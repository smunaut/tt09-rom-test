magic
tech sky130A
magscale 1 2
timestamp 1730749471
<< nwell >>
rect 27265 4520 27773 22220
<< locali >>
rect 27111 22140 27145 22156
rect 27111 22090 27145 22106
rect 27111 22000 27145 22016
rect 27111 21950 27145 21966
rect 27111 21860 27145 21876
rect 27111 21810 27145 21826
rect 27111 21720 27145 21736
rect 27111 21670 27145 21686
rect 27111 21580 27145 21596
rect 27111 21530 27145 21546
rect 27111 21440 27145 21456
rect 27111 21390 27145 21406
rect 27111 21300 27145 21316
rect 27111 21250 27145 21266
rect 27111 21160 27145 21176
rect 27111 21110 27145 21126
rect 27111 20930 27145 20946
rect 27111 20880 27145 20896
rect 27111 20790 27145 20806
rect 27111 20740 27145 20756
rect 27111 20650 27145 20666
rect 27111 20600 27145 20616
rect 27111 20510 27145 20526
rect 27111 20460 27145 20476
rect 27111 20370 27145 20386
rect 27111 20320 27145 20336
rect 27111 20230 27145 20246
rect 27111 20180 27145 20196
rect 27111 20090 27145 20106
rect 27111 20040 27145 20056
rect 27111 19950 27145 19966
rect 27111 19900 27145 19916
rect 27111 19720 27145 19736
rect 27111 19670 27145 19686
rect 27111 19580 27145 19596
rect 27111 19530 27145 19546
rect 27111 19440 27145 19456
rect 27111 19390 27145 19406
rect 27111 19300 27145 19316
rect 27111 19250 27145 19266
rect 27111 19160 27145 19176
rect 27111 19110 27145 19126
rect 27111 19020 27145 19036
rect 27111 18970 27145 18986
rect 27111 18880 27145 18896
rect 27111 18830 27145 18846
rect 27111 18740 27145 18756
rect 27111 18690 27145 18706
rect 27111 18510 27145 18526
rect 27111 18460 27145 18476
rect 27111 18370 27145 18386
rect 27111 18320 27145 18336
rect 27111 18230 27145 18246
rect 27111 18180 27145 18196
rect 27111 18090 27145 18106
rect 27111 18040 27145 18056
rect 27111 17950 27145 17966
rect 27111 17900 27145 17916
rect 27111 17810 27145 17826
rect 27111 17760 27145 17776
rect 27111 17670 27145 17686
rect 27111 17620 27145 17636
rect 27111 17530 27145 17546
rect 27111 17480 27145 17496
rect 27111 17160 27145 17176
rect 27111 17110 27145 17126
rect 27111 17020 27145 17036
rect 27111 16970 27145 16986
rect 27111 16880 27145 16896
rect 27111 16830 27145 16846
rect 27111 16740 27145 16756
rect 27111 16690 27145 16706
rect 27111 16600 27145 16616
rect 27111 16550 27145 16566
rect 27111 16460 27145 16476
rect 27111 16410 27145 16426
rect 27111 16320 27145 16336
rect 27111 16270 27145 16286
rect 27111 16180 27145 16196
rect 27111 16130 27145 16146
rect 27111 15950 27145 15966
rect 27111 15900 27145 15916
rect 27111 15810 27145 15826
rect 27111 15760 27145 15776
rect 27111 15670 27145 15686
rect 27111 15620 27145 15636
rect 27111 15530 27145 15546
rect 27111 15480 27145 15496
rect 27111 15390 27145 15406
rect 27111 15340 27145 15356
rect 27111 15250 27145 15266
rect 27111 15200 27145 15216
rect 27111 15110 27145 15126
rect 27111 15060 27145 15076
rect 27111 14970 27145 14986
rect 27111 14920 27145 14936
rect 27111 14740 27145 14756
rect 27111 14690 27145 14706
rect 27111 14600 27145 14616
rect 27111 14550 27145 14566
rect 27111 14460 27145 14476
rect 27111 14410 27145 14426
rect 27111 14320 27145 14336
rect 27111 14270 27145 14286
rect 27111 14180 27145 14196
rect 27111 14130 27145 14146
rect 27111 14040 27145 14056
rect 27111 13990 27145 14006
rect 27111 13900 27145 13916
rect 27111 13850 27145 13866
rect 27111 13760 27145 13776
rect 27111 13710 27145 13726
rect 27111 13530 27145 13546
rect 27111 13480 27145 13496
rect 27111 13390 27145 13406
rect 27111 13340 27145 13356
rect 27111 13250 27145 13266
rect 27111 13200 27145 13216
rect 27111 13110 27145 13126
rect 27111 13060 27145 13076
rect 27111 12970 27145 12986
rect 27111 12920 27145 12936
rect 27111 12830 27145 12846
rect 27111 12780 27145 12796
rect 27111 12690 27145 12706
rect 27111 12640 27145 12656
rect 27111 12550 27145 12566
rect 27111 12500 27145 12516
rect 27111 12180 27145 12196
rect 27111 12130 27145 12146
rect 27111 12040 27145 12056
rect 27111 11990 27145 12006
rect 27111 11900 27145 11916
rect 27111 11850 27145 11866
rect 27111 11760 27145 11776
rect 27111 11710 27145 11726
rect 27111 11620 27145 11636
rect 27111 11570 27145 11586
rect 27111 11480 27145 11496
rect 27111 11430 27145 11446
rect 27111 11340 27145 11356
rect 27111 11290 27145 11306
rect 27111 11200 27145 11216
rect 27111 11150 27145 11166
rect 27111 10970 27145 10986
rect 27111 10920 27145 10936
rect 27111 10830 27145 10846
rect 27111 10780 27145 10796
rect 27111 10690 27145 10706
rect 27111 10640 27145 10656
rect 27111 10550 27145 10566
rect 27111 10500 27145 10516
rect 27111 10410 27145 10426
rect 27111 10360 27145 10376
rect 27111 10270 27145 10286
rect 27111 10220 27145 10236
rect 27111 10130 27145 10146
rect 27111 10080 27145 10096
rect 27111 9990 27145 10006
rect 27111 9940 27145 9956
rect 27111 9760 27145 9776
rect 27111 9710 27145 9726
rect 27111 9620 27145 9636
rect 27111 9570 27145 9586
rect 27111 9480 27145 9496
rect 27111 9430 27145 9446
rect 27111 9340 27145 9356
rect 27111 9290 27145 9306
rect 27111 9200 27145 9216
rect 27111 9150 27145 9166
rect 27111 9060 27145 9076
rect 27111 9010 27145 9026
rect 27111 8920 27145 8936
rect 27111 8870 27145 8886
rect 27111 8780 27145 8796
rect 27111 8730 27145 8746
rect 27111 8550 27145 8566
rect 27111 8500 27145 8516
rect 27111 8410 27145 8426
rect 27111 8360 27145 8376
rect 27111 8270 27145 8286
rect 27111 8220 27145 8236
rect 27111 8130 27145 8146
rect 27111 8080 27145 8096
rect 27111 7990 27145 8006
rect 27111 7940 27145 7956
rect 27111 7850 27145 7866
rect 27111 7800 27145 7816
rect 27111 7710 27145 7726
rect 27111 7660 27145 7676
rect 27111 7570 27145 7586
rect 27111 7520 27145 7536
rect 27111 7200 27145 7216
rect 27111 7150 27145 7166
rect 27111 7060 27145 7076
rect 27111 7010 27145 7026
rect 27111 6920 27145 6936
rect 27111 6870 27145 6886
rect 27111 6780 27145 6796
rect 27111 6730 27145 6746
rect 27111 6640 27145 6656
rect 27111 6590 27145 6606
rect 27111 6500 27145 6516
rect 27111 6450 27145 6466
rect 27111 6360 27145 6376
rect 27111 6310 27145 6326
rect 27111 6220 27145 6236
rect 27111 6170 27145 6186
rect 27111 5990 27145 6006
rect 27111 5940 27145 5956
rect 27111 5850 27145 5866
rect 27111 5800 27145 5816
rect 27111 5710 27145 5726
rect 27111 5660 27145 5676
rect 27111 5570 27145 5586
rect 27111 5520 27145 5536
rect 27111 5430 27145 5446
rect 27111 5380 27145 5396
rect 27111 5290 27145 5306
rect 27111 5240 27145 5256
rect 27111 5150 27145 5166
rect 27111 5100 27145 5116
rect 27111 5010 27145 5026
rect 27111 4960 27145 4976
rect 27111 4780 27145 4796
rect 27111 4730 27145 4746
rect 27111 4640 27145 4656
rect 27111 4590 27145 4606
rect 27111 4500 27145 4516
rect 27111 4450 27145 4466
rect 27111 4360 27145 4376
rect 27111 4310 27145 4326
rect 27111 4220 27145 4236
rect 27111 4170 27145 4186
rect 27111 4080 27145 4096
rect 27111 4030 27145 4046
rect 27111 3940 27145 3956
rect 27111 3890 27145 3906
rect 27111 3800 27145 3816
rect 27111 3750 27145 3766
rect 27111 3570 27145 3586
rect 27111 3520 27145 3536
rect 27111 3430 27145 3446
rect 27111 3380 27145 3396
rect 27111 3290 27145 3306
rect 27111 3240 27145 3256
rect 27111 3150 27145 3166
rect 27111 3100 27145 3116
rect 27111 3010 27145 3026
rect 27111 2960 27145 2976
rect 27111 2870 27145 2886
rect 27111 2820 27145 2836
rect 27111 2730 27145 2746
rect 27111 2680 27145 2696
rect 27111 2590 27145 2606
rect 27111 2540 27145 2556
<< viali >>
rect 27111 22106 27145 22140
rect 27111 21966 27145 22000
rect 27111 21826 27145 21860
rect 27111 21686 27145 21720
rect 27111 21546 27145 21580
rect 27111 21406 27145 21440
rect 27111 21266 27145 21300
rect 27111 21126 27145 21160
rect 27111 20896 27145 20930
rect 27111 20756 27145 20790
rect 27111 20616 27145 20650
rect 27111 20476 27145 20510
rect 27111 20336 27145 20370
rect 27111 20196 27145 20230
rect 27111 20056 27145 20090
rect 27111 19916 27145 19950
rect 27111 19686 27145 19720
rect 27111 19546 27145 19580
rect 27111 19406 27145 19440
rect 27111 19266 27145 19300
rect 27111 19126 27145 19160
rect 27111 18986 27145 19020
rect 27111 18846 27145 18880
rect 27111 18706 27145 18740
rect 27111 18476 27145 18510
rect 27111 18336 27145 18370
rect 27111 18196 27145 18230
rect 27111 18056 27145 18090
rect 27111 17916 27145 17950
rect 27111 17776 27145 17810
rect 27111 17636 27145 17670
rect 27111 17496 27145 17530
rect 27111 17126 27145 17160
rect 27111 16986 27145 17020
rect 27111 16846 27145 16880
rect 27111 16706 27145 16740
rect 27111 16566 27145 16600
rect 27111 16426 27145 16460
rect 27111 16286 27145 16320
rect 27111 16146 27145 16180
rect 27111 15916 27145 15950
rect 27111 15776 27145 15810
rect 27111 15636 27145 15670
rect 27111 15496 27145 15530
rect 27111 15356 27145 15390
rect 27111 15216 27145 15250
rect 27111 15076 27145 15110
rect 27111 14936 27145 14970
rect 27111 14706 27145 14740
rect 27111 14566 27145 14600
rect 27111 14426 27145 14460
rect 27111 14286 27145 14320
rect 27111 14146 27145 14180
rect 27111 14006 27145 14040
rect 27111 13866 27145 13900
rect 27111 13726 27145 13760
rect 27111 13496 27145 13530
rect 27111 13356 27145 13390
rect 27111 13216 27145 13250
rect 27111 13076 27145 13110
rect 27111 12936 27145 12970
rect 27111 12796 27145 12830
rect 27111 12656 27145 12690
rect 27111 12516 27145 12550
rect 27111 12146 27145 12180
rect 27111 12006 27145 12040
rect 27111 11866 27145 11900
rect 27111 11726 27145 11760
rect 27111 11586 27145 11620
rect 27111 11446 27145 11480
rect 27111 11306 27145 11340
rect 27111 11166 27145 11200
rect 27111 10936 27145 10970
rect 27111 10796 27145 10830
rect 27111 10656 27145 10690
rect 27111 10516 27145 10550
rect 27111 10376 27145 10410
rect 27111 10236 27145 10270
rect 27111 10096 27145 10130
rect 27111 9956 27145 9990
rect 27111 9726 27145 9760
rect 27111 9586 27145 9620
rect 27111 9446 27145 9480
rect 27111 9306 27145 9340
rect 27111 9166 27145 9200
rect 27111 9026 27145 9060
rect 27111 8886 27145 8920
rect 27111 8746 27145 8780
rect 27111 8516 27145 8550
rect 27111 8376 27145 8410
rect 27111 8236 27145 8270
rect 27111 8096 27145 8130
rect 27111 7956 27145 7990
rect 27111 7816 27145 7850
rect 27111 7676 27145 7710
rect 27111 7536 27145 7570
rect 27111 7166 27145 7200
rect 27111 7026 27145 7060
rect 27111 6886 27145 6920
rect 27111 6746 27145 6780
rect 27111 6606 27145 6640
rect 27111 6466 27145 6500
rect 27111 6326 27145 6360
rect 27111 6186 27145 6220
rect 27111 5956 27145 5990
rect 27111 5816 27145 5850
rect 27111 5676 27145 5710
rect 27111 5536 27145 5570
rect 27111 5396 27145 5430
rect 27111 5256 27145 5290
rect 27111 5116 27145 5150
rect 27111 4976 27145 5010
rect 27111 4746 27145 4780
rect 27111 4606 27145 4640
rect 27111 4466 27145 4500
rect 27111 4326 27145 4360
rect 27111 4186 27145 4220
rect 27111 4046 27145 4080
rect 27111 3906 27145 3940
rect 27111 3766 27145 3800
rect 27111 3536 27145 3570
rect 27111 3396 27145 3430
rect 27111 3256 27145 3290
rect 27111 3116 27145 3150
rect 27111 2976 27145 3010
rect 27111 2836 27145 2870
rect 27111 2696 27145 2730
rect 27111 2556 27145 2590
<< metal1 >>
rect 27111 22155 27145 22163
rect 27102 22149 27154 22155
rect 27102 22091 27154 22097
rect 27111 22012 27145 22091
rect 27105 22000 27151 22012
rect 27105 21966 27111 22000
rect 27145 21966 27151 22000
rect 27105 21954 27151 21966
rect 27111 21872 27145 21954
rect 27105 21860 27151 21872
rect 27105 21826 27111 21860
rect 27145 21826 27151 21860
rect 27105 21814 27151 21826
rect 27111 21732 27145 21814
rect 27105 21720 27151 21732
rect 27105 21686 27111 21720
rect 27145 21686 27151 21720
rect 27105 21674 27151 21686
rect 27111 21592 27145 21674
rect 27105 21580 27151 21592
rect 27105 21546 27111 21580
rect 27145 21546 27151 21580
rect 27105 21534 27151 21546
rect 27111 21452 27145 21534
rect 27105 21440 27151 21452
rect 27105 21406 27111 21440
rect 27145 21406 27151 21440
rect 27105 21394 27151 21406
rect 27111 21312 27145 21394
rect 27105 21300 27151 21312
rect 27105 21266 27111 21300
rect 27145 21266 27151 21300
rect 27105 21254 27151 21266
rect 27111 21172 27145 21254
rect 27105 21160 27151 21172
rect 27105 21126 27111 21160
rect 27145 21126 27151 21160
rect 27105 21114 27151 21126
rect 27111 20942 27145 21114
rect 27105 20930 27151 20942
rect 27105 20896 27111 20930
rect 27145 20896 27151 20930
rect 27105 20884 27151 20896
rect 27111 20802 27145 20884
rect 27105 20790 27151 20802
rect 27105 20756 27111 20790
rect 27145 20756 27151 20790
rect 27105 20744 27151 20756
rect 27111 20662 27145 20744
rect 27105 20650 27151 20662
rect 27105 20616 27111 20650
rect 27145 20616 27151 20650
rect 27105 20604 27151 20616
rect 27111 20522 27145 20604
rect 27105 20510 27151 20522
rect 27105 20476 27111 20510
rect 27145 20476 27151 20510
rect 27105 20464 27151 20476
rect 27111 20382 27145 20464
rect 27105 20370 27151 20382
rect 27105 20336 27111 20370
rect 27145 20336 27151 20370
rect 27105 20324 27151 20336
rect 27111 20242 27145 20324
rect 27105 20230 27151 20242
rect 27105 20196 27111 20230
rect 27145 20196 27151 20230
rect 27105 20184 27151 20196
rect 27111 20102 27145 20184
rect 27105 20090 27151 20102
rect 27105 20056 27111 20090
rect 27145 20056 27151 20090
rect 27105 20044 27151 20056
rect 27111 19962 27145 20044
rect 27105 19950 27151 19962
rect 27105 19916 27111 19950
rect 27145 19916 27151 19950
rect 27105 19904 27151 19916
rect 27111 19894 27145 19904
rect 27111 19735 27145 19743
rect 27102 19729 27154 19735
rect 27102 19671 27154 19677
rect 27111 19592 27145 19671
rect 27105 19580 27151 19592
rect 27105 19546 27111 19580
rect 27145 19546 27151 19580
rect 27105 19534 27151 19546
rect 27111 19452 27145 19534
rect 27105 19440 27151 19452
rect 27105 19406 27111 19440
rect 27145 19406 27151 19440
rect 27105 19394 27151 19406
rect 27111 19312 27145 19394
rect 27105 19300 27151 19312
rect 27105 19266 27111 19300
rect 27145 19266 27151 19300
rect 27105 19254 27151 19266
rect 27111 19172 27145 19254
rect 27105 19160 27151 19172
rect 27105 19126 27111 19160
rect 27145 19126 27151 19160
rect 27105 19114 27151 19126
rect 27111 19032 27145 19114
rect 27105 19020 27151 19032
rect 27105 18986 27111 19020
rect 27145 18986 27151 19020
rect 27105 18974 27151 18986
rect 27111 18892 27145 18974
rect 27105 18880 27151 18892
rect 27105 18846 27111 18880
rect 27145 18846 27151 18880
rect 27105 18834 27151 18846
rect 27111 18752 27145 18834
rect 27105 18740 27151 18752
rect 27105 18706 27111 18740
rect 27145 18706 27151 18740
rect 27105 18694 27151 18706
rect 27111 18522 27145 18694
rect 27105 18510 27151 18522
rect 27105 18476 27111 18510
rect 27145 18476 27151 18510
rect 27105 18464 27151 18476
rect 27111 18382 27145 18464
rect 27105 18370 27151 18382
rect 27105 18336 27111 18370
rect 27145 18336 27151 18370
rect 27105 18324 27151 18336
rect 27111 18242 27145 18324
rect 27105 18230 27151 18242
rect 27105 18196 27111 18230
rect 27145 18196 27151 18230
rect 27105 18184 27151 18196
rect 27111 18102 27145 18184
rect 27105 18090 27151 18102
rect 27105 18056 27111 18090
rect 27145 18056 27151 18090
rect 27105 18044 27151 18056
rect 27111 17962 27145 18044
rect 27105 17950 27151 17962
rect 27105 17916 27111 17950
rect 27145 17916 27151 17950
rect 27105 17904 27151 17916
rect 27111 17822 27145 17904
rect 27105 17810 27151 17822
rect 27105 17776 27111 17810
rect 27145 17776 27151 17810
rect 27105 17764 27151 17776
rect 27111 17682 27145 17764
rect 27105 17670 27151 17682
rect 27105 17636 27111 17670
rect 27145 17636 27151 17670
rect 27105 17624 27151 17636
rect 27111 17542 27145 17624
rect 27105 17530 27151 17542
rect 27105 17496 27111 17530
rect 27145 17496 27151 17530
rect 27105 17484 27151 17496
rect 27111 17474 27145 17484
rect 27111 17175 27145 17183
rect 27102 17169 27154 17175
rect 27102 17111 27154 17117
rect 27111 17032 27145 17111
rect 27105 17020 27151 17032
rect 27105 16986 27111 17020
rect 27145 16986 27151 17020
rect 27105 16974 27151 16986
rect 27111 16892 27145 16974
rect 27105 16880 27151 16892
rect 27105 16846 27111 16880
rect 27145 16846 27151 16880
rect 27105 16834 27151 16846
rect 27111 16752 27145 16834
rect 27105 16740 27151 16752
rect 27105 16706 27111 16740
rect 27145 16706 27151 16740
rect 27105 16694 27151 16706
rect 27111 16612 27145 16694
rect 27105 16600 27151 16612
rect 27105 16566 27111 16600
rect 27145 16566 27151 16600
rect 27105 16554 27151 16566
rect 27111 16472 27145 16554
rect 27105 16460 27151 16472
rect 27105 16426 27111 16460
rect 27145 16426 27151 16460
rect 27105 16414 27151 16426
rect 27111 16332 27145 16414
rect 27105 16320 27151 16332
rect 27105 16286 27111 16320
rect 27145 16286 27151 16320
rect 27105 16274 27151 16286
rect 27111 16192 27145 16274
rect 27105 16180 27151 16192
rect 27105 16146 27111 16180
rect 27145 16146 27151 16180
rect 27105 16134 27151 16146
rect 27111 15962 27145 16134
rect 27105 15950 27151 15962
rect 27105 15916 27111 15950
rect 27145 15916 27151 15950
rect 27105 15904 27151 15916
rect 27111 15822 27145 15904
rect 27105 15810 27151 15822
rect 27105 15776 27111 15810
rect 27145 15776 27151 15810
rect 27105 15764 27151 15776
rect 27111 15682 27145 15764
rect 27105 15670 27151 15682
rect 27105 15636 27111 15670
rect 27145 15636 27151 15670
rect 27105 15624 27151 15636
rect 27111 15542 27145 15624
rect 27105 15530 27151 15542
rect 27105 15496 27111 15530
rect 27145 15496 27151 15530
rect 27105 15484 27151 15496
rect 27111 15402 27145 15484
rect 27105 15390 27151 15402
rect 27105 15356 27111 15390
rect 27145 15356 27151 15390
rect 27105 15344 27151 15356
rect 27111 15262 27145 15344
rect 27105 15250 27151 15262
rect 27105 15216 27111 15250
rect 27145 15216 27151 15250
rect 27105 15204 27151 15216
rect 27111 15122 27145 15204
rect 27105 15110 27151 15122
rect 27105 15076 27111 15110
rect 27145 15076 27151 15110
rect 27105 15064 27151 15076
rect 27111 14982 27145 15064
rect 27105 14970 27151 14982
rect 27105 14936 27111 14970
rect 27145 14936 27151 14970
rect 27105 14924 27151 14936
rect 27111 14914 27145 14924
rect 27111 14755 27145 14763
rect 27102 14749 27154 14755
rect 27102 14691 27154 14697
rect 27111 14612 27145 14691
rect 27105 14600 27151 14612
rect 27105 14566 27111 14600
rect 27145 14566 27151 14600
rect 27105 14554 27151 14566
rect 27111 14472 27145 14554
rect 27105 14460 27151 14472
rect 27105 14426 27111 14460
rect 27145 14426 27151 14460
rect 27105 14414 27151 14426
rect 27111 14332 27145 14414
rect 27105 14320 27151 14332
rect 27105 14286 27111 14320
rect 27145 14286 27151 14320
rect 27105 14274 27151 14286
rect 27111 14192 27145 14274
rect 27105 14180 27151 14192
rect 27105 14146 27111 14180
rect 27145 14146 27151 14180
rect 27105 14134 27151 14146
rect 27111 14052 27145 14134
rect 27105 14040 27151 14052
rect 27105 14006 27111 14040
rect 27145 14006 27151 14040
rect 27105 13994 27151 14006
rect 27111 13912 27145 13994
rect 27105 13900 27151 13912
rect 27105 13866 27111 13900
rect 27145 13866 27151 13900
rect 27105 13854 27151 13866
rect 27111 13772 27145 13854
rect 27105 13760 27151 13772
rect 27105 13726 27111 13760
rect 27145 13726 27151 13760
rect 27105 13714 27151 13726
rect 27111 13542 27145 13714
rect 27105 13530 27151 13542
rect 27105 13496 27111 13530
rect 27145 13496 27151 13530
rect 27105 13484 27151 13496
rect 27111 13402 27145 13484
rect 27105 13390 27151 13402
rect 27105 13356 27111 13390
rect 27145 13356 27151 13390
rect 27105 13344 27151 13356
rect 27111 13262 27145 13344
rect 27105 13250 27151 13262
rect 27105 13216 27111 13250
rect 27145 13216 27151 13250
rect 27105 13204 27151 13216
rect 27111 13122 27145 13204
rect 27105 13110 27151 13122
rect 27105 13076 27111 13110
rect 27145 13076 27151 13110
rect 27105 13064 27151 13076
rect 27111 12982 27145 13064
rect 27105 12970 27151 12982
rect 27105 12936 27111 12970
rect 27145 12936 27151 12970
rect 27105 12924 27151 12936
rect 27111 12842 27145 12924
rect 27105 12830 27151 12842
rect 27105 12796 27111 12830
rect 27145 12796 27151 12830
rect 27105 12784 27151 12796
rect 27111 12702 27145 12784
rect 27105 12690 27151 12702
rect 27105 12656 27111 12690
rect 27145 12656 27151 12690
rect 27105 12644 27151 12656
rect 27111 12562 27145 12644
rect 27105 12550 27151 12562
rect 27105 12516 27111 12550
rect 27145 12516 27151 12550
rect 27105 12504 27151 12516
rect 27111 12494 27145 12504
rect 27111 12195 27145 12203
rect 27102 12189 27154 12195
rect 27102 12131 27154 12137
rect 27111 12052 27145 12131
rect 27105 12040 27151 12052
rect 27105 12006 27111 12040
rect 27145 12006 27151 12040
rect 27105 11994 27151 12006
rect 27111 11912 27145 11994
rect 27105 11900 27151 11912
rect 27105 11866 27111 11900
rect 27145 11866 27151 11900
rect 27105 11854 27151 11866
rect 27111 11772 27145 11854
rect 27105 11760 27151 11772
rect 27105 11726 27111 11760
rect 27145 11726 27151 11760
rect 27105 11714 27151 11726
rect 27111 11632 27145 11714
rect 27105 11620 27151 11632
rect 27105 11586 27111 11620
rect 27145 11586 27151 11620
rect 27105 11574 27151 11586
rect 27111 11492 27145 11574
rect 27105 11480 27151 11492
rect 27105 11446 27111 11480
rect 27145 11446 27151 11480
rect 27105 11434 27151 11446
rect 27111 11352 27145 11434
rect 27105 11340 27151 11352
rect 27105 11306 27111 11340
rect 27145 11306 27151 11340
rect 27105 11294 27151 11306
rect 27111 11212 27145 11294
rect 27105 11200 27151 11212
rect 27105 11166 27111 11200
rect 27145 11166 27151 11200
rect 27105 11154 27151 11166
rect 27111 10982 27145 11154
rect 27105 10970 27151 10982
rect 27105 10936 27111 10970
rect 27145 10936 27151 10970
rect 27105 10924 27151 10936
rect 27111 10842 27145 10924
rect 27105 10830 27151 10842
rect 27105 10796 27111 10830
rect 27145 10796 27151 10830
rect 27105 10784 27151 10796
rect 27111 10702 27145 10784
rect 27105 10690 27151 10702
rect 27105 10656 27111 10690
rect 27145 10656 27151 10690
rect 27105 10644 27151 10656
rect 27111 10562 27145 10644
rect 27105 10550 27151 10562
rect 27105 10516 27111 10550
rect 27145 10516 27151 10550
rect 27105 10504 27151 10516
rect 27111 10422 27145 10504
rect 27105 10410 27151 10422
rect 27105 10376 27111 10410
rect 27145 10376 27151 10410
rect 27105 10364 27151 10376
rect 27111 10282 27145 10364
rect 27105 10270 27151 10282
rect 27105 10236 27111 10270
rect 27145 10236 27151 10270
rect 27105 10224 27151 10236
rect 27111 10142 27145 10224
rect 27105 10130 27151 10142
rect 27105 10096 27111 10130
rect 27145 10096 27151 10130
rect 27105 10084 27151 10096
rect 27111 10002 27145 10084
rect 27105 9990 27151 10002
rect 27105 9956 27111 9990
rect 27145 9956 27151 9990
rect 27105 9944 27151 9956
rect 27111 9934 27145 9944
rect 27111 9775 27145 9783
rect 27102 9769 27154 9775
rect 27102 9711 27154 9717
rect 27111 9632 27145 9711
rect 27105 9620 27151 9632
rect 27105 9586 27111 9620
rect 27145 9586 27151 9620
rect 27105 9574 27151 9586
rect 27111 9492 27145 9574
rect 27105 9480 27151 9492
rect 27105 9446 27111 9480
rect 27145 9446 27151 9480
rect 27105 9434 27151 9446
rect 27111 9352 27145 9434
rect 27105 9340 27151 9352
rect 27105 9306 27111 9340
rect 27145 9306 27151 9340
rect 27105 9294 27151 9306
rect 27111 9212 27145 9294
rect 27105 9200 27151 9212
rect 27105 9166 27111 9200
rect 27145 9166 27151 9200
rect 27105 9154 27151 9166
rect 27111 9072 27145 9154
rect 27105 9060 27151 9072
rect 27105 9026 27111 9060
rect 27145 9026 27151 9060
rect 27105 9014 27151 9026
rect 27111 8932 27145 9014
rect 27105 8920 27151 8932
rect 27105 8886 27111 8920
rect 27145 8886 27151 8920
rect 27105 8874 27151 8886
rect 27111 8792 27145 8874
rect 27105 8780 27151 8792
rect 27105 8746 27111 8780
rect 27145 8746 27151 8780
rect 27105 8734 27151 8746
rect 27111 8562 27145 8734
rect 27105 8550 27151 8562
rect 27105 8516 27111 8550
rect 27145 8516 27151 8550
rect 27105 8504 27151 8516
rect 27111 8422 27145 8504
rect 27105 8410 27151 8422
rect 27105 8376 27111 8410
rect 27145 8376 27151 8410
rect 27105 8364 27151 8376
rect 27111 8282 27145 8364
rect 27105 8270 27151 8282
rect 27105 8236 27111 8270
rect 27145 8236 27151 8270
rect 27105 8224 27151 8236
rect 27111 8142 27145 8224
rect 27105 8130 27151 8142
rect 27105 8096 27111 8130
rect 27145 8096 27151 8130
rect 27105 8084 27151 8096
rect 27111 8002 27145 8084
rect 27105 7990 27151 8002
rect 27105 7956 27111 7990
rect 27145 7956 27151 7990
rect 27105 7944 27151 7956
rect 27111 7862 27145 7944
rect 27105 7850 27151 7862
rect 27105 7816 27111 7850
rect 27145 7816 27151 7850
rect 27105 7804 27151 7816
rect 27111 7722 27145 7804
rect 27105 7710 27151 7722
rect 27105 7676 27111 7710
rect 27145 7676 27151 7710
rect 27105 7664 27151 7676
rect 27111 7582 27145 7664
rect 27105 7570 27151 7582
rect 27105 7536 27111 7570
rect 27145 7536 27151 7570
rect 27105 7524 27151 7536
rect 27111 7514 27145 7524
rect 27111 7215 27145 7223
rect 27102 7209 27154 7215
rect 27102 7151 27154 7157
rect 27111 7072 27145 7151
rect 27105 7060 27151 7072
rect 27105 7026 27111 7060
rect 27145 7026 27151 7060
rect 27105 7014 27151 7026
rect 27111 6932 27145 7014
rect 27105 6920 27151 6932
rect 27105 6886 27111 6920
rect 27145 6886 27151 6920
rect 27105 6874 27151 6886
rect 27111 6792 27145 6874
rect 27105 6780 27151 6792
rect 27105 6746 27111 6780
rect 27145 6746 27151 6780
rect 27105 6734 27151 6746
rect 27111 6652 27145 6734
rect 27105 6640 27151 6652
rect 27105 6606 27111 6640
rect 27145 6606 27151 6640
rect 27105 6594 27151 6606
rect 27111 6512 27145 6594
rect 27105 6500 27151 6512
rect 27105 6466 27111 6500
rect 27145 6466 27151 6500
rect 27105 6454 27151 6466
rect 27111 6372 27145 6454
rect 27105 6360 27151 6372
rect 27105 6326 27111 6360
rect 27145 6326 27151 6360
rect 27105 6314 27151 6326
rect 27111 6232 27145 6314
rect 27105 6220 27151 6232
rect 27105 6186 27111 6220
rect 27145 6186 27151 6220
rect 27105 6174 27151 6186
rect 27111 6002 27145 6174
rect 27105 5990 27151 6002
rect 27105 5956 27111 5990
rect 27145 5956 27151 5990
rect 27105 5944 27151 5956
rect 27111 5862 27145 5944
rect 27105 5850 27151 5862
rect 27105 5816 27111 5850
rect 27145 5816 27151 5850
rect 27105 5804 27151 5816
rect 27111 5722 27145 5804
rect 27105 5710 27151 5722
rect 27105 5676 27111 5710
rect 27145 5676 27151 5710
rect 27105 5664 27151 5676
rect 27111 5582 27145 5664
rect 27105 5570 27151 5582
rect 27105 5536 27111 5570
rect 27145 5536 27151 5570
rect 27105 5524 27151 5536
rect 27111 5442 27145 5524
rect 27105 5430 27151 5442
rect 27105 5396 27111 5430
rect 27145 5396 27151 5430
rect 27105 5384 27151 5396
rect 27111 5302 27145 5384
rect 27105 5290 27151 5302
rect 27105 5256 27111 5290
rect 27145 5256 27151 5290
rect 27105 5244 27151 5256
rect 27111 5162 27145 5244
rect 27105 5150 27151 5162
rect 27105 5116 27111 5150
rect 27145 5116 27151 5150
rect 27105 5104 27151 5116
rect 27111 5022 27145 5104
rect 27105 5010 27151 5022
rect 27105 4976 27111 5010
rect 27145 4976 27151 5010
rect 27105 4964 27151 4976
rect 27111 4954 27145 4964
rect 27111 4795 27145 4803
rect 27102 4789 27154 4795
rect 27102 4731 27154 4737
rect 27111 4652 27145 4731
rect 27105 4640 27151 4652
rect 27105 4606 27111 4640
rect 27145 4606 27151 4640
rect 27105 4594 27151 4606
rect 27111 4512 27145 4594
rect 27220 4553 27254 22193
rect 28000 22027 28006 22079
rect 28074 22027 28080 22079
rect 28000 19607 28006 19659
rect 28074 19607 28080 19659
rect 28000 17047 28006 17099
rect 28074 17047 28080 17099
rect 28000 14627 28006 14679
rect 28074 14627 28080 14679
rect 28000 12067 28006 12119
rect 28074 12067 28080 12119
rect 28000 9647 28006 9699
rect 28074 9647 28080 9699
rect 28000 7087 28006 7139
rect 28074 7087 28080 7139
rect 28000 4667 28006 4719
rect 28074 4667 28080 4719
rect 27105 4500 27151 4512
rect 27105 4466 27111 4500
rect 27145 4466 27151 4500
rect 27105 4454 27151 4466
rect 27111 4372 27145 4454
rect 27105 4360 27151 4372
rect 27105 4326 27111 4360
rect 27145 4326 27151 4360
rect 27105 4314 27151 4326
rect 27111 4232 27145 4314
rect 27105 4220 27151 4232
rect 27105 4186 27111 4220
rect 27145 4186 27151 4220
rect 27105 4174 27151 4186
rect 27111 4092 27145 4174
rect 27105 4080 27151 4092
rect 27105 4046 27111 4080
rect 27145 4046 27151 4080
rect 27105 4034 27151 4046
rect 27111 3952 27145 4034
rect 27105 3940 27151 3952
rect 27105 3906 27111 3940
rect 27145 3906 27151 3940
rect 27105 3894 27151 3906
rect 27111 3812 27145 3894
rect 27105 3800 27151 3812
rect 27105 3766 27111 3800
rect 27145 3766 27151 3800
rect 27105 3754 27151 3766
rect 27111 3582 27145 3754
rect 27105 3570 27151 3582
rect 27105 3536 27111 3570
rect 27145 3536 27151 3570
rect 27105 3524 27151 3536
rect 27111 3442 27145 3524
rect 27105 3430 27151 3442
rect 27105 3396 27111 3430
rect 27145 3396 27151 3430
rect 27105 3384 27151 3396
rect 27111 3302 27145 3384
rect 27105 3290 27151 3302
rect 27105 3256 27111 3290
rect 27145 3256 27151 3290
rect 27105 3244 27151 3256
rect 27111 3162 27145 3244
rect 27105 3150 27151 3162
rect 27105 3116 27111 3150
rect 27145 3116 27151 3150
rect 27105 3104 27151 3116
rect 27111 3022 27145 3104
rect 27105 3010 27151 3022
rect 27105 2976 27111 3010
rect 27145 2976 27151 3010
rect 27105 2964 27151 2976
rect 27111 2882 27145 2964
rect 27105 2870 27151 2882
rect 27105 2836 27111 2870
rect 27145 2836 27151 2870
rect 27105 2824 27151 2836
rect 27111 2742 27145 2824
rect 27105 2730 27151 2742
rect 27105 2696 27111 2730
rect 27145 2696 27151 2730
rect 27105 2684 27151 2696
rect 27111 2602 27145 2684
rect 27105 2590 27151 2602
rect 27105 2556 27111 2590
rect 27145 2556 27151 2590
rect 27105 2544 27151 2556
rect 27111 2534 27145 2544
rect 27270 2473 27449 2503
rect 41 2203 157 2233
rect 25811 2203 25927 2233
rect 41 1781 71 2203
rect 25897 1781 25927 2203
rect 41 1751 101 1781
rect 25867 1751 25927 1781
rect 26039 1603 26069 2413
rect 26099 1703 26129 2413
rect 26329 1803 26359 2413
rect 26429 1903 26459 2413
rect 26529 2003 26559 2413
rect 26629 2103 26659 2413
rect 26729 2203 26759 2413
rect 26829 2287 26859 2413
rect 26929 2347 26959 2413
rect 27029 2407 27059 2413
rect 27270 2407 27300 2473
rect 27029 2377 27300 2407
rect 27330 2373 27449 2403
rect 27330 2347 27360 2373
rect 26929 2317 27360 2347
rect 27390 2287 27449 2303
rect 26829 2273 27449 2287
rect 26829 2257 27420 2273
rect 26729 2173 27449 2203
rect 26629 2073 27449 2103
rect 26529 1973 27449 2003
rect 26429 1873 27449 1903
rect 26329 1773 27449 1803
rect 26099 1673 27449 1703
rect 26039 1573 27449 1603
rect 25825 1473 27449 1503
rect 25825 1373 27449 1403
rect 25825 1273 27449 1303
rect 25825 1173 27449 1203
rect 25825 1073 27449 1103
rect 25825 973 27449 1003
rect 25825 873 27449 903
rect 25825 773 27449 803
rect 25825 673 27449 703
rect 25825 573 27449 603
rect 25825 473 27449 503
rect 25825 373 27449 403
rect 25825 273 27449 303
rect 25825 173 27449 203
rect 11 90 211 96
rect 11 32 17 90
rect 205 32 211 90
rect 11 26 211 32
rect 25757 90 25957 96
rect 25757 32 25763 90
rect 25951 32 25957 90
rect 25757 26 25957 32
<< via1 >>
rect 27102 22140 27154 22149
rect 27102 22106 27111 22140
rect 27111 22106 27145 22140
rect 27145 22106 27154 22140
rect 27102 22097 27154 22106
rect 27102 19720 27154 19729
rect 27102 19686 27111 19720
rect 27111 19686 27145 19720
rect 27145 19686 27154 19720
rect 27102 19677 27154 19686
rect 27102 17160 27154 17169
rect 27102 17126 27111 17160
rect 27111 17126 27145 17160
rect 27145 17126 27154 17160
rect 27102 17117 27154 17126
rect 27102 14740 27154 14749
rect 27102 14706 27111 14740
rect 27111 14706 27145 14740
rect 27145 14706 27154 14740
rect 27102 14697 27154 14706
rect 27102 12180 27154 12189
rect 27102 12146 27111 12180
rect 27111 12146 27145 12180
rect 27145 12146 27154 12180
rect 27102 12137 27154 12146
rect 27102 9760 27154 9769
rect 27102 9726 27111 9760
rect 27111 9726 27145 9760
rect 27145 9726 27154 9760
rect 27102 9717 27154 9726
rect 27102 7200 27154 7209
rect 27102 7166 27111 7200
rect 27111 7166 27145 7200
rect 27145 7166 27154 7200
rect 27102 7157 27154 7166
rect 27102 4780 27154 4789
rect 27102 4746 27111 4780
rect 27111 4746 27145 4780
rect 27145 4746 27154 4780
rect 27102 4737 27154 4746
rect 28006 22027 28074 22079
rect 28006 19607 28074 19659
rect 28006 17047 28074 17099
rect 28006 14627 28074 14679
rect 28006 12067 28074 12119
rect 28006 9647 28074 9699
rect 28006 7087 28074 7139
rect 28006 4667 28074 4719
rect 17 32 205 90
rect 25763 32 25951 90
<< metal2 >>
rect 27102 22149 27154 22155
rect 27102 22076 27154 22097
rect 27102 22030 27200 22076
rect 28000 22027 28006 22079
rect 28074 22027 28980 22079
rect 27102 19729 27154 19735
rect 27102 19656 27154 19677
rect 27102 19610 27200 19656
rect 28000 19607 28006 19659
rect 28074 19607 28980 19659
rect 27102 17169 27154 17175
rect 27102 17096 27154 17117
rect 27102 17050 27200 17096
rect 28000 17047 28006 17099
rect 28074 17047 28980 17099
rect 27102 14749 27154 14755
rect 27102 14676 27154 14697
rect 27102 14630 27200 14676
rect 28000 14627 28006 14679
rect 28074 14627 28980 14679
rect 27102 12189 27154 12195
rect 27102 12116 27154 12137
rect 27102 12070 27200 12116
rect 28000 12067 28006 12119
rect 28074 12067 28980 12119
rect 27102 9769 27154 9775
rect 27102 9696 27154 9717
rect 27102 9650 27200 9696
rect 28000 9647 28006 9699
rect 28074 9647 28980 9699
rect 27102 7209 27154 7215
rect 27102 7136 27154 7157
rect 27102 7090 27200 7136
rect 28000 7087 28006 7139
rect 28074 7087 28980 7139
rect 27102 4789 27154 4795
rect 27102 4716 27154 4737
rect 27102 4670 27200 4716
rect 28000 4667 28006 4719
rect 28074 4667 28980 4719
rect 27217 2703 27226 2853
rect 27465 2848 28595 2853
rect 27465 2708 27854 2848
rect 28586 2708 28595 2848
rect 27465 2703 28595 2708
rect 28889 2462 28980 2514
rect 11 1734 111 2303
rect 11 1494 16 1734
rect 106 1494 111 1734
rect 11 96 111 1494
rect 25857 2268 26057 2303
rect 25857 2178 25876 2268
rect 26052 2178 26057 2268
rect 28889 2262 28980 2314
rect 25857 1734 26057 2178
rect 28889 2062 28980 2114
rect 28889 1862 28980 1914
rect 25857 1494 25862 1734
rect 26052 1494 26057 1734
rect 28889 1662 28980 1714
rect 25857 1485 26057 1494
rect 25857 96 25957 1485
rect 28889 1462 28980 1514
rect 28889 1262 28980 1314
rect 28889 1062 28980 1114
rect 28889 862 28980 914
rect 28889 662 28980 714
rect 28889 462 28980 514
rect 28889 262 28980 314
rect 11 90 211 96
rect 11 32 17 90
rect 205 32 211 90
rect 11 26 211 32
rect 25757 90 25957 96
rect 25757 32 25763 90
rect 25951 32 25957 90
rect 25757 26 25957 32
<< via2 >>
rect 27226 2703 27465 2853
rect 27854 2708 28586 2848
rect 16 1494 106 1734
rect 25876 2178 26052 2268
rect 25862 1494 26052 1734
<< metal3 >>
rect 27475 3502 27743 22193
rect 27221 3253 27743 3502
rect 27221 2853 27470 3253
rect 27859 3153 27969 22193
rect 27221 2703 27226 2853
rect 27465 2703 27470 2853
rect 111 2268 26057 2273
rect 111 2178 25876 2268
rect 26052 2178 26057 2268
rect 111 2173 26057 2178
rect 27221 2089 27470 2703
rect 27570 2953 28870 3153
rect 27570 2653 27751 2953
rect 27849 2848 28591 2853
rect 27849 2708 27854 2848
rect 28586 2708 28591 2848
rect 27849 2653 28591 2708
rect 28689 2653 28870 2953
rect 151 1839 27470 2089
rect 11 1734 27570 1739
rect 11 1494 16 1734
rect 106 1494 25862 1734
rect 26052 1494 27570 1734
rect 11 1489 27570 1494
use out_drive  out_drive_0
timestamp 1728730538
transform 1 0 22500 0 1 21773
box 4700 -55 5500 474
use out_drive  out_drive_1
timestamp 1728730538
transform 1 0 22500 0 1 4413
box 4700 -55 5500 474
use out_drive  out_drive_2
timestamp 1728730538
transform 1 0 22500 0 1 6833
box 4700 -55 5500 474
use out_drive  out_drive_3
timestamp 1728730538
transform 1 0 22500 0 1 9393
box 4700 -55 5500 474
use out_drive  out_drive_4
timestamp 1728730538
transform 1 0 22500 0 1 11813
box 4700 -55 5500 474
use out_drive  out_drive_5
timestamp 1728730538
transform 1 0 22500 0 1 14373
box 4700 -55 5500 474
use out_drive  out_drive_6
timestamp 1728730538
transform 1 0 22500 0 1 16793
box 4700 -55 5500 474
use out_drive  out_drive_7
timestamp 1728730538
transform 1 0 22500 0 1 19353
box 4700 -55 5500 474
use rom_32k_core  rom_32k_core_0
timestamp 1730660059
transform 1 0 249 0 1 2413
box -169 -2413 28640 20010
<< labels >>
flabel metal3 s 151 1839 27470 2089 0 FreeSans 400 0 0 0 VPWR
port 21 nsew power bidirectional
flabel metal3 s 111 2173 26057 2273 0 FreeSans 400 0 0 0 VGND
port 20 nsew ground bidirectional
flabel metal3 s 11 1489 27751 1739 0 FreeSans 400 0 0 0 VGND
port 20 nsew ground bidirectional
flabel metal2 s 28920 22027 28980 22079 0 FreeSans 160 0 0 0 q[7]
port 19 nsew signal output
flabel metal2 s 28920 19607 28980 19659 0 FreeSans 160 0 0 0 q[6]
port 18 nsew signal output
flabel metal2 s 28920 17047 28980 17099 0 FreeSans 160 0 0 0 q[5]
port 17 nsew signal output
flabel metal2 s 28920 14627 28980 14679 0 FreeSans 160 0 0 0 q[4]
port 16 nsew signal output
flabel metal2 s 28920 12067 28980 12119 0 FreeSans 160 0 0 0 q[3]
port 15 nsew signal output
flabel metal2 s 28920 9647 28980 9699 0 FreeSans 160 0 0 0 q[2]
port 14 nsew signal output
flabel metal2 s 28920 7087 28980 7139 0 FreeSans 160 0 0 0 q[1]
port 13 nsew signal output
flabel metal2 s 28920 4667 28980 4719 0 FreeSans 160 0 0 0 q[0]
port 12 nsew signal output
flabel metal2 s 28920 262 28980 314 0 FreeSans 160 0 0 0 addr[11]
port 11 nsew signal input
flabel metal2 s 28920 462 28980 514 0 FreeSans 160 0 0 0 addr[10]
port 10 nsew signal input
flabel metal2 s 28920 662 28980 714 0 FreeSans 160 0 0 0 addr[9]
port 9 nsew signal input
flabel metal2 s 28920 862 28980 914 0 FreeSans 160 0 0 0 addr[8]
port 8 nsew signal input
flabel metal2 s 28920 1062 28980 1114 0 FreeSans 160 0 0 0 addr[7]
port 7 nsew signal input
flabel metal2 s 28920 1262 28980 1314 0 FreeSans 160 0 0 0 addr[6]
port 6 nsew signal input
flabel metal2 s 28920 1462 28980 1514 0 FreeSans 160 0 0 0 addr[5]
port 5 nsew signal input
flabel metal2 s 28920 2462 28980 2514 0 FreeSans 160 0 0 0 addr[4]
port 4 nsew signal input
flabel metal2 s 28920 2262 28980 2314 0 FreeSans 160 0 0 0 addr[3]
port 3 nsew signal input
flabel metal2 s 28920 2062 28980 2114 0 FreeSans 160 0 0 0 addr[2]
port 2 nsew signal input
flabel metal2 s 28920 1862 28980 1914 0 FreeSans 160 0 0 0 addr[1]
port 1 nsew signal input
flabel metal2 s 28920 1662 28980 1714 0 FreeSans 160 0 0 0 addr[0]
port 0 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 28980 22460
<< end >>
