magic
tech sky130A
magscale 1 2
timestamp 1730654005
<< viali >>
rect 2881 8517 2915 8551
rect 7665 8517 7699 8551
rect 9045 8517 9079 8551
rect 11069 8517 11103 8551
rect 2053 8449 2087 8483
rect 8401 8449 8435 8483
rect 9873 8449 9907 8483
rect 10241 8449 10275 8483
rect 6009 7837 6043 7871
rect 6101 7837 6135 7871
rect 6837 7837 6871 7871
rect 8148 7837 8182 7871
rect 8401 7837 8435 7871
rect 9712 7837 9746 7871
rect 9965 7837 9999 7871
rect 7044 7701 7078 7735
rect 8608 7701 8642 7735
rect 7044 7497 7078 7531
rect 8608 7497 8642 7531
rect 6009 7361 6043 7395
rect 6101 7361 6135 7395
rect 6837 7361 6871 7395
rect 8148 7361 8182 7395
rect 8401 7361 8435 7395
rect 9712 7361 9746 7395
rect 9965 7361 9999 7395
rect 857 6749 891 6783
rect 949 6749 983 6783
rect 2053 6749 2087 6783
rect 6009 6749 6043 6783
rect 6101 6749 6135 6783
rect 6837 6749 6871 6783
rect 8148 6749 8182 6783
rect 8401 6749 8435 6783
rect 9712 6749 9746 6783
rect 9965 6749 9999 6783
rect 1317 6681 1351 6715
rect 1685 6681 1719 6715
rect 2306 6681 2340 6715
rect 581 6613 615 6647
rect 1869 6613 1903 6647
rect 3410 6613 3444 6647
rect 7044 6613 7078 6647
rect 8608 6613 8642 6647
rect 581 6409 615 6443
rect 1869 6409 1903 6443
rect 3410 6409 3444 6443
rect 7044 6409 7078 6443
rect 8608 6409 8642 6443
rect 1317 6341 1351 6375
rect 1685 6341 1719 6375
rect 2306 6341 2340 6375
rect 857 6273 891 6307
rect 949 6273 983 6307
rect 2053 6273 2087 6307
rect 6009 6273 6043 6307
rect 6101 6273 6135 6307
rect 6837 6273 6871 6307
rect 8148 6273 8182 6307
rect 8401 6273 8435 6307
rect 9712 6273 9746 6307
rect 9965 6273 9999 6307
rect 857 5661 891 5695
rect 949 5661 983 5695
rect 2053 5661 2087 5695
rect 6009 5661 6043 5695
rect 6101 5661 6135 5695
rect 6837 5661 6871 5695
rect 8148 5661 8182 5695
rect 8401 5661 8435 5695
rect 9712 5661 9746 5695
rect 9965 5661 9999 5695
rect 1317 5593 1351 5627
rect 1685 5593 1719 5627
rect 2306 5593 2340 5627
rect 581 5525 615 5559
rect 1869 5525 1903 5559
rect 3410 5525 3444 5559
rect 7044 5525 7078 5559
rect 8608 5525 8642 5559
rect 581 5321 615 5355
rect 1869 5321 1903 5355
rect 3410 5321 3444 5355
rect 7044 5321 7078 5355
rect 8608 5321 8642 5355
rect 1317 5253 1351 5287
rect 1685 5253 1719 5287
rect 2306 5253 2340 5287
rect 857 5185 891 5219
rect 949 5185 983 5219
rect 2053 5185 2087 5219
rect 6009 5185 6043 5219
rect 6101 5185 6135 5219
rect 6837 5185 6871 5219
rect 8148 5185 8182 5219
rect 8401 5185 8435 5219
rect 9712 5185 9746 5219
rect 9965 5185 9999 5219
rect 857 4573 891 4607
rect 949 4573 983 4607
rect 2053 4573 2087 4607
rect 6009 4573 6043 4607
rect 6101 4573 6135 4607
rect 6837 4573 6871 4607
rect 8148 4573 8182 4607
rect 8401 4573 8435 4607
rect 9712 4573 9746 4607
rect 9965 4573 9999 4607
rect 1317 4505 1351 4539
rect 1685 4505 1719 4539
rect 2306 4505 2340 4539
rect 581 4437 615 4471
rect 1869 4437 1903 4471
rect 3410 4437 3444 4471
rect 7044 4437 7078 4471
rect 8608 4437 8642 4471
rect 581 4233 615 4267
rect 1869 4233 1903 4267
rect 3410 4233 3444 4267
rect 7044 4233 7078 4267
rect 8608 4233 8642 4267
rect 1317 4165 1351 4199
rect 1685 4165 1719 4199
rect 2306 4165 2340 4199
rect 857 4097 891 4131
rect 949 4097 983 4131
rect 2053 4097 2087 4131
rect 6009 4097 6043 4131
rect 6101 4097 6135 4131
rect 6837 4097 6871 4131
rect 8148 4097 8182 4131
rect 8401 4097 8435 4131
rect 9712 4097 9746 4131
rect 9965 4097 9999 4131
rect 857 3485 891 3519
rect 949 3485 983 3519
rect 2053 3485 2087 3519
rect 6009 3485 6043 3519
rect 6101 3485 6135 3519
rect 6837 3485 6871 3519
rect 8148 3485 8182 3519
rect 8401 3485 8435 3519
rect 9712 3485 9746 3519
rect 9965 3485 9999 3519
rect 1317 3417 1351 3451
rect 1685 3417 1719 3451
rect 2306 3417 2340 3451
rect 581 3349 615 3383
rect 1869 3349 1903 3383
rect 3410 3349 3444 3383
rect 7044 3349 7078 3383
rect 8608 3349 8642 3383
rect 581 3145 615 3179
rect 1869 3145 1903 3179
rect 3410 3145 3444 3179
rect 7044 3145 7078 3179
rect 8608 3145 8642 3179
rect 1317 3077 1351 3111
rect 1685 3077 1719 3111
rect 2306 3077 2340 3111
rect 857 3009 891 3043
rect 949 3009 983 3043
rect 2053 3009 2087 3043
rect 6009 3009 6043 3043
rect 6101 3009 6135 3043
rect 6837 3009 6871 3043
rect 8148 3009 8182 3043
rect 8401 3009 8435 3043
rect 9712 3009 9746 3043
rect 9965 3009 9999 3043
rect 857 2397 891 2431
rect 949 2397 983 2431
rect 2053 2397 2087 2431
rect 6009 2397 6043 2431
rect 6101 2397 6135 2431
rect 6837 2397 6871 2431
rect 8148 2397 8182 2431
rect 8401 2397 8435 2431
rect 9712 2397 9746 2431
rect 9965 2397 9999 2431
rect 1317 2329 1351 2363
rect 1685 2329 1719 2363
rect 2306 2329 2340 2363
rect 581 2261 615 2295
rect 1869 2261 1903 2295
rect 3410 2261 3444 2295
rect 7044 2261 7078 2295
rect 8608 2261 8642 2295
rect 581 2057 615 2091
rect 1869 2057 1903 2091
rect 3410 2057 3444 2091
rect 7044 2057 7078 2091
rect 8608 2057 8642 2091
rect 1317 1989 1351 2023
rect 1685 1989 1719 2023
rect 2306 1989 2340 2023
rect 857 1921 891 1955
rect 949 1921 983 1955
rect 2053 1921 2087 1955
rect 6009 1921 6043 1955
rect 6101 1921 6135 1955
rect 6837 1921 6871 1955
rect 8148 1921 8182 1955
rect 8401 1921 8435 1955
rect 9712 1921 9746 1955
rect 9965 1921 9999 1955
rect 6009 1309 6043 1343
rect 6101 1309 6135 1343
rect 6837 1309 6871 1343
rect 8148 1309 8182 1343
rect 8401 1309 8435 1343
rect 9712 1309 9746 1343
rect 9965 1309 9999 1343
rect 7044 1173 7078 1207
rect 8608 1173 8642 1207
rect 7044 969 7078 1003
rect 8608 969 8642 1003
rect 6009 833 6043 867
rect 6101 833 6135 867
rect 6837 833 6871 867
rect 8148 833 8182 867
rect 8401 833 8435 867
rect 9712 833 9746 867
rect 9965 833 9999 867
<< metal1 >>
rect 2866 8508 2872 8560
rect 2924 8508 2930 8560
rect 7650 8508 7656 8560
rect 7708 8508 7714 8560
rect 9030 8508 9036 8560
rect 9088 8508 9094 8560
rect 11054 8508 11060 8560
rect 11112 8508 11118 8560
rect 2038 8440 2044 8492
rect 2096 8440 2102 8492
rect 8386 8440 8392 8492
rect 8444 8440 8450 8492
rect 9858 8440 9864 8492
rect 9916 8440 9922 8492
rect 10226 8440 10232 8492
rect 10284 8440 10290 8492
rect 4706 7828 4712 7880
rect 4764 7868 4770 7880
rect 5997 7871 6055 7877
rect 5997 7868 6009 7871
rect 4764 7840 6009 7868
rect 4764 7828 4770 7840
rect 5997 7837 6009 7840
rect 6043 7868 6055 7871
rect 6089 7871 6147 7877
rect 6089 7868 6101 7871
rect 6043 7840 6101 7868
rect 6043 7837 6055 7840
rect 5997 7831 6055 7837
rect 6089 7837 6101 7840
rect 6135 7837 6147 7871
rect 6089 7831 6147 7837
rect 6825 7871 6883 7877
rect 6825 7837 6837 7871
rect 6871 7868 6883 7871
rect 8136 7871 8194 7877
rect 6871 7840 6960 7868
rect 6871 7837 6883 7840
rect 6825 7831 6883 7837
rect 6932 7732 6960 7840
rect 8136 7837 8148 7871
rect 8182 7868 8194 7871
rect 8182 7840 8340 7868
rect 8182 7837 8194 7840
rect 8136 7831 8194 7837
rect 7032 7735 7090 7741
rect 7032 7732 7044 7735
rect 6932 7704 7044 7732
rect 7032 7701 7044 7704
rect 7078 7701 7090 7735
rect 8312 7732 8340 7840
rect 8386 7828 8392 7880
rect 8444 7828 8450 7880
rect 9700 7871 9758 7877
rect 9700 7837 9712 7871
rect 9746 7868 9758 7871
rect 9746 7840 9858 7868
rect 9746 7837 9758 7840
rect 9700 7831 9758 7837
rect 9830 7800 9858 7840
rect 9950 7828 9956 7880
rect 10008 7828 10014 7880
rect 10410 7800 10416 7812
rect 9830 7772 10416 7800
rect 10410 7760 10416 7772
rect 10468 7760 10474 7812
rect 8596 7735 8654 7741
rect 8596 7732 8608 7735
rect 8312 7704 8608 7732
rect 7032 7695 7090 7701
rect 8596 7701 8608 7704
rect 8642 7701 8654 7735
rect 8596 7695 8654 7701
rect 7032 7531 7090 7537
rect 7032 7528 7044 7531
rect 6932 7500 7044 7528
rect 4798 7352 4804 7404
rect 4856 7392 4862 7404
rect 5997 7395 6055 7401
rect 5997 7392 6009 7395
rect 4856 7364 6009 7392
rect 4856 7352 4862 7364
rect 5997 7361 6009 7364
rect 6043 7392 6055 7395
rect 6089 7395 6147 7401
rect 6089 7392 6101 7395
rect 6043 7364 6101 7392
rect 6043 7361 6055 7364
rect 5997 7355 6055 7361
rect 6089 7361 6101 7364
rect 6135 7361 6147 7395
rect 6089 7355 6147 7361
rect 6825 7395 6883 7401
rect 6825 7361 6837 7395
rect 6871 7392 6883 7395
rect 6932 7392 6960 7500
rect 7032 7497 7044 7500
rect 7078 7497 7090 7531
rect 8596 7531 8654 7537
rect 8596 7528 8608 7531
rect 7032 7491 7090 7497
rect 8312 7500 8608 7528
rect 6871 7364 6960 7392
rect 8136 7395 8194 7401
rect 6871 7361 6883 7364
rect 6825 7355 6883 7361
rect 8136 7361 8148 7395
rect 8182 7392 8194 7395
rect 8312 7392 8340 7500
rect 8596 7497 8608 7500
rect 8642 7497 8654 7531
rect 8596 7491 8654 7497
rect 10502 7460 10508 7472
rect 9830 7432 10508 7460
rect 8182 7364 8340 7392
rect 8182 7361 8194 7364
rect 8136 7355 8194 7361
rect 8386 7352 8392 7404
rect 8444 7352 8450 7404
rect 9700 7395 9758 7401
rect 9700 7361 9712 7395
rect 9746 7392 9758 7395
rect 9830 7392 9858 7432
rect 10502 7420 10508 7432
rect 10560 7420 10566 7472
rect 9746 7364 9858 7392
rect 9746 7361 9758 7364
rect 9700 7355 9758 7361
rect 9950 7352 9956 7404
rect 10008 7352 10014 7404
rect 1780 6956 6776 6984
rect 1578 6808 1584 6860
rect 1636 6808 1642 6860
rect -906 6740 -900 6792
rect -848 6780 -842 6792
rect 845 6783 903 6789
rect 845 6780 857 6783
rect -848 6752 857 6780
rect -848 6740 -842 6752
rect 845 6749 857 6752
rect 891 6749 903 6783
rect 845 6743 903 6749
rect 934 6740 940 6792
rect 992 6740 998 6792
rect -2746 6672 -2740 6724
rect -2688 6712 -2682 6724
rect 1305 6715 1363 6721
rect 1305 6712 1317 6715
rect -2688 6684 1317 6712
rect -2688 6672 -2682 6684
rect 1305 6681 1317 6684
rect 1351 6681 1363 6715
rect 1305 6675 1363 6681
rect 1673 6715 1731 6721
rect 1673 6681 1685 6715
rect 1719 6712 1731 6715
rect 1780 6712 1808 6956
rect 2038 6740 2044 6792
rect 2096 6740 2102 6792
rect 4890 6740 4896 6792
rect 4948 6780 4954 6792
rect 5997 6783 6055 6789
rect 5997 6780 6009 6783
rect 4948 6752 6009 6780
rect 4948 6740 4954 6752
rect 5997 6749 6009 6752
rect 6043 6780 6055 6783
rect 6089 6783 6147 6789
rect 6089 6780 6101 6783
rect 6043 6752 6101 6780
rect 6043 6749 6055 6752
rect 5997 6743 6055 6749
rect 6089 6749 6101 6752
rect 6135 6749 6147 6783
rect 6748 6780 6776 6956
rect 6825 6783 6883 6789
rect 6825 6780 6837 6783
rect 6748 6752 6837 6780
rect 6089 6743 6147 6749
rect 6825 6749 6837 6752
rect 6871 6780 6883 6783
rect 8136 6783 8194 6789
rect 6871 6752 6960 6780
rect 6871 6749 6883 6752
rect 6825 6743 6883 6749
rect 2294 6715 2352 6721
rect 2294 6712 2306 6715
rect 1719 6684 1808 6712
rect 2148 6684 2306 6712
rect 1719 6681 1731 6684
rect 1673 6675 1731 6681
rect -1826 6604 -1820 6656
rect -1768 6644 -1762 6656
rect 569 6647 627 6653
rect 569 6644 581 6647
rect -1768 6616 581 6644
rect -1768 6604 -1762 6616
rect 569 6613 581 6616
rect 615 6613 627 6647
rect 569 6607 627 6613
rect 1857 6647 1915 6653
rect 1857 6613 1869 6647
rect 1903 6644 1915 6647
rect 2148 6644 2176 6684
rect 2294 6681 2306 6684
rect 2340 6681 2352 6715
rect 2294 6675 2352 6681
rect 1903 6616 2176 6644
rect 3398 6647 3456 6653
rect 1903 6613 1915 6616
rect 1857 6607 1915 6613
rect 3398 6613 3410 6647
rect 3444 6644 3456 6647
rect 3510 6644 3516 6656
rect 3444 6616 3516 6644
rect 3444 6613 3456 6616
rect 3398 6607 3456 6613
rect 3510 6604 3516 6616
rect 3568 6604 3574 6656
rect 6932 6644 6960 6752
rect 8136 6749 8148 6783
rect 8182 6780 8194 6783
rect 8182 6752 8340 6780
rect 8182 6749 8194 6752
rect 8136 6743 8194 6749
rect 7032 6647 7090 6653
rect 7032 6644 7044 6647
rect 6932 6616 7044 6644
rect 7032 6613 7044 6616
rect 7078 6613 7090 6647
rect 8312 6644 8340 6752
rect 8386 6740 8392 6792
rect 8444 6740 8450 6792
rect 9700 6783 9758 6789
rect 9700 6749 9712 6783
rect 9746 6780 9758 6783
rect 9746 6752 9858 6780
rect 9746 6749 9758 6752
rect 9700 6743 9758 6749
rect 9830 6712 9858 6752
rect 9950 6740 9956 6792
rect 10008 6740 10014 6792
rect 10594 6712 10600 6724
rect 9830 6684 10600 6712
rect 10594 6672 10600 6684
rect 10652 6672 10658 6724
rect 8596 6647 8654 6653
rect 8596 6644 8608 6647
rect 8312 6616 8608 6644
rect 7032 6607 7090 6613
rect 8596 6613 8608 6616
rect 8642 6613 8654 6647
rect 8596 6607 8654 6613
rect -1734 6400 -1728 6452
rect -1676 6440 -1670 6452
rect 569 6443 627 6449
rect 569 6440 581 6443
rect -1676 6412 581 6440
rect -1676 6400 -1670 6412
rect 569 6409 581 6412
rect 615 6409 627 6443
rect 569 6403 627 6409
rect 1857 6443 1915 6449
rect 1857 6409 1869 6443
rect 1903 6440 1915 6443
rect 3398 6443 3456 6449
rect 1903 6412 2176 6440
rect 1903 6409 1915 6412
rect 1857 6403 1915 6409
rect -2654 6332 -2648 6384
rect -2596 6372 -2590 6384
rect 1305 6375 1363 6381
rect 1305 6372 1317 6375
rect -2596 6344 1317 6372
rect -2596 6332 -2590 6344
rect 1305 6341 1317 6344
rect 1351 6341 1363 6375
rect 1305 6335 1363 6341
rect 1673 6375 1731 6381
rect 1673 6341 1685 6375
rect 1719 6372 1731 6375
rect 2148 6372 2176 6412
rect 3398 6409 3410 6443
rect 3444 6440 3456 6443
rect 3602 6440 3608 6452
rect 3444 6412 3608 6440
rect 3444 6409 3456 6412
rect 3398 6403 3456 6409
rect 3602 6400 3608 6412
rect 3660 6400 3666 6452
rect 7032 6443 7090 6449
rect 7032 6440 7044 6443
rect 6932 6412 7044 6440
rect 2294 6375 2352 6381
rect 2294 6372 2306 6375
rect 1719 6344 1808 6372
rect 2148 6344 2306 6372
rect 1719 6341 1731 6344
rect 1673 6335 1731 6341
rect -814 6264 -808 6316
rect -756 6304 -750 6316
rect 845 6307 903 6313
rect 845 6304 857 6307
rect -756 6276 857 6304
rect -756 6264 -750 6276
rect 845 6273 857 6276
rect 891 6273 903 6307
rect 845 6267 903 6273
rect 934 6264 940 6316
rect 992 6264 998 6316
rect 1578 6196 1584 6248
rect 1636 6196 1642 6248
rect 1780 6100 1808 6344
rect 2294 6341 2306 6344
rect 2340 6341 2352 6375
rect 2294 6335 2352 6341
rect 2038 6264 2044 6316
rect 2096 6264 2102 6316
rect 4982 6264 4988 6316
rect 5040 6304 5046 6316
rect 5997 6307 6055 6313
rect 5997 6304 6009 6307
rect 5040 6276 6009 6304
rect 5040 6264 5046 6276
rect 5997 6273 6009 6276
rect 6043 6304 6055 6307
rect 6089 6307 6147 6313
rect 6089 6304 6101 6307
rect 6043 6276 6101 6304
rect 6043 6273 6055 6276
rect 5997 6267 6055 6273
rect 6089 6273 6101 6276
rect 6135 6273 6147 6307
rect 6825 6307 6883 6313
rect 6825 6304 6837 6307
rect 6089 6267 6147 6273
rect 6748 6276 6837 6304
rect 6748 6100 6776 6276
rect 6825 6273 6837 6276
rect 6871 6304 6883 6307
rect 6932 6304 6960 6412
rect 7032 6409 7044 6412
rect 7078 6409 7090 6443
rect 8596 6443 8654 6449
rect 8596 6440 8608 6443
rect 7032 6403 7090 6409
rect 8312 6412 8608 6440
rect 6871 6276 6960 6304
rect 8136 6307 8194 6313
rect 6871 6273 6883 6276
rect 6825 6267 6883 6273
rect 8136 6273 8148 6307
rect 8182 6304 8194 6307
rect 8312 6304 8340 6412
rect 8596 6409 8608 6412
rect 8642 6409 8654 6443
rect 8596 6403 8654 6409
rect 10686 6372 10692 6384
rect 9830 6344 10692 6372
rect 8182 6276 8340 6304
rect 8182 6273 8194 6276
rect 8136 6267 8194 6273
rect 8386 6264 8392 6316
rect 8444 6264 8450 6316
rect 9700 6307 9758 6313
rect 9700 6273 9712 6307
rect 9746 6304 9758 6307
rect 9830 6304 9858 6344
rect 10686 6332 10692 6344
rect 10744 6332 10750 6384
rect 9746 6276 9858 6304
rect 9746 6273 9758 6276
rect 9700 6267 9758 6273
rect 9950 6264 9956 6316
rect 10008 6264 10014 6316
rect 1780 6072 6776 6100
rect 1780 5868 6776 5896
rect 1578 5720 1584 5772
rect 1636 5720 1642 5772
rect -722 5652 -716 5704
rect -664 5692 -658 5704
rect 845 5695 903 5701
rect 845 5692 857 5695
rect -664 5664 857 5692
rect -664 5652 -658 5664
rect 845 5661 857 5664
rect 891 5661 903 5695
rect 845 5655 903 5661
rect 934 5652 940 5704
rect 992 5652 998 5704
rect -2562 5584 -2556 5636
rect -2504 5624 -2498 5636
rect 1305 5627 1363 5633
rect 1305 5624 1317 5627
rect -2504 5596 1317 5624
rect -2504 5584 -2498 5596
rect 1305 5593 1317 5596
rect 1351 5593 1363 5627
rect 1305 5587 1363 5593
rect 1673 5627 1731 5633
rect 1673 5593 1685 5627
rect 1719 5624 1731 5627
rect 1780 5624 1808 5868
rect 2038 5652 2044 5704
rect 2096 5652 2102 5704
rect 5074 5652 5080 5704
rect 5132 5692 5138 5704
rect 5997 5695 6055 5701
rect 5997 5692 6009 5695
rect 5132 5664 6009 5692
rect 5132 5652 5138 5664
rect 5997 5661 6009 5664
rect 6043 5692 6055 5695
rect 6089 5695 6147 5701
rect 6089 5692 6101 5695
rect 6043 5664 6101 5692
rect 6043 5661 6055 5664
rect 5997 5655 6055 5661
rect 6089 5661 6101 5664
rect 6135 5661 6147 5695
rect 6748 5692 6776 5868
rect 6825 5695 6883 5701
rect 6825 5692 6837 5695
rect 6748 5664 6837 5692
rect 6089 5655 6147 5661
rect 6825 5661 6837 5664
rect 6871 5692 6883 5695
rect 8136 5695 8194 5701
rect 6871 5664 6960 5692
rect 6871 5661 6883 5664
rect 6825 5655 6883 5661
rect 2294 5627 2352 5633
rect 2294 5624 2306 5627
rect 1719 5596 1808 5624
rect 2148 5596 2306 5624
rect 1719 5593 1731 5596
rect 1673 5587 1731 5593
rect -1642 5516 -1636 5568
rect -1584 5556 -1578 5568
rect 569 5559 627 5565
rect 569 5556 581 5559
rect -1584 5528 581 5556
rect -1584 5516 -1578 5528
rect 569 5525 581 5528
rect 615 5525 627 5559
rect 569 5519 627 5525
rect 1857 5559 1915 5565
rect 1857 5525 1869 5559
rect 1903 5556 1915 5559
rect 2148 5556 2176 5596
rect 2294 5593 2306 5596
rect 2340 5593 2352 5627
rect 2294 5587 2352 5593
rect 1903 5528 2176 5556
rect 3398 5559 3456 5565
rect 1903 5525 1915 5528
rect 1857 5519 1915 5525
rect 3398 5525 3410 5559
rect 3444 5556 3456 5559
rect 3694 5556 3700 5568
rect 3444 5528 3700 5556
rect 3444 5525 3456 5528
rect 3398 5519 3456 5525
rect 3694 5516 3700 5528
rect 3752 5516 3758 5568
rect 6932 5556 6960 5664
rect 8136 5661 8148 5695
rect 8182 5692 8194 5695
rect 8182 5664 8340 5692
rect 8182 5661 8194 5664
rect 8136 5655 8194 5661
rect 7032 5559 7090 5565
rect 7032 5556 7044 5559
rect 6932 5528 7044 5556
rect 7032 5525 7044 5528
rect 7078 5525 7090 5559
rect 8312 5556 8340 5664
rect 8386 5652 8392 5704
rect 8444 5652 8450 5704
rect 9700 5695 9758 5701
rect 9700 5661 9712 5695
rect 9746 5692 9758 5695
rect 9746 5664 9858 5692
rect 9746 5661 9758 5664
rect 9700 5655 9758 5661
rect 9830 5624 9858 5664
rect 9950 5652 9956 5704
rect 10008 5652 10014 5704
rect 10778 5624 10784 5636
rect 9830 5596 10784 5624
rect 10778 5584 10784 5596
rect 10836 5584 10842 5636
rect 8596 5559 8654 5565
rect 8596 5556 8608 5559
rect 8312 5528 8608 5556
rect 7032 5519 7090 5525
rect 8596 5525 8608 5528
rect 8642 5525 8654 5559
rect 8596 5519 8654 5525
rect -1550 5312 -1544 5364
rect -1492 5352 -1486 5364
rect 569 5355 627 5361
rect 569 5352 581 5355
rect -1492 5324 581 5352
rect -1492 5312 -1486 5324
rect 569 5321 581 5324
rect 615 5321 627 5355
rect 569 5315 627 5321
rect 1857 5355 1915 5361
rect 1857 5321 1869 5355
rect 1903 5352 1915 5355
rect 3398 5355 3456 5361
rect 1903 5324 2176 5352
rect 1903 5321 1915 5324
rect 1857 5315 1915 5321
rect -2470 5244 -2464 5296
rect -2412 5284 -2406 5296
rect 1305 5287 1363 5293
rect 1305 5284 1317 5287
rect -2412 5256 1317 5284
rect -2412 5244 -2406 5256
rect 1305 5253 1317 5256
rect 1351 5253 1363 5287
rect 1305 5247 1363 5253
rect 1673 5287 1731 5293
rect 1673 5253 1685 5287
rect 1719 5284 1731 5287
rect 2148 5284 2176 5324
rect 3398 5321 3410 5355
rect 3444 5352 3456 5355
rect 3786 5352 3792 5364
rect 3444 5324 3792 5352
rect 3444 5321 3456 5324
rect 3398 5315 3456 5321
rect 3786 5312 3792 5324
rect 3844 5312 3850 5364
rect 7032 5355 7090 5361
rect 7032 5352 7044 5355
rect 6932 5324 7044 5352
rect 2294 5287 2352 5293
rect 2294 5284 2306 5287
rect 1719 5256 1808 5284
rect 2148 5256 2306 5284
rect 1719 5253 1731 5256
rect 1673 5247 1731 5253
rect -630 5176 -624 5228
rect -572 5216 -566 5228
rect 845 5219 903 5225
rect 845 5216 857 5219
rect -572 5188 857 5216
rect -572 5176 -566 5188
rect 845 5185 857 5188
rect 891 5185 903 5219
rect 845 5179 903 5185
rect 934 5176 940 5228
rect 992 5176 998 5228
rect 1578 5108 1584 5160
rect 1636 5108 1642 5160
rect 1780 5012 1808 5256
rect 2294 5253 2306 5256
rect 2340 5253 2352 5287
rect 2294 5247 2352 5253
rect 2038 5176 2044 5228
rect 2096 5176 2102 5228
rect 5166 5176 5172 5228
rect 5224 5216 5230 5228
rect 5997 5219 6055 5225
rect 5997 5216 6009 5219
rect 5224 5188 6009 5216
rect 5224 5176 5230 5188
rect 5997 5185 6009 5188
rect 6043 5216 6055 5219
rect 6089 5219 6147 5225
rect 6089 5216 6101 5219
rect 6043 5188 6101 5216
rect 6043 5185 6055 5188
rect 5997 5179 6055 5185
rect 6089 5185 6101 5188
rect 6135 5185 6147 5219
rect 6825 5219 6883 5225
rect 6825 5216 6837 5219
rect 6089 5179 6147 5185
rect 6748 5188 6837 5216
rect 6748 5012 6776 5188
rect 6825 5185 6837 5188
rect 6871 5216 6883 5219
rect 6932 5216 6960 5324
rect 7032 5321 7044 5324
rect 7078 5321 7090 5355
rect 8596 5355 8654 5361
rect 8596 5352 8608 5355
rect 7032 5315 7090 5321
rect 8312 5324 8608 5352
rect 6871 5188 6960 5216
rect 8136 5219 8194 5225
rect 6871 5185 6883 5188
rect 6825 5179 6883 5185
rect 8136 5185 8148 5219
rect 8182 5216 8194 5219
rect 8312 5216 8340 5324
rect 8596 5321 8608 5324
rect 8642 5321 8654 5355
rect 8596 5315 8654 5321
rect 10870 5284 10876 5296
rect 9830 5256 10876 5284
rect 8182 5188 8340 5216
rect 8182 5185 8194 5188
rect 8136 5179 8194 5185
rect 8386 5176 8392 5228
rect 8444 5176 8450 5228
rect 9700 5219 9758 5225
rect 9700 5185 9712 5219
rect 9746 5216 9758 5219
rect 9830 5216 9858 5256
rect 10870 5244 10876 5256
rect 10928 5244 10934 5296
rect 9746 5188 9858 5216
rect 9746 5185 9758 5188
rect 9700 5179 9758 5185
rect 9950 5176 9956 5228
rect 10008 5176 10014 5228
rect 1780 4984 6776 5012
rect 1780 4780 6776 4808
rect 1578 4632 1584 4684
rect 1636 4632 1642 4684
rect -538 4564 -532 4616
rect -480 4604 -474 4616
rect 845 4607 903 4613
rect 845 4604 857 4607
rect -480 4576 857 4604
rect -480 4564 -474 4576
rect 845 4573 857 4576
rect 891 4573 903 4607
rect 845 4567 903 4573
rect 934 4564 940 4616
rect 992 4564 998 4616
rect -2378 4496 -2372 4548
rect -2320 4536 -2314 4548
rect 1305 4539 1363 4545
rect 1305 4536 1317 4539
rect -2320 4508 1317 4536
rect -2320 4496 -2314 4508
rect 1305 4505 1317 4508
rect 1351 4505 1363 4539
rect 1305 4499 1363 4505
rect 1673 4539 1731 4545
rect 1673 4505 1685 4539
rect 1719 4536 1731 4539
rect 1780 4536 1808 4780
rect 2038 4564 2044 4616
rect 2096 4564 2102 4616
rect 5258 4564 5264 4616
rect 5316 4604 5322 4616
rect 5997 4607 6055 4613
rect 5997 4604 6009 4607
rect 5316 4576 6009 4604
rect 5316 4564 5322 4576
rect 5997 4573 6009 4576
rect 6043 4604 6055 4607
rect 6089 4607 6147 4613
rect 6089 4604 6101 4607
rect 6043 4576 6101 4604
rect 6043 4573 6055 4576
rect 5997 4567 6055 4573
rect 6089 4573 6101 4576
rect 6135 4573 6147 4607
rect 6748 4604 6776 4780
rect 6825 4607 6883 4613
rect 6825 4604 6837 4607
rect 6748 4576 6837 4604
rect 6089 4567 6147 4573
rect 6825 4573 6837 4576
rect 6871 4604 6883 4607
rect 8136 4607 8194 4613
rect 6871 4576 6960 4604
rect 6871 4573 6883 4576
rect 6825 4567 6883 4573
rect 2294 4539 2352 4545
rect 2294 4536 2306 4539
rect 1719 4508 1808 4536
rect 2148 4508 2306 4536
rect 1719 4505 1731 4508
rect 1673 4499 1731 4505
rect -1458 4428 -1452 4480
rect -1400 4468 -1394 4480
rect 569 4471 627 4477
rect 569 4468 581 4471
rect -1400 4440 581 4468
rect -1400 4428 -1394 4440
rect 569 4437 581 4440
rect 615 4437 627 4471
rect 569 4431 627 4437
rect 1857 4471 1915 4477
rect 1857 4437 1869 4471
rect 1903 4468 1915 4471
rect 2148 4468 2176 4508
rect 2294 4505 2306 4508
rect 2340 4505 2352 4539
rect 2294 4499 2352 4505
rect 1903 4440 2176 4468
rect 3398 4471 3456 4477
rect 1903 4437 1915 4440
rect 1857 4431 1915 4437
rect 3398 4437 3410 4471
rect 3444 4468 3456 4471
rect 3878 4468 3884 4480
rect 3444 4440 3884 4468
rect 3444 4437 3456 4440
rect 3398 4431 3456 4437
rect 3878 4428 3884 4440
rect 3936 4428 3942 4480
rect 6932 4468 6960 4576
rect 8136 4573 8148 4607
rect 8182 4604 8194 4607
rect 8182 4576 8340 4604
rect 8182 4573 8194 4576
rect 8136 4567 8194 4573
rect 7032 4471 7090 4477
rect 7032 4468 7044 4471
rect 6932 4440 7044 4468
rect 7032 4437 7044 4440
rect 7078 4437 7090 4471
rect 8312 4468 8340 4576
rect 8386 4564 8392 4616
rect 8444 4564 8450 4616
rect 9700 4607 9758 4613
rect 9700 4573 9712 4607
rect 9746 4604 9758 4607
rect 9746 4576 9858 4604
rect 9746 4573 9758 4576
rect 9700 4567 9758 4573
rect 9830 4536 9858 4576
rect 9950 4564 9956 4616
rect 10008 4564 10014 4616
rect 10962 4536 10968 4548
rect 9830 4508 10968 4536
rect 10962 4496 10968 4508
rect 11020 4496 11026 4548
rect 8596 4471 8654 4477
rect 8596 4468 8608 4471
rect 8312 4440 8608 4468
rect 7032 4431 7090 4437
rect 8596 4437 8608 4440
rect 8642 4437 8654 4471
rect 8596 4431 8654 4437
rect -1366 4224 -1360 4276
rect -1308 4264 -1302 4276
rect 569 4267 627 4273
rect 569 4264 581 4267
rect -1308 4236 581 4264
rect -1308 4224 -1302 4236
rect 569 4233 581 4236
rect 615 4233 627 4267
rect 569 4227 627 4233
rect 1857 4267 1915 4273
rect 1857 4233 1869 4267
rect 1903 4264 1915 4267
rect 3398 4267 3456 4273
rect 1903 4236 2176 4264
rect 1903 4233 1915 4236
rect 1857 4227 1915 4233
rect -2286 4156 -2280 4208
rect -2228 4196 -2222 4208
rect 1305 4199 1363 4205
rect 1305 4196 1317 4199
rect -2228 4168 1317 4196
rect -2228 4156 -2222 4168
rect 1305 4165 1317 4168
rect 1351 4165 1363 4199
rect 1305 4159 1363 4165
rect 1673 4199 1731 4205
rect 1673 4165 1685 4199
rect 1719 4196 1731 4199
rect 2148 4196 2176 4236
rect 3398 4233 3410 4267
rect 3444 4264 3456 4267
rect 3970 4264 3976 4276
rect 3444 4236 3976 4264
rect 3444 4233 3456 4236
rect 3398 4227 3456 4233
rect 3970 4224 3976 4236
rect 4028 4224 4034 4276
rect 7032 4267 7090 4273
rect 7032 4264 7044 4267
rect 6932 4236 7044 4264
rect 2294 4199 2352 4205
rect 2294 4196 2306 4199
rect 1719 4168 1808 4196
rect 2148 4168 2306 4196
rect 1719 4165 1731 4168
rect 1673 4159 1731 4165
rect -446 4088 -440 4140
rect -388 4128 -382 4140
rect 845 4131 903 4137
rect 845 4128 857 4131
rect -388 4100 857 4128
rect -388 4088 -382 4100
rect 845 4097 857 4100
rect 891 4097 903 4131
rect 845 4091 903 4097
rect 934 4088 940 4140
rect 992 4088 998 4140
rect 1578 4020 1584 4072
rect 1636 4020 1642 4072
rect 1780 3924 1808 4168
rect 2294 4165 2306 4168
rect 2340 4165 2352 4199
rect 2294 4159 2352 4165
rect 2038 4088 2044 4140
rect 2096 4088 2102 4140
rect 5350 4088 5356 4140
rect 5408 4128 5414 4140
rect 5997 4131 6055 4137
rect 5997 4128 6009 4131
rect 5408 4100 6009 4128
rect 5408 4088 5414 4100
rect 5997 4097 6009 4100
rect 6043 4128 6055 4131
rect 6089 4131 6147 4137
rect 6089 4128 6101 4131
rect 6043 4100 6101 4128
rect 6043 4097 6055 4100
rect 5997 4091 6055 4097
rect 6089 4097 6101 4100
rect 6135 4097 6147 4131
rect 6825 4131 6883 4137
rect 6825 4128 6837 4131
rect 6089 4091 6147 4097
rect 6748 4100 6837 4128
rect 6748 3924 6776 4100
rect 6825 4097 6837 4100
rect 6871 4128 6883 4131
rect 6932 4128 6960 4236
rect 7032 4233 7044 4236
rect 7078 4233 7090 4267
rect 8596 4267 8654 4273
rect 8596 4264 8608 4267
rect 7032 4227 7090 4233
rect 8312 4236 8608 4264
rect 6871 4100 6960 4128
rect 8136 4131 8194 4137
rect 6871 4097 6883 4100
rect 6825 4091 6883 4097
rect 8136 4097 8148 4131
rect 8182 4128 8194 4131
rect 8312 4128 8340 4236
rect 8596 4233 8608 4236
rect 8642 4233 8654 4267
rect 8596 4227 8654 4233
rect 10410 4196 10416 4208
rect 9830 4168 10416 4196
rect 8182 4100 8340 4128
rect 8182 4097 8194 4100
rect 8136 4091 8194 4097
rect 8386 4088 8392 4140
rect 8444 4088 8450 4140
rect 9700 4131 9758 4137
rect 9700 4097 9712 4131
rect 9746 4128 9758 4131
rect 9830 4128 9858 4168
rect 10410 4156 10416 4168
rect 10468 4156 10474 4208
rect 9746 4100 9858 4128
rect 9746 4097 9758 4100
rect 9700 4091 9758 4097
rect 9950 4088 9956 4140
rect 10008 4088 10014 4140
rect 1780 3896 6776 3924
rect 1780 3692 6776 3720
rect 1578 3544 1584 3596
rect 1636 3544 1642 3596
rect -354 3476 -348 3528
rect -296 3516 -290 3528
rect 845 3519 903 3525
rect 845 3516 857 3519
rect -296 3488 857 3516
rect -296 3476 -290 3488
rect 845 3485 857 3488
rect 891 3485 903 3519
rect 845 3479 903 3485
rect 934 3476 940 3528
rect 992 3476 998 3528
rect -2194 3408 -2188 3460
rect -2136 3448 -2130 3460
rect 1305 3451 1363 3457
rect 1305 3448 1317 3451
rect -2136 3420 1317 3448
rect -2136 3408 -2130 3420
rect 1305 3417 1317 3420
rect 1351 3417 1363 3451
rect 1305 3411 1363 3417
rect 1673 3451 1731 3457
rect 1673 3417 1685 3451
rect 1719 3448 1731 3451
rect 1780 3448 1808 3692
rect 2038 3476 2044 3528
rect 2096 3476 2102 3528
rect 5442 3476 5448 3528
rect 5500 3516 5506 3528
rect 5997 3519 6055 3525
rect 5997 3516 6009 3519
rect 5500 3488 6009 3516
rect 5500 3476 5506 3488
rect 5997 3485 6009 3488
rect 6043 3516 6055 3519
rect 6089 3519 6147 3525
rect 6089 3516 6101 3519
rect 6043 3488 6101 3516
rect 6043 3485 6055 3488
rect 5997 3479 6055 3485
rect 6089 3485 6101 3488
rect 6135 3485 6147 3519
rect 6748 3516 6776 3692
rect 6825 3519 6883 3525
rect 6825 3516 6837 3519
rect 6748 3488 6837 3516
rect 6089 3479 6147 3485
rect 6825 3485 6837 3488
rect 6871 3516 6883 3519
rect 8136 3519 8194 3525
rect 6871 3488 6960 3516
rect 6871 3485 6883 3488
rect 6825 3479 6883 3485
rect 2294 3451 2352 3457
rect 2294 3448 2306 3451
rect 1719 3420 1808 3448
rect 2148 3420 2306 3448
rect 1719 3417 1731 3420
rect 1673 3411 1731 3417
rect -1274 3340 -1268 3392
rect -1216 3380 -1210 3392
rect 569 3383 627 3389
rect 569 3380 581 3383
rect -1216 3352 581 3380
rect -1216 3340 -1210 3352
rect 569 3349 581 3352
rect 615 3349 627 3383
rect 569 3343 627 3349
rect 1857 3383 1915 3389
rect 1857 3349 1869 3383
rect 1903 3380 1915 3383
rect 2148 3380 2176 3420
rect 2294 3417 2306 3420
rect 2340 3417 2352 3451
rect 2294 3411 2352 3417
rect 1903 3352 2176 3380
rect 3398 3383 3456 3389
rect 1903 3349 1915 3352
rect 1857 3343 1915 3349
rect 3398 3349 3410 3383
rect 3444 3380 3456 3383
rect 4062 3380 4068 3392
rect 3444 3352 4068 3380
rect 3444 3349 3456 3352
rect 3398 3343 3456 3349
rect 4062 3340 4068 3352
rect 4120 3340 4126 3392
rect 6932 3380 6960 3488
rect 8136 3485 8148 3519
rect 8182 3516 8194 3519
rect 8182 3488 8340 3516
rect 8182 3485 8194 3488
rect 8136 3479 8194 3485
rect 7032 3383 7090 3389
rect 7032 3380 7044 3383
rect 6932 3352 7044 3380
rect 7032 3349 7044 3352
rect 7078 3349 7090 3383
rect 8312 3380 8340 3488
rect 8386 3476 8392 3528
rect 8444 3476 8450 3528
rect 9700 3519 9758 3525
rect 9700 3485 9712 3519
rect 9746 3516 9758 3519
rect 9746 3488 9858 3516
rect 9746 3485 9758 3488
rect 9700 3479 9758 3485
rect 9830 3448 9858 3488
rect 9950 3476 9956 3528
rect 10008 3476 10014 3528
rect 10502 3448 10508 3460
rect 9830 3420 10508 3448
rect 10502 3408 10508 3420
rect 10560 3408 10566 3460
rect 8596 3383 8654 3389
rect 8596 3380 8608 3383
rect 8312 3352 8608 3380
rect 7032 3343 7090 3349
rect 8596 3349 8608 3352
rect 8642 3349 8654 3383
rect 8596 3343 8654 3349
rect -1182 3136 -1176 3188
rect -1124 3176 -1118 3188
rect 569 3179 627 3185
rect 569 3176 581 3179
rect -1124 3148 581 3176
rect -1124 3136 -1118 3148
rect 569 3145 581 3148
rect 615 3145 627 3179
rect 569 3139 627 3145
rect 1857 3179 1915 3185
rect 1857 3145 1869 3179
rect 1903 3176 1915 3179
rect 3398 3179 3456 3185
rect 1903 3148 2176 3176
rect 1903 3145 1915 3148
rect 1857 3139 1915 3145
rect -2102 3068 -2096 3120
rect -2044 3108 -2038 3120
rect 1305 3111 1363 3117
rect 1305 3108 1317 3111
rect -2044 3080 1317 3108
rect -2044 3068 -2038 3080
rect 1305 3077 1317 3080
rect 1351 3077 1363 3111
rect 1305 3071 1363 3077
rect 1673 3111 1731 3117
rect 1673 3077 1685 3111
rect 1719 3108 1731 3111
rect 2148 3108 2176 3148
rect 3398 3145 3410 3179
rect 3444 3176 3456 3179
rect 4154 3176 4160 3188
rect 3444 3148 4160 3176
rect 3444 3145 3456 3148
rect 3398 3139 3456 3145
rect 4154 3136 4160 3148
rect 4212 3136 4218 3188
rect 7032 3179 7090 3185
rect 7032 3176 7044 3179
rect 6932 3148 7044 3176
rect 2294 3111 2352 3117
rect 2294 3108 2306 3111
rect 1719 3080 1808 3108
rect 2148 3080 2306 3108
rect 1719 3077 1731 3080
rect 1673 3071 1731 3077
rect -262 3000 -256 3052
rect -204 3040 -198 3052
rect 845 3043 903 3049
rect 845 3040 857 3043
rect -204 3012 857 3040
rect -204 3000 -198 3012
rect 845 3009 857 3012
rect 891 3009 903 3043
rect 845 3003 903 3009
rect 934 3000 940 3052
rect 992 3000 998 3052
rect 1578 2932 1584 2984
rect 1636 2932 1642 2984
rect 1780 2836 1808 3080
rect 2294 3077 2306 3080
rect 2340 3077 2352 3111
rect 2294 3071 2352 3077
rect 2038 3000 2044 3052
rect 2096 3000 2102 3052
rect 5534 3000 5540 3052
rect 5592 3040 5598 3052
rect 5997 3043 6055 3049
rect 5997 3040 6009 3043
rect 5592 3012 6009 3040
rect 5592 3000 5598 3012
rect 5997 3009 6009 3012
rect 6043 3040 6055 3043
rect 6089 3043 6147 3049
rect 6089 3040 6101 3043
rect 6043 3012 6101 3040
rect 6043 3009 6055 3012
rect 5997 3003 6055 3009
rect 6089 3009 6101 3012
rect 6135 3009 6147 3043
rect 6825 3043 6883 3049
rect 6825 3040 6837 3043
rect 6089 3003 6147 3009
rect 6748 3012 6837 3040
rect 6748 2836 6776 3012
rect 6825 3009 6837 3012
rect 6871 3040 6883 3043
rect 6932 3040 6960 3148
rect 7032 3145 7044 3148
rect 7078 3145 7090 3179
rect 8596 3179 8654 3185
rect 8596 3176 8608 3179
rect 7032 3139 7090 3145
rect 8312 3148 8608 3176
rect 6871 3012 6960 3040
rect 8136 3043 8194 3049
rect 6871 3009 6883 3012
rect 6825 3003 6883 3009
rect 8136 3009 8148 3043
rect 8182 3040 8194 3043
rect 8312 3040 8340 3148
rect 8596 3145 8608 3148
rect 8642 3145 8654 3179
rect 8596 3139 8654 3145
rect 10594 3108 10600 3120
rect 9830 3080 10600 3108
rect 8182 3012 8340 3040
rect 8182 3009 8194 3012
rect 8136 3003 8194 3009
rect 8386 3000 8392 3052
rect 8444 3000 8450 3052
rect 9700 3043 9758 3049
rect 9700 3009 9712 3043
rect 9746 3040 9758 3043
rect 9830 3040 9858 3080
rect 10594 3068 10600 3080
rect 10652 3068 10658 3120
rect 9746 3012 9858 3040
rect 9746 3009 9758 3012
rect 9700 3003 9758 3009
rect 9950 3000 9956 3052
rect 10008 3000 10014 3052
rect 1780 2808 6776 2836
rect 1780 2604 6776 2632
rect 1578 2456 1584 2508
rect 1636 2456 1642 2508
rect -170 2388 -164 2440
rect -112 2428 -106 2440
rect 845 2431 903 2437
rect 845 2428 857 2431
rect -112 2400 857 2428
rect -112 2388 -106 2400
rect 845 2397 857 2400
rect 891 2397 903 2431
rect 845 2391 903 2397
rect 934 2388 940 2440
rect 992 2388 998 2440
rect -2010 2320 -2004 2372
rect -1952 2360 -1946 2372
rect 1305 2363 1363 2369
rect 1305 2360 1317 2363
rect -1952 2332 1317 2360
rect -1952 2320 -1946 2332
rect 1305 2329 1317 2332
rect 1351 2329 1363 2363
rect 1305 2323 1363 2329
rect 1673 2363 1731 2369
rect 1673 2329 1685 2363
rect 1719 2360 1731 2363
rect 1780 2360 1808 2604
rect 2038 2388 2044 2440
rect 2096 2388 2102 2440
rect 5626 2388 5632 2440
rect 5684 2428 5690 2440
rect 5997 2431 6055 2437
rect 5997 2428 6009 2431
rect 5684 2400 6009 2428
rect 5684 2388 5690 2400
rect 5997 2397 6009 2400
rect 6043 2428 6055 2431
rect 6089 2431 6147 2437
rect 6089 2428 6101 2431
rect 6043 2400 6101 2428
rect 6043 2397 6055 2400
rect 5997 2391 6055 2397
rect 6089 2397 6101 2400
rect 6135 2397 6147 2431
rect 6748 2428 6776 2604
rect 6825 2431 6883 2437
rect 6825 2428 6837 2431
rect 6748 2400 6837 2428
rect 6089 2391 6147 2397
rect 6825 2397 6837 2400
rect 6871 2428 6883 2431
rect 8136 2431 8194 2437
rect 6871 2400 6960 2428
rect 6871 2397 6883 2400
rect 6825 2391 6883 2397
rect 2294 2363 2352 2369
rect 2294 2360 2306 2363
rect 1719 2332 1808 2360
rect 2148 2332 2306 2360
rect 1719 2329 1731 2332
rect 1673 2323 1731 2329
rect -1090 2252 -1084 2304
rect -1032 2292 -1026 2304
rect 569 2295 627 2301
rect 569 2292 581 2295
rect -1032 2264 581 2292
rect -1032 2252 -1026 2264
rect 569 2261 581 2264
rect 615 2261 627 2295
rect 569 2255 627 2261
rect 1857 2295 1915 2301
rect 1857 2261 1869 2295
rect 1903 2292 1915 2295
rect 2148 2292 2176 2332
rect 2294 2329 2306 2332
rect 2340 2329 2352 2363
rect 2294 2323 2352 2329
rect 1903 2264 2176 2292
rect 3398 2295 3456 2301
rect 1903 2261 1915 2264
rect 1857 2255 1915 2261
rect 3398 2261 3410 2295
rect 3444 2292 3456 2295
rect 4246 2292 4252 2304
rect 3444 2264 4252 2292
rect 3444 2261 3456 2264
rect 3398 2255 3456 2261
rect 4246 2252 4252 2264
rect 4304 2252 4310 2304
rect 6932 2292 6960 2400
rect 8136 2397 8148 2431
rect 8182 2428 8194 2431
rect 8182 2400 8340 2428
rect 8182 2397 8194 2400
rect 8136 2391 8194 2397
rect 7032 2295 7090 2301
rect 7032 2292 7044 2295
rect 6932 2264 7044 2292
rect 7032 2261 7044 2264
rect 7078 2261 7090 2295
rect 8312 2292 8340 2400
rect 8386 2388 8392 2440
rect 8444 2388 8450 2440
rect 9700 2431 9758 2437
rect 9700 2397 9712 2431
rect 9746 2428 9758 2431
rect 9746 2400 9858 2428
rect 9746 2397 9758 2400
rect 9700 2391 9758 2397
rect 9830 2360 9858 2400
rect 9950 2388 9956 2440
rect 10008 2388 10014 2440
rect 10686 2360 10692 2372
rect 9830 2332 10692 2360
rect 10686 2320 10692 2332
rect 10744 2320 10750 2372
rect 8596 2295 8654 2301
rect 8596 2292 8608 2295
rect 8312 2264 8608 2292
rect 7032 2255 7090 2261
rect 8596 2261 8608 2264
rect 8642 2261 8654 2295
rect 8596 2255 8654 2261
rect -998 2048 -992 2100
rect -940 2088 -934 2100
rect 569 2091 627 2097
rect 569 2088 581 2091
rect -940 2060 581 2088
rect -940 2048 -934 2060
rect 569 2057 581 2060
rect 615 2057 627 2091
rect 569 2051 627 2057
rect 1857 2091 1915 2097
rect 1857 2057 1869 2091
rect 1903 2088 1915 2091
rect 3398 2091 3456 2097
rect 1903 2060 2176 2088
rect 1903 2057 1915 2060
rect 1857 2051 1915 2057
rect -1918 1980 -1912 2032
rect -1860 2020 -1854 2032
rect 1305 2023 1363 2029
rect 1305 2020 1317 2023
rect -1860 1992 1317 2020
rect -1860 1980 -1854 1992
rect 1305 1989 1317 1992
rect 1351 1989 1363 2023
rect 1305 1983 1363 1989
rect 1673 2023 1731 2029
rect 1673 1989 1685 2023
rect 1719 2020 1731 2023
rect 2148 2020 2176 2060
rect 3398 2057 3410 2091
rect 3444 2088 3456 2091
rect 4338 2088 4344 2100
rect 3444 2060 4344 2088
rect 3444 2057 3456 2060
rect 3398 2051 3456 2057
rect 4338 2048 4344 2060
rect 4396 2048 4402 2100
rect 7032 2091 7090 2097
rect 7032 2088 7044 2091
rect 6932 2060 7044 2088
rect 2294 2023 2352 2029
rect 2294 2020 2306 2023
rect 1719 1992 1808 2020
rect 2148 1992 2306 2020
rect 1719 1989 1731 1992
rect 1673 1983 1731 1989
rect -78 1912 -72 1964
rect -20 1952 -14 1964
rect 845 1955 903 1961
rect 845 1952 857 1955
rect -20 1924 857 1952
rect -20 1912 -14 1924
rect 845 1921 857 1924
rect 891 1921 903 1955
rect 845 1915 903 1921
rect 934 1912 940 1964
rect 992 1912 998 1964
rect 1578 1844 1584 1896
rect 1636 1844 1642 1896
rect 1780 1748 1808 1992
rect 2294 1989 2306 1992
rect 2340 1989 2352 2023
rect 2294 1983 2352 1989
rect 2038 1912 2044 1964
rect 2096 1912 2102 1964
rect 5718 1912 5724 1964
rect 5776 1952 5782 1964
rect 5997 1955 6055 1961
rect 5997 1952 6009 1955
rect 5776 1924 6009 1952
rect 5776 1912 5782 1924
rect 5997 1921 6009 1924
rect 6043 1952 6055 1955
rect 6089 1955 6147 1961
rect 6089 1952 6101 1955
rect 6043 1924 6101 1952
rect 6043 1921 6055 1924
rect 5997 1915 6055 1921
rect 6089 1921 6101 1924
rect 6135 1921 6147 1955
rect 6825 1955 6883 1961
rect 6825 1952 6837 1955
rect 6089 1915 6147 1921
rect 6748 1924 6837 1952
rect 6748 1748 6776 1924
rect 6825 1921 6837 1924
rect 6871 1952 6883 1955
rect 6932 1952 6960 2060
rect 7032 2057 7044 2060
rect 7078 2057 7090 2091
rect 8596 2091 8654 2097
rect 8596 2088 8608 2091
rect 7032 2051 7090 2057
rect 8312 2060 8608 2088
rect 6871 1924 6960 1952
rect 8136 1955 8194 1961
rect 6871 1921 6883 1924
rect 6825 1915 6883 1921
rect 8136 1921 8148 1955
rect 8182 1952 8194 1955
rect 8312 1952 8340 2060
rect 8596 2057 8608 2060
rect 8642 2057 8654 2091
rect 8596 2051 8654 2057
rect 10778 2020 10784 2032
rect 9830 1992 10784 2020
rect 8182 1924 8340 1952
rect 8182 1921 8194 1924
rect 8136 1915 8194 1921
rect 8386 1912 8392 1964
rect 8444 1912 8450 1964
rect 9700 1955 9758 1961
rect 9700 1921 9712 1955
rect 9746 1952 9758 1955
rect 9830 1952 9858 1992
rect 10778 1980 10784 1992
rect 10836 1980 10842 2032
rect 9746 1924 9858 1952
rect 9746 1921 9758 1924
rect 9700 1915 9758 1921
rect 9950 1912 9956 1964
rect 10008 1912 10014 1964
rect 1780 1720 6776 1748
rect 5810 1300 5816 1352
rect 5868 1340 5874 1352
rect 5997 1343 6055 1349
rect 5997 1340 6009 1343
rect 5868 1312 6009 1340
rect 5868 1300 5874 1312
rect 5997 1309 6009 1312
rect 6043 1340 6055 1343
rect 6089 1343 6147 1349
rect 6089 1340 6101 1343
rect 6043 1312 6101 1340
rect 6043 1309 6055 1312
rect 5997 1303 6055 1309
rect 6089 1309 6101 1312
rect 6135 1309 6147 1343
rect 6089 1303 6147 1309
rect 6825 1343 6883 1349
rect 6825 1309 6837 1343
rect 6871 1340 6883 1343
rect 8136 1343 8194 1349
rect 6871 1312 6960 1340
rect 6871 1309 6883 1312
rect 6825 1303 6883 1309
rect 6932 1204 6960 1312
rect 8136 1309 8148 1343
rect 8182 1340 8194 1343
rect 8182 1312 8340 1340
rect 8182 1309 8194 1312
rect 8136 1303 8194 1309
rect 7032 1207 7090 1213
rect 7032 1204 7044 1207
rect 6932 1176 7044 1204
rect 7032 1173 7044 1176
rect 7078 1173 7090 1207
rect 8312 1204 8340 1312
rect 8386 1300 8392 1352
rect 8444 1300 8450 1352
rect 9700 1343 9758 1349
rect 9700 1309 9712 1343
rect 9746 1340 9758 1343
rect 9746 1312 9858 1340
rect 9746 1309 9758 1312
rect 9700 1303 9758 1309
rect 9830 1272 9858 1312
rect 9950 1300 9956 1352
rect 10008 1300 10014 1352
rect 10870 1272 10876 1284
rect 9830 1244 10876 1272
rect 10870 1232 10876 1244
rect 10928 1232 10934 1284
rect 8596 1207 8654 1213
rect 8596 1204 8608 1207
rect 8312 1176 8608 1204
rect 7032 1167 7090 1173
rect 8596 1173 8608 1176
rect 8642 1173 8654 1207
rect 8596 1167 8654 1173
rect 7032 1003 7090 1009
rect 7032 1000 7044 1003
rect 6932 972 7044 1000
rect 5902 824 5908 876
rect 5960 864 5966 876
rect 5997 867 6055 873
rect 5997 864 6009 867
rect 5960 836 6009 864
rect 5960 824 5966 836
rect 5997 833 6009 836
rect 6043 864 6055 867
rect 6089 867 6147 873
rect 6089 864 6101 867
rect 6043 836 6101 864
rect 6043 833 6055 836
rect 5997 827 6055 833
rect 6089 833 6101 836
rect 6135 833 6147 867
rect 6089 827 6147 833
rect 6825 867 6883 873
rect 6825 833 6837 867
rect 6871 864 6883 867
rect 6932 864 6960 972
rect 7032 969 7044 972
rect 7078 969 7090 1003
rect 8596 1003 8654 1009
rect 8596 1000 8608 1003
rect 7032 963 7090 969
rect 8312 972 8608 1000
rect 6871 836 6960 864
rect 8136 867 8194 873
rect 6871 833 6883 836
rect 6825 827 6883 833
rect 8136 833 8148 867
rect 8182 864 8194 867
rect 8312 864 8340 972
rect 8596 969 8608 972
rect 8642 969 8654 1003
rect 8596 963 8654 969
rect 10962 932 10968 944
rect 9830 904 10968 932
rect 8182 836 8340 864
rect 8182 833 8194 836
rect 8136 827 8194 833
rect 8386 824 8392 876
rect 8444 824 8450 876
rect 9700 867 9758 873
rect 9700 833 9712 867
rect 9746 864 9758 867
rect 9830 864 9858 904
rect 10962 892 10968 904
rect 11020 892 11026 944
rect 9746 836 9858 864
rect 9746 833 9758 836
rect 9700 827 9758 833
rect 9950 824 9956 876
rect 10008 824 10014 876
<< via1 >>
rect 0 8662 250 8746
rect 11176 8662 11426 8746
rect 2872 8551 2924 8560
rect 2872 8517 2881 8551
rect 2881 8517 2915 8551
rect 2915 8517 2924 8551
rect 2872 8508 2924 8517
rect 7656 8551 7708 8560
rect 7656 8517 7665 8551
rect 7665 8517 7699 8551
rect 7699 8517 7708 8551
rect 7656 8508 7708 8517
rect 9036 8551 9088 8560
rect 9036 8517 9045 8551
rect 9045 8517 9079 8551
rect 9079 8517 9088 8551
rect 9036 8508 9088 8517
rect 11060 8551 11112 8560
rect 11060 8517 11069 8551
rect 11069 8517 11103 8551
rect 11103 8517 11112 8551
rect 11060 8508 11112 8517
rect 2044 8483 2096 8492
rect 2044 8449 2053 8483
rect 2053 8449 2087 8483
rect 2087 8449 2096 8483
rect 2044 8440 2096 8449
rect 8392 8483 8444 8492
rect 8392 8449 8401 8483
rect 8401 8449 8435 8483
rect 8435 8449 8444 8483
rect 8392 8440 8444 8449
rect 9864 8483 9916 8492
rect 9864 8449 9873 8483
rect 9873 8449 9907 8483
rect 9907 8449 9916 8483
rect 9864 8440 9916 8449
rect 10232 8483 10284 8492
rect 10232 8449 10241 8483
rect 10241 8449 10275 8483
rect 10275 8449 10284 8483
rect 10232 8440 10284 8449
rect 350 8118 600 8202
rect 11526 8118 11776 8202
rect 4712 7828 4764 7880
rect 8392 7871 8444 7880
rect 8392 7837 8401 7871
rect 8401 7837 8435 7871
rect 8435 7837 8444 7871
rect 8392 7828 8444 7837
rect 9956 7871 10008 7880
rect 9956 7837 9965 7871
rect 9965 7837 9999 7871
rect 9999 7837 10008 7871
rect 9956 7828 10008 7837
rect 10416 7760 10468 7812
rect 0 7574 250 7658
rect 11176 7574 11426 7658
rect 4804 7352 4856 7404
rect 8392 7395 8444 7404
rect 8392 7361 8401 7395
rect 8401 7361 8435 7395
rect 8435 7361 8444 7395
rect 8392 7352 8444 7361
rect 10508 7420 10560 7472
rect 9956 7395 10008 7404
rect 9956 7361 9965 7395
rect 9965 7361 9999 7395
rect 9999 7361 10008 7395
rect 9956 7352 10008 7361
rect 350 7030 600 7114
rect 11526 7030 11776 7114
rect 1584 6808 1636 6860
rect -900 6740 -848 6792
rect 940 6783 992 6792
rect 940 6749 949 6783
rect 949 6749 983 6783
rect 983 6749 992 6783
rect 940 6740 992 6749
rect -2740 6672 -2688 6724
rect 2044 6783 2096 6792
rect 2044 6749 2053 6783
rect 2053 6749 2087 6783
rect 2087 6749 2096 6783
rect 2044 6740 2096 6749
rect 4896 6740 4948 6792
rect -1820 6604 -1768 6656
rect 3516 6604 3568 6656
rect 8392 6783 8444 6792
rect 8392 6749 8401 6783
rect 8401 6749 8435 6783
rect 8435 6749 8444 6783
rect 8392 6740 8444 6749
rect 9956 6783 10008 6792
rect 9956 6749 9965 6783
rect 9965 6749 9999 6783
rect 9999 6749 10008 6783
rect 9956 6740 10008 6749
rect 10600 6672 10652 6724
rect 0 6486 250 6570
rect 11176 6486 11426 6570
rect -1728 6400 -1676 6452
rect -2648 6332 -2596 6384
rect 3608 6400 3660 6452
rect -808 6264 -756 6316
rect 940 6307 992 6316
rect 940 6273 949 6307
rect 949 6273 983 6307
rect 983 6273 992 6307
rect 940 6264 992 6273
rect 1584 6196 1636 6248
rect 2044 6307 2096 6316
rect 2044 6273 2053 6307
rect 2053 6273 2087 6307
rect 2087 6273 2096 6307
rect 2044 6264 2096 6273
rect 4988 6264 5040 6316
rect 8392 6307 8444 6316
rect 8392 6273 8401 6307
rect 8401 6273 8435 6307
rect 8435 6273 8444 6307
rect 8392 6264 8444 6273
rect 10692 6332 10744 6384
rect 9956 6307 10008 6316
rect 9956 6273 9965 6307
rect 9965 6273 9999 6307
rect 9999 6273 10008 6307
rect 9956 6264 10008 6273
rect 350 5942 600 6026
rect 11526 5942 11776 6026
rect 1584 5720 1636 5772
rect -716 5652 -664 5704
rect 940 5695 992 5704
rect 940 5661 949 5695
rect 949 5661 983 5695
rect 983 5661 992 5695
rect 940 5652 992 5661
rect -2556 5584 -2504 5636
rect 2044 5695 2096 5704
rect 2044 5661 2053 5695
rect 2053 5661 2087 5695
rect 2087 5661 2096 5695
rect 2044 5652 2096 5661
rect 5080 5652 5132 5704
rect -1636 5516 -1584 5568
rect 3700 5516 3752 5568
rect 8392 5695 8444 5704
rect 8392 5661 8401 5695
rect 8401 5661 8435 5695
rect 8435 5661 8444 5695
rect 8392 5652 8444 5661
rect 9956 5695 10008 5704
rect 9956 5661 9965 5695
rect 9965 5661 9999 5695
rect 9999 5661 10008 5695
rect 9956 5652 10008 5661
rect 10784 5584 10836 5636
rect 0 5398 250 5482
rect 11176 5398 11426 5482
rect -1544 5312 -1492 5364
rect -2464 5244 -2412 5296
rect 3792 5312 3844 5364
rect -624 5176 -572 5228
rect 940 5219 992 5228
rect 940 5185 949 5219
rect 949 5185 983 5219
rect 983 5185 992 5219
rect 940 5176 992 5185
rect 1584 5108 1636 5160
rect 2044 5219 2096 5228
rect 2044 5185 2053 5219
rect 2053 5185 2087 5219
rect 2087 5185 2096 5219
rect 2044 5176 2096 5185
rect 5172 5176 5224 5228
rect 8392 5219 8444 5228
rect 8392 5185 8401 5219
rect 8401 5185 8435 5219
rect 8435 5185 8444 5219
rect 8392 5176 8444 5185
rect 10876 5244 10928 5296
rect 9956 5219 10008 5228
rect 9956 5185 9965 5219
rect 9965 5185 9999 5219
rect 9999 5185 10008 5219
rect 9956 5176 10008 5185
rect 350 4854 600 4938
rect 11526 4854 11776 4938
rect 1584 4632 1636 4684
rect -532 4564 -480 4616
rect 940 4607 992 4616
rect 940 4573 949 4607
rect 949 4573 983 4607
rect 983 4573 992 4607
rect 940 4564 992 4573
rect -2372 4496 -2320 4548
rect 2044 4607 2096 4616
rect 2044 4573 2053 4607
rect 2053 4573 2087 4607
rect 2087 4573 2096 4607
rect 2044 4564 2096 4573
rect 5264 4564 5316 4616
rect -1452 4428 -1400 4480
rect 3884 4428 3936 4480
rect 8392 4607 8444 4616
rect 8392 4573 8401 4607
rect 8401 4573 8435 4607
rect 8435 4573 8444 4607
rect 8392 4564 8444 4573
rect 9956 4607 10008 4616
rect 9956 4573 9965 4607
rect 9965 4573 9999 4607
rect 9999 4573 10008 4607
rect 9956 4564 10008 4573
rect 10968 4496 11020 4548
rect 0 4310 250 4394
rect 11176 4310 11426 4394
rect -1360 4224 -1308 4276
rect -2280 4156 -2228 4208
rect 3976 4224 4028 4276
rect -440 4088 -388 4140
rect 940 4131 992 4140
rect 940 4097 949 4131
rect 949 4097 983 4131
rect 983 4097 992 4131
rect 940 4088 992 4097
rect 1584 4020 1636 4072
rect 2044 4131 2096 4140
rect 2044 4097 2053 4131
rect 2053 4097 2087 4131
rect 2087 4097 2096 4131
rect 2044 4088 2096 4097
rect 5356 4088 5408 4140
rect 8392 4131 8444 4140
rect 8392 4097 8401 4131
rect 8401 4097 8435 4131
rect 8435 4097 8444 4131
rect 8392 4088 8444 4097
rect 10416 4156 10468 4208
rect 9956 4131 10008 4140
rect 9956 4097 9965 4131
rect 9965 4097 9999 4131
rect 9999 4097 10008 4131
rect 9956 4088 10008 4097
rect 350 3766 600 3850
rect 11526 3766 11776 3850
rect 1584 3544 1636 3596
rect -348 3476 -296 3528
rect 940 3519 992 3528
rect 940 3485 949 3519
rect 949 3485 983 3519
rect 983 3485 992 3519
rect 940 3476 992 3485
rect -2188 3408 -2136 3460
rect 2044 3519 2096 3528
rect 2044 3485 2053 3519
rect 2053 3485 2087 3519
rect 2087 3485 2096 3519
rect 2044 3476 2096 3485
rect 5448 3476 5500 3528
rect -1268 3340 -1216 3392
rect 4068 3340 4120 3392
rect 8392 3519 8444 3528
rect 8392 3485 8401 3519
rect 8401 3485 8435 3519
rect 8435 3485 8444 3519
rect 8392 3476 8444 3485
rect 9956 3519 10008 3528
rect 9956 3485 9965 3519
rect 9965 3485 9999 3519
rect 9999 3485 10008 3519
rect 9956 3476 10008 3485
rect 10508 3408 10560 3460
rect 0 3222 250 3306
rect 11176 3222 11426 3306
rect -1176 3136 -1124 3188
rect -2096 3068 -2044 3120
rect 4160 3136 4212 3188
rect -256 3000 -204 3052
rect 940 3043 992 3052
rect 940 3009 949 3043
rect 949 3009 983 3043
rect 983 3009 992 3043
rect 940 3000 992 3009
rect 1584 2932 1636 2984
rect 2044 3043 2096 3052
rect 2044 3009 2053 3043
rect 2053 3009 2087 3043
rect 2087 3009 2096 3043
rect 2044 3000 2096 3009
rect 5540 3000 5592 3052
rect 8392 3043 8444 3052
rect 8392 3009 8401 3043
rect 8401 3009 8435 3043
rect 8435 3009 8444 3043
rect 8392 3000 8444 3009
rect 10600 3068 10652 3120
rect 9956 3043 10008 3052
rect 9956 3009 9965 3043
rect 9965 3009 9999 3043
rect 9999 3009 10008 3043
rect 9956 3000 10008 3009
rect 350 2678 600 2762
rect 11526 2678 11776 2762
rect 1584 2456 1636 2508
rect -164 2388 -112 2440
rect 940 2431 992 2440
rect 940 2397 949 2431
rect 949 2397 983 2431
rect 983 2397 992 2431
rect 940 2388 992 2397
rect -2004 2320 -1952 2372
rect 2044 2431 2096 2440
rect 2044 2397 2053 2431
rect 2053 2397 2087 2431
rect 2087 2397 2096 2431
rect 2044 2388 2096 2397
rect 5632 2388 5684 2440
rect -1084 2252 -1032 2304
rect 4252 2252 4304 2304
rect 8392 2431 8444 2440
rect 8392 2397 8401 2431
rect 8401 2397 8435 2431
rect 8435 2397 8444 2431
rect 8392 2388 8444 2397
rect 9956 2431 10008 2440
rect 9956 2397 9965 2431
rect 9965 2397 9999 2431
rect 9999 2397 10008 2431
rect 9956 2388 10008 2397
rect 10692 2320 10744 2372
rect 0 2134 250 2218
rect 11176 2134 11426 2218
rect -992 2048 -940 2100
rect -1912 1980 -1860 2032
rect 4344 2048 4396 2100
rect -72 1912 -20 1964
rect 940 1955 992 1964
rect 940 1921 949 1955
rect 949 1921 983 1955
rect 983 1921 992 1955
rect 940 1912 992 1921
rect 1584 1844 1636 1896
rect 2044 1955 2096 1964
rect 2044 1921 2053 1955
rect 2053 1921 2087 1955
rect 2087 1921 2096 1955
rect 2044 1912 2096 1921
rect 5724 1912 5776 1964
rect 8392 1955 8444 1964
rect 8392 1921 8401 1955
rect 8401 1921 8435 1955
rect 8435 1921 8444 1955
rect 8392 1912 8444 1921
rect 10784 1980 10836 2032
rect 9956 1955 10008 1964
rect 9956 1921 9965 1955
rect 9965 1921 9999 1955
rect 9999 1921 10008 1955
rect 9956 1912 10008 1921
rect 350 1590 600 1674
rect 11526 1590 11776 1674
rect 5816 1300 5868 1352
rect 8392 1343 8444 1352
rect 8392 1309 8401 1343
rect 8401 1309 8435 1343
rect 8435 1309 8444 1343
rect 8392 1300 8444 1309
rect 9956 1343 10008 1352
rect 9956 1309 9965 1343
rect 9965 1309 9999 1343
rect 9999 1309 10008 1343
rect 9956 1300 10008 1309
rect 10876 1232 10928 1284
rect 0 1046 250 1130
rect 11176 1046 11426 1130
rect 5908 824 5960 876
rect 8392 867 8444 876
rect 8392 833 8401 867
rect 8401 833 8435 867
rect 8435 833 8444 867
rect 8392 824 8444 833
rect 10968 892 11020 944
rect 9956 867 10008 876
rect 9956 833 9965 867
rect 9965 833 9999 867
rect 9999 833 10008 867
rect 9956 824 10008 833
rect 350 502 600 586
rect 11526 502 11776 586
rect 0 -42 250 42
rect 11176 -42 11426 42
<< metal2 >>
rect 0 8746 250 8752
rect 0 8656 250 8662
rect 350 8202 600 8208
rect 350 8112 600 8118
rect 0 7658 250 7664
rect 0 7568 250 7574
rect 350 7114 600 7120
rect 350 7024 600 7030
rect 952 6798 980 8820
rect 1596 6866 1624 8820
rect 2884 8566 2912 8820
rect 2872 8560 2924 8566
rect 2872 8502 2924 8508
rect 2044 8492 2096 8498
rect 2044 8434 2096 8440
rect 1584 6860 1636 6866
rect 1584 6802 1636 6808
rect -900 6792 -848 6798
rect -900 6734 -848 6740
rect 940 6792 992 6798
rect 940 6734 992 6740
rect -2740 6724 -2688 6730
rect -2740 6666 -2688 6672
rect -2728 -116 -2700 6666
rect -1820 6656 -1768 6662
rect -1820 6598 -1768 6604
rect -2648 6384 -2596 6390
rect -2648 6326 -2596 6332
rect -2636 -116 -2608 6326
rect -2556 5636 -2504 5642
rect -2556 5578 -2504 5584
rect -2544 -116 -2516 5578
rect -2464 5296 -2412 5302
rect -2464 5238 -2412 5244
rect -2452 -116 -2424 5238
rect -2372 4548 -2320 4554
rect -2372 4490 -2320 4496
rect -2360 -116 -2332 4490
rect -2280 4208 -2228 4214
rect -2280 4150 -2228 4156
rect -2268 -116 -2240 4150
rect -2188 3460 -2136 3466
rect -2188 3402 -2136 3408
rect -2176 -116 -2148 3402
rect -2096 3120 -2044 3126
rect -2096 3062 -2044 3068
rect -2084 -116 -2056 3062
rect -2004 2372 -1952 2378
rect -2004 2314 -1952 2320
rect -1992 -116 -1964 2314
rect -1912 2032 -1860 2038
rect -1912 1974 -1860 1980
rect -1900 -116 -1872 1974
rect -1808 -116 -1780 6598
rect -1728 6452 -1676 6458
rect -1728 6394 -1676 6400
rect -1716 -116 -1688 6394
rect -1636 5568 -1584 5574
rect -1636 5510 -1584 5516
rect -1624 -116 -1596 5510
rect -1544 5364 -1492 5370
rect -1544 5306 -1492 5312
rect -1532 -116 -1504 5306
rect -1452 4480 -1400 4486
rect -1452 4422 -1400 4428
rect -1440 -116 -1412 4422
rect -1360 4276 -1308 4282
rect -1360 4218 -1308 4224
rect -1348 -116 -1320 4218
rect -1268 3392 -1216 3398
rect -1268 3334 -1216 3340
rect -1256 -116 -1228 3334
rect -1176 3188 -1124 3194
rect -1176 3130 -1124 3136
rect -1164 -116 -1136 3130
rect -1084 2304 -1032 2310
rect -1084 2246 -1032 2252
rect -1072 -116 -1044 2246
rect -992 2100 -940 2106
rect -992 2042 -940 2048
rect -980 -116 -952 2042
rect -888 -116 -860 6734
rect 0 6570 250 6576
rect 0 6480 250 6486
rect 952 6322 980 6734
rect -808 6316 -756 6322
rect -808 6258 -756 6264
rect 940 6316 992 6322
rect 940 6258 992 6264
rect -796 -116 -768 6258
rect 350 6026 600 6032
rect 350 5936 600 5942
rect 952 5710 980 6258
rect 1596 6254 1624 6802
rect 2056 6798 2084 8434
rect 2044 6792 2096 6798
rect 2044 6734 2096 6740
rect 2056 6322 2084 6734
rect 3528 6662 3556 8820
rect 3516 6656 3568 6662
rect 3516 6598 3568 6604
rect 3620 6458 3648 8820
rect 3608 6452 3660 6458
rect 3608 6394 3660 6400
rect 2044 6316 2096 6322
rect 2044 6258 2096 6264
rect 1584 6248 1636 6254
rect 1584 6190 1636 6196
rect 1596 5778 1624 6190
rect 1584 5772 1636 5778
rect 1584 5714 1636 5720
rect -716 5704 -664 5710
rect -716 5646 -664 5652
rect 940 5704 992 5710
rect 940 5646 992 5652
rect -704 -116 -676 5646
rect 0 5482 250 5488
rect 0 5392 250 5398
rect 952 5234 980 5646
rect -624 5228 -572 5234
rect -624 5170 -572 5176
rect 940 5228 992 5234
rect 940 5170 992 5176
rect -612 -116 -584 5170
rect 350 4938 600 4944
rect 350 4848 600 4854
rect 952 4622 980 5170
rect 1596 5166 1624 5714
rect 2056 5710 2084 6258
rect 2044 5704 2096 5710
rect 2044 5646 2096 5652
rect 2056 5234 2084 5646
rect 3712 5574 3740 8820
rect 3700 5568 3752 5574
rect 3700 5510 3752 5516
rect 3804 5370 3832 8820
rect 3792 5364 3844 5370
rect 3792 5306 3844 5312
rect 2044 5228 2096 5234
rect 2044 5170 2096 5176
rect 1584 5160 1636 5166
rect 1584 5102 1636 5108
rect 1596 4690 1624 5102
rect 1584 4684 1636 4690
rect 1584 4626 1636 4632
rect -532 4616 -480 4622
rect -532 4558 -480 4564
rect 940 4616 992 4622
rect 940 4558 992 4564
rect -520 -116 -492 4558
rect 0 4394 250 4400
rect 0 4304 250 4310
rect 952 4146 980 4558
rect -440 4140 -388 4146
rect -440 4082 -388 4088
rect 940 4140 992 4146
rect 940 4082 992 4088
rect -428 -116 -400 4082
rect 350 3850 600 3856
rect 350 3760 600 3766
rect 952 3534 980 4082
rect 1596 4078 1624 4626
rect 2056 4622 2084 5170
rect 2044 4616 2096 4622
rect 2044 4558 2096 4564
rect 2056 4146 2084 4558
rect 3896 4486 3924 8820
rect 3884 4480 3936 4486
rect 3884 4422 3936 4428
rect 3988 4282 4016 8820
rect 3976 4276 4028 4282
rect 3976 4218 4028 4224
rect 2044 4140 2096 4146
rect 2044 4082 2096 4088
rect 1584 4072 1636 4078
rect 1584 4014 1636 4020
rect 1596 3602 1624 4014
rect 1584 3596 1636 3602
rect 1584 3538 1636 3544
rect -348 3528 -296 3534
rect -348 3470 -296 3476
rect 940 3528 992 3534
rect 940 3470 992 3476
rect -336 -116 -308 3470
rect 0 3306 250 3312
rect 0 3216 250 3222
rect 952 3058 980 3470
rect -256 3052 -204 3058
rect -256 2994 -204 3000
rect 940 3052 992 3058
rect 940 2994 992 3000
rect -244 -116 -216 2994
rect 350 2762 600 2768
rect 350 2672 600 2678
rect 952 2446 980 2994
rect 1596 2990 1624 3538
rect 2056 3534 2084 4082
rect 2044 3528 2096 3534
rect 2044 3470 2096 3476
rect 2056 3058 2084 3470
rect 4080 3398 4108 8820
rect 4068 3392 4120 3398
rect 4068 3334 4120 3340
rect 4172 3194 4200 8820
rect 4160 3188 4212 3194
rect 4160 3130 4212 3136
rect 2044 3052 2096 3058
rect 2044 2994 2096 3000
rect 1584 2984 1636 2990
rect 1584 2926 1636 2932
rect 1596 2514 1624 2926
rect 1584 2508 1636 2514
rect 1584 2450 1636 2456
rect -164 2440 -112 2446
rect -164 2382 -112 2388
rect 940 2440 992 2446
rect 940 2382 992 2388
rect -152 -116 -124 2382
rect 0 2218 250 2224
rect 0 2128 250 2134
rect 952 1970 980 2382
rect -72 1964 -20 1970
rect -72 1906 -20 1912
rect 940 1964 992 1970
rect 940 1906 992 1912
rect -60 -116 -32 1906
rect 1596 1902 1624 2450
rect 2056 2446 2084 2994
rect 2044 2440 2096 2446
rect 2044 2382 2096 2388
rect 2056 1970 2084 2382
rect 4264 2310 4292 8820
rect 4252 2304 4304 2310
rect 4252 2246 4304 2252
rect 4356 2106 4384 8820
rect 7668 8566 7696 8820
rect 9048 8566 9076 8820
rect 7656 8560 7708 8566
rect 7656 8502 7708 8508
rect 9036 8560 9088 8566
rect 9036 8502 9088 8508
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 9864 8492 9916 8498
rect 9864 8434 9916 8440
rect 10232 8492 10284 8498
rect 10232 8434 10284 8440
rect 8404 7886 8432 8434
rect 4712 7880 4764 7886
rect 4712 7822 4764 7828
rect 8392 7880 8444 7886
rect 8392 7822 8444 7828
rect 9876 7868 9904 8434
rect 9950 7868 9956 7880
rect 9876 7840 9956 7868
rect 4344 2100 4396 2106
rect 4344 2042 4396 2048
rect 2044 1964 2096 1970
rect 2044 1906 2096 1912
rect 1584 1896 1636 1902
rect 1584 1838 1636 1844
rect 350 1674 600 1680
rect 350 1584 600 1590
rect 0 1130 250 1136
rect 0 1040 250 1046
rect 350 586 600 592
rect 350 496 600 502
rect 0 42 250 48
rect 0 -48 250 -42
rect 4724 -116 4752 7822
rect 8404 7410 8432 7822
rect 4804 7404 4856 7410
rect 4804 7346 4856 7352
rect 8392 7404 8444 7410
rect 8392 7346 8444 7352
rect 9876 7392 9904 7840
rect 9950 7828 9956 7840
rect 10008 7828 10014 7880
rect 9950 7392 9956 7404
rect 9876 7364 9956 7392
rect 4816 -116 4844 7346
rect 8404 6798 8432 7346
rect 4896 6792 4948 6798
rect 4896 6734 4948 6740
rect 8392 6792 8444 6798
rect 8392 6734 8444 6740
rect 9876 6780 9904 7364
rect 9950 7352 9956 7364
rect 10008 7352 10014 7404
rect 9950 6780 9956 6792
rect 9876 6752 9956 6780
rect 4908 -116 4936 6734
rect 8404 6322 8432 6734
rect 4988 6316 5040 6322
rect 4988 6258 5040 6264
rect 8392 6316 8444 6322
rect 8392 6258 8444 6264
rect 9876 6304 9904 6752
rect 9950 6740 9956 6752
rect 10008 6740 10014 6792
rect 9950 6304 9956 6316
rect 9876 6276 9956 6304
rect 5000 -116 5028 6258
rect 8404 5710 8432 6258
rect 5080 5704 5132 5710
rect 5080 5646 5132 5652
rect 8392 5704 8444 5710
rect 8392 5646 8444 5652
rect 9876 5692 9904 6276
rect 9950 6264 9956 6276
rect 10008 6264 10014 6316
rect 9950 5692 9956 5704
rect 9876 5664 9956 5692
rect 5092 -116 5120 5646
rect 8404 5234 8432 5646
rect 5172 5228 5224 5234
rect 5172 5170 5224 5176
rect 8392 5228 8444 5234
rect 8392 5170 8444 5176
rect 9876 5216 9904 5664
rect 9950 5652 9956 5664
rect 10008 5652 10014 5704
rect 9950 5216 9956 5228
rect 9876 5188 9956 5216
rect 5184 -116 5212 5170
rect 8404 4622 8432 5170
rect 5264 4616 5316 4622
rect 5264 4558 5316 4564
rect 8392 4616 8444 4622
rect 9876 4604 9904 5188
rect 9950 5176 9956 5188
rect 10008 5176 10014 5228
rect 9950 4604 9956 4616
rect 9876 4576 9956 4604
rect 9950 4564 9956 4576
rect 10008 4564 10014 4616
rect 8392 4558 8444 4564
rect 5276 -116 5304 4558
rect 8404 4146 8432 4558
rect 5356 4140 5408 4146
rect 5356 4082 5408 4088
rect 8392 4140 8444 4146
rect 9950 4088 9956 4140
rect 10008 4128 10014 4140
rect 10244 4128 10272 8434
rect 10428 7818 10456 8820
rect 10416 7812 10468 7818
rect 10416 7754 10468 7760
rect 10428 4214 10456 7754
rect 10520 7478 10548 8820
rect 10508 7472 10560 7478
rect 10508 7414 10560 7420
rect 10416 4208 10468 4214
rect 10416 4150 10468 4156
rect 10008 4100 10272 4128
rect 10008 4088 10014 4100
rect 8392 4082 8444 4088
rect 5368 -116 5396 4082
rect 8404 3534 8432 4082
rect 5448 3528 5500 3534
rect 5448 3470 5500 3476
rect 8392 3528 8444 3534
rect 9950 3476 9956 3528
rect 10008 3516 10014 3528
rect 10244 3516 10272 4100
rect 10008 3488 10272 3516
rect 10008 3476 10014 3488
rect 8392 3470 8444 3476
rect 5460 -116 5488 3470
rect 8404 3058 8432 3470
rect 5540 3052 5592 3058
rect 5540 2994 5592 3000
rect 8392 3052 8444 3058
rect 9950 3000 9956 3052
rect 10008 3040 10014 3052
rect 10244 3040 10272 3488
rect 10520 3466 10548 7414
rect 10612 6730 10640 8820
rect 10600 6724 10652 6730
rect 10600 6666 10652 6672
rect 10508 3460 10560 3466
rect 10508 3402 10560 3408
rect 10612 3126 10640 6666
rect 10704 6390 10732 8820
rect 10692 6384 10744 6390
rect 10692 6326 10744 6332
rect 10600 3120 10652 3126
rect 10600 3062 10652 3068
rect 10008 3012 10272 3040
rect 10008 3000 10014 3012
rect 8392 2994 8444 3000
rect 5552 -116 5580 2994
rect 8404 2446 8432 2994
rect 5632 2440 5684 2446
rect 5632 2382 5684 2388
rect 8392 2440 8444 2446
rect 9950 2388 9956 2440
rect 10008 2428 10014 2440
rect 10244 2428 10272 3012
rect 10008 2400 10272 2428
rect 10008 2388 10014 2400
rect 8392 2382 8444 2388
rect 5644 -116 5672 2382
rect 8404 1970 8432 2382
rect 5724 1964 5776 1970
rect 5724 1906 5776 1912
rect 8392 1964 8444 1970
rect 9950 1912 9956 1964
rect 10008 1952 10014 1964
rect 10244 1952 10272 2400
rect 10704 2378 10732 6326
rect 10796 5642 10824 8820
rect 10784 5636 10836 5642
rect 10784 5578 10836 5584
rect 10692 2372 10744 2378
rect 10692 2314 10744 2320
rect 10796 2038 10824 5578
rect 10888 5302 10916 8820
rect 10876 5296 10928 5302
rect 10876 5238 10928 5244
rect 10784 2032 10836 2038
rect 10784 1974 10836 1980
rect 10008 1924 10272 1952
rect 10008 1912 10014 1924
rect 8392 1906 8444 1912
rect 5736 -116 5764 1906
rect 8404 1358 8432 1906
rect 5816 1352 5868 1358
rect 5816 1294 5868 1300
rect 8392 1352 8444 1358
rect 9950 1300 9956 1352
rect 10008 1340 10014 1352
rect 10244 1340 10272 1924
rect 10008 1312 10272 1340
rect 10008 1300 10014 1312
rect 8392 1294 8444 1300
rect 5828 -116 5856 1294
rect 8404 882 8432 1294
rect 5908 876 5960 882
rect 5908 818 5960 824
rect 8392 876 8444 882
rect 9950 824 9956 876
rect 10008 864 10014 876
rect 10244 864 10272 1312
rect 10888 1290 10916 5238
rect 10980 4554 11008 8820
rect 11072 8566 11100 8820
rect 11176 8746 11426 8752
rect 11176 8656 11426 8662
rect 11060 8560 11112 8566
rect 11060 8502 11112 8508
rect 11526 8202 11776 8208
rect 11526 8112 11776 8118
rect 11176 7658 11426 7664
rect 11176 7568 11426 7574
rect 11526 7114 11776 7120
rect 11526 7024 11776 7030
rect 11176 6570 11426 6576
rect 11176 6480 11426 6486
rect 11526 6026 11776 6032
rect 11526 5936 11776 5942
rect 11176 5482 11426 5488
rect 11176 5392 11426 5398
rect 11526 4938 11776 4944
rect 11526 4848 11776 4854
rect 10968 4548 11020 4554
rect 10968 4490 11020 4496
rect 10876 1284 10928 1290
rect 10876 1226 10928 1232
rect 10980 950 11008 4490
rect 11176 4394 11426 4400
rect 11176 4304 11426 4310
rect 11526 3850 11776 3856
rect 11526 3760 11776 3766
rect 11176 3306 11426 3312
rect 11176 3216 11426 3222
rect 11526 2762 11776 2768
rect 11526 2672 11776 2678
rect 11176 2218 11426 2224
rect 11176 2128 11426 2134
rect 11526 1674 11776 1680
rect 11526 1584 11776 1590
rect 11176 1130 11426 1136
rect 11176 1040 11426 1046
rect 10968 944 11020 950
rect 10968 886 11020 892
rect 10008 836 10272 864
rect 10008 824 10014 836
rect 8392 818 8444 824
rect 5920 -116 5948 818
rect 11526 586 11776 592
rect 11526 496 11776 502
rect 11176 42 11426 48
rect 11176 -48 11426 -42
<< via2 >>
rect 5 8665 245 8743
rect 355 8121 595 8199
rect 5 7577 245 7655
rect 355 7033 595 7111
rect 5 6489 245 6567
rect 355 5945 595 6023
rect 5 5401 245 5479
rect 355 4857 595 4935
rect 5 4313 245 4391
rect 355 3769 595 3847
rect 5 3225 245 3303
rect 355 2681 595 2759
rect 5 2137 245 2215
rect 355 1593 595 1671
rect 5 1049 245 1127
rect 355 505 595 583
rect 5 -39 245 39
rect 11181 8665 11421 8743
rect 11531 8121 11771 8199
rect 11181 7577 11421 7655
rect 11531 7033 11771 7111
rect 11181 6489 11421 6567
rect 11531 5945 11771 6023
rect 11181 5401 11421 5479
rect 11531 4857 11771 4935
rect 11181 4313 11421 4391
rect 11531 3769 11771 3847
rect 11181 3225 11421 3303
rect 11531 2681 11771 2759
rect 11181 2137 11421 2215
rect 11531 1593 11771 1671
rect 11181 1049 11421 1127
rect 11531 505 11771 583
rect 11181 -39 11421 39
<< metal3 >>
rect 0 8746 250 8752
rect 0 8662 1 8746
rect 249 8662 250 8746
rect 0 8656 250 8662
rect 11176 8746 11426 8752
rect 11176 8662 11177 8746
rect 11425 8662 11426 8746
rect 11176 8656 11426 8662
rect 350 8202 600 8208
rect 350 8118 351 8202
rect 599 8118 600 8202
rect 350 8112 600 8118
rect 11526 8202 11776 8208
rect 11526 8118 11527 8202
rect 11775 8118 11776 8202
rect 11526 8112 11776 8118
rect 0 7658 250 7664
rect 0 7574 1 7658
rect 249 7574 250 7658
rect 0 7568 250 7574
rect 11176 7658 11426 7664
rect 11176 7574 11177 7658
rect 11425 7574 11426 7658
rect 11176 7568 11426 7574
rect 350 7114 600 7120
rect 350 7030 351 7114
rect 599 7030 600 7114
rect 350 7024 600 7030
rect 11526 7114 11776 7120
rect 11526 7030 11527 7114
rect 11775 7030 11776 7114
rect 11526 7024 11776 7030
rect 0 6570 250 6576
rect 0 6486 1 6570
rect 249 6486 250 6570
rect 0 6480 250 6486
rect 11176 6570 11426 6576
rect 11176 6486 11177 6570
rect 11425 6486 11426 6570
rect 11176 6480 11426 6486
rect 350 6026 600 6032
rect 350 5942 351 6026
rect 599 5942 600 6026
rect 350 5936 600 5942
rect 11526 6026 11776 6032
rect 11526 5942 11527 6026
rect 11775 5942 11776 6026
rect 11526 5936 11776 5942
rect 0 5482 250 5488
rect 0 5398 1 5482
rect 249 5398 250 5482
rect 0 5392 250 5398
rect 11176 5482 11426 5488
rect 11176 5398 11177 5482
rect 11425 5398 11426 5482
rect 11176 5392 11426 5398
rect 350 4938 600 4944
rect 350 4854 351 4938
rect 599 4854 600 4938
rect 350 4848 600 4854
rect 11526 4938 11776 4944
rect 11526 4854 11527 4938
rect 11775 4854 11776 4938
rect 11526 4848 11776 4854
rect 0 4394 250 4400
rect 0 4310 1 4394
rect 249 4310 250 4394
rect 0 4304 250 4310
rect 11176 4394 11426 4400
rect 11176 4310 11177 4394
rect 11425 4310 11426 4394
rect 11176 4304 11426 4310
rect 350 3850 600 3856
rect 350 3766 351 3850
rect 599 3766 600 3850
rect 350 3760 600 3766
rect 11526 3850 11776 3856
rect 11526 3766 11527 3850
rect 11775 3766 11776 3850
rect 11526 3760 11776 3766
rect 0 3306 250 3312
rect 0 3222 1 3306
rect 249 3222 250 3306
rect 0 3216 250 3222
rect 11176 3306 11426 3312
rect 11176 3222 11177 3306
rect 11425 3222 11426 3306
rect 11176 3216 11426 3222
rect 350 2762 600 2768
rect 350 2678 351 2762
rect 599 2678 600 2762
rect 350 2672 600 2678
rect 11526 2762 11776 2768
rect 11526 2678 11527 2762
rect 11775 2678 11776 2762
rect 11526 2672 11776 2678
rect 0 2218 250 2224
rect 0 2134 1 2218
rect 249 2134 250 2218
rect 0 2128 250 2134
rect 11176 2218 11426 2224
rect 11176 2134 11177 2218
rect 11425 2134 11426 2218
rect 11176 2128 11426 2134
rect 350 1674 600 1680
rect 350 1590 351 1674
rect 599 1590 600 1674
rect 350 1584 600 1590
rect 11526 1674 11776 1680
rect 11526 1590 11527 1674
rect 11775 1590 11776 1674
rect 11526 1584 11776 1590
rect 0 1130 250 1136
rect 0 1046 1 1130
rect 249 1046 250 1130
rect 0 1040 250 1046
rect 11176 1130 11426 1136
rect 11176 1046 11177 1130
rect 11425 1046 11426 1130
rect 11176 1040 11426 1046
rect 350 586 600 592
rect 350 502 351 586
rect 599 502 600 586
rect 350 496 600 502
rect 11526 586 11776 592
rect 11526 502 11527 586
rect 11775 502 11776 586
rect 11526 496 11776 502
rect 0 42 250 48
rect 0 -42 1 42
rect 249 -42 250 42
rect 0 -48 250 -42
rect 11176 42 11426 48
rect 11176 -42 11177 42
rect 11425 -42 11426 42
rect 11176 -48 11426 -42
<< via3 >>
rect 1 8743 249 8746
rect 1 8665 5 8743
rect 5 8665 245 8743
rect 245 8665 249 8743
rect 1 8662 249 8665
rect 11177 8743 11425 8746
rect 11177 8665 11181 8743
rect 11181 8665 11421 8743
rect 11421 8665 11425 8743
rect 11177 8662 11425 8665
rect 351 8199 599 8202
rect 351 8121 355 8199
rect 355 8121 595 8199
rect 595 8121 599 8199
rect 351 8118 599 8121
rect 11527 8199 11775 8202
rect 11527 8121 11531 8199
rect 11531 8121 11771 8199
rect 11771 8121 11775 8199
rect 11527 8118 11775 8121
rect 1 7655 249 7658
rect 1 7577 5 7655
rect 5 7577 245 7655
rect 245 7577 249 7655
rect 1 7574 249 7577
rect 11177 7655 11425 7658
rect 11177 7577 11181 7655
rect 11181 7577 11421 7655
rect 11421 7577 11425 7655
rect 11177 7574 11425 7577
rect 351 7111 599 7114
rect 351 7033 355 7111
rect 355 7033 595 7111
rect 595 7033 599 7111
rect 351 7030 599 7033
rect 11527 7111 11775 7114
rect 11527 7033 11531 7111
rect 11531 7033 11771 7111
rect 11771 7033 11775 7111
rect 11527 7030 11775 7033
rect 1 6567 249 6570
rect 1 6489 5 6567
rect 5 6489 245 6567
rect 245 6489 249 6567
rect 1 6486 249 6489
rect 11177 6567 11425 6570
rect 11177 6489 11181 6567
rect 11181 6489 11421 6567
rect 11421 6489 11425 6567
rect 11177 6486 11425 6489
rect 351 6023 599 6026
rect 351 5945 355 6023
rect 355 5945 595 6023
rect 595 5945 599 6023
rect 351 5942 599 5945
rect 11527 6023 11775 6026
rect 11527 5945 11531 6023
rect 11531 5945 11771 6023
rect 11771 5945 11775 6023
rect 11527 5942 11775 5945
rect 1 5479 249 5482
rect 1 5401 5 5479
rect 5 5401 245 5479
rect 245 5401 249 5479
rect 1 5398 249 5401
rect 11177 5479 11425 5482
rect 11177 5401 11181 5479
rect 11181 5401 11421 5479
rect 11421 5401 11425 5479
rect 11177 5398 11425 5401
rect 351 4935 599 4938
rect 351 4857 355 4935
rect 355 4857 595 4935
rect 595 4857 599 4935
rect 351 4854 599 4857
rect 11527 4935 11775 4938
rect 11527 4857 11531 4935
rect 11531 4857 11771 4935
rect 11771 4857 11775 4935
rect 11527 4854 11775 4857
rect 1 4391 249 4394
rect 1 4313 5 4391
rect 5 4313 245 4391
rect 245 4313 249 4391
rect 1 4310 249 4313
rect 11177 4391 11425 4394
rect 11177 4313 11181 4391
rect 11181 4313 11421 4391
rect 11421 4313 11425 4391
rect 11177 4310 11425 4313
rect 351 3847 599 3850
rect 351 3769 355 3847
rect 355 3769 595 3847
rect 595 3769 599 3847
rect 351 3766 599 3769
rect 11527 3847 11775 3850
rect 11527 3769 11531 3847
rect 11531 3769 11771 3847
rect 11771 3769 11775 3847
rect 11527 3766 11775 3769
rect 1 3303 249 3306
rect 1 3225 5 3303
rect 5 3225 245 3303
rect 245 3225 249 3303
rect 1 3222 249 3225
rect 11177 3303 11425 3306
rect 11177 3225 11181 3303
rect 11181 3225 11421 3303
rect 11421 3225 11425 3303
rect 11177 3222 11425 3225
rect 351 2759 599 2762
rect 351 2681 355 2759
rect 355 2681 595 2759
rect 595 2681 599 2759
rect 351 2678 599 2681
rect 11527 2759 11775 2762
rect 11527 2681 11531 2759
rect 11531 2681 11771 2759
rect 11771 2681 11775 2759
rect 11527 2678 11775 2681
rect 1 2215 249 2218
rect 1 2137 5 2215
rect 5 2137 245 2215
rect 245 2137 249 2215
rect 1 2134 249 2137
rect 11177 2215 11425 2218
rect 11177 2137 11181 2215
rect 11181 2137 11421 2215
rect 11421 2137 11425 2215
rect 11177 2134 11425 2137
rect 351 1671 599 1674
rect 351 1593 355 1671
rect 355 1593 595 1671
rect 595 1593 599 1671
rect 351 1590 599 1593
rect 11527 1671 11775 1674
rect 11527 1593 11531 1671
rect 11531 1593 11771 1671
rect 11771 1593 11775 1671
rect 11527 1590 11775 1593
rect 1 1127 249 1130
rect 1 1049 5 1127
rect 5 1049 245 1127
rect 245 1049 249 1127
rect 1 1046 249 1049
rect 11177 1127 11425 1130
rect 11177 1049 11181 1127
rect 11181 1049 11421 1127
rect 11421 1049 11425 1127
rect 11177 1046 11425 1049
rect 351 583 599 586
rect 351 505 355 583
rect 355 505 595 583
rect 595 505 599 583
rect 351 502 599 505
rect 11527 583 11775 586
rect 11527 505 11531 583
rect 11531 505 11771 583
rect 11771 505 11775 583
rect 11527 502 11775 505
rect 1 39 249 42
rect 1 -39 5 39
rect 5 -39 245 39
rect 245 -39 249 39
rect 1 -42 249 -39
rect 11177 39 11425 42
rect 11177 -39 11181 39
rect 11181 -39 11421 39
rect 11421 -39 11425 39
rect 11177 -42 11425 -39
<< metal4 >>
rect 0 8746 250 8752
rect 0 8662 1 8746
rect 249 8662 250 8746
rect 0 7658 250 8662
rect 0 7574 1 7658
rect 249 7574 250 7658
rect 0 6570 250 7574
rect 0 6486 1 6570
rect 249 6486 250 6570
rect 0 5482 250 6486
rect 0 5398 1 5482
rect 249 5398 250 5482
rect 0 4394 250 5398
rect 0 4310 1 4394
rect 249 4310 250 4394
rect 0 3306 250 4310
rect 0 3222 1 3306
rect 249 3222 250 3306
rect 0 2218 250 3222
rect 0 2134 1 2218
rect 249 2134 250 2218
rect 0 1130 250 2134
rect 0 1046 1 1130
rect 249 1046 250 1130
rect 0 42 250 1046
rect 0 -42 1 42
rect 249 -42 250 42
rect 0 -48 250 -42
rect 350 8202 600 8752
rect 350 8118 351 8202
rect 599 8118 600 8202
rect 350 7114 600 8118
rect 350 7030 351 7114
rect 599 7030 600 7114
rect 350 6026 600 7030
rect 350 5942 351 6026
rect 599 5942 600 6026
rect 350 4938 600 5942
rect 350 4854 351 4938
rect 599 4854 600 4938
rect 350 3850 600 4854
rect 350 3766 351 3850
rect 599 3766 600 3850
rect 350 2762 600 3766
rect 350 2678 351 2762
rect 599 2678 600 2762
rect 350 1674 600 2678
rect 350 1590 351 1674
rect 599 1590 600 1674
rect 350 586 600 1590
rect 350 502 351 586
rect 599 502 600 586
rect 350 -48 600 502
rect 11176 8746 11426 8752
rect 11176 8662 11177 8746
rect 11425 8662 11426 8746
rect 11176 7658 11426 8662
rect 11176 7574 11177 7658
rect 11425 7574 11426 7658
rect 11176 6570 11426 7574
rect 11176 6486 11177 6570
rect 11425 6486 11426 6570
rect 11176 5482 11426 6486
rect 11176 5398 11177 5482
rect 11425 5398 11426 5482
rect 11176 4394 11426 5398
rect 11176 4310 11177 4394
rect 11425 4310 11426 4394
rect 11176 3306 11426 4310
rect 11176 3222 11177 3306
rect 11425 3222 11426 3306
rect 11176 2218 11426 3222
rect 11176 2134 11177 2218
rect 11425 2134 11426 2218
rect 11176 1130 11426 2134
rect 11176 1046 11177 1130
rect 11425 1046 11426 1130
rect 11176 42 11426 1046
rect 11176 -42 11177 42
rect 11425 -42 11426 42
rect 11176 -48 11426 -42
rect 11526 8202 11776 8752
rect 11526 8118 11527 8202
rect 11775 8118 11776 8202
rect 11526 7114 11776 8118
rect 11526 7030 11527 7114
rect 11775 7030 11776 7114
rect 11526 6026 11776 7030
rect 11526 5942 11527 6026
rect 11775 5942 11776 6026
rect 11526 4938 11776 5942
rect 11526 4854 11527 4938
rect 11775 4854 11776 4938
rect 11526 3850 11776 4854
rect 11526 3766 11527 3850
rect 11775 3766 11776 3850
rect 11526 2762 11776 3766
rect 11526 2678 11527 2762
rect 11775 2678 11776 2762
rect 11526 1674 11776 2678
rect 11526 1590 11527 1674
rect 11775 1590 11776 1674
rect 11526 586 11776 1590
rect 11526 502 11527 586
rect 11775 502 11776 586
rect 11526 -48 11776 502
use sky130_fd_sc_hd__clkbuf_8  sky130_fd_sc_hd__clkbuf_8_0 $PDK_ROOT/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 6900 0 -1 1088
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  sky130_fd_sc_hd__clkbuf_8_1
timestamp 1707688321
transform -1 0 6900 0 1 1088
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  sky130_fd_sc_hd__clkbuf_8_2
timestamp 1707688321
transform -1 0 6900 0 -1 2176
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  sky130_fd_sc_hd__clkbuf_8_3
timestamp 1707688321
transform -1 0 6900 0 1 2176
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  sky130_fd_sc_hd__clkbuf_8_4
timestamp 1707688321
transform -1 0 6900 0 -1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  sky130_fd_sc_hd__clkbuf_8_5
timestamp 1707688321
transform -1 0 6900 0 1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  sky130_fd_sc_hd__clkbuf_8_6
timestamp 1707688321
transform -1 0 6900 0 -1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  sky130_fd_sc_hd__clkbuf_8_7
timestamp 1707688321
transform -1 0 6900 0 1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  sky130_fd_sc_hd__clkbuf_8_8
timestamp 1707688321
transform -1 0 6900 0 -1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  sky130_fd_sc_hd__clkbuf_8_9
timestamp 1707688321
transform -1 0 6900 0 1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  sky130_fd_sc_hd__clkbuf_8_10
timestamp 1707688321
transform -1 0 6900 0 -1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  sky130_fd_sc_hd__clkbuf_8_11
timestamp 1707688321
transform -1 0 6900 0 1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  sky130_fd_sc_hd__clkbuf_8_12
timestamp 1707688321
transform -1 0 6900 0 -1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  sky130_fd_sc_hd__clkbuf_8_13
timestamp 1707688321
transform -1 0 6900 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  sky130_fd_sc_hd__clkbuf_8_14
timestamp 1707688321
transform -1 0 2944 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  sky130_fd_sc_hd__clkbuf_8_15
timestamp 1707688321
transform 1 0 7636 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  sky130_fd_sc_hd__clkbuf_8_16
timestamp 1707688321
transform 1 0 9016 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  sky130_fd_sc_hd__clkbuf_8_17
timestamp 1707688321
transform -1 0 11132 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_0 $PDK_ROOT/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 0 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_1
timestamp 1707688321
transform 1 0 3312 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_2
timestamp 1707688321
transform 1 0 5520 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_3
timestamp 1707688321
transform 1 0 0 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_4
timestamp 1707688321
transform 1 0 3312 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_5
timestamp 1707688321
transform 1 0 5520 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_6
timestamp 1707688321
transform 1 0 0 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_7
timestamp 1707688321
transform 1 0 3312 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_8
timestamp 1707688321
transform 1 0 5520 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_9
timestamp 1707688321
transform 1 0 0 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_10
timestamp 1707688321
transform 1 0 5520 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_11
timestamp 1707688321
transform 1 0 0 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_12
timestamp 1707688321
transform 1 0 5520 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_13
timestamp 1707688321
transform 1 0 0 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_14
timestamp 1707688321
transform 1 0 5520 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_15
timestamp 1707688321
transform 1 0 0 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_16
timestamp 1707688321
transform 1 0 5520 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_17
timestamp 1707688321
transform 1 0 0 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_18
timestamp 1707688321
transform 1 0 5520 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_19
timestamp 1707688321
transform 1 0 0 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_20
timestamp 1707688321
transform 1 0 5520 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_21
timestamp 1707688321
transform 1 0 0 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_22
timestamp 1707688321
transform 1 0 5520 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_23
timestamp 1707688321
transform 1 0 0 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_24
timestamp 1707688321
transform 1 0 5520 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_25
timestamp 1707688321
transform 1 0 0 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_26
timestamp 1707688321
transform 1 0 5520 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_27
timestamp 1707688321
transform 1 0 0 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_28
timestamp 1707688321
transform 1 0 5520 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_29
timestamp 1707688321
transform 1 0 0 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_30
timestamp 1707688321
transform 1 0 3312 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_31
timestamp 1707688321
transform 1 0 5520 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_32
timestamp 1707688321
transform 1 0 0 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_33
timestamp 1707688321
transform 1 0 3312 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_34
timestamp 1707688321
transform 1 0 5520 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_35
timestamp 1707688321
transform 1 0 0 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_36
timestamp 1707688321
transform 1 0 5520 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_0 $PDK_ROOT/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 1472 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_1
timestamp 1707688321
transform 1 0 8648 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_0 $PDK_ROOT/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 11224 0 1 0
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_1
timestamp 1707688321
transform 1 0 11224 0 -1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_2
timestamp 1707688321
transform 1 0 11224 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_3
timestamp 1707688321
transform 1 0 11224 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_4
timestamp 1707688321
transform 1 0 11224 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_5
timestamp 1707688321
transform 1 0 11224 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_6
timestamp 1707688321
transform 1 0 11224 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_7
timestamp 1707688321
transform 1 0 11224 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_8
timestamp 1707688321
transform 1 0 11224 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_9
timestamp 1707688321
transform 1 0 11224 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_10
timestamp 1707688321
transform 1 0 11224 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_11
timestamp 1707688321
transform 1 0 11224 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_12
timestamp 1707688321
transform 1 0 11224 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_13
timestamp 1707688321
transform 1 0 11224 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_14
timestamp 1707688321
transform 1 0 11224 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_15
timestamp 1707688321
transform 1 0 2944 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_16
timestamp 1707688321
transform 1 0 6992 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_17
timestamp 1707688321
transform 1 0 11132 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_0 $PDK_ROOT/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 2576 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_1
timestamp 1707688321
transform 1 0 4784 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_2
timestamp 1707688321
transform 1 0 9200 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_3
timestamp 1707688321
transform 1 0 2576 0 -1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_4
timestamp 1707688321
transform 1 0 4784 0 -1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_5
timestamp 1707688321
transform 1 0 2576 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_6
timestamp 1707688321
transform 1 0 4784 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_7
timestamp 1707688321
transform 1 0 4784 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_8
timestamp 1707688321
transform 1 0 4784 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_9
timestamp 1707688321
transform 1 0 4784 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_10
timestamp 1707688321
transform 1 0 4784 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_11
timestamp 1707688321
transform 1 0 4784 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_12
timestamp 1707688321
transform 1 0 4784 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_13
timestamp 1707688321
transform 1 0 4784 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_14
timestamp 1707688321
transform 1 0 4784 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_15
timestamp 1707688321
transform 1 0 4784 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_16
timestamp 1707688321
transform 1 0 4784 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_17
timestamp 1707688321
transform 1 0 2576 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_18
timestamp 1707688321
transform 1 0 4784 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_19
timestamp 1707688321
transform 1 0 2576 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_20
timestamp 1707688321
transform 1 0 4784 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_21
timestamp 1707688321
transform 1 0 4784 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_0 $PDK_ROOT/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 368 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_1
timestamp 1707688321
transform 1 0 1472 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_2
timestamp 1707688321
transform 1 0 3680 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_3
timestamp 1707688321
transform 1 0 5888 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_4
timestamp 1707688321
transform 1 0 6992 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_5
timestamp 1707688321
transform 1 0 8096 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_6
timestamp 1707688321
transform 1 0 10120 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_7
timestamp 1707688321
transform 1 0 368 0 -1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_8
timestamp 1707688321
transform 1 0 1472 0 -1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_9
timestamp 1707688321
transform 1 0 3680 0 -1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_10
timestamp 1707688321
transform 1 0 10120 0 -1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_11
timestamp 1707688321
transform 1 0 368 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_12
timestamp 1707688321
transform 1 0 1472 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_13
timestamp 1707688321
transform 1 0 3680 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_14
timestamp 1707688321
transform 1 0 10120 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_15
timestamp 1707688321
transform 1 0 3680 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_16
timestamp 1707688321
transform 1 0 10120 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_17
timestamp 1707688321
transform 1 0 3680 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_18
timestamp 1707688321
transform 1 0 10120 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_19
timestamp 1707688321
transform 1 0 3680 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_20
timestamp 1707688321
transform 1 0 10120 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_21
timestamp 1707688321
transform 1 0 3680 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_22
timestamp 1707688321
transform 1 0 10120 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_23
timestamp 1707688321
transform 1 0 3680 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_24
timestamp 1707688321
transform 1 0 10120 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_25
timestamp 1707688321
transform 1 0 3680 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_26
timestamp 1707688321
transform 1 0 10120 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_27
timestamp 1707688321
transform 1 0 3680 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_28
timestamp 1707688321
transform 1 0 10120 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_29
timestamp 1707688321
transform 1 0 3680 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_30
timestamp 1707688321
transform 1 0 10120 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_31
timestamp 1707688321
transform 1 0 3680 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_32
timestamp 1707688321
transform 1 0 10120 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_33
timestamp 1707688321
transform 1 0 3680 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_34
timestamp 1707688321
transform 1 0 10120 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_35
timestamp 1707688321
transform 1 0 368 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_36
timestamp 1707688321
transform 1 0 1472 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_37
timestamp 1707688321
transform 1 0 3680 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_38
timestamp 1707688321
transform 1 0 10120 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_39
timestamp 1707688321
transform 1 0 368 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_40
timestamp 1707688321
transform 1 0 1472 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_41
timestamp 1707688321
transform 1 0 3680 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_42
timestamp 1707688321
transform 1 0 10120 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_43
timestamp 1707688321
transform 1 0 368 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_44
timestamp 1707688321
transform 1 0 3680 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_45
timestamp 1707688321
transform 1 0 5888 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_2  sky130_fd_sc_hd__dfxtp_2_0 $PDK_ROOT/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 8464 0 -1 1088
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  sky130_fd_sc_hd__dfxtp_2_1
timestamp 1707688321
transform -1 0 10028 0 -1 1088
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  sky130_fd_sc_hd__dfxtp_2_2
timestamp 1707688321
transform -1 0 8464 0 1 1088
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  sky130_fd_sc_hd__dfxtp_2_3
timestamp 1707688321
transform -1 0 10028 0 1 1088
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  sky130_fd_sc_hd__dfxtp_2_4
timestamp 1707688321
transform 1 0 2024 0 -1 2176
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  sky130_fd_sc_hd__dfxtp_2_5
timestamp 1707688321
transform -1 0 8464 0 -1 2176
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  sky130_fd_sc_hd__dfxtp_2_6
timestamp 1707688321
transform -1 0 10028 0 -1 2176
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  sky130_fd_sc_hd__dfxtp_2_7
timestamp 1707688321
transform 1 0 2024 0 1 2176
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  sky130_fd_sc_hd__dfxtp_2_8
timestamp 1707688321
transform -1 0 8464 0 1 2176
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  sky130_fd_sc_hd__dfxtp_2_9
timestamp 1707688321
transform -1 0 10028 0 1 2176
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  sky130_fd_sc_hd__dfxtp_2_10
timestamp 1707688321
transform 1 0 2024 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  sky130_fd_sc_hd__dfxtp_2_11
timestamp 1707688321
transform -1 0 8464 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  sky130_fd_sc_hd__dfxtp_2_12
timestamp 1707688321
transform -1 0 10028 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  sky130_fd_sc_hd__dfxtp_2_13
timestamp 1707688321
transform 1 0 2024 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  sky130_fd_sc_hd__dfxtp_2_14
timestamp 1707688321
transform -1 0 8464 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  sky130_fd_sc_hd__dfxtp_2_15
timestamp 1707688321
transform -1 0 10028 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  sky130_fd_sc_hd__dfxtp_2_16
timestamp 1707688321
transform 1 0 2024 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  sky130_fd_sc_hd__dfxtp_2_17
timestamp 1707688321
transform -1 0 8464 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  sky130_fd_sc_hd__dfxtp_2_18
timestamp 1707688321
transform -1 0 10028 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  sky130_fd_sc_hd__dfxtp_2_19
timestamp 1707688321
transform 1 0 2024 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  sky130_fd_sc_hd__dfxtp_2_20
timestamp 1707688321
transform -1 0 8464 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  sky130_fd_sc_hd__dfxtp_2_21
timestamp 1707688321
transform -1 0 10028 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  sky130_fd_sc_hd__dfxtp_2_22
timestamp 1707688321
transform 1 0 2024 0 -1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  sky130_fd_sc_hd__dfxtp_2_23
timestamp 1707688321
transform -1 0 8464 0 -1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  sky130_fd_sc_hd__dfxtp_2_24
timestamp 1707688321
transform -1 0 10028 0 -1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  sky130_fd_sc_hd__dfxtp_2_25
timestamp 1707688321
transform 1 0 2024 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  sky130_fd_sc_hd__dfxtp_2_26
timestamp 1707688321
transform -1 0 8464 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  sky130_fd_sc_hd__dfxtp_2_27
timestamp 1707688321
transform -1 0 10028 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  sky130_fd_sc_hd__dfxtp_2_28
timestamp 1707688321
transform 1 0 2024 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  sky130_fd_sc_hd__dfxtp_2_29
timestamp 1707688321
transform -1 0 8464 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  sky130_fd_sc_hd__dfxtp_2_30
timestamp 1707688321
transform -1 0 10028 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  sky130_fd_sc_hd__dfxtp_2_31
timestamp 1707688321
transform 1 0 2024 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  sky130_fd_sc_hd__dfxtp_2_32
timestamp 1707688321
transform -1 0 8464 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  sky130_fd_sc_hd__dfxtp_2_33
timestamp 1707688321
transform -1 0 10028 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  sky130_fd_sc_hd__dfxtp_2_34
timestamp 1707688321
transform -1 0 8464 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  sky130_fd_sc_hd__dfxtp_2_35
timestamp 1707688321
transform -1 0 10028 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  sky130_fd_sc_hd__dfxtp_2_36
timestamp 1707688321
transform -1 0 8464 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  sky130_fd_sc_hd__dfxtp_2_37
timestamp 1707688321
transform -1 0 10028 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_0 $PDK_ROOT/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 9936 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_1
timestamp 1707688321
transform 1 0 1840 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_2
timestamp 1707688321
transform 1 0 3496 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_3
timestamp 1707688321
transform 1 0 7544 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_4
timestamp 1707688321
transform 1 0 11684 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__mux4_2  sky130_fd_sc_hd__mux4_2_0 $PDK_ROOT/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 368 0 -1 2176
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  sky130_fd_sc_hd__mux4_2_1
timestamp 1707688321
transform 1 0 368 0 1 2176
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  sky130_fd_sc_hd__mux4_2_2
timestamp 1707688321
transform 1 0 368 0 -1 3264
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  sky130_fd_sc_hd__mux4_2_3
timestamp 1707688321
transform 1 0 368 0 1 3264
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  sky130_fd_sc_hd__mux4_2_4
timestamp 1707688321
transform 1 0 368 0 -1 4352
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  sky130_fd_sc_hd__mux4_2_5
timestamp 1707688321
transform 1 0 368 0 1 4352
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  sky130_fd_sc_hd__mux4_2_6
timestamp 1707688321
transform 1 0 368 0 -1 5440
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  sky130_fd_sc_hd__mux4_2_7
timestamp 1707688321
transform 1 0 368 0 1 5440
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  sky130_fd_sc_hd__mux4_2_8
timestamp 1707688321
transform 1 0 368 0 -1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  sky130_fd_sc_hd__mux4_2_9
timestamp 1707688321
transform 1 0 368 0 1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDK_ROOT/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 276 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1707688321
transform 1 0 3588 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1707688321
transform 1 0 5796 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1707688321
transform 1 0 10028 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1707688321
transform 1 0 276 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1707688321
transform 1 0 3588 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_6
timestamp 1707688321
transform 1 0 5796 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_7
timestamp 1707688321
transform 1 0 10028 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_8
timestamp 1707688321
transform 1 0 276 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_9
timestamp 1707688321
transform 1 0 3588 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_10
timestamp 1707688321
transform 1 0 5796 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_11
timestamp 1707688321
transform 1 0 10028 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_12
timestamp 1707688321
transform 1 0 276 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_13
timestamp 1707688321
transform 1 0 3588 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_14
timestamp 1707688321
transform 1 0 5796 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_15
timestamp 1707688321
transform 1 0 10028 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_16
timestamp 1707688321
transform 1 0 276 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_17
timestamp 1707688321
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_18
timestamp 1707688321
transform 1 0 5796 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_19
timestamp 1707688321
transform 1 0 10028 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_20
timestamp 1707688321
transform 1 0 276 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_21
timestamp 1707688321
transform 1 0 3588 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_22
timestamp 1707688321
transform 1 0 5796 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_23
timestamp 1707688321
transform 1 0 10028 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_24
timestamp 1707688321
transform 1 0 276 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_25
timestamp 1707688321
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_26
timestamp 1707688321
transform 1 0 5796 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_27
timestamp 1707688321
transform 1 0 10028 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_28
timestamp 1707688321
transform 1 0 276 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_29
timestamp 1707688321
transform 1 0 3588 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_30
timestamp 1707688321
transform 1 0 5796 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_31
timestamp 1707688321
transform 1 0 10028 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_32
timestamp 1707688321
transform 1 0 276 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_33
timestamp 1707688321
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_34
timestamp 1707688321
transform 1 0 5796 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_35
timestamp 1707688321
transform 1 0 10028 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_36
timestamp 1707688321
transform 1 0 276 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_37
timestamp 1707688321
transform 1 0 3588 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_38
timestamp 1707688321
transform 1 0 5796 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_39
timestamp 1707688321
transform 1 0 10028 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_40
timestamp 1707688321
transform 1 0 276 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_41
timestamp 1707688321
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_42
timestamp 1707688321
transform 1 0 5796 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_43
timestamp 1707688321
transform 1 0 10028 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_44
timestamp 1707688321
transform 1 0 276 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_45
timestamp 1707688321
transform 1 0 3588 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_46
timestamp 1707688321
transform 1 0 5796 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_47
timestamp 1707688321
transform 1 0 10028 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_48
timestamp 1707688321
transform 1 0 276 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_49
timestamp 1707688321
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_50
timestamp 1707688321
transform 1 0 5796 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_51
timestamp 1707688321
transform 1 0 10028 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_52
timestamp 1707688321
transform 1 0 276 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_53
timestamp 1707688321
transform 1 0 3588 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_54
timestamp 1707688321
transform 1 0 5796 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_55
timestamp 1707688321
transform 1 0 10028 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_56
timestamp 1707688321
transform 1 0 276 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_57
timestamp 1707688321
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_58
timestamp 1707688321
transform 1 0 5796 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_59
timestamp 1707688321
transform 1 0 10028 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_60
timestamp 1707688321
transform 1 0 276 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_61
timestamp 1707688321
transform 1 0 3588 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_62
timestamp 1707688321
transform 1 0 5796 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_63
timestamp 1707688321
transform 1 0 10028 0 -1 8704
box -38 -48 130 592
<< labels >>
flabel metal4 0 -48 250 8752 1 FreeSans 160 0 0 0 VGND
port 0 n ground input
flabel metal4 350 -48 600 8752 1 FreeSans 160 0 0 0 VDPWR
port 1 n power input
flabel metal4 11176 -48 11426 8752 1 FreeSans 160 0 0 0 VGND
port 0 n ground input
flabel metal4 11526 -48 11776 8752 1 FreeSans 160 0 0 0 VDPWR
port 1 n power input
flabel metal2 2884 8792 2912 8820 1 FreeSans 40 0 0 0 usr_data_clk
port 12 n signal input
flabel metal2 7668 8792 7696 8820 1 FreeSans 40 0 0 0 usr_addr_clk
port 11 n signal input
flabel metal2 9048 8792 9076 8820 1 FreeSans 40 0 0 0 usr_addr_hi_clk
port 9 n signal input
flabel metal2 11072 8792 11100 8820 1 FreeSans 40 0 0 0 usr_addr_lo_clk
port 10 n signal input
flabel metal2 -1900 -116 -1872 -88 1 FreeSans 40 0 0 0 rom_data0_in[0]
port 48 n signal input
flabel metal2 -1992 -116 -1964 -88 1 FreeSans 40 0 0 0 rom_data0_in[1]
port 47 n signal input
flabel metal2 -2084 -116 -2056 -88 1 FreeSans 40 0 0 0 rom_data0_in[2]
port 46 n signal input
flabel metal2 -2176 -116 -2148 -88 1 FreeSans 40 0 0 0 rom_data0_in[3]
port 45 n signal input
flabel metal2 -2268 -116 -2240 -88 1 FreeSans 40 0 0 0 rom_data0_in[4]
port 44 n signal input
flabel metal2 -2360 -116 -2332 -88 1 FreeSans 40 0 0 0 rom_data0_in[5]
port 43 n signal input
flabel metal2 -2452 -116 -2424 -88 1 FreeSans 40 0 0 0 rom_data0_in[6]
port 42 n signal input
flabel metal2 -2544 -116 -2516 -88 1 FreeSans 40 0 0 0 rom_data0_in[7]
port 41 n signal input
flabel metal2 -2636 -116 -2608 -88 1 FreeSans 40 0 0 0 rom_data0_in[8]
port 40 n signal input
flabel metal2 -2728 -116 -2700 -88 1 FreeSans 40 0 0 0 rom_data0_in[9]
port 39 n signal input
flabel metal2 -980 -116 -952 -88 1 FreeSans 40 0 0 0 rom_data1_in[0]
port 58 n signal input
flabel metal2 -1072 -116 -1044 -88 1 FreeSans 40 0 0 0 rom_data1_in[1]
port 57 n signal input
flabel metal2 -1164 -116 -1136 -88 1 FreeSans 40 0 0 0 rom_data1_in[2]
port 56 n signal input
flabel metal2 -1256 -116 -1228 -88 1 FreeSans 40 0 0 0 rom_data1_in[3]
port 55 n signal input
flabel metal2 -1348 -116 -1320 -88 1 FreeSans 40 0 0 0 rom_data1_in[4]
port 54 n signal input
flabel metal2 -1440 -116 -1412 -88 1 FreeSans 40 0 0 0 rom_data1_in[5]
port 53 n signal input
flabel metal2 -1532 -116 -1504 -88 1 FreeSans 40 0 0 0 rom_data1_in[6]
port 52 n signal input
flabel metal2 -1624 -116 -1596 -88 1 FreeSans 40 0 0 0 rom_data1_in[7]
port 51 n signal input
flabel metal2 -1716 -116 -1688 -88 1 FreeSans 40 0 0 0 rom_data1_in[8]
port 50 n signal input
flabel metal2 -1808 -116 -1780 -88 1 FreeSans 40 0 0 0 rom_data1_in[9]
port 49 n signal input
flabel metal2 -60 -116 -32 -88 1 FreeSans 40 0 0 0 rom_data2_in[0]
port 68 n signal input
flabel metal2 -152 -116 -124 -88 1 FreeSans 40 0 0 0 rom_data2_in[1]
port 67 n signal input
flabel metal2 -244 -116 -216 -88 1 FreeSans 40 0 0 0 rom_data2_in[2]
port 66 n signal input
flabel metal2 -336 -116 -308 -88 1 FreeSans 40 0 0 0 rom_data2_in[3]
port 65 n signal input
flabel metal2 -428 -116 -400 -88 1 FreeSans 40 0 0 0 rom_data2_in[4]
port 64 n signal input
flabel metal2 -520 -116 -492 -88 1 FreeSans 40 0 0 0 rom_data2_in[5]
port 63 n signal input
flabel metal2 -612 -116 -584 -88 1 FreeSans 40 0 0 0 rom_data2_in[6]
port 62 n signal input
flabel metal2 -704 -116 -676 -88 1 FreeSans 40 0 0 0 rom_data2_in[7]
port 61 n signal input
flabel metal2 -796 -116 -768 -88 1 FreeSans 40 0 0 0 rom_data2_in[8]
port 60 n signal input
flabel metal2 -888 -116 -860 -88 1 FreeSans 40 0 0 0 rom_data2_in[9]
port 59 n signal input
flabel metal2 1596 8792 1624 8820 1 FreeSans 40 0 0 0 usr_data_sel[0]
port 24 n signal input
flabel metal2 952 8792 980 8820 1 FreeSans 40 0 0 0 usr_data_sel[1]
port 23 n signal input
flabel metal2 4356 8792 4384 8820 1 FreeSans 40 0 0 0 usr_data_out[0]
port 22 n signal output
flabel metal2 4264 8792 4292 8820 1 FreeSans 40 0 0 0 usr_data_out[1]
port 21 n signal output
flabel metal2 4172 8792 4200 8820 1 FreeSans 40 0 0 0 usr_data_out[2]
port 20 n signal output
flabel metal2 4080 8792 4108 8820 1 FreeSans 40 0 0 0 usr_data_out[3]
port 19 n signal output
flabel metal2 3988 8792 4016 8820 1 FreeSans 40 0 0 0 usr_data_out[4]
port 18 n signal output
flabel metal2 3896 8792 3924 8820 1 FreeSans 40 0 0 0 usr_data_out[5]
port 17 n signal output
flabel metal2 3804 8792 3832 8820 1 FreeSans 40 0 0 0 usr_data_out[6]
port 16 n signal output
flabel metal2 3712 8792 3740 8820 1 FreeSans 40 0 0 0 usr_data_out[7]
port 15 n signal output
flabel metal2 3620 8792 3648 8820 1 FreeSans 40 0 0 0 usr_data_out[8]
port 14 n signal output
flabel metal2 3528 8792 3556 8820 1 FreeSans 40 0 0 0 usr_data_out[9]
port 13 n signal output
flabel metal2 10980 8792 11008 8820 1 FreeSans 40 0 0 0 usr_addr_in[0]
port 8 n signal input
flabel metal2 10888 8792 10916 8820 1 FreeSans 40 0 0 0 usr_addr_in[1]
port 7 n signal input
flabel metal2 10796 8792 10824 8820 1 FreeSans 40 0 0 0 usr_addr_in[2]
port 6 n signal input
flabel metal2 10704 8792 10732 8820 1 FreeSans 40 0 0 0 usr_addr_in[3]
port 5 n signal input
flabel metal2 10612 8792 10640 8820 1 FreeSans 40 0 0 0 usr_addr_in[4]
port 4 n signal input
flabel metal2 10520 8792 10548 8820 1 FreeSans 40 0 0 0 usr_addr_in[5]
port 3 n signal input
flabel metal2 10428 8792 10456 8820 1 FreeSans 40 0 0 0 usr_addr_in[6]
port 2 n signal input
flabel metal2 5920 -116 5948 -88 1 FreeSans 40 0 0 0 rom_addr_out[0]
port 38 n signal output
flabel metal2 5828 -116 5856 -88 1 FreeSans 40 0 0 0 rom_addr_out[1]
port 37 n signal output
flabel metal2 5736 -116 5764 -88 1 FreeSans 40 0 0 0 rom_addr_out[2]
port 36 n signal output
flabel metal2 5644 -116 5672 -88 1 FreeSans 40 0 0 0 rom_addr_out[3]
port 35 n signal output
flabel metal2 5552 -116 5580 -88 1 FreeSans 40 0 0 0 rom_addr_out[4]
port 34 n signal output
flabel metal2 5460 -116 5488 -88 1 FreeSans 40 0 0 0 rom_addr_out[5]
port 33 n signal output
flabel metal2 5368 -116 5396 -88 1 FreeSans 40 0 0 0 rom_addr_out[6]
port 32 n signal output
flabel metal2 5276 -116 5304 -88 1 FreeSans 40 0 0 0 rom_addr_out[7]
port 31 n signal output
flabel metal2 5184 -116 5212 -88 1 FreeSans 40 0 0 0 rom_addr_out[8]
port 30 n signal output
flabel metal2 5092 -116 5120 -88 1 FreeSans 40 0 0 0 rom_addr_out[9]
port 29 n signal output
flabel metal2 5000 -116 5028 -88 1 FreeSans 40 0 0 0 rom_addr_out[10]
port 28 n signal output
flabel metal2 4908 -116 4936 -88 1 FreeSans 40 0 0 0 rom_addr_out[11]
port 27 n signal output
flabel metal2 4816 -116 4844 -88 1 FreeSans 40 0 0 0 rom_addr_out[12]
port 26 n signal output
flabel metal2 4724 -116 4752 -88 1 FreeSans 40 0 0 0 rom_addr_out[13]
port 25 n signal output
<< end >>
