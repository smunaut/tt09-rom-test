magic
tech sky130A
magscale 1 2
timestamp 1730764879
<< metal1 >>
rect 3324 28506 3376 28512
rect 3324 24881 3376 28454
rect 4234 27726 4286 27732
rect 4234 27301 4286 27674
rect 4234 27243 4286 27249
rect 3324 24823 3376 24829
<< via1 >>
rect 3324 28454 3376 28506
rect 4234 27674 4286 27726
rect 4234 27249 4286 27301
rect 3324 24829 3376 24881
<< metal2 >>
rect 3866 44788 3922 44797
rect 3866 44723 3922 44732
rect 3880 41936 3908 44723
rect 4510 44658 4566 44667
rect 4510 44593 4566 44602
rect 4524 41936 4552 44593
rect 7270 44528 7326 44537
rect 7270 44463 7326 44472
rect 7178 44398 7234 44407
rect 7178 44333 7234 44342
rect 7086 44268 7142 44277
rect 7086 44203 7142 44212
rect 6994 44138 7050 44147
rect 6994 44073 7050 44082
rect 6902 44008 6958 44017
rect 6902 43943 6958 43952
rect 6810 43878 6866 43887
rect 6810 43813 6866 43822
rect 6718 43748 6774 43757
rect 6718 43683 6774 43692
rect 6626 43618 6682 43627
rect 6626 43553 6682 43562
rect 6534 43488 6590 43497
rect 6534 43423 6590 43432
rect 6442 43358 6498 43367
rect 6442 43293 6498 43302
rect 5798 42448 5854 42457
rect 5798 42383 5854 42392
rect 5812 41936 5840 42383
rect 6456 41936 6484 43293
rect 6548 41936 6576 43423
rect 6640 41936 6668 43553
rect 6732 41936 6760 43683
rect 6824 41936 6852 43813
rect 6916 41936 6944 43943
rect 7008 41936 7036 44073
rect 7100 41936 7128 44203
rect 7192 41936 7220 44333
rect 7284 41936 7312 44463
rect 13895 43488 13951 43497
rect 13895 43423 13951 43432
rect 13908 43407 13937 43423
rect 13802 43358 13858 43367
rect 13802 43293 13858 43302
rect 13710 43228 13766 43237
rect 13710 43163 13766 43172
rect 13618 43098 13674 43107
rect 13618 43033 13674 43042
rect 13526 42968 13582 42977
rect 13526 42903 13582 42912
rect 13434 42838 13490 42847
rect 13434 42773 13490 42782
rect 13342 42708 13398 42717
rect 13342 42643 13398 42652
rect 10582 42318 10638 42327
rect 10582 42253 10638 42262
rect 10596 41936 10624 42253
rect 11962 42188 12018 42197
rect 11962 42123 12018 42132
rect 11976 41936 12004 42123
rect 13356 41936 13384 42643
rect 13448 41936 13476 42773
rect 13540 41936 13568 42903
rect 13632 41936 13660 43033
rect 13724 41936 13752 43163
rect 13816 41936 13844 43293
rect 13908 41936 13936 43407
rect 13986 42058 14042 42067
rect 13986 41993 14042 42002
rect 14000 41936 14028 41993
rect 19373 34747 19382 34803
rect 19438 34801 19447 34803
rect 19438 34749 22200 34801
rect 19438 34747 19447 34749
rect 19503 34547 19512 34603
rect 19568 34601 19577 34603
rect 19568 34549 22200 34601
rect 19568 34547 19577 34549
rect 19763 34347 19772 34403
rect 19828 34401 19837 34403
rect 19828 34349 22200 34401
rect 19828 34347 19837 34349
rect 19893 34147 19902 34203
rect 19958 34201 19967 34203
rect 19958 34149 22200 34201
rect 19958 34147 19967 34149
rect 20283 33947 20292 34003
rect 20348 34001 20357 34003
rect 20348 33949 22200 34001
rect 20348 33947 20357 33949
rect 20933 33747 20942 33803
rect 20998 33801 21007 33803
rect 20998 33749 22200 33801
rect 20998 33747 21007 33749
rect 20803 33547 20812 33603
rect 20868 33601 20877 33603
rect 20868 33549 22200 33601
rect 20868 33547 20877 33549
rect 20673 33347 20682 33403
rect 20738 33401 20747 33403
rect 20738 33349 22200 33401
rect 20738 33347 20747 33349
rect 20413 33147 20422 33203
rect 20478 33201 20487 33203
rect 20478 33149 22200 33201
rect 20478 33147 20487 33149
rect 200 436 228 33000
rect 292 2856 320 33000
rect 384 4084 412 33000
rect 476 5416 504 33000
rect 568 7836 596 33000
rect 660 10396 688 33000
rect 752 12816 780 33000
rect 844 14096 872 33000
rect 936 15376 964 33000
rect 1028 17796 1056 33000
rect 1120 22628 1148 33000
rect 1212 22720 1240 33000
rect 1304 22812 1332 33000
rect 1396 22904 1424 33000
rect 1488 22996 1516 33000
rect 1580 23088 1608 33000
rect 1672 23180 1700 33000
rect 1764 23272 1792 33000
rect 1856 23364 1884 33000
rect 1948 23456 1976 33000
rect 2040 23996 2068 33000
rect 2132 24556 2160 33000
rect 2224 24881 2252 33000
rect 2316 25206 2344 33000
rect 2408 25766 2436 33000
rect 2500 26416 2528 33000
rect 2592 26976 2620 33000
rect 2684 27301 2712 33000
rect 2776 27626 2804 33000
rect 2868 28186 2896 33000
rect 7652 32797 7680 33000
rect 7638 32788 7694 32797
rect 7638 32723 7694 32732
rect 7744 32667 7772 33000
rect 7730 32658 7786 32667
rect 7730 32593 7786 32602
rect 7836 32537 7864 33000
rect 7822 32528 7878 32537
rect 7822 32463 7878 32472
rect 7928 32431 7956 33000
rect 7927 32407 7956 32431
rect 7913 32398 7969 32407
rect 7913 32333 7969 32342
rect 8020 32277 8048 33000
rect 8006 32268 8062 32277
rect 8006 32203 8062 32212
rect 8112 32147 8140 33000
rect 8098 32138 8154 32147
rect 8098 32073 8154 32082
rect 8204 32017 8232 33000
rect 8190 32008 8246 32017
rect 8190 31943 8246 31952
rect 8296 31887 8324 33000
rect 8282 31878 8338 31887
rect 8282 31813 8338 31822
rect 8388 31781 8416 33000
rect 8388 31757 8417 31781
rect 8375 31748 8431 31757
rect 8375 31683 8431 31692
rect 8480 31627 8508 33000
rect 8466 31618 8522 31627
rect 8466 31553 8522 31562
rect 8572 31497 8600 33000
rect 8558 31488 8614 31497
rect 8558 31423 8614 31432
rect 8664 31367 8692 33000
rect 8650 31358 8706 31367
rect 8650 31293 8706 31302
rect 8756 31237 8784 33000
rect 8742 31228 8798 31237
rect 8742 31163 8798 31172
rect 8848 31107 8876 33000
rect 21144 31954 22200 32006
rect 8834 31098 8890 31107
rect 8834 31033 8890 31042
rect 3053 30567 3062 30623
rect 3118 30621 3127 30623
rect 3118 30569 4800 30621
rect 3118 30567 3127 30569
rect 3183 30367 3192 30423
rect 3248 30421 3257 30423
rect 3248 30369 4800 30421
rect 3248 30367 3257 30369
rect 3443 30167 3452 30223
rect 3508 30221 3517 30223
rect 3508 30169 4800 30221
rect 3508 30167 3517 30169
rect 3573 29967 3582 30023
rect 3638 30021 3647 30023
rect 3638 29969 4800 30021
rect 3638 29967 3647 29969
rect 3963 29767 3972 29823
rect 4028 29821 4037 29823
rect 4028 29769 4800 29821
rect 4028 29767 4037 29769
rect 4093 29567 4102 29623
rect 4158 29621 4167 29623
rect 4158 29569 4800 29621
rect 4158 29567 4167 29569
rect 4613 29367 4622 29423
rect 4678 29421 4687 29423
rect 4678 29369 4800 29421
rect 4678 29367 4687 29369
rect 4483 29167 4492 29223
rect 4548 29221 4557 29223
rect 4548 29169 4800 29221
rect 4548 29167 4557 29169
rect 4353 28967 4362 29023
rect 4418 29021 4427 29023
rect 4418 28969 4800 29021
rect 4418 28967 4427 28969
rect 3313 28452 3322 28508
rect 3378 28452 3387 28508
rect 2868 28134 4800 28186
rect 4223 27672 4232 27728
rect 4288 27672 4297 27728
rect 2776 27574 4800 27626
rect 2684 27249 4234 27301
rect 4286 27249 4292 27301
rect 2592 26924 4800 26976
rect 2500 26364 4800 26416
rect 2408 25714 4800 25766
rect 2316 25154 4800 25206
rect 2224 24829 3324 24881
rect 3376 24829 3382 24881
rect 2132 24504 4800 24556
rect 2040 23944 4800 23996
rect 21144 23456 21172 31954
rect 1948 23428 21172 23456
rect 21236 30744 22200 30796
rect 21236 23364 21264 30744
rect 21314 29729 21370 29738
rect 21314 29664 21370 29673
rect 1856 23336 21264 23364
rect 21328 23272 21356 29664
rect 1764 23244 21356 23272
rect 21420 29534 22200 29586
rect 21420 23180 21448 29534
rect 1672 23152 21448 23180
rect 21512 28324 22200 28376
rect 21512 23088 21540 28324
rect 1580 23060 21540 23088
rect 21604 26974 22200 27026
rect 21604 22996 21632 26974
rect 1488 22968 21632 22996
rect 21696 25764 22200 25816
rect 21696 22904 21724 25764
rect 21774 24739 21830 24748
rect 21774 24674 21830 24683
rect 1396 22876 21724 22904
rect 21788 22812 21816 24674
rect 1304 22784 21816 22812
rect 21880 24554 22200 24606
rect 21880 22720 21908 24554
rect 1212 22692 21908 22720
rect 21972 23344 22200 23396
rect 21972 22628 22000 23344
rect 1120 22600 22000 22628
rect 1123 22147 1132 22203
rect 1188 22201 1197 22203
rect 1188 22149 3000 22201
rect 1188 22147 1197 22149
rect 1253 21947 1262 22003
rect 1318 22001 1327 22003
rect 1318 21949 3000 22001
rect 1318 21947 1327 21949
rect 1383 21747 1392 21803
rect 1448 21801 1457 21803
rect 1448 21749 3000 21801
rect 1448 21747 1457 21749
rect 1643 21547 1652 21603
rect 1708 21601 1717 21603
rect 1708 21549 3000 21601
rect 1708 21547 1717 21549
rect 1773 21347 1782 21403
rect 1838 21401 1847 21403
rect 1838 21349 3000 21401
rect 1838 21347 1847 21349
rect 1903 21147 1912 21203
rect 1968 21201 1977 21203
rect 1968 21149 3000 21201
rect 1968 21147 1977 21149
rect 2033 20947 2042 21003
rect 2098 21001 2107 21003
rect 2098 20949 3000 21001
rect 2098 20947 2107 20949
rect 2813 20747 2822 20803
rect 2878 20801 2887 20803
rect 2878 20749 3000 20801
rect 2878 20747 2887 20749
rect 2683 20547 2692 20603
rect 2748 20601 2757 20603
rect 2748 20549 3000 20601
rect 2748 20547 2757 20549
rect 2553 20347 2562 20403
rect 2618 20401 2627 20403
rect 2618 20349 3000 20401
rect 2618 20347 2627 20349
rect 2293 20147 2302 20203
rect 2358 20201 2367 20203
rect 2358 20149 3000 20201
rect 2358 20147 2367 20149
rect 2163 19947 2172 20003
rect 2228 20001 2237 20003
rect 2228 19949 3000 20001
rect 2228 19947 2237 19949
rect 1028 17744 3000 17796
rect 936 15324 3000 15376
rect 2423 14097 2432 14099
rect 2417 14096 2432 14097
rect 844 14044 2432 14096
rect 2423 14043 2432 14044
rect 2488 14043 2497 14099
rect 752 12764 3000 12816
rect 660 10344 3000 10396
rect 568 7784 3000 7836
rect 476 5364 3000 5416
rect 1513 4085 1522 4087
rect 1507 4084 1522 4085
rect 384 4032 1522 4084
rect 1513 4031 1522 4032
rect 1578 4031 1587 4087
rect 292 2804 3000 2856
rect 200 384 3000 436
<< via2 >>
rect 3866 44732 3922 44788
rect 4510 44602 4566 44658
rect 7270 44472 7326 44528
rect 7178 44342 7234 44398
rect 7086 44212 7142 44268
rect 6994 44082 7050 44138
rect 6902 43952 6958 44008
rect 6810 43822 6866 43878
rect 6718 43692 6774 43748
rect 6626 43562 6682 43618
rect 6534 43432 6590 43488
rect 6442 43302 6498 43358
rect 5798 42392 5854 42448
rect 13895 43432 13951 43488
rect 13802 43302 13858 43358
rect 13710 43172 13766 43228
rect 13618 43042 13674 43098
rect 13526 42912 13582 42968
rect 13434 42782 13490 42838
rect 13342 42652 13398 42708
rect 10582 42262 10638 42318
rect 11962 42132 12018 42188
rect 13986 42002 14042 42058
rect 19382 34747 19438 34803
rect 19512 34547 19568 34603
rect 19772 34347 19828 34403
rect 19902 34147 19958 34203
rect 20292 33947 20348 34003
rect 20942 33747 20998 33803
rect 20812 33547 20868 33603
rect 20682 33347 20738 33403
rect 20422 33147 20478 33203
rect 7638 32732 7694 32788
rect 7730 32602 7786 32658
rect 7822 32472 7878 32528
rect 7913 32342 7969 32398
rect 8006 32212 8062 32268
rect 8098 32082 8154 32138
rect 8190 31952 8246 32008
rect 8282 31822 8338 31878
rect 8375 31692 8431 31748
rect 8466 31562 8522 31618
rect 8558 31432 8614 31488
rect 8650 31302 8706 31358
rect 8742 31172 8798 31228
rect 8834 31042 8890 31098
rect 3062 30567 3118 30623
rect 3192 30367 3248 30423
rect 3452 30167 3508 30223
rect 3582 29967 3638 30023
rect 3972 29767 4028 29823
rect 4102 29567 4158 29623
rect 4622 29367 4678 29423
rect 4492 29167 4548 29223
rect 4362 28967 4418 29023
rect 3322 28506 3378 28508
rect 3322 28454 3324 28506
rect 3324 28454 3376 28506
rect 3376 28454 3378 28506
rect 3322 28452 3378 28454
rect 4232 27726 4288 27728
rect 4232 27674 4234 27726
rect 4234 27674 4286 27726
rect 4286 27674 4288 27726
rect 4232 27672 4288 27674
rect 21314 29673 21370 29729
rect 21774 24683 21830 24739
rect 1132 22147 1188 22203
rect 1262 21947 1318 22003
rect 1392 21747 1448 21803
rect 1652 21547 1708 21603
rect 1782 21347 1838 21403
rect 1912 21147 1968 21203
rect 2042 20947 2098 21003
rect 2822 20747 2878 20803
rect 2692 20547 2748 20603
rect 2562 20347 2618 20403
rect 2302 20147 2358 20203
rect 2172 19947 2228 20003
rect 2432 14043 2488 14099
rect 1522 4031 1578 4087
<< metal3 >>
rect 7230 44950 7236 45014
rect 7300 45012 7306 45014
rect 11094 45012 11100 45014
rect 7300 44952 11100 45012
rect 7300 44950 7306 44952
rect 11094 44950 11100 44952
rect 11164 45012 11170 45014
rect 14958 45012 14964 45014
rect 11164 44952 14964 45012
rect 11164 44950 11170 44952
rect 14958 44950 14964 44952
rect 15028 44950 15034 45014
rect 3861 44790 3927 44793
rect 28758 44790 28764 44792
rect 3861 44788 28764 44790
rect 3861 44732 3866 44788
rect 3922 44732 28764 44788
rect 3861 44730 28764 44732
rect 3861 44727 3927 44730
rect 28758 44728 28764 44730
rect 28828 44728 28834 44792
rect 4505 44660 4571 44663
rect 28206 44660 28212 44662
rect 4505 44658 28212 44660
rect 4505 44602 4510 44658
rect 4566 44602 28212 44658
rect 4505 44600 28212 44602
rect 4505 44597 4571 44600
rect 28206 44598 28212 44600
rect 28276 44598 28282 44662
rect 7265 44530 7331 44533
rect 18822 44530 18828 44532
rect 7265 44528 18828 44530
rect 7265 44472 7270 44528
rect 7326 44472 18828 44528
rect 7265 44470 18828 44472
rect 7265 44467 7331 44470
rect 18822 44468 18828 44470
rect 18892 44468 18898 44532
rect 27654 44530 27660 44532
rect 19120 44470 27660 44530
rect 7173 44400 7239 44403
rect 18270 44400 18276 44402
rect 7173 44398 18276 44400
rect 7173 44342 7178 44398
rect 7234 44342 18276 44398
rect 7173 44340 18276 44342
rect 7173 44337 7239 44340
rect 18270 44338 18276 44340
rect 18340 44338 18346 44402
rect 7081 44270 7147 44273
rect 17718 44270 17724 44272
rect 7081 44268 17724 44270
rect 7081 44212 7086 44268
rect 7142 44212 17724 44268
rect 7081 44210 17724 44212
rect 7081 44207 7147 44210
rect 17718 44208 17724 44210
rect 17788 44208 17794 44272
rect 6989 44140 7055 44143
rect 17166 44140 17172 44142
rect 6989 44138 17172 44140
rect 6989 44082 6994 44138
rect 7050 44082 17172 44138
rect 6989 44080 17172 44082
rect 6989 44077 7055 44080
rect 17166 44078 17172 44080
rect 17236 44078 17242 44142
rect 6897 44010 6963 44013
rect 16614 44010 16620 44012
rect 6897 44008 16620 44010
rect 6897 43952 6902 44008
rect 6958 43952 16620 44008
rect 6897 43950 16620 43952
rect 6897 43947 6963 43950
rect 16614 43948 16620 43950
rect 16684 44010 16690 44012
rect 16684 43950 16705 44010
rect 16684 43948 16690 43950
rect 6805 43880 6871 43883
rect 14406 43880 14412 43882
rect 6805 43878 14412 43880
rect 6805 43822 6810 43878
rect 6866 43822 14412 43878
rect 6805 43820 14412 43822
rect 6805 43817 6871 43820
rect 14406 43818 14412 43820
rect 14476 43818 14482 43882
rect 6713 43750 6779 43753
rect 13854 43750 13860 43752
rect 6713 43748 13860 43750
rect 6713 43692 6718 43748
rect 6774 43692 13860 43748
rect 6713 43690 13860 43692
rect 6713 43687 6779 43690
rect 13854 43688 13860 43690
rect 13924 43688 13930 43752
rect 6621 43620 6687 43623
rect 13302 43620 13308 43622
rect 6621 43618 13308 43620
rect 6621 43562 6626 43618
rect 6682 43562 13308 43618
rect 6621 43560 13308 43562
rect 6621 43557 6687 43560
rect 13302 43558 13308 43560
rect 13372 43558 13378 43622
rect 6529 43490 6595 43493
rect 12750 43490 12756 43492
rect 6529 43488 12756 43490
rect 6529 43432 6534 43488
rect 6590 43432 12756 43488
rect 6529 43430 12756 43432
rect 6529 43427 6595 43430
rect 12750 43428 12756 43430
rect 12820 43428 12826 43492
rect 13890 43490 13956 43493
rect 19120 43490 19180 44470
rect 27654 44468 27660 44470
rect 27724 44468 27730 44532
rect 27102 44400 27108 44402
rect 13890 43488 19180 43490
rect 13890 43432 13895 43488
rect 13951 43432 19180 43488
rect 13890 43430 19180 43432
rect 19250 44340 27108 44400
rect 13890 43427 13956 43430
rect 6437 43360 6503 43363
rect 12198 43360 12204 43362
rect 6437 43358 12204 43360
rect 6437 43302 6442 43358
rect 6498 43302 12204 43358
rect 6437 43300 12204 43302
rect 6437 43297 6503 43300
rect 12198 43298 12204 43300
rect 12268 43298 12274 43362
rect 13797 43360 13863 43363
rect 19250 43360 19310 44340
rect 27102 44338 27108 44340
rect 27172 44338 27178 44402
rect 26550 44270 26556 44272
rect 13797 43358 19310 43360
rect 13797 43302 13802 43358
rect 13858 43302 19310 43358
rect 13797 43300 19310 43302
rect 19380 44210 26556 44270
rect 13797 43297 13863 43300
rect 13705 43230 13771 43233
rect 19380 43230 19440 44210
rect 26550 44208 26556 44210
rect 26620 44208 26626 44272
rect 25998 44140 26004 44142
rect 13705 43228 19440 43230
rect 13705 43172 13710 43228
rect 13766 43172 19440 43228
rect 13705 43170 19440 43172
rect 19510 44080 26004 44140
rect 13705 43167 13771 43170
rect 13613 43100 13679 43103
rect 19510 43100 19570 44080
rect 25998 44078 26004 44080
rect 26068 44078 26074 44142
rect 25446 44010 25452 44012
rect 13613 43098 19570 43100
rect 13613 43042 13618 43098
rect 13674 43042 19570 43098
rect 13613 43040 19570 43042
rect 19640 43950 25452 44010
rect 13613 43037 13679 43040
rect 13521 42970 13587 42973
rect 19640 42970 19700 43950
rect 25446 43948 25452 43950
rect 25516 43948 25522 44012
rect 24894 43880 24900 43882
rect 13521 42968 19700 42970
rect 13521 42912 13526 42968
rect 13582 42912 19700 42968
rect 13521 42910 19700 42912
rect 19770 43820 24900 43880
rect 13521 42907 13587 42910
rect 13429 42840 13495 42843
rect 19770 42840 19830 43820
rect 24894 43818 24900 43820
rect 24964 43818 24970 43882
rect 24342 43750 24348 43752
rect 13429 42838 19830 42840
rect 13429 42782 13434 42838
rect 13490 42782 19830 42838
rect 13429 42780 19830 42782
rect 19900 43690 24348 43750
rect 13429 42777 13495 42780
rect 13337 42710 13403 42713
rect 19900 42710 19960 43690
rect 24342 43688 24348 43690
rect 24412 43688 24418 43752
rect 23790 43490 23796 43492
rect 13337 42708 19960 42710
rect 13337 42652 13342 42708
rect 13398 42652 19960 42708
rect 13337 42650 19960 42652
rect 20658 43430 23796 43490
rect 13337 42647 13403 42650
rect 5793 42450 5859 42453
rect 20478 42450 20484 42452
rect 5793 42448 20484 42450
rect 5793 42392 5798 42448
rect 5854 42392 20484 42448
rect 5793 42390 20484 42392
rect 5793 42387 5859 42390
rect 20478 42388 20484 42390
rect 20548 42388 20554 42452
rect 10577 42320 10643 42323
rect 19926 42320 19932 42322
rect 10577 42318 19932 42320
rect 10577 42262 10582 42318
rect 10638 42262 19932 42318
rect 10577 42260 19932 42262
rect 10577 42257 10643 42260
rect 19926 42258 19932 42260
rect 19996 42258 20002 42322
rect 11957 42190 12023 42193
rect 20658 42190 20718 43430
rect 23790 43428 23796 43430
rect 23860 43428 23866 43492
rect 11957 42188 20718 42190
rect 11957 42132 11962 42188
rect 12018 42132 20718 42188
rect 11957 42130 20718 42132
rect 11957 42127 12023 42130
rect 13981 42060 14047 42063
rect 19374 42060 19380 42062
rect 13981 42058 19380 42060
rect 13981 42002 13986 42058
rect 14042 42002 19380 42058
rect 13981 42000 19380 42002
rect 13981 41997 14047 42000
rect 19374 41998 19380 42000
rect 19444 41998 19450 42062
rect 19640 35050 21832 35110
rect 7633 32790 7699 32793
rect 19250 32790 19310 34808
rect 19377 34803 19443 34808
rect 19377 34747 19382 34803
rect 19438 34747 19443 34803
rect 19377 34742 19443 34747
rect 2930 32788 19310 32790
rect 2930 32732 7638 32788
rect 7694 32732 19310 32788
rect 2930 32730 19310 32732
rect 2930 28900 2990 32730
rect 7633 32727 7699 32730
rect 7725 32660 7791 32663
rect 19380 32660 19440 34742
rect 19510 34608 19570 34808
rect 19507 34603 19573 34608
rect 19507 34547 19512 34603
rect 19568 34547 19573 34603
rect 19507 34542 19573 34547
rect 3060 32658 19440 32660
rect 3060 32602 7730 32658
rect 7786 32602 19440 32658
rect 3060 32600 19440 32602
rect 3060 30628 3120 32600
rect 7725 32597 7791 32600
rect 7817 32530 7883 32533
rect 19510 32530 19570 34542
rect 3190 32528 19570 32530
rect 3190 32472 7822 32528
rect 7878 32472 19570 32528
rect 3190 32470 19570 32472
rect 3057 30623 3123 30628
rect 3057 30567 3062 30623
rect 3118 30567 3123 30623
rect 3057 30562 3123 30567
rect 1130 28840 2990 28900
rect 1130 22208 1190 28840
rect 3060 28770 3120 30562
rect 3190 30428 3250 32470
rect 7817 32467 7883 32470
rect 7908 32400 7974 32403
rect 19640 32400 19700 35050
rect 20550 34920 21372 34980
rect 19770 34408 19830 34808
rect 19767 34403 19833 34408
rect 19767 34347 19772 34403
rect 19828 34347 19833 34403
rect 19767 34342 19833 34347
rect 3320 32398 19700 32400
rect 3320 32342 7913 32398
rect 7969 32342 19700 32398
rect 3320 32340 19700 32342
rect 3187 30423 3253 30428
rect 3187 30367 3192 30423
rect 3248 30367 3253 30423
rect 3187 30362 3253 30367
rect 1260 28710 3120 28770
rect 1127 22203 1193 22208
rect 1127 22147 1132 22203
rect 1188 22147 1193 22203
rect 1127 22142 1193 22147
rect 1130 19942 1190 22142
rect 1260 22008 1320 28710
rect 3190 28640 3250 30362
rect 1390 28580 3250 28640
rect 1257 22003 1323 22008
rect 1257 21947 1262 22003
rect 1318 21947 1323 22003
rect 1257 21942 1323 21947
rect 1260 19942 1320 21942
rect 1390 21808 1450 28580
rect 3320 28513 3380 32340
rect 7908 32337 7974 32340
rect 8001 32270 8067 32273
rect 19770 32270 19830 34342
rect 19900 34208 19960 34808
rect 19897 34203 19963 34208
rect 19897 34147 19902 34203
rect 19958 34147 19963 34203
rect 19897 34142 19963 34147
rect 3450 32268 19830 32270
rect 3450 32212 8006 32268
rect 8062 32212 19830 32268
rect 3450 32210 19830 32212
rect 3450 30228 3510 32210
rect 8001 32207 8067 32210
rect 8093 32140 8159 32143
rect 19900 32140 19960 34142
rect 3580 32138 19960 32140
rect 3580 32082 8098 32138
rect 8154 32082 19960 32138
rect 3580 32080 19960 32082
rect 3447 30223 3513 30228
rect 3447 30167 3452 30223
rect 3508 30167 3513 30223
rect 3447 30162 3513 30167
rect 3317 28510 3383 28513
rect 1520 28508 3383 28510
rect 1520 28452 3322 28508
rect 3378 28452 3383 28508
rect 1520 28450 3383 28452
rect 1387 21803 1453 21808
rect 1387 21747 1392 21803
rect 1448 21747 1453 21803
rect 1387 21742 1453 21747
rect 1390 19942 1450 21742
rect 1520 4092 1580 28450
rect 3317 28447 3383 28450
rect 3450 28380 3510 30162
rect 3580 30028 3640 32080
rect 8093 32077 8159 32080
rect 8185 32010 8251 32013
rect 20030 32010 20090 34808
rect 3710 32008 20090 32010
rect 3710 31952 8190 32008
rect 8246 31952 20090 32008
rect 3710 31950 20090 31952
rect 3577 30023 3643 30028
rect 3577 29967 3582 30023
rect 3638 29967 3643 30023
rect 3577 29962 3643 29967
rect 1650 28320 3510 28380
rect 1650 21608 1710 28320
rect 3580 28250 3640 29962
rect 1780 28190 3640 28250
rect 1647 21603 1713 21608
rect 1647 21547 1652 21603
rect 1708 21547 1713 21603
rect 1647 21542 1713 21547
rect 1650 19942 1710 21542
rect 1780 21408 1840 28190
rect 3710 28120 3770 31950
rect 8185 31947 8251 31950
rect 8277 31880 8343 31883
rect 20160 31880 20220 34808
rect 20290 34008 20350 34808
rect 20287 34003 20353 34008
rect 20287 33947 20292 34003
rect 20348 33947 20353 34003
rect 20287 33942 20353 33947
rect 1910 28060 3770 28120
rect 3840 31878 20220 31880
rect 3840 31822 8282 31878
rect 8338 31822 20220 31878
rect 3840 31820 20220 31822
rect 1777 21403 1843 21408
rect 1777 21347 1782 21403
rect 1838 21347 1843 21403
rect 1777 21342 1843 21347
rect 1780 19942 1840 21342
rect 1910 21208 1970 28060
rect 3840 27990 3900 31820
rect 8277 31817 8343 31820
rect 8370 31750 8436 31753
rect 20290 31750 20350 33942
rect 20420 33208 20480 34808
rect 20417 33203 20483 33208
rect 20417 33147 20422 33203
rect 20478 33147 20483 33203
rect 20417 33142 20483 33147
rect 3970 31748 20350 31750
rect 3970 31692 8375 31748
rect 8431 31692 20350 31748
rect 3970 31690 20350 31692
rect 3970 29828 4030 31690
rect 8370 31687 8436 31690
rect 8461 31620 8527 31623
rect 20420 31620 20480 33142
rect 4100 31618 20480 31620
rect 4100 31562 8466 31618
rect 8522 31562 20480 31618
rect 4100 31560 20480 31562
rect 3967 29823 4033 29828
rect 3967 29767 3972 29823
rect 4028 29767 4033 29823
rect 3967 29762 4033 29767
rect 2040 27930 3900 27990
rect 1907 21203 1973 21208
rect 1907 21147 1912 21203
rect 1968 21147 1973 21203
rect 1907 21142 1973 21147
rect 1910 19942 1970 21142
rect 2040 21008 2100 27930
rect 3970 27860 4030 29762
rect 4100 29628 4160 31560
rect 8461 31557 8527 31560
rect 8553 31490 8619 31493
rect 20550 31490 20610 34920
rect 20680 33408 20740 34808
rect 20810 33608 20870 34808
rect 20940 33808 21000 34808
rect 20937 33803 21003 33808
rect 20937 33747 20942 33803
rect 20998 33747 21003 33803
rect 20937 33742 21003 33747
rect 20807 33603 20873 33608
rect 20807 33547 20812 33603
rect 20868 33547 20873 33603
rect 20807 33542 20873 33547
rect 20677 33403 20743 33408
rect 20677 33347 20682 33403
rect 20738 33347 20743 33403
rect 20677 33342 20743 33347
rect 4230 31488 20610 31490
rect 4230 31432 8558 31488
rect 8614 31432 20610 31488
rect 4230 31430 20610 31432
rect 4097 29623 4163 29628
rect 4097 29567 4102 29623
rect 4158 29567 4163 29623
rect 4097 29562 4163 29567
rect 2170 27800 4030 27860
rect 2037 21003 2103 21008
rect 2037 20947 2042 21003
rect 2098 20947 2103 21003
rect 2037 20942 2103 20947
rect 2040 19942 2100 20942
rect 2170 20008 2230 27800
rect 4100 27730 4160 29562
rect 4230 27733 4290 31430
rect 8553 31427 8619 31430
rect 8645 31360 8711 31363
rect 20680 31360 20740 33342
rect 4360 31358 20740 31360
rect 4360 31302 8650 31358
rect 8706 31302 20740 31358
rect 4360 31300 20740 31302
rect 4360 29028 4420 31300
rect 8645 31297 8711 31300
rect 8737 31230 8803 31233
rect 20810 31230 20870 33542
rect 4490 31228 20870 31230
rect 4490 31172 8742 31228
rect 8798 31172 20870 31228
rect 4490 31170 20870 31172
rect 4490 29228 4550 31170
rect 8737 31167 8803 31170
rect 8829 31100 8895 31103
rect 20940 31100 21000 33742
rect 4620 31098 21000 31100
rect 4620 31042 8834 31098
rect 8890 31042 21000 31098
rect 4620 31040 21000 31042
rect 4620 29428 4680 31040
rect 8829 31037 8895 31040
rect 21312 29734 21372 34920
rect 21309 29729 21375 29734
rect 21309 29673 21314 29729
rect 21370 29673 21375 29729
rect 21309 29668 21375 29673
rect 4617 29423 4683 29428
rect 4617 29367 4622 29423
rect 4678 29367 4683 29423
rect 4617 29362 4683 29367
rect 4487 29223 4553 29228
rect 4487 29167 4492 29223
rect 4548 29167 4553 29223
rect 4487 29162 4553 29167
rect 4357 29023 4423 29028
rect 4357 28967 4362 29023
rect 4418 28967 4423 29023
rect 4357 28962 4423 28967
rect 2300 27670 4160 27730
rect 4227 27728 4293 27733
rect 4227 27672 4232 27728
rect 4288 27672 4293 27728
rect 2300 20208 2360 27670
rect 4227 27667 4293 27672
rect 4230 27600 4290 27667
rect 2430 27540 4290 27600
rect 2297 20203 2363 20208
rect 2297 20147 2302 20203
rect 2358 20147 2363 20203
rect 2297 20142 2363 20147
rect 2167 20003 2233 20008
rect 2167 19947 2172 20003
rect 2228 19947 2233 20003
rect 2167 19942 2233 19947
rect 2300 19942 2360 20142
rect 2430 14104 2490 27540
rect 4360 27470 4420 28962
rect 2560 27410 4420 27470
rect 2560 20408 2620 27410
rect 4490 27340 4550 29162
rect 2690 27280 4550 27340
rect 2690 20608 2750 27280
rect 4620 27210 4680 29362
rect 2820 27150 4680 27210
rect 2820 20808 2880 27150
rect 21772 24744 21832 35050
rect 21769 24739 21835 24744
rect 21769 24683 21774 24739
rect 21830 24683 21835 24739
rect 21769 24678 21835 24683
rect 2817 20803 2883 20808
rect 2817 20747 2822 20803
rect 2878 20747 2883 20803
rect 2817 20742 2883 20747
rect 2687 20603 2753 20608
rect 2687 20547 2692 20603
rect 2748 20547 2753 20603
rect 2687 20542 2753 20547
rect 2557 20403 2623 20408
rect 2557 20347 2562 20403
rect 2618 20347 2623 20403
rect 2557 20342 2623 20347
rect 2560 19942 2620 20342
rect 2690 19942 2750 20542
rect 2820 19942 2880 20742
rect 2427 14099 2493 14104
rect 2427 14043 2432 14099
rect 2488 14043 2493 14099
rect 2427 14038 2493 14043
rect 2430 14029 2490 14038
rect 1517 4087 1583 4092
rect 1517 4031 1522 4087
rect 1578 4031 1583 4087
rect 1517 4026 1583 4031
rect 1520 4017 1580 4026
<< via3 >>
rect 7236 44950 7300 45014
rect 11100 44950 11164 45014
rect 14964 44950 15028 45014
rect 28764 44728 28828 44792
rect 28212 44598 28276 44662
rect 18828 44468 18892 44532
rect 18276 44338 18340 44402
rect 17724 44208 17788 44272
rect 17172 44078 17236 44142
rect 16620 43948 16684 44012
rect 14412 43818 14476 43882
rect 13860 43688 13924 43752
rect 13308 43558 13372 43622
rect 12756 43428 12820 43492
rect 27660 44468 27724 44532
rect 12204 43298 12268 43362
rect 27108 44338 27172 44402
rect 26556 44208 26620 44272
rect 26004 44078 26068 44142
rect 25452 43948 25516 44012
rect 24900 43818 24964 43882
rect 24348 43688 24412 43752
rect 20484 42388 20548 42452
rect 19932 42258 19996 42322
rect 23796 43428 23860 43492
rect 19380 41998 19444 42062
rect 8001 29345 8249 29593
rect 14105 29345 14353 29593
rect 8351 28995 8599 29243
rect 14455 28995 14703 29243
rect 8001 28811 8249 28909
rect 14105 28811 14353 28909
rect 25351 33725 25599 33973
rect 30351 33725 30599 33973
rect 25001 33375 25249 33623
rect 30001 33375 30249 33623
rect 25351 33191 25599 33289
rect 30351 33191 30599 33289
rect 8001 20725 8249 20973
rect 14105 20725 14353 20973
rect 25351 20725 25599 20973
rect 30351 20725 30599 20973
rect 8351 20375 8599 20623
rect 14455 20375 14703 20623
rect 25001 20375 25249 20623
rect 30001 20375 30249 20623
rect 8001 20191 8249 20289
rect 14105 20191 14353 20289
rect 25351 20191 25599 20289
rect 30351 20191 30599 20289
<< metal4 >>
rect 6134 45012 6194 45152
rect 6686 45012 6746 45152
rect 7238 45015 7298 45152
rect 7235 45014 7301 45015
rect 7235 45012 7236 45014
rect 6134 44952 7236 45012
rect 7235 44950 7236 44952
rect 7300 44950 7301 45014
rect 7790 45012 7850 45152
rect 8342 45012 8402 45152
rect 8894 45012 8954 45152
rect 9446 45012 9506 45152
rect 9998 45012 10058 45152
rect 7790 44952 10058 45012
rect 10550 45012 10610 45152
rect 11102 45015 11162 45152
rect 11099 45014 11165 45015
rect 11099 45012 11100 45014
rect 10550 44952 11100 45012
rect 7235 44949 7301 44950
rect 7238 44840 7298 44949
rect 7238 44780 8060 44840
rect 8000 43152 8060 44780
rect 8350 43152 8410 44952
rect 11099 44950 11100 44952
rect 11164 45012 11165 45014
rect 11654 45012 11714 45152
rect 11164 44952 11714 45012
rect 11164 44950 11165 44952
rect 11099 44949 11165 44950
rect 12206 43363 12266 45152
rect 12758 43493 12818 45152
rect 13310 43623 13370 45152
rect 13862 43753 13922 45152
rect 14414 43883 14474 45152
rect 14966 45015 15026 45152
rect 14963 45014 15029 45015
rect 14963 44950 14964 45014
rect 15028 45012 15029 45014
rect 15518 45012 15578 45152
rect 16070 45012 16130 45152
rect 15028 44952 16130 45012
rect 15028 44950 15029 44952
rect 14963 44949 15029 44950
rect 16622 44013 16682 45152
rect 17174 44143 17234 45152
rect 17726 44273 17786 45152
rect 18278 44403 18338 45152
rect 18830 44533 18890 45152
rect 18827 44532 18893 44533
rect 18827 44468 18828 44532
rect 18892 44468 18893 44532
rect 18827 44467 18893 44468
rect 18275 44402 18341 44403
rect 18275 44338 18276 44402
rect 18340 44338 18341 44402
rect 18275 44337 18341 44338
rect 17723 44272 17789 44273
rect 17723 44208 17724 44272
rect 17788 44208 17789 44272
rect 17723 44207 17789 44208
rect 17171 44142 17237 44143
rect 17171 44078 17172 44142
rect 17236 44078 17237 44142
rect 17171 44077 17237 44078
rect 16619 44012 16685 44013
rect 16619 43948 16620 44012
rect 16684 43948 16685 44012
rect 16619 43947 16685 43948
rect 14411 43882 14477 43883
rect 14411 43818 14412 43882
rect 14476 43818 14477 43882
rect 14411 43817 14477 43818
rect 13859 43752 13925 43753
rect 13859 43688 13860 43752
rect 13924 43688 13925 43752
rect 13859 43687 13925 43688
rect 13307 43622 13373 43623
rect 13307 43558 13308 43622
rect 13372 43558 13373 43622
rect 13307 43557 13373 43558
rect 12755 43492 12821 43493
rect 12755 43428 12756 43492
rect 12820 43428 12821 43492
rect 12755 43427 12821 43428
rect 12203 43362 12269 43363
rect 12203 43298 12204 43362
rect 12268 43298 12269 43362
rect 12203 43297 12269 43298
rect 2928 2000 3178 43152
rect 3278 2000 3528 43152
rect 8000 29593 8250 43152
rect 8000 29345 8001 29593
rect 8249 29345 8250 29593
rect 8000 28909 8250 29345
rect 8000 28811 8001 28909
rect 8249 28811 8250 28909
rect 8000 20973 8250 28811
rect 8000 20725 8001 20973
rect 8249 20725 8250 20973
rect 8000 20289 8250 20725
rect 8000 20191 8001 20289
rect 8249 20191 8250 20289
rect 8000 2000 8250 20191
rect 8350 29243 8600 43152
rect 8350 28995 8351 29243
rect 8599 28995 8600 29243
rect 8350 20623 8600 28995
rect 8350 20375 8351 20623
rect 8599 20375 8600 20623
rect 8350 2000 8600 20375
rect 14104 29593 14354 43152
rect 14104 29345 14105 29593
rect 14353 29345 14354 29593
rect 14104 28909 14354 29345
rect 14104 28811 14105 28909
rect 14353 28811 14354 28909
rect 14104 20973 14354 28811
rect 14104 20725 14105 20973
rect 14353 20725 14354 20973
rect 14104 20289 14354 20725
rect 14104 20191 14105 20289
rect 14353 20191 14354 20289
rect 14104 2000 14354 20191
rect 14454 29243 14704 43152
rect 19382 42063 19442 45152
rect 19934 42323 19994 45152
rect 20486 42453 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 43493 23858 45152
rect 24350 43753 24410 45152
rect 24902 43883 24962 45152
rect 25454 44013 25514 45152
rect 26006 44143 26066 45152
rect 26558 44273 26618 45152
rect 27110 44403 27170 45152
rect 27662 44533 27722 45152
rect 28214 44663 28274 45152
rect 28766 44793 28826 45152
rect 29318 44952 29378 45152
rect 28763 44792 28829 44793
rect 28763 44728 28764 44792
rect 28828 44728 28829 44792
rect 28763 44727 28829 44728
rect 28211 44662 28277 44663
rect 28211 44598 28212 44662
rect 28276 44598 28277 44662
rect 28211 44597 28277 44598
rect 27659 44532 27725 44533
rect 27659 44468 27660 44532
rect 27724 44468 27725 44532
rect 27659 44467 27725 44468
rect 27107 44402 27173 44403
rect 27107 44338 27108 44402
rect 27172 44338 27173 44402
rect 27107 44337 27173 44338
rect 26555 44272 26621 44273
rect 26555 44208 26556 44272
rect 26620 44208 26621 44272
rect 26555 44207 26621 44208
rect 26003 44142 26069 44143
rect 26003 44078 26004 44142
rect 26068 44078 26069 44142
rect 26003 44077 26069 44078
rect 25451 44012 25517 44013
rect 25451 43948 25452 44012
rect 25516 43948 25517 44012
rect 25451 43947 25517 43948
rect 24899 43882 24965 43883
rect 24899 43818 24900 43882
rect 24964 43818 24965 43882
rect 24899 43817 24965 43818
rect 24347 43752 24413 43753
rect 24347 43688 24348 43752
rect 24412 43688 24413 43752
rect 24347 43687 24413 43688
rect 23795 43492 23861 43493
rect 23795 43428 23796 43492
rect 23860 43428 23861 43492
rect 23795 43427 23861 43428
rect 20483 42452 20549 42453
rect 20483 42388 20484 42452
rect 20548 42388 20549 42452
rect 20483 42387 20549 42388
rect 19931 42322 19997 42323
rect 19931 42258 19932 42322
rect 19996 42258 19997 42322
rect 19931 42257 19997 42258
rect 19379 42062 19445 42063
rect 19379 41998 19380 42062
rect 19444 41998 19445 42062
rect 19379 41997 19445 41998
rect 14454 28995 14455 29243
rect 14703 28995 14704 29243
rect 14454 20623 14704 28995
rect 14454 20375 14455 20623
rect 14703 20375 14704 20623
rect 14454 2000 14704 20375
rect 25000 33623 25250 43152
rect 25000 33375 25001 33623
rect 25249 33375 25250 33623
rect 25000 20623 25250 33375
rect 25000 20375 25001 20623
rect 25249 20375 25250 20623
rect 25000 2000 25250 20375
rect 25350 33973 25600 43152
rect 25350 33725 25351 33973
rect 25599 33725 25600 33973
rect 25350 33289 25600 33725
rect 25350 33191 25351 33289
rect 25599 33191 25600 33289
rect 25350 20973 25600 33191
rect 25350 20725 25351 20973
rect 25599 20725 25600 20973
rect 25350 20289 25600 20725
rect 25350 20191 25351 20289
rect 25599 20191 25600 20289
rect 25350 2000 25600 20191
rect 30000 33623 30250 43152
rect 30000 33375 30001 33623
rect 30249 33375 30250 33623
rect 30000 20623 30250 33375
rect 30000 20375 30001 20623
rect 30249 20375 30250 20623
rect 30000 2000 30250 20375
rect 30350 33973 30600 43152
rect 30350 33725 30351 33973
rect 30599 33725 30600 33973
rect 30350 33289 30600 33725
rect 30350 33191 30351 33289
rect 30599 33191 30600 33289
rect 30350 20973 30600 33191
rect 30350 20725 30351 20973
rect 30599 20725 30600 20973
rect 30350 20289 30600 20725
rect 30350 20191 30351 20289
rect 30599 20191 30600 20289
rect 30350 2000 30600 20191
use control  control_0
timestamp 1730654005
transform 1 0 2928 0 1 33116
box -2746 -116 11814 8820
use rom_4k_0  rom_4k_0_0
timestamp 1730749399
transform -1 0 31980 0 -1 35063
box 11 0 9780 12063
use rom_4k_1  rom_4k_1_0
timestamp 1730748763
transform -1 0 20980 0 -1 30883
box 11 0 16180 7283
use rom_32k  rom_32k_0
timestamp 1730749471
transform -1 0 31980 0 -1 22463
box 11 0 28980 22423
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 3 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 4 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 5 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 6 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 7 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 8 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 9 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 10 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 11 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 12 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 13 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 14 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 15 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 16 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 17 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 18 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 19 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 20 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 21 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 22 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 23 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 24 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 25 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 26 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 27 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 28 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 29 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 30 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 31 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 32 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 33 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 34 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 35 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 36 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 37 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 38 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 39 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 40 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 41 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 42 nsew signal output
flabel metal4 2928 2000 3178 43152 1 FreeSans 160 0 0 0 VGND
port 43 n ground input
flabel metal4 14104 2000 14354 43152 1 FreeSans 160 0 0 0 VGND
port 43 n
flabel metal4 8000 2000 8250 43152 1 FreeSans 160 0 0 0 VGND
port 43 n
flabel metal4 25350 2000 25600 43152 1 FreeSans 160 0 0 0 VGND
port 43 n
flabel metal4 30350 2000 30600 43152 1 FreeSans 160 0 0 0 VGND
port 43 n
flabel metal4 3278 2000 3528 43152 1 FreeSans 160 0 0 0 VDPWR
port 44 n power input
flabel metal4 8350 2000 8600 43152 1 FreeSans 160 0 0 0 VDPWR
port 44 n
flabel metal4 14454 2000 14704 43152 1 FreeSans 160 0 0 0 VDPWR
port 44 n
flabel metal4 25000 2000 25250 43152 1 FreeSans 160 0 0 0 VDPWR
port 44 n
flabel metal4 30000 2000 30250 43152 1 FreeSans 160 0 0 0 VDPWR
port 44 n
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
