magic
tech sky130A
magscale 1 2
timestamp 1730660070
<< nwell >>
rect -169 -778 6439 -294
rect 8380 -1973 9162 123
<< pwell >>
rect 90 9819 6380 10047
rect -10 5071 7496 9819
rect 90 4839 6380 5071
rect -10 91 7496 4839
rect -10 -1 6436 91
rect -166 -87 6436 -1
rect -120 -236 6390 -87
rect -36 -2013 6306 -820
rect 8114 -1963 8316 113
rect 9226 -1963 9428 113
<< nmos >>
rect 8140 -90 8290 -60
rect 9252 -90 9402 -60
rect -30 -210 0 -126
rect 70 -210 100 -126
rect 170 -210 200 -126
rect 270 -210 300 -126
rect 370 -210 400 -126
rect 470 -210 500 -126
rect 570 -210 600 -126
rect 670 -210 700 -126
rect 770 -210 800 -126
rect 870 -210 900 -126
rect 970 -210 1000 -126
rect 1070 -210 1100 -126
rect 1170 -210 1200 -126
rect 1270 -210 1300 -126
rect 1370 -210 1400 -126
rect 1470 -210 1500 -126
rect 1570 -210 1600 -126
rect 1670 -210 1700 -126
rect 1770 -210 1800 -126
rect 1870 -210 1900 -126
rect 1970 -210 2000 -126
rect 2070 -210 2100 -126
rect 2170 -210 2200 -126
rect 2270 -210 2300 -126
rect 2370 -210 2400 -126
rect 2470 -210 2500 -126
rect 2570 -210 2600 -126
rect 2670 -210 2700 -126
rect 2770 -210 2800 -126
rect 2870 -210 2900 -126
rect 2970 -210 3000 -126
rect 3070 -210 3100 -126
rect 3170 -210 3200 -126
rect 3270 -210 3300 -126
rect 3370 -210 3400 -126
rect 3470 -210 3500 -126
rect 3570 -210 3600 -126
rect 3670 -210 3700 -126
rect 3770 -210 3800 -126
rect 3870 -210 3900 -126
rect 3970 -210 4000 -126
rect 4070 -210 4100 -126
rect 4170 -210 4200 -126
rect 4270 -210 4300 -126
rect 4370 -210 4400 -126
rect 4470 -210 4500 -126
rect 4570 -210 4600 -126
rect 4670 -210 4700 -126
rect 4770 -210 4800 -126
rect 4870 -210 4900 -126
rect 4970 -210 5000 -126
rect 5070 -210 5100 -126
rect 5170 -210 5200 -126
rect 5270 -210 5300 -126
rect 5370 -210 5400 -126
rect 5470 -210 5500 -126
rect 5570 -210 5600 -126
rect 5670 -210 5700 -126
rect 5770 -210 5800 -126
rect 5870 -210 5900 -126
rect 5970 -210 6000 -126
rect 6070 -210 6100 -126
rect 6170 -210 6200 -126
rect 6270 -210 6300 -126
rect 8140 -190 8290 -160
rect 9252 -190 9402 -160
rect 8140 -290 8290 -260
rect 9252 -290 9402 -260
rect 8140 -390 8290 -360
rect 9252 -390 9402 -360
rect 8140 -490 8290 -460
rect 9252 -490 9402 -460
rect 8140 -590 8290 -560
rect 9252 -590 9402 -560
rect 8140 -690 8290 -660
rect 9252 -690 9402 -660
rect 8140 -790 8290 -760
rect 9252 -790 9402 -760
rect 8140 -890 8290 -860
rect 9252 -890 9402 -860
rect 8140 -990 8290 -960
rect 9252 -990 9402 -960
rect 8140 -1090 8290 -1060
rect 9252 -1090 9402 -1060
rect 8140 -1190 8290 -1160
rect 9252 -1190 9402 -1160
rect 8140 -1290 8290 -1260
rect 9252 -1290 9402 -1260
rect 8140 -1390 8290 -1360
rect 9252 -1390 9402 -1360
rect 8140 -1490 8290 -1460
rect 9252 -1490 9402 -1460
rect 8140 -1590 8290 -1560
rect 9252 -1590 9402 -1560
rect 8140 -1690 8290 -1660
rect 9252 -1690 9402 -1660
rect 8140 -1790 8290 -1760
rect 9252 -1790 9402 -1760
<< pmos >>
rect 8416 -90 8716 -60
rect 8826 -90 9126 -60
rect 8416 -190 8716 -160
rect 8826 -190 9126 -160
rect 8416 -290 8716 -260
rect 8826 -290 9126 -260
rect 8416 -390 8716 -360
rect 8826 -390 9126 -360
rect 8416 -490 8716 -460
rect 8826 -490 9126 -460
rect 8416 -590 8716 -560
rect 8826 -590 9126 -560
rect 15 -742 107 -658
rect 163 -742 255 -658
rect 415 -742 507 -658
rect 563 -742 655 -658
rect 815 -742 907 -658
rect 963 -742 1055 -658
rect 1215 -742 1307 -658
rect 1363 -742 1455 -658
rect 1615 -742 1707 -658
rect 1763 -742 1855 -658
rect 2015 -742 2107 -658
rect 2163 -742 2255 -658
rect 2415 -742 2507 -658
rect 2563 -742 2655 -658
rect 2815 -742 2907 -658
rect 2963 -742 3055 -658
rect 3215 -742 3307 -658
rect 3363 -742 3455 -658
rect 3615 -742 3707 -658
rect 3763 -742 3855 -658
rect 4015 -742 4107 -658
rect 4163 -742 4255 -658
rect 4415 -742 4507 -658
rect 4563 -742 4655 -658
rect 4815 -742 4907 -658
rect 4963 -742 5055 -658
rect 5215 -742 5307 -658
rect 5363 -742 5455 -658
rect 5615 -742 5707 -658
rect 5763 -742 5855 -658
rect 6015 -742 6107 -658
rect 6163 -742 6255 -658
rect 8416 -690 8716 -660
rect 8826 -690 9126 -660
rect 8416 -790 8716 -760
rect 8826 -790 9126 -760
rect 8416 -890 8716 -860
rect 8826 -890 9126 -860
rect 8416 -990 8716 -960
rect 8826 -990 9126 -960
rect 8416 -1090 8716 -1060
rect 8826 -1090 9126 -1060
rect 8416 -1190 8716 -1160
rect 8826 -1190 9126 -1160
rect 8416 -1290 8716 -1260
rect 8826 -1290 9126 -1260
rect 8416 -1390 8716 -1360
rect 8826 -1390 9126 -1360
rect 8416 -1490 8716 -1460
rect 8826 -1490 9126 -1460
rect 8416 -1590 8716 -1560
rect 8826 -1590 9126 -1560
rect 8416 -1690 8716 -1660
rect 8826 -1690 9126 -1660
rect 8416 -1790 8716 -1760
rect 8826 -1790 9126 -1760
<< pmoshvt >>
rect -30 -498 0 -330
rect 70 -498 100 -330
rect 170 -498 200 -330
rect 270 -498 300 -330
rect 370 -498 400 -330
rect 470 -498 500 -330
rect 570 -498 600 -330
rect 670 -498 700 -330
rect 770 -498 800 -330
rect 870 -498 900 -330
rect 970 -498 1000 -330
rect 1070 -498 1100 -330
rect 1170 -498 1200 -330
rect 1270 -498 1300 -330
rect 1370 -498 1400 -330
rect 1470 -498 1500 -330
rect 1570 -498 1600 -330
rect 1670 -498 1700 -330
rect 1770 -498 1800 -330
rect 1870 -498 1900 -330
rect 1970 -498 2000 -330
rect 2070 -498 2100 -330
rect 2170 -498 2200 -330
rect 2270 -498 2300 -330
rect 2370 -498 2400 -330
rect 2470 -498 2500 -330
rect 2570 -498 2600 -330
rect 2670 -498 2700 -330
rect 2770 -498 2800 -330
rect 2870 -498 2900 -330
rect 2970 -498 3000 -330
rect 3070 -498 3100 -330
rect 3170 -498 3200 -330
rect 3270 -498 3300 -330
rect 3370 -498 3400 -330
rect 3470 -498 3500 -330
rect 3570 -498 3600 -330
rect 3670 -498 3700 -330
rect 3770 -498 3800 -330
rect 3870 -498 3900 -330
rect 3970 -498 4000 -330
rect 4070 -498 4100 -330
rect 4170 -498 4200 -330
rect 4270 -498 4300 -330
rect 4370 -498 4400 -330
rect 4470 -498 4500 -330
rect 4570 -498 4600 -330
rect 4670 -498 4700 -330
rect 4770 -498 4800 -330
rect 4870 -498 4900 -330
rect 4970 -498 5000 -330
rect 5070 -498 5100 -330
rect 5170 -498 5200 -330
rect 5270 -498 5300 -330
rect 5370 -498 5400 -330
rect 5470 -498 5500 -330
rect 5570 -498 5600 -330
rect 5670 -498 5700 -330
rect 5770 -498 5800 -330
rect 5870 -498 5900 -330
rect 5970 -498 6000 -330
rect 6070 -498 6100 -330
rect 6170 -498 6200 -330
rect 6270 -498 6300 -330
<< nmoslvt >>
rect 70 9707 100 9793
rect 170 9707 200 9793
rect 270 9707 300 9793
rect 370 9707 400 9793
rect 470 9707 500 9793
rect 570 9707 600 9793
rect 670 9707 700 9793
rect 770 9707 800 9793
rect 870 9707 900 9793
rect 970 9707 1000 9793
rect 1070 9707 1100 9793
rect 1170 9707 1200 9793
rect 1270 9707 1300 9793
rect 1370 9707 1400 9793
rect 1470 9707 1500 9793
rect 70 9567 100 9653
rect 170 9567 200 9653
rect 270 9567 300 9653
rect 370 9567 400 9653
rect 470 9567 500 9653
rect 570 9567 600 9653
rect 70 9427 100 9513
rect 170 9427 200 9513
rect 270 9427 300 9513
rect 370 9427 400 9513
rect 1670 9707 1700 9793
rect 1770 9707 1800 9793
rect 1870 9707 1900 9793
rect 1970 9707 2000 9793
rect 2070 9707 2100 9793
rect 770 9567 800 9653
rect 870 9567 900 9653
rect 970 9567 1000 9653
rect 1070 9567 1100 9653
rect 1170 9567 1200 9653
rect 1270 9567 1300 9653
rect 1370 9567 1400 9653
rect 1470 9567 1500 9653
rect 1570 9567 1600 9653
rect 1670 9567 1700 9653
rect 1770 9567 1800 9653
rect 1870 9567 1900 9653
rect 1970 9567 2000 9653
rect 2070 9567 2100 9653
rect 570 9427 600 9513
rect 670 9427 700 9513
rect 770 9427 800 9513
rect 870 9427 900 9513
rect 1070 9427 1100 9513
rect 1270 9427 1300 9513
rect 1370 9427 1400 9513
rect 1470 9427 1500 9513
rect 1570 9427 1600 9513
rect 1670 9427 1700 9513
rect 70 9287 100 9373
rect 170 9287 200 9373
rect 270 9287 300 9373
rect 370 9287 400 9373
rect 470 9287 500 9373
rect 570 9287 600 9373
rect 670 9287 700 9373
rect 770 9287 800 9373
rect 870 9287 900 9373
rect 970 9287 1000 9373
rect 1070 9287 1100 9373
rect 1170 9287 1200 9373
rect 1270 9287 1300 9373
rect 1370 9287 1400 9373
rect 1470 9287 1500 9373
rect 1570 9287 1600 9373
rect 1670 9287 1700 9373
rect 70 9147 100 9233
rect 170 9147 200 9233
rect 270 9147 300 9233
rect 370 9147 400 9233
rect 470 9147 500 9233
rect 570 9147 600 9233
rect 670 9147 700 9233
rect 770 9147 800 9233
rect 870 9147 900 9233
rect 970 9147 1000 9233
rect 1070 9147 1100 9233
rect 1170 9147 1200 9233
rect 1270 9147 1300 9233
rect 1370 9147 1400 9233
rect 1470 9147 1500 9233
rect 70 9007 100 9093
rect 170 9007 200 9093
rect 270 9007 300 9093
rect 370 9007 400 9093
rect 470 9007 500 9093
rect 570 9007 600 9093
rect 1870 9427 1900 9513
rect 1970 9427 2000 9513
rect 2270 9707 2300 9793
rect 2370 9707 2400 9793
rect 2470 9707 2500 9793
rect 2570 9707 2600 9793
rect 2670 9707 2700 9793
rect 2270 9567 2300 9653
rect 2170 9427 2200 9513
rect 2270 9427 2300 9513
rect 2870 9707 2900 9793
rect 2970 9707 3000 9793
rect 3070 9707 3100 9793
rect 3170 9707 3200 9793
rect 2470 9567 2500 9653
rect 2570 9567 2600 9653
rect 2670 9567 2700 9653
rect 2770 9567 2800 9653
rect 2870 9567 2900 9653
rect 2470 9427 2500 9513
rect 2670 9427 2700 9513
rect 3370 9707 3400 9793
rect 3470 9707 3500 9793
rect 3670 9707 3700 9793
rect 3770 9707 3800 9793
rect 3870 9707 3900 9793
rect 3970 9707 4000 9793
rect 4070 9707 4100 9793
rect 4170 9707 4200 9793
rect 4270 9707 4300 9793
rect 4370 9707 4400 9793
rect 4470 9707 4500 9793
rect 4570 9707 4600 9793
rect 4670 9707 4700 9793
rect 4770 9707 4800 9793
rect 4870 9707 4900 9793
rect 4970 9707 5000 9793
rect 5070 9707 5100 9793
rect 5170 9707 5200 9793
rect 5270 9707 5300 9793
rect 5370 9707 5400 9793
rect 3070 9567 3100 9653
rect 3170 9567 3200 9653
rect 3270 9567 3300 9653
rect 3370 9567 3400 9653
rect 3470 9567 3500 9653
rect 3570 9567 3600 9653
rect 3670 9567 3700 9653
rect 3770 9567 3800 9653
rect 3870 9567 3900 9653
rect 3970 9567 4000 9653
rect 2870 9427 2900 9513
rect 2970 9427 3000 9513
rect 3070 9427 3100 9513
rect 3170 9427 3200 9513
rect 3270 9427 3300 9513
rect 3370 9427 3400 9513
rect 3470 9427 3500 9513
rect 3570 9427 3600 9513
rect 3670 9427 3700 9513
rect 3770 9427 3800 9513
rect 3870 9427 3900 9513
rect 3970 9427 4000 9513
rect 5570 9707 5600 9793
rect 5670 9707 5700 9793
rect 5870 9707 5900 9793
rect 4170 9567 4200 9653
rect 4270 9567 4300 9653
rect 4370 9567 4400 9653
rect 4470 9567 4500 9653
rect 4570 9567 4600 9653
rect 4670 9567 4700 9653
rect 4770 9567 4800 9653
rect 4870 9567 4900 9653
rect 4970 9567 5000 9653
rect 5070 9567 5100 9653
rect 5170 9567 5200 9653
rect 5270 9567 5300 9653
rect 5370 9567 5400 9653
rect 5470 9567 5500 9653
rect 5570 9567 5600 9653
rect 5670 9567 5700 9653
rect 5770 9567 5800 9653
rect 5870 9567 5900 9653
rect 4170 9427 4200 9513
rect 4270 9427 4300 9513
rect 4370 9427 4400 9513
rect 4470 9427 4500 9513
rect 1870 9287 1900 9373
rect 1970 9287 2000 9373
rect 2070 9287 2100 9373
rect 2170 9287 2200 9373
rect 2270 9287 2300 9373
rect 2370 9287 2400 9373
rect 2470 9287 2500 9373
rect 2570 9287 2600 9373
rect 2670 9287 2700 9373
rect 2770 9287 2800 9373
rect 2870 9287 2900 9373
rect 2970 9287 3000 9373
rect 3070 9287 3100 9373
rect 3170 9287 3200 9373
rect 3270 9287 3300 9373
rect 3370 9287 3400 9373
rect 3470 9287 3500 9373
rect 3570 9287 3600 9373
rect 3670 9287 3700 9373
rect 3770 9287 3800 9373
rect 3870 9287 3900 9373
rect 3970 9287 4000 9373
rect 4070 9287 4100 9373
rect 1670 9147 1700 9233
rect 1770 9147 1800 9233
rect 1870 9147 1900 9233
rect 1970 9147 2000 9233
rect 2070 9147 2100 9233
rect 2170 9147 2200 9233
rect 2270 9147 2300 9233
rect 2370 9147 2400 9233
rect 770 9007 800 9093
rect 870 9007 900 9093
rect 970 9007 1000 9093
rect 1070 9007 1100 9093
rect 1170 9007 1200 9093
rect 1270 9007 1300 9093
rect 1370 9007 1400 9093
rect 1470 9007 1500 9093
rect 1570 9007 1600 9093
rect 1670 9007 1700 9093
rect 1870 9007 1900 9093
rect 2570 9147 2600 9233
rect 2670 9147 2700 9233
rect 2770 9147 2800 9233
rect 2870 9147 2900 9233
rect 2970 9147 3000 9233
rect 3070 9147 3100 9233
rect 3170 9147 3200 9233
rect 3270 9147 3300 9233
rect 3370 9147 3400 9233
rect 3470 9147 3500 9233
rect 3570 9147 3600 9233
rect 3670 9147 3700 9233
rect 3770 9147 3800 9233
rect 3870 9147 3900 9233
rect 3970 9147 4000 9233
rect 2070 9007 2100 9093
rect 2170 9007 2200 9093
rect 2270 9007 2300 9093
rect 2370 9007 2400 9093
rect 2470 9007 2500 9093
rect 2570 9007 2600 9093
rect 70 8867 100 8953
rect 170 8867 200 8953
rect 270 8867 300 8953
rect 370 8867 400 8953
rect 470 8867 500 8953
rect 570 8867 600 8953
rect 670 8867 700 8953
rect 770 8867 800 8953
rect 870 8867 900 8953
rect 970 8867 1000 8953
rect 1070 8867 1100 8953
rect 1170 8867 1200 8953
rect 1270 8867 1300 8953
rect 1370 8867 1400 8953
rect 1470 8867 1500 8953
rect 1570 8867 1600 8953
rect 1670 8867 1700 8953
rect 1770 8867 1800 8953
rect 1870 8867 1900 8953
rect 1970 8867 2000 8953
rect 2070 8867 2100 8953
rect 2170 8867 2200 8953
rect 2270 8867 2300 8953
rect 2370 8867 2400 8953
rect 2470 8867 2500 8953
rect 2570 8867 2600 8953
rect 70 8727 100 8813
rect 170 8727 200 8813
rect 370 8727 400 8813
rect 470 8727 500 8813
rect 570 8727 600 8813
rect 670 8727 700 8813
rect 770 8727 800 8813
rect 870 8727 900 8813
rect 970 8727 1000 8813
rect 1070 8727 1100 8813
rect 1170 8727 1200 8813
rect 1270 8727 1300 8813
rect 1370 8727 1400 8813
rect 1470 8727 1500 8813
rect 1570 8727 1600 8813
rect 1670 8727 1700 8813
rect 1770 8727 1800 8813
rect 1870 8727 1900 8813
rect 1970 8727 2000 8813
rect 2070 8727 2100 8813
rect 2170 8727 2200 8813
rect 2270 8727 2300 8813
rect 2370 8727 2400 8813
rect 2470 8727 2500 8813
rect 2570 8727 2600 8813
rect 70 8497 100 8583
rect 170 8497 200 8583
rect 270 8497 300 8583
rect 370 8497 400 8583
rect 470 8497 500 8583
rect 570 8497 600 8583
rect 670 8497 700 8583
rect 770 8497 800 8583
rect 970 8497 1000 8583
rect 2770 9007 2800 9093
rect 2970 9007 3000 9093
rect 3070 9007 3100 9093
rect 3170 9007 3200 9093
rect 4670 9427 4700 9513
rect 4770 9427 4800 9513
rect 4970 9427 5000 9513
rect 5170 9427 5200 9513
rect 5370 9427 5400 9513
rect 5470 9427 5500 9513
rect 5570 9427 5600 9513
rect 5770 9427 5800 9513
rect 6070 9707 6100 9793
rect 6170 9707 6200 9793
rect 6270 9707 6300 9793
rect 6370 9707 6400 9793
rect 6570 9707 6600 9793
rect 6670 9707 6700 9793
rect 6880 9707 6910 9793
rect 6980 9707 7010 9793
rect 7080 9707 7110 9793
rect 7180 9707 7210 9793
rect 7280 9707 7310 9793
rect 7380 9707 7410 9793
rect 6070 9567 6100 9653
rect 6170 9567 6200 9653
rect 6270 9567 6300 9653
rect 6370 9567 6400 9653
rect 6570 9567 6600 9653
rect 6670 9567 6700 9653
rect 6880 9567 6910 9653
rect 6980 9567 7010 9653
rect 7080 9567 7110 9653
rect 7180 9567 7210 9653
rect 7280 9567 7310 9653
rect 7380 9567 7410 9653
rect 5970 9427 6000 9513
rect 6070 9427 6100 9513
rect 6270 9427 6300 9513
rect 6370 9427 6400 9513
rect 6570 9427 6600 9513
rect 6670 9427 6700 9513
rect 6880 9427 6910 9513
rect 6980 9427 7010 9513
rect 7080 9427 7110 9513
rect 7180 9427 7210 9513
rect 7280 9427 7310 9513
rect 7380 9427 7410 9513
rect 4270 9287 4300 9373
rect 4370 9287 4400 9373
rect 4470 9287 4500 9373
rect 4570 9287 4600 9373
rect 4670 9287 4700 9373
rect 4770 9287 4800 9373
rect 4870 9287 4900 9373
rect 4970 9287 5000 9373
rect 5070 9287 5100 9373
rect 5170 9287 5200 9373
rect 5270 9287 5300 9373
rect 5370 9287 5400 9373
rect 5470 9287 5500 9373
rect 5570 9287 5600 9373
rect 5670 9287 5700 9373
rect 5770 9287 5800 9373
rect 5870 9287 5900 9373
rect 5970 9287 6000 9373
rect 6070 9287 6100 9373
rect 6170 9287 6200 9373
rect 6270 9287 6300 9373
rect 6370 9287 6400 9373
rect 6570 9287 6600 9373
rect 6670 9287 6700 9373
rect 6880 9287 6910 9373
rect 6980 9287 7010 9373
rect 7080 9287 7110 9373
rect 7180 9287 7210 9373
rect 7280 9287 7310 9373
rect 7380 9287 7410 9373
rect 4170 9147 4200 9233
rect 4270 9147 4300 9233
rect 4370 9147 4400 9233
rect 4470 9147 4500 9233
rect 4570 9147 4600 9233
rect 4670 9147 4700 9233
rect 4770 9147 4800 9233
rect 4870 9147 4900 9233
rect 4970 9147 5000 9233
rect 3370 9007 3400 9093
rect 3470 9007 3500 9093
rect 3570 9007 3600 9093
rect 3670 9007 3700 9093
rect 3770 9007 3800 9093
rect 3870 9007 3900 9093
rect 3970 9007 4000 9093
rect 4070 9007 4100 9093
rect 4170 9007 4200 9093
rect 4270 9007 4300 9093
rect 4370 9007 4400 9093
rect 4470 9007 4500 9093
rect 2770 8867 2800 8953
rect 2870 8867 2900 8953
rect 2970 8867 3000 8953
rect 3070 8867 3100 8953
rect 3170 8867 3200 8953
rect 3270 8867 3300 8953
rect 3370 8867 3400 8953
rect 3470 8867 3500 8953
rect 3570 8867 3600 8953
rect 3670 8867 3700 8953
rect 3770 8867 3800 8953
rect 3870 8867 3900 8953
rect 3970 8867 4000 8953
rect 4070 8867 4100 8953
rect 4170 8867 4200 8953
rect 4270 8867 4300 8953
rect 4370 8867 4400 8953
rect 2770 8727 2800 8813
rect 2870 8727 2900 8813
rect 2970 8727 3000 8813
rect 3070 8727 3100 8813
rect 1170 8497 1200 8583
rect 1270 8497 1300 8583
rect 1370 8497 1400 8583
rect 1470 8497 1500 8583
rect 1570 8497 1600 8583
rect 1670 8497 1700 8583
rect 1770 8497 1800 8583
rect 1870 8497 1900 8583
rect 1970 8497 2000 8583
rect 2070 8497 2100 8583
rect 2170 8497 2200 8583
rect 2270 8497 2300 8583
rect 2370 8497 2400 8583
rect 2470 8497 2500 8583
rect 2570 8497 2600 8583
rect 2670 8497 2700 8583
rect 70 8357 100 8443
rect 170 8357 200 8443
rect 270 8357 300 8443
rect 370 8357 400 8443
rect 470 8357 500 8443
rect 570 8357 600 8443
rect 670 8357 700 8443
rect 770 8357 800 8443
rect 870 8357 900 8443
rect 970 8357 1000 8443
rect 1070 8357 1100 8443
rect 1170 8357 1200 8443
rect 1270 8357 1300 8443
rect 70 8217 100 8303
rect 170 8217 200 8303
rect 270 8217 300 8303
rect 370 8217 400 8303
rect 470 8217 500 8303
rect 570 8217 600 8303
rect 770 8217 800 8303
rect 1470 8357 1500 8443
rect 1570 8357 1600 8443
rect 1670 8357 1700 8443
rect 1770 8357 1800 8443
rect 1970 8357 2000 8443
rect 970 8217 1000 8303
rect 1070 8217 1100 8303
rect 1170 8217 1200 8303
rect 1270 8217 1300 8303
rect 1370 8217 1400 8303
rect 1470 8217 1500 8303
rect 1570 8217 1600 8303
rect 1670 8217 1700 8303
rect 1770 8217 1800 8303
rect 1870 8217 1900 8303
rect 70 8077 100 8163
rect 170 8077 200 8163
rect 270 8077 300 8163
rect 370 8077 400 8163
rect 470 8077 500 8163
rect 570 8077 600 8163
rect 670 8077 700 8163
rect 770 8077 800 8163
rect 870 8077 900 8163
rect 970 8077 1000 8163
rect 1070 8077 1100 8163
rect 1170 8077 1200 8163
rect 70 7937 100 8023
rect 170 7937 200 8023
rect 370 7937 400 8023
rect 470 7937 500 8023
rect 570 7937 600 8023
rect 670 7937 700 8023
rect 770 7937 800 8023
rect 870 7937 900 8023
rect 970 7937 1000 8023
rect 70 7797 100 7883
rect 170 7797 200 7883
rect 270 7797 300 7883
rect 370 7797 400 7883
rect 470 7797 500 7883
rect 570 7797 600 7883
rect 770 7797 800 7883
rect 2170 8357 2200 8443
rect 2270 8357 2300 8443
rect 2070 8217 2100 8303
rect 2170 8217 2200 8303
rect 2270 8217 2300 8303
rect 4670 9007 4700 9093
rect 4570 8867 4600 8953
rect 5170 9147 5200 9233
rect 5270 9147 5300 9233
rect 5370 9147 5400 9233
rect 4870 9007 4900 9093
rect 4970 9007 5000 9093
rect 5070 9007 5100 9093
rect 5170 9007 5200 9093
rect 4770 8867 4800 8953
rect 5570 9147 5600 9233
rect 5670 9147 5700 9233
rect 5870 9147 5900 9233
rect 5970 9147 6000 9233
rect 6070 9147 6100 9233
rect 6170 9147 6200 9233
rect 6270 9147 6300 9233
rect 6370 9147 6400 9233
rect 6570 9147 6600 9233
rect 6670 9147 6700 9233
rect 6880 9147 6910 9233
rect 6980 9147 7010 9233
rect 7080 9147 7110 9233
rect 7180 9147 7210 9233
rect 7280 9147 7310 9233
rect 7380 9147 7410 9233
rect 5370 9007 5400 9093
rect 5470 9007 5500 9093
rect 5570 9007 5600 9093
rect 5670 9007 5700 9093
rect 5770 9007 5800 9093
rect 5870 9007 5900 9093
rect 5970 9007 6000 9093
rect 6070 9007 6100 9093
rect 6170 9007 6200 9093
rect 6270 9007 6300 9093
rect 6370 9007 6400 9093
rect 6570 9007 6600 9093
rect 6670 9007 6700 9093
rect 6880 9007 6910 9093
rect 6980 9007 7010 9093
rect 7080 9007 7110 9093
rect 7180 9007 7210 9093
rect 7280 9007 7310 9093
rect 7380 9007 7410 9093
rect 4970 8867 5000 8953
rect 5070 8867 5100 8953
rect 5170 8867 5200 8953
rect 5270 8867 5300 8953
rect 5370 8867 5400 8953
rect 5470 8867 5500 8953
rect 5570 8867 5600 8953
rect 3270 8727 3300 8813
rect 3370 8727 3400 8813
rect 3470 8727 3500 8813
rect 3570 8727 3600 8813
rect 3670 8727 3700 8813
rect 3770 8727 3800 8813
rect 3870 8727 3900 8813
rect 3970 8727 4000 8813
rect 4070 8727 4100 8813
rect 4170 8727 4200 8813
rect 4270 8727 4300 8813
rect 4370 8727 4400 8813
rect 4470 8727 4500 8813
rect 4570 8727 4600 8813
rect 4670 8727 4700 8813
rect 4770 8727 4800 8813
rect 4870 8727 4900 8813
rect 4970 8727 5000 8813
rect 5070 8727 5100 8813
rect 5170 8727 5200 8813
rect 5270 8727 5300 8813
rect 5370 8727 5400 8813
rect 5470 8727 5500 8813
rect 2870 8497 2900 8583
rect 2970 8497 3000 8583
rect 3070 8497 3100 8583
rect 3170 8497 3200 8583
rect 3270 8497 3300 8583
rect 3470 8497 3500 8583
rect 3670 8497 3700 8583
rect 3770 8497 3800 8583
rect 3870 8497 3900 8583
rect 3970 8497 4000 8583
rect 2470 8357 2500 8443
rect 2570 8357 2600 8443
rect 2670 8357 2700 8443
rect 2770 8357 2800 8443
rect 2870 8357 2900 8443
rect 2970 8357 3000 8443
rect 3070 8357 3100 8443
rect 3170 8357 3200 8443
rect 3270 8357 3300 8443
rect 3370 8357 3400 8443
rect 3470 8357 3500 8443
rect 3570 8357 3600 8443
rect 3670 8357 3700 8443
rect 3770 8357 3800 8443
rect 2470 8217 2500 8303
rect 2670 8217 2700 8303
rect 2770 8217 2800 8303
rect 2870 8217 2900 8303
rect 2970 8217 3000 8303
rect 3070 8217 3100 8303
rect 1370 8077 1400 8163
rect 1470 8077 1500 8163
rect 1570 8077 1600 8163
rect 1670 8077 1700 8163
rect 1770 8077 1800 8163
rect 1870 8077 1900 8163
rect 1970 8077 2000 8163
rect 2070 8077 2100 8163
rect 2170 8077 2200 8163
rect 2270 8077 2300 8163
rect 2370 8077 2400 8163
rect 2470 8077 2500 8163
rect 2570 8077 2600 8163
rect 1170 7937 1200 8023
rect 1270 7937 1300 8023
rect 1470 7937 1500 8023
rect 1570 7937 1600 8023
rect 1670 7937 1700 8023
rect 970 7797 1000 7883
rect 1070 7797 1100 7883
rect 1170 7797 1200 7883
rect 1270 7797 1300 7883
rect 1370 7797 1400 7883
rect 1570 7797 1600 7883
rect 70 7657 100 7743
rect 170 7657 200 7743
rect 270 7657 300 7743
rect 370 7657 400 7743
rect 470 7657 500 7743
rect 570 7657 600 7743
rect 670 7657 700 7743
rect 770 7657 800 7743
rect 870 7657 900 7743
rect 970 7657 1000 7743
rect 1070 7657 1100 7743
rect 1170 7657 1200 7743
rect 1270 7657 1300 7743
rect 1370 7657 1400 7743
rect 1470 7657 1500 7743
rect 70 7517 100 7603
rect 170 7517 200 7603
rect 270 7517 300 7603
rect 370 7517 400 7603
rect 470 7517 500 7603
rect 570 7517 600 7603
rect 670 7517 700 7603
rect 770 7517 800 7603
rect 870 7517 900 7603
rect 970 7517 1000 7603
rect 1170 7517 1200 7603
rect 1270 7517 1300 7603
rect 1870 7937 1900 8023
rect 1970 7937 2000 8023
rect 2770 8077 2800 8163
rect 2170 7937 2200 8023
rect 2270 7937 2300 8023
rect 2370 7937 2400 8023
rect 2470 7937 2500 8023
rect 2570 7937 2600 8023
rect 2670 7937 2700 8023
rect 1770 7797 1800 7883
rect 1870 7797 1900 7883
rect 1970 7797 2000 7883
rect 2070 7797 2100 7883
rect 2170 7797 2200 7883
rect 2270 7797 2300 7883
rect 2370 7797 2400 7883
rect 2470 7797 2500 7883
rect 1670 7657 1700 7743
rect 3270 8217 3300 8303
rect 3370 8217 3400 8303
rect 3470 8217 3500 8303
rect 4170 8497 4200 8583
rect 4270 8497 4300 8583
rect 4470 8497 4500 8583
rect 4570 8497 4600 8583
rect 4670 8497 4700 8583
rect 3970 8357 4000 8443
rect 4070 8357 4100 8443
rect 4170 8357 4200 8443
rect 4270 8357 4300 8443
rect 4370 8357 4400 8443
rect 4470 8357 4500 8443
rect 4570 8357 4600 8443
rect 4670 8357 4700 8443
rect 5770 8867 5800 8953
rect 5870 8867 5900 8953
rect 5970 8867 6000 8953
rect 6070 8867 6100 8953
rect 5670 8727 5700 8813
rect 5770 8727 5800 8813
rect 5870 8727 5900 8813
rect 4870 8497 4900 8583
rect 4970 8497 5000 8583
rect 5070 8497 5100 8583
rect 5170 8497 5200 8583
rect 5270 8497 5300 8583
rect 5370 8497 5400 8583
rect 5470 8497 5500 8583
rect 5570 8497 5600 8583
rect 4870 8357 4900 8443
rect 6270 8867 6300 8953
rect 6370 8867 6400 8953
rect 6570 8867 6600 8953
rect 6670 8867 6700 8953
rect 6880 8867 6910 8953
rect 6980 8867 7010 8953
rect 7080 8867 7110 8953
rect 7180 8867 7210 8953
rect 7280 8867 7310 8953
rect 7380 8867 7410 8953
rect 6070 8727 6100 8813
rect 6170 8727 6200 8813
rect 6270 8727 6300 8813
rect 6370 8727 6400 8813
rect 6570 8727 6600 8813
rect 6670 8727 6700 8813
rect 6880 8727 6910 8813
rect 6980 8727 7010 8813
rect 7080 8727 7110 8813
rect 7180 8727 7210 8813
rect 7280 8727 7310 8813
rect 7380 8727 7410 8813
rect 5770 8497 5800 8583
rect 5870 8497 5900 8583
rect 5970 8497 6000 8583
rect 6070 8497 6100 8583
rect 6170 8497 6200 8583
rect 6270 8497 6300 8583
rect 6370 8497 6400 8583
rect 6570 8497 6600 8583
rect 6670 8497 6700 8583
rect 6880 8497 6910 8583
rect 6980 8497 7010 8583
rect 7080 8497 7110 8583
rect 7180 8497 7210 8583
rect 7280 8497 7310 8583
rect 7380 8497 7410 8583
rect 5070 8357 5100 8443
rect 5170 8357 5200 8443
rect 5270 8357 5300 8443
rect 5370 8357 5400 8443
rect 5470 8357 5500 8443
rect 5570 8357 5600 8443
rect 5670 8357 5700 8443
rect 5770 8357 5800 8443
rect 5970 8357 6000 8443
rect 6070 8357 6100 8443
rect 6170 8357 6200 8443
rect 6270 8357 6300 8443
rect 6370 8357 6400 8443
rect 6570 8357 6600 8443
rect 6670 8357 6700 8443
rect 6880 8357 6910 8443
rect 6980 8357 7010 8443
rect 7080 8357 7110 8443
rect 7180 8357 7210 8443
rect 7280 8357 7310 8443
rect 7380 8357 7410 8443
rect 3670 8217 3700 8303
rect 3770 8217 3800 8303
rect 3870 8217 3900 8303
rect 3970 8217 4000 8303
rect 4070 8217 4100 8303
rect 4170 8217 4200 8303
rect 4270 8217 4300 8303
rect 4370 8217 4400 8303
rect 4470 8217 4500 8303
rect 4570 8217 4600 8303
rect 4670 8217 4700 8303
rect 4770 8217 4800 8303
rect 4870 8217 4900 8303
rect 4970 8217 5000 8303
rect 5070 8217 5100 8303
rect 5170 8217 5200 8303
rect 5270 8217 5300 8303
rect 5370 8217 5400 8303
rect 5470 8217 5500 8303
rect 5570 8217 5600 8303
rect 5670 8217 5700 8303
rect 5770 8217 5800 8303
rect 5870 8217 5900 8303
rect 5970 8217 6000 8303
rect 6070 8217 6100 8303
rect 6170 8217 6200 8303
rect 6270 8217 6300 8303
rect 6370 8217 6400 8303
rect 6570 8217 6600 8303
rect 6670 8217 6700 8303
rect 6880 8217 6910 8303
rect 6980 8217 7010 8303
rect 7080 8217 7110 8303
rect 7180 8217 7210 8303
rect 7280 8217 7310 8303
rect 7380 8217 7410 8303
rect 2970 8077 3000 8163
rect 3070 8077 3100 8163
rect 3170 8077 3200 8163
rect 3270 8077 3300 8163
rect 3370 8077 3400 8163
rect 3470 8077 3500 8163
rect 3570 8077 3600 8163
rect 3670 8077 3700 8163
rect 2870 7937 2900 8023
rect 3870 8077 3900 8163
rect 3970 8077 4000 8163
rect 4070 8077 4100 8163
rect 4170 8077 4200 8163
rect 4270 8077 4300 8163
rect 4370 8077 4400 8163
rect 4470 8077 4500 8163
rect 4570 8077 4600 8163
rect 4670 8077 4700 8163
rect 4770 8077 4800 8163
rect 4870 8077 4900 8163
rect 4970 8077 5000 8163
rect 5070 8077 5100 8163
rect 5170 8077 5200 8163
rect 5270 8077 5300 8163
rect 5370 8077 5400 8163
rect 5470 8077 5500 8163
rect 5570 8077 5600 8163
rect 5670 8077 5700 8163
rect 5770 8077 5800 8163
rect 5870 8077 5900 8163
rect 5970 8077 6000 8163
rect 6070 8077 6100 8163
rect 6170 8077 6200 8163
rect 6270 8077 6300 8163
rect 6370 8077 6400 8163
rect 6570 8077 6600 8163
rect 6670 8077 6700 8163
rect 6880 8077 6910 8163
rect 6980 8077 7010 8163
rect 7080 8077 7110 8163
rect 7180 8077 7210 8163
rect 7280 8077 7310 8163
rect 7380 8077 7410 8163
rect 3070 7937 3100 8023
rect 3170 7937 3200 8023
rect 3270 7937 3300 8023
rect 3370 7937 3400 8023
rect 3470 7937 3500 8023
rect 3570 7937 3600 8023
rect 3670 7937 3700 8023
rect 3770 7937 3800 8023
rect 3870 7937 3900 8023
rect 3970 7937 4000 8023
rect 4070 7937 4100 8023
rect 4170 7937 4200 8023
rect 4270 7937 4300 8023
rect 4370 7937 4400 8023
rect 4470 7937 4500 8023
rect 4570 7937 4600 8023
rect 4670 7937 4700 8023
rect 4770 7937 4800 8023
rect 4870 7937 4900 8023
rect 2670 7797 2700 7883
rect 2770 7797 2800 7883
rect 2870 7797 2900 7883
rect 2970 7797 3000 7883
rect 3070 7797 3100 7883
rect 3170 7797 3200 7883
rect 3270 7797 3300 7883
rect 1870 7657 1900 7743
rect 1970 7657 2000 7743
rect 2070 7657 2100 7743
rect 2170 7657 2200 7743
rect 2270 7657 2300 7743
rect 2370 7657 2400 7743
rect 2470 7657 2500 7743
rect 2570 7657 2600 7743
rect 2670 7657 2700 7743
rect 1470 7517 1500 7603
rect 1570 7517 1600 7603
rect 1670 7517 1700 7603
rect 1770 7517 1800 7603
rect 1870 7517 1900 7603
rect 1970 7517 2000 7603
rect 2070 7517 2100 7603
rect 2170 7517 2200 7603
rect 2270 7517 2300 7603
rect 2370 7517 2400 7603
rect 2470 7517 2500 7603
rect 2570 7517 2600 7603
rect 2670 7517 2700 7603
rect 70 7287 100 7373
rect 170 7287 200 7373
rect 270 7287 300 7373
rect 370 7287 400 7373
rect 470 7287 500 7373
rect 570 7287 600 7373
rect 670 7287 700 7373
rect 770 7287 800 7373
rect 870 7287 900 7373
rect 970 7287 1000 7373
rect 1070 7287 1100 7373
rect 1170 7287 1200 7373
rect 70 7147 100 7233
rect 170 7147 200 7233
rect 270 7147 300 7233
rect 70 7007 100 7093
rect 170 7007 200 7093
rect 270 7007 300 7093
rect 1370 7287 1400 7373
rect 1470 7287 1500 7373
rect 1670 7287 1700 7373
rect 1770 7287 1800 7373
rect 1870 7287 1900 7373
rect 1970 7287 2000 7373
rect 2070 7287 2100 7373
rect 2270 7287 2300 7373
rect 2470 7287 2500 7373
rect 470 7147 500 7233
rect 570 7147 600 7233
rect 670 7147 700 7233
rect 770 7147 800 7233
rect 870 7147 900 7233
rect 970 7147 1000 7233
rect 1070 7147 1100 7233
rect 1170 7147 1200 7233
rect 1270 7147 1300 7233
rect 1370 7147 1400 7233
rect 1470 7147 1500 7233
rect 1570 7147 1600 7233
rect 1670 7147 1700 7233
rect 1770 7147 1800 7233
rect 1870 7147 1900 7233
rect 1970 7147 2000 7233
rect 2070 7147 2100 7233
rect 2170 7147 2200 7233
rect 2270 7147 2300 7233
rect 2370 7147 2400 7233
rect 2470 7147 2500 7233
rect 470 7007 500 7093
rect 570 7007 600 7093
rect 670 7007 700 7093
rect 770 7007 800 7093
rect 870 7007 900 7093
rect 970 7007 1000 7093
rect 1070 7007 1100 7093
rect 1170 7007 1200 7093
rect 1370 7007 1400 7093
rect 1470 7007 1500 7093
rect 1570 7007 1600 7093
rect 1670 7007 1700 7093
rect 1770 7007 1800 7093
rect 1870 7007 1900 7093
rect 1970 7007 2000 7093
rect 2070 7007 2100 7093
rect 2170 7007 2200 7093
rect 70 6867 100 6953
rect 170 6867 200 6953
rect 270 6867 300 6953
rect 370 6867 400 6953
rect 470 6867 500 6953
rect 570 6867 600 6953
rect 670 6867 700 6953
rect 770 6867 800 6953
rect 870 6867 900 6953
rect 970 6867 1000 6953
rect 1070 6867 1100 6953
rect 1170 6867 1200 6953
rect 1270 6867 1300 6953
rect 1370 6867 1400 6953
rect 70 6727 100 6813
rect 170 6727 200 6813
rect 270 6727 300 6813
rect 370 6727 400 6813
rect 470 6727 500 6813
rect 570 6727 600 6813
rect 670 6727 700 6813
rect 770 6727 800 6813
rect 870 6727 900 6813
rect 970 6727 1000 6813
rect 1070 6727 1100 6813
rect 1170 6727 1200 6813
rect 1270 6727 1300 6813
rect 70 6587 100 6673
rect 170 6587 200 6673
rect 370 6587 400 6673
rect 470 6587 500 6673
rect 570 6587 600 6673
rect 670 6587 700 6673
rect 770 6587 800 6673
rect 870 6587 900 6673
rect 970 6587 1000 6673
rect 70 6447 100 6533
rect 170 6447 200 6533
rect 270 6447 300 6533
rect 370 6447 400 6533
rect 470 6447 500 6533
rect 70 6307 100 6393
rect 1170 6587 1200 6673
rect 1570 6867 1600 6953
rect 1670 6867 1700 6953
rect 1770 6867 1800 6953
rect 1870 6867 1900 6953
rect 1970 6867 2000 6953
rect 1470 6727 1500 6813
rect 3470 7797 3500 7883
rect 3570 7797 3600 7883
rect 3670 7797 3700 7883
rect 3870 7797 3900 7883
rect 4070 7797 4100 7883
rect 2870 7657 2900 7743
rect 2970 7657 3000 7743
rect 3070 7657 3100 7743
rect 3170 7657 3200 7743
rect 3270 7657 3300 7743
rect 3370 7657 3400 7743
rect 3470 7657 3500 7743
rect 3570 7657 3600 7743
rect 3670 7657 3700 7743
rect 3770 7657 3800 7743
rect 3870 7657 3900 7743
rect 3970 7657 4000 7743
rect 4070 7657 4100 7743
rect 2870 7517 2900 7603
rect 2970 7517 3000 7603
rect 3170 7517 3200 7603
rect 3370 7517 3400 7603
rect 3470 7517 3500 7603
rect 3570 7517 3600 7603
rect 3670 7517 3700 7603
rect 3770 7517 3800 7603
rect 3870 7517 3900 7603
rect 4270 7797 4300 7883
rect 4370 7797 4400 7883
rect 4470 7797 4500 7883
rect 4270 7657 4300 7743
rect 4670 7797 4700 7883
rect 4870 7797 4900 7883
rect 5070 7937 5100 8023
rect 5170 7937 5200 8023
rect 5270 7937 5300 8023
rect 5370 7937 5400 8023
rect 5470 7937 5500 8023
rect 5570 7937 5600 8023
rect 5670 7937 5700 8023
rect 5770 7937 5800 8023
rect 5870 7937 5900 8023
rect 5970 7937 6000 8023
rect 6070 7937 6100 8023
rect 6170 7937 6200 8023
rect 6270 7937 6300 8023
rect 6370 7937 6400 8023
rect 6570 7937 6600 8023
rect 6670 7937 6700 8023
rect 6880 7937 6910 8023
rect 6980 7937 7010 8023
rect 7080 7937 7110 8023
rect 7180 7937 7210 8023
rect 7280 7937 7310 8023
rect 7380 7937 7410 8023
rect 5070 7797 5100 7883
rect 5170 7797 5200 7883
rect 5270 7797 5300 7883
rect 5370 7797 5400 7883
rect 5470 7797 5500 7883
rect 4470 7657 4500 7743
rect 4570 7657 4600 7743
rect 4670 7657 4700 7743
rect 4770 7657 4800 7743
rect 4870 7657 4900 7743
rect 4970 7657 5000 7743
rect 5070 7657 5100 7743
rect 5170 7657 5200 7743
rect 5270 7657 5300 7743
rect 5370 7657 5400 7743
rect 5470 7657 5500 7743
rect 4070 7517 4100 7603
rect 4170 7517 4200 7603
rect 4270 7517 4300 7603
rect 4370 7517 4400 7603
rect 4470 7517 4500 7603
rect 4570 7517 4600 7603
rect 4670 7517 4700 7603
rect 4770 7517 4800 7603
rect 4870 7517 4900 7603
rect 5070 7517 5100 7603
rect 5670 7797 5700 7883
rect 5670 7657 5700 7743
rect 5870 7797 5900 7883
rect 5970 7797 6000 7883
rect 6070 7797 6100 7883
rect 6170 7797 6200 7883
rect 6270 7797 6300 7883
rect 6370 7797 6400 7883
rect 6570 7797 6600 7883
rect 6670 7797 6700 7883
rect 6880 7797 6910 7883
rect 6980 7797 7010 7883
rect 7080 7797 7110 7883
rect 7180 7797 7210 7883
rect 7280 7797 7310 7883
rect 7380 7797 7410 7883
rect 5870 7657 5900 7743
rect 5970 7657 6000 7743
rect 6070 7657 6100 7743
rect 6170 7657 6200 7743
rect 6270 7657 6300 7743
rect 6370 7657 6400 7743
rect 6570 7657 6600 7743
rect 6670 7657 6700 7743
rect 6880 7657 6910 7743
rect 6980 7657 7010 7743
rect 7080 7657 7110 7743
rect 7180 7657 7210 7743
rect 7280 7657 7310 7743
rect 7380 7657 7410 7743
rect 5270 7517 5300 7603
rect 5370 7517 5400 7603
rect 5470 7517 5500 7603
rect 5570 7517 5600 7603
rect 5670 7517 5700 7603
rect 5770 7517 5800 7603
rect 5870 7517 5900 7603
rect 5970 7517 6000 7603
rect 6070 7517 6100 7603
rect 6170 7517 6200 7603
rect 6270 7517 6300 7603
rect 6370 7517 6400 7603
rect 6570 7517 6600 7603
rect 6670 7517 6700 7603
rect 6880 7517 6910 7603
rect 6980 7517 7010 7603
rect 7080 7517 7110 7603
rect 7180 7517 7210 7603
rect 7280 7517 7310 7603
rect 7380 7517 7410 7603
rect 2670 7287 2700 7373
rect 2770 7287 2800 7373
rect 2870 7287 2900 7373
rect 2970 7287 3000 7373
rect 3070 7287 3100 7373
rect 3170 7287 3200 7373
rect 3270 7287 3300 7373
rect 3370 7287 3400 7373
rect 3470 7287 3500 7373
rect 3570 7287 3600 7373
rect 3670 7287 3700 7373
rect 3770 7287 3800 7373
rect 3870 7287 3900 7373
rect 3970 7287 4000 7373
rect 4070 7287 4100 7373
rect 4170 7287 4200 7373
rect 4270 7287 4300 7373
rect 4370 7287 4400 7373
rect 4470 7287 4500 7373
rect 4570 7287 4600 7373
rect 4670 7287 4700 7373
rect 4770 7287 4800 7373
rect 4870 7287 4900 7373
rect 4970 7287 5000 7373
rect 5070 7287 5100 7373
rect 5170 7287 5200 7373
rect 5270 7287 5300 7373
rect 5370 7287 5400 7373
rect 5470 7287 5500 7373
rect 5570 7287 5600 7373
rect 5670 7287 5700 7373
rect 5770 7287 5800 7373
rect 5870 7287 5900 7373
rect 5970 7287 6000 7373
rect 6070 7287 6100 7373
rect 6170 7287 6200 7373
rect 6270 7287 6300 7373
rect 6370 7287 6400 7373
rect 6570 7287 6600 7373
rect 6670 7287 6700 7373
rect 6880 7287 6910 7373
rect 6980 7287 7010 7373
rect 7080 7287 7110 7373
rect 7180 7287 7210 7373
rect 7280 7287 7310 7373
rect 7380 7287 7410 7373
rect 2670 7147 2700 7233
rect 2770 7147 2800 7233
rect 2870 7147 2900 7233
rect 3070 7147 3100 7233
rect 3170 7147 3200 7233
rect 2370 7007 2400 7093
rect 2470 7007 2500 7093
rect 2570 7007 2600 7093
rect 2670 7007 2700 7093
rect 2770 7007 2800 7093
rect 2870 7007 2900 7093
rect 2970 7007 3000 7093
rect 2170 6867 2200 6953
rect 2270 6867 2300 6953
rect 2370 6867 2400 6953
rect 2470 6867 2500 6953
rect 2570 6867 2600 6953
rect 2670 6867 2700 6953
rect 2770 6867 2800 6953
rect 2870 6867 2900 6953
rect 1670 6727 1700 6813
rect 1770 6727 1800 6813
rect 1870 6727 1900 6813
rect 1970 6727 2000 6813
rect 2070 6727 2100 6813
rect 3370 7147 3400 7233
rect 3470 7147 3500 7233
rect 3570 7147 3600 7233
rect 3670 7147 3700 7233
rect 3770 7147 3800 7233
rect 3870 7147 3900 7233
rect 3970 7147 4000 7233
rect 4070 7147 4100 7233
rect 4170 7147 4200 7233
rect 4270 7147 4300 7233
rect 3170 7007 3200 7093
rect 3270 7007 3300 7093
rect 3370 7007 3400 7093
rect 3070 6867 3100 6953
rect 3270 6867 3300 6953
rect 3370 6867 3400 6953
rect 3570 7007 3600 7093
rect 3670 7007 3700 7093
rect 3770 7007 3800 7093
rect 3870 7007 3900 7093
rect 3970 7007 4000 7093
rect 4470 7147 4500 7233
rect 4570 7147 4600 7233
rect 4770 7147 4800 7233
rect 4870 7147 4900 7233
rect 4970 7147 5000 7233
rect 5170 7147 5200 7233
rect 5270 7147 5300 7233
rect 5370 7147 5400 7233
rect 5470 7147 5500 7233
rect 5570 7147 5600 7233
rect 5670 7147 5700 7233
rect 5770 7147 5800 7233
rect 5870 7147 5900 7233
rect 5970 7147 6000 7233
rect 4170 7007 4200 7093
rect 4270 7007 4300 7093
rect 4370 7007 4400 7093
rect 4470 7007 4500 7093
rect 4570 7007 4600 7093
rect 4670 7007 4700 7093
rect 4770 7007 4800 7093
rect 4870 7007 4900 7093
rect 4970 7007 5000 7093
rect 5070 7007 5100 7093
rect 3570 6867 3600 6953
rect 3670 6867 3700 6953
rect 3770 6867 3800 6953
rect 3870 6867 3900 6953
rect 3970 6867 4000 6953
rect 4070 6867 4100 6953
rect 4170 6867 4200 6953
rect 4370 6867 4400 6953
rect 4470 6867 4500 6953
rect 4570 6867 4600 6953
rect 4670 6867 4700 6953
rect 4770 6867 4800 6953
rect 4970 6867 5000 6953
rect 5070 6867 5100 6953
rect 6170 7147 6200 7233
rect 6270 7147 6300 7233
rect 6370 7147 6400 7233
rect 6570 7147 6600 7233
rect 6670 7147 6700 7233
rect 6880 7147 6910 7233
rect 6980 7147 7010 7233
rect 7080 7147 7110 7233
rect 7180 7147 7210 7233
rect 7280 7147 7310 7233
rect 7380 7147 7410 7233
rect 5270 7007 5300 7093
rect 5370 7007 5400 7093
rect 5470 7007 5500 7093
rect 5570 7007 5600 7093
rect 5670 7007 5700 7093
rect 5770 7007 5800 7093
rect 5870 7007 5900 7093
rect 5970 7007 6000 7093
rect 6070 7007 6100 7093
rect 5270 6867 5300 6953
rect 5470 6867 5500 6953
rect 5570 6867 5600 6953
rect 5670 6867 5700 6953
rect 5770 6867 5800 6953
rect 5870 6867 5900 6953
rect 5970 6867 6000 6953
rect 6070 6867 6100 6953
rect 2270 6727 2300 6813
rect 2370 6727 2400 6813
rect 2470 6727 2500 6813
rect 2570 6727 2600 6813
rect 2670 6727 2700 6813
rect 2770 6727 2800 6813
rect 2870 6727 2900 6813
rect 2970 6727 3000 6813
rect 3070 6727 3100 6813
rect 3170 6727 3200 6813
rect 3270 6727 3300 6813
rect 3370 6727 3400 6813
rect 3470 6727 3500 6813
rect 3570 6727 3600 6813
rect 3670 6727 3700 6813
rect 3770 6727 3800 6813
rect 3870 6727 3900 6813
rect 3970 6727 4000 6813
rect 4070 6727 4100 6813
rect 4170 6727 4200 6813
rect 4270 6727 4300 6813
rect 4370 6727 4400 6813
rect 4470 6727 4500 6813
rect 4570 6727 4600 6813
rect 4670 6727 4700 6813
rect 4770 6727 4800 6813
rect 4870 6727 4900 6813
rect 4970 6727 5000 6813
rect 5070 6727 5100 6813
rect 5170 6727 5200 6813
rect 5270 6727 5300 6813
rect 5370 6727 5400 6813
rect 1370 6587 1400 6673
rect 1470 6587 1500 6673
rect 1570 6587 1600 6673
rect 1670 6587 1700 6673
rect 1770 6587 1800 6673
rect 1870 6587 1900 6673
rect 1970 6587 2000 6673
rect 2070 6587 2100 6673
rect 2170 6587 2200 6673
rect 2270 6587 2300 6673
rect 2370 6587 2400 6673
rect 2470 6587 2500 6673
rect 2570 6587 2600 6673
rect 2670 6587 2700 6673
rect 2770 6587 2800 6673
rect 2870 6587 2900 6673
rect 2970 6587 3000 6673
rect 3070 6587 3100 6673
rect 3170 6587 3200 6673
rect 3270 6587 3300 6673
rect 3370 6587 3400 6673
rect 670 6447 700 6533
rect 770 6447 800 6533
rect 870 6447 900 6533
rect 970 6447 1000 6533
rect 1070 6447 1100 6533
rect 1170 6447 1200 6533
rect 1270 6447 1300 6533
rect 1370 6447 1400 6533
rect 1470 6447 1500 6533
rect 1570 6447 1600 6533
rect 270 6307 300 6393
rect 370 6307 400 6393
rect 470 6307 500 6393
rect 570 6307 600 6393
rect 670 6307 700 6393
rect 770 6307 800 6393
rect 970 6307 1000 6393
rect 1170 6307 1200 6393
rect 1270 6307 1300 6393
rect 1370 6307 1400 6393
rect 1470 6307 1500 6393
rect 1570 6307 1600 6393
rect 3570 6587 3600 6673
rect 3770 6587 3800 6673
rect 3870 6587 3900 6673
rect 3970 6587 4000 6673
rect 4070 6587 4100 6673
rect 4170 6587 4200 6673
rect 4270 6587 4300 6673
rect 4370 6587 4400 6673
rect 1770 6447 1800 6533
rect 1870 6447 1900 6533
rect 1970 6447 2000 6533
rect 2070 6447 2100 6533
rect 2170 6447 2200 6533
rect 2270 6447 2300 6533
rect 2370 6447 2400 6533
rect 2470 6447 2500 6533
rect 2570 6447 2600 6533
rect 2670 6447 2700 6533
rect 2770 6447 2800 6533
rect 2870 6447 2900 6533
rect 2970 6447 3000 6533
rect 3070 6447 3100 6533
rect 3170 6447 3200 6533
rect 3270 6447 3300 6533
rect 3370 6447 3400 6533
rect 3470 6447 3500 6533
rect 3570 6447 3600 6533
rect 3670 6447 3700 6533
rect 1770 6307 1800 6393
rect 1870 6307 1900 6393
rect 2070 6307 2100 6393
rect 2170 6307 2200 6393
rect 2270 6307 2300 6393
rect 2370 6307 2400 6393
rect 2470 6307 2500 6393
rect 2570 6307 2600 6393
rect 2670 6307 2700 6393
rect 2770 6307 2800 6393
rect 70 6077 100 6163
rect 170 6077 200 6163
rect 270 6077 300 6163
rect 370 6077 400 6163
rect 470 6077 500 6163
rect 570 6077 600 6163
rect 670 6077 700 6163
rect 770 6077 800 6163
rect 870 6077 900 6163
rect 970 6077 1000 6163
rect 1070 6077 1100 6163
rect 1170 6077 1200 6163
rect 1270 6077 1300 6163
rect 1370 6077 1400 6163
rect 1470 6077 1500 6163
rect 1570 6077 1600 6163
rect 1670 6077 1700 6163
rect 1770 6077 1800 6163
rect 1870 6077 1900 6163
rect 1970 6077 2000 6163
rect 2070 6077 2100 6163
rect 2170 6077 2200 6163
rect 2270 6077 2300 6163
rect 2370 6077 2400 6163
rect 70 5937 100 6023
rect 170 5937 200 6023
rect 270 5937 300 6023
rect 370 5937 400 6023
rect 570 5937 600 6023
rect 670 5937 700 6023
rect 770 5937 800 6023
rect 870 5937 900 6023
rect 970 5937 1000 6023
rect 1070 5937 1100 6023
rect 1170 5937 1200 6023
rect 1270 5937 1300 6023
rect 2970 6307 3000 6393
rect 3070 6307 3100 6393
rect 3170 6307 3200 6393
rect 3270 6307 3300 6393
rect 5570 6727 5600 6813
rect 5770 6727 5800 6813
rect 4570 6587 4600 6673
rect 4670 6587 4700 6673
rect 4770 6587 4800 6673
rect 4870 6587 4900 6673
rect 4970 6587 5000 6673
rect 5070 6587 5100 6673
rect 5170 6587 5200 6673
rect 5270 6587 5300 6673
rect 5370 6587 5400 6673
rect 5470 6587 5500 6673
rect 5570 6587 5600 6673
rect 5670 6587 5700 6673
rect 5770 6587 5800 6673
rect 3870 6447 3900 6533
rect 3970 6447 4000 6533
rect 4070 6447 4100 6533
rect 4170 6447 4200 6533
rect 4270 6447 4300 6533
rect 4370 6447 4400 6533
rect 4470 6447 4500 6533
rect 4570 6447 4600 6533
rect 4670 6447 4700 6533
rect 4770 6447 4800 6533
rect 4870 6447 4900 6533
rect 4970 6447 5000 6533
rect 5070 6447 5100 6533
rect 3470 6307 3500 6393
rect 3570 6307 3600 6393
rect 3670 6307 3700 6393
rect 3770 6307 3800 6393
rect 3870 6307 3900 6393
rect 3970 6307 4000 6393
rect 4070 6307 4100 6393
rect 4170 6307 4200 6393
rect 4270 6307 4300 6393
rect 4370 6307 4400 6393
rect 4470 6307 4500 6393
rect 4570 6307 4600 6393
rect 4670 6307 4700 6393
rect 4770 6307 4800 6393
rect 4870 6307 4900 6393
rect 4970 6307 5000 6393
rect 2570 6077 2600 6163
rect 2670 6077 2700 6163
rect 2770 6077 2800 6163
rect 2870 6077 2900 6163
rect 2970 6077 3000 6163
rect 3070 6077 3100 6163
rect 3170 6077 3200 6163
rect 3270 6077 3300 6163
rect 3370 6077 3400 6163
rect 3470 6077 3500 6163
rect 3570 6077 3600 6163
rect 3670 6077 3700 6163
rect 1470 5937 1500 6023
rect 1570 5937 1600 6023
rect 1670 5937 1700 6023
rect 1770 5937 1800 6023
rect 1870 5937 1900 6023
rect 1970 5937 2000 6023
rect 2070 5937 2100 6023
rect 2170 5937 2200 6023
rect 2270 5937 2300 6023
rect 2370 5937 2400 6023
rect 2470 5937 2500 6023
rect 2570 5937 2600 6023
rect 2670 5937 2700 6023
rect 2770 5937 2800 6023
rect 2870 5937 2900 6023
rect 2970 5937 3000 6023
rect 3070 5937 3100 6023
rect 3170 5937 3200 6023
rect 3270 5937 3300 6023
rect 70 5797 100 5883
rect 170 5797 200 5883
rect 270 5797 300 5883
rect 370 5797 400 5883
rect 470 5797 500 5883
rect 570 5797 600 5883
rect 670 5797 700 5883
rect 770 5797 800 5883
rect 870 5797 900 5883
rect 970 5797 1000 5883
rect 1070 5797 1100 5883
rect 1170 5797 1200 5883
rect 1270 5797 1300 5883
rect 1370 5797 1400 5883
rect 1470 5797 1500 5883
rect 1570 5797 1600 5883
rect 1670 5797 1700 5883
rect 1770 5797 1800 5883
rect 1870 5797 1900 5883
rect 1970 5797 2000 5883
rect 70 5657 100 5743
rect 170 5657 200 5743
rect 270 5657 300 5743
rect 470 5657 500 5743
rect 570 5657 600 5743
rect 670 5657 700 5743
rect 770 5657 800 5743
rect 870 5657 900 5743
rect 970 5657 1000 5743
rect 3870 6077 3900 6163
rect 3970 6077 4000 6163
rect 4170 6077 4200 6163
rect 4270 6077 4300 6163
rect 4370 6077 4400 6163
rect 4570 6077 4600 6163
rect 5270 6447 5300 6533
rect 5170 6307 5200 6393
rect 5270 6307 5300 6393
rect 6270 7007 6300 7093
rect 6370 7007 6400 7093
rect 6570 7007 6600 7093
rect 6670 7007 6700 7093
rect 6880 7007 6910 7093
rect 6980 7007 7010 7093
rect 7080 7007 7110 7093
rect 7180 7007 7210 7093
rect 7280 7007 7310 7093
rect 7380 7007 7410 7093
rect 6270 6867 6300 6953
rect 6370 6867 6400 6953
rect 6570 6867 6600 6953
rect 6670 6867 6700 6953
rect 6880 6867 6910 6953
rect 6980 6867 7010 6953
rect 7080 6867 7110 6953
rect 7180 6867 7210 6953
rect 7280 6867 7310 6953
rect 7380 6867 7410 6953
rect 5970 6727 6000 6813
rect 6070 6727 6100 6813
rect 6170 6727 6200 6813
rect 6270 6727 6300 6813
rect 6370 6727 6400 6813
rect 6570 6727 6600 6813
rect 6670 6727 6700 6813
rect 6880 6727 6910 6813
rect 6980 6727 7010 6813
rect 7080 6727 7110 6813
rect 7180 6727 7210 6813
rect 7280 6727 7310 6813
rect 7380 6727 7410 6813
rect 5970 6587 6000 6673
rect 6070 6587 6100 6673
rect 6170 6587 6200 6673
rect 6270 6587 6300 6673
rect 6370 6587 6400 6673
rect 6570 6587 6600 6673
rect 6670 6587 6700 6673
rect 6880 6587 6910 6673
rect 6980 6587 7010 6673
rect 7080 6587 7110 6673
rect 7180 6587 7210 6673
rect 7280 6587 7310 6673
rect 7380 6587 7410 6673
rect 5470 6447 5500 6533
rect 5570 6447 5600 6533
rect 5670 6447 5700 6533
rect 5770 6447 5800 6533
rect 5870 6447 5900 6533
rect 5970 6447 6000 6533
rect 6070 6447 6100 6533
rect 6170 6447 6200 6533
rect 6270 6447 6300 6533
rect 6370 6447 6400 6533
rect 6570 6447 6600 6533
rect 6670 6447 6700 6533
rect 6880 6447 6910 6533
rect 6980 6447 7010 6533
rect 7080 6447 7110 6533
rect 7180 6447 7210 6533
rect 7280 6447 7310 6533
rect 7380 6447 7410 6533
rect 5470 6307 5500 6393
rect 5570 6307 5600 6393
rect 5670 6307 5700 6393
rect 5770 6307 5800 6393
rect 5870 6307 5900 6393
rect 5970 6307 6000 6393
rect 6070 6307 6100 6393
rect 6270 6307 6300 6393
rect 6370 6307 6400 6393
rect 6570 6307 6600 6393
rect 6670 6307 6700 6393
rect 6880 6307 6910 6393
rect 6980 6307 7010 6393
rect 7080 6307 7110 6393
rect 7180 6307 7210 6393
rect 7280 6307 7310 6393
rect 7380 6307 7410 6393
rect 4770 6077 4800 6163
rect 4870 6077 4900 6163
rect 4970 6077 5000 6163
rect 5070 6077 5100 6163
rect 5170 6077 5200 6163
rect 5270 6077 5300 6163
rect 5370 6077 5400 6163
rect 5470 6077 5500 6163
rect 5570 6077 5600 6163
rect 5670 6077 5700 6163
rect 5770 6077 5800 6163
rect 5870 6077 5900 6163
rect 5970 6077 6000 6163
rect 3470 5937 3500 6023
rect 3570 5937 3600 6023
rect 3670 5937 3700 6023
rect 3770 5937 3800 6023
rect 3870 5937 3900 6023
rect 3970 5937 4000 6023
rect 4070 5937 4100 6023
rect 4170 5937 4200 6023
rect 4270 5937 4300 6023
rect 4370 5937 4400 6023
rect 4470 5937 4500 6023
rect 4570 5937 4600 6023
rect 4670 5937 4700 6023
rect 4770 5937 4800 6023
rect 4870 5937 4900 6023
rect 4970 5937 5000 6023
rect 5070 5937 5100 6023
rect 5170 5937 5200 6023
rect 2170 5797 2200 5883
rect 2270 5797 2300 5883
rect 2370 5797 2400 5883
rect 2470 5797 2500 5883
rect 2570 5797 2600 5883
rect 2670 5797 2700 5883
rect 2770 5797 2800 5883
rect 2870 5797 2900 5883
rect 2970 5797 3000 5883
rect 3070 5797 3100 5883
rect 3170 5797 3200 5883
rect 3270 5797 3300 5883
rect 3370 5797 3400 5883
rect 1170 5657 1200 5743
rect 1270 5657 1300 5743
rect 1370 5657 1400 5743
rect 1470 5657 1500 5743
rect 1570 5657 1600 5743
rect 1670 5657 1700 5743
rect 1770 5657 1800 5743
rect 1870 5657 1900 5743
rect 1970 5657 2000 5743
rect 2070 5657 2100 5743
rect 2170 5657 2200 5743
rect 2270 5657 2300 5743
rect 2370 5657 2400 5743
rect 2470 5657 2500 5743
rect 2570 5657 2600 5743
rect 2670 5657 2700 5743
rect 2770 5657 2800 5743
rect 70 5517 100 5603
rect 170 5517 200 5603
rect 270 5517 300 5603
rect 370 5517 400 5603
rect 470 5517 500 5603
rect 570 5517 600 5603
rect 670 5517 700 5603
rect 770 5517 800 5603
rect 870 5517 900 5603
rect 970 5517 1000 5603
rect 1070 5517 1100 5603
rect 70 5377 100 5463
rect 170 5377 200 5463
rect 270 5377 300 5463
rect 370 5377 400 5463
rect 1270 5517 1300 5603
rect 1470 5517 1500 5603
rect 1570 5517 1600 5603
rect 1670 5517 1700 5603
rect 1770 5517 1800 5603
rect 1870 5517 1900 5603
rect 570 5377 600 5463
rect 670 5377 700 5463
rect 770 5377 800 5463
rect 870 5377 900 5463
rect 970 5377 1000 5463
rect 1070 5377 1100 5463
rect 1170 5377 1200 5463
rect 1270 5377 1300 5463
rect 1370 5377 1400 5463
rect 1570 5377 1600 5463
rect 1670 5377 1700 5463
rect 2070 5517 2100 5603
rect 2170 5517 2200 5603
rect 1870 5377 1900 5463
rect 1970 5377 2000 5463
rect 2070 5377 2100 5463
rect 2170 5377 2200 5463
rect 70 5237 100 5323
rect 170 5237 200 5323
rect 270 5237 300 5323
rect 370 5237 400 5323
rect 470 5237 500 5323
rect 570 5237 600 5323
rect 670 5237 700 5323
rect 770 5237 800 5323
rect 870 5237 900 5323
rect 970 5237 1000 5323
rect 1070 5237 1100 5323
rect 1170 5237 1200 5323
rect 1270 5237 1300 5323
rect 1370 5237 1400 5323
rect 1470 5237 1500 5323
rect 1570 5237 1600 5323
rect 1670 5237 1700 5323
rect 1770 5237 1800 5323
rect 1870 5237 1900 5323
rect 1970 5237 2000 5323
rect 2070 5237 2100 5323
rect 70 5097 100 5183
rect 170 5097 200 5183
rect 270 5097 300 5183
rect 370 5097 400 5183
rect 470 5097 500 5183
rect 570 5097 600 5183
rect 670 5097 700 5183
rect 770 5097 800 5183
rect 870 5097 900 5183
rect 970 5097 1000 5183
rect 1070 5097 1100 5183
rect 1170 5097 1200 5183
rect 1270 5097 1300 5183
rect 70 4727 100 4813
rect 170 4727 200 4813
rect 370 4727 400 4813
rect 470 4727 500 4813
rect 570 4727 600 4813
rect 670 4727 700 4813
rect 770 4727 800 4813
rect 870 4727 900 4813
rect 970 4727 1000 4813
rect 1070 4727 1100 4813
rect 1470 5097 1500 5183
rect 1570 5097 1600 5183
rect 1670 5097 1700 5183
rect 1770 5097 1800 5183
rect 1870 5097 1900 5183
rect 1970 5097 2000 5183
rect 2070 5097 2100 5183
rect 2970 5657 3000 5743
rect 3170 5657 3200 5743
rect 3370 5657 3400 5743
rect 3570 5797 3600 5883
rect 3670 5797 3700 5883
rect 3770 5797 3800 5883
rect 3870 5797 3900 5883
rect 3970 5797 4000 5883
rect 4070 5797 4100 5883
rect 3570 5657 3600 5743
rect 3770 5657 3800 5743
rect 3870 5657 3900 5743
rect 3970 5657 4000 5743
rect 4070 5657 4100 5743
rect 2370 5517 2400 5603
rect 2470 5517 2500 5603
rect 2570 5517 2600 5603
rect 2670 5517 2700 5603
rect 2770 5517 2800 5603
rect 2870 5517 2900 5603
rect 2970 5517 3000 5603
rect 3070 5517 3100 5603
rect 3170 5517 3200 5603
rect 3270 5517 3300 5603
rect 3370 5517 3400 5603
rect 3470 5517 3500 5603
rect 3570 5517 3600 5603
rect 3670 5517 3700 5603
rect 3770 5517 3800 5603
rect 3870 5517 3900 5603
rect 3970 5517 4000 5603
rect 2370 5377 2400 5463
rect 2470 5377 2500 5463
rect 2570 5377 2600 5463
rect 2670 5377 2700 5463
rect 2770 5377 2800 5463
rect 2870 5377 2900 5463
rect 2970 5377 3000 5463
rect 3070 5377 3100 5463
rect 3170 5377 3200 5463
rect 3270 5377 3300 5463
rect 3370 5377 3400 5463
rect 3470 5377 3500 5463
rect 3570 5377 3600 5463
rect 3670 5377 3700 5463
rect 2270 5237 2300 5323
rect 2470 5237 2500 5323
rect 2570 5237 2600 5323
rect 2770 5237 2800 5323
rect 2870 5237 2900 5323
rect 3070 5237 3100 5323
rect 5370 5937 5400 6023
rect 5470 5937 5500 6023
rect 5570 5937 5600 6023
rect 5670 5937 5700 6023
rect 5770 5937 5800 6023
rect 4270 5797 4300 5883
rect 4370 5797 4400 5883
rect 4470 5797 4500 5883
rect 4570 5797 4600 5883
rect 4670 5797 4700 5883
rect 4770 5797 4800 5883
rect 4870 5797 4900 5883
rect 4970 5797 5000 5883
rect 5070 5797 5100 5883
rect 5170 5797 5200 5883
rect 5270 5797 5300 5883
rect 5370 5797 5400 5883
rect 5470 5797 5500 5883
rect 5570 5797 5600 5883
rect 5670 5797 5700 5883
rect 4270 5657 4300 5743
rect 4470 5657 4500 5743
rect 4670 5657 4700 5743
rect 4770 5657 4800 5743
rect 4870 5657 4900 5743
rect 4970 5657 5000 5743
rect 5070 5657 5100 5743
rect 5170 5657 5200 5743
rect 5270 5657 5300 5743
rect 5370 5657 5400 5743
rect 5470 5657 5500 5743
rect 6170 6077 6200 6163
rect 6370 6077 6400 6163
rect 6570 6077 6600 6163
rect 6670 6077 6700 6163
rect 6880 6077 6910 6163
rect 6980 6077 7010 6163
rect 7080 6077 7110 6163
rect 7180 6077 7210 6163
rect 7280 6077 7310 6163
rect 7380 6077 7410 6163
rect 5970 5937 6000 6023
rect 6070 5937 6100 6023
rect 6170 5937 6200 6023
rect 6270 5937 6300 6023
rect 6370 5937 6400 6023
rect 6570 5937 6600 6023
rect 6670 5937 6700 6023
rect 6880 5937 6910 6023
rect 6980 5937 7010 6023
rect 7080 5937 7110 6023
rect 7180 5937 7210 6023
rect 7280 5937 7310 6023
rect 7380 5937 7410 6023
rect 5870 5797 5900 5883
rect 6070 5797 6100 5883
rect 6170 5797 6200 5883
rect 6270 5797 6300 5883
rect 6370 5797 6400 5883
rect 6570 5797 6600 5883
rect 6670 5797 6700 5883
rect 6880 5797 6910 5883
rect 6980 5797 7010 5883
rect 7080 5797 7110 5883
rect 7180 5797 7210 5883
rect 7280 5797 7310 5883
rect 7380 5797 7410 5883
rect 5670 5657 5700 5743
rect 5770 5657 5800 5743
rect 5870 5657 5900 5743
rect 5970 5657 6000 5743
rect 6070 5657 6100 5743
rect 6170 5657 6200 5743
rect 6270 5657 6300 5743
rect 6370 5657 6400 5743
rect 6570 5657 6600 5743
rect 6670 5657 6700 5743
rect 6880 5657 6910 5743
rect 6980 5657 7010 5743
rect 7080 5657 7110 5743
rect 7180 5657 7210 5743
rect 7280 5657 7310 5743
rect 7380 5657 7410 5743
rect 4170 5517 4200 5603
rect 4270 5517 4300 5603
rect 4370 5517 4400 5603
rect 4470 5517 4500 5603
rect 4570 5517 4600 5603
rect 4670 5517 4700 5603
rect 4770 5517 4800 5603
rect 4870 5517 4900 5603
rect 4970 5517 5000 5603
rect 5070 5517 5100 5603
rect 5170 5517 5200 5603
rect 5270 5517 5300 5603
rect 5370 5517 5400 5603
rect 5470 5517 5500 5603
rect 5570 5517 5600 5603
rect 5670 5517 5700 5603
rect 5770 5517 5800 5603
rect 5870 5517 5900 5603
rect 5970 5517 6000 5603
rect 6070 5517 6100 5603
rect 6170 5517 6200 5603
rect 6270 5517 6300 5603
rect 6370 5517 6400 5603
rect 6570 5517 6600 5603
rect 6670 5517 6700 5603
rect 6880 5517 6910 5603
rect 6980 5517 7010 5603
rect 7080 5517 7110 5603
rect 7180 5517 7210 5603
rect 7280 5517 7310 5603
rect 7380 5517 7410 5603
rect 3870 5377 3900 5463
rect 3970 5377 4000 5463
rect 4070 5377 4100 5463
rect 4170 5377 4200 5463
rect 4270 5377 4300 5463
rect 4370 5377 4400 5463
rect 4470 5377 4500 5463
rect 4570 5377 4600 5463
rect 4670 5377 4700 5463
rect 4770 5377 4800 5463
rect 4870 5377 4900 5463
rect 4970 5377 5000 5463
rect 5070 5377 5100 5463
rect 5270 5377 5300 5463
rect 3270 5237 3300 5323
rect 3370 5237 3400 5323
rect 3470 5237 3500 5323
rect 3570 5237 3600 5323
rect 3670 5237 3700 5323
rect 3770 5237 3800 5323
rect 3870 5237 3900 5323
rect 3970 5237 4000 5323
rect 4070 5237 4100 5323
rect 4170 5237 4200 5323
rect 4270 5237 4300 5323
rect 4370 5237 4400 5323
rect 4470 5237 4500 5323
rect 4570 5237 4600 5323
rect 4670 5237 4700 5323
rect 4770 5237 4800 5323
rect 4870 5237 4900 5323
rect 4970 5237 5000 5323
rect 5070 5237 5100 5323
rect 5170 5237 5200 5323
rect 2270 5097 2300 5183
rect 2370 5097 2400 5183
rect 2470 5097 2500 5183
rect 2570 5097 2600 5183
rect 2670 5097 2700 5183
rect 2770 5097 2800 5183
rect 2870 5097 2900 5183
rect 2970 5097 3000 5183
rect 3070 5097 3100 5183
rect 3170 5097 3200 5183
rect 3270 5097 3300 5183
rect 3370 5097 3400 5183
rect 3470 5097 3500 5183
rect 3570 5097 3600 5183
rect 3670 5097 3700 5183
rect 3770 5097 3800 5183
rect 3870 5097 3900 5183
rect 3970 5097 4000 5183
rect 4070 5097 4100 5183
rect 4170 5097 4200 5183
rect 4270 5097 4300 5183
rect 1270 4727 1300 4813
rect 1370 4727 1400 4813
rect 1470 4727 1500 4813
rect 1570 4727 1600 4813
rect 1670 4727 1700 4813
rect 1770 4727 1800 4813
rect 1870 4727 1900 4813
rect 1970 4727 2000 4813
rect 2070 4727 2100 4813
rect 2170 4727 2200 4813
rect 2270 4727 2300 4813
rect 2370 4727 2400 4813
rect 2470 4727 2500 4813
rect 2570 4727 2600 4813
rect 2670 4727 2700 4813
rect 2770 4727 2800 4813
rect 70 4587 100 4673
rect 170 4587 200 4673
rect 270 4587 300 4673
rect 370 4587 400 4673
rect 470 4587 500 4673
rect 570 4587 600 4673
rect 670 4587 700 4673
rect 770 4587 800 4673
rect 870 4587 900 4673
rect 970 4587 1000 4673
rect 1070 4587 1100 4673
rect 1170 4587 1200 4673
rect 1270 4587 1300 4673
rect 1370 4587 1400 4673
rect 1470 4587 1500 4673
rect 1570 4587 1600 4673
rect 1670 4587 1700 4673
rect 1770 4587 1800 4673
rect 70 4447 100 4533
rect 270 4447 300 4533
rect 370 4447 400 4533
rect 470 4447 500 4533
rect 570 4447 600 4533
rect 670 4447 700 4533
rect 770 4447 800 4533
rect 870 4447 900 4533
rect 970 4447 1000 4533
rect 1070 4447 1100 4533
rect 1170 4447 1200 4533
rect 1270 4447 1300 4533
rect 1370 4447 1400 4533
rect 1470 4447 1500 4533
rect 1570 4447 1600 4533
rect 70 4307 100 4393
rect 170 4307 200 4393
rect 270 4307 300 4393
rect 370 4307 400 4393
rect 70 4167 100 4253
rect 270 4167 300 4253
rect 570 4307 600 4393
rect 670 4307 700 4393
rect 1970 4587 2000 4673
rect 4470 5097 4500 5183
rect 4570 5097 4600 5183
rect 4670 5097 4700 5183
rect 5470 5377 5500 5463
rect 5370 5237 5400 5323
rect 5670 5377 5700 5463
rect 5870 5377 5900 5463
rect 5970 5377 6000 5463
rect 6070 5377 6100 5463
rect 6170 5377 6200 5463
rect 6270 5377 6300 5463
rect 6370 5377 6400 5463
rect 6570 5377 6600 5463
rect 6670 5377 6700 5463
rect 6880 5377 6910 5463
rect 6980 5377 7010 5463
rect 7080 5377 7110 5463
rect 7180 5377 7210 5463
rect 7280 5377 7310 5463
rect 7380 5377 7410 5463
rect 5570 5237 5600 5323
rect 5670 5237 5700 5323
rect 5770 5237 5800 5323
rect 5870 5237 5900 5323
rect 5970 5237 6000 5323
rect 6070 5237 6100 5323
rect 6170 5237 6200 5323
rect 6270 5237 6300 5323
rect 6370 5237 6400 5323
rect 6570 5237 6600 5323
rect 6670 5237 6700 5323
rect 6880 5237 6910 5323
rect 6980 5237 7010 5323
rect 7080 5237 7110 5323
rect 7180 5237 7210 5323
rect 7280 5237 7310 5323
rect 7380 5237 7410 5323
rect 4870 5097 4900 5183
rect 4970 5097 5000 5183
rect 5070 5097 5100 5183
rect 5170 5097 5200 5183
rect 5270 5097 5300 5183
rect 5370 5097 5400 5183
rect 5470 5097 5500 5183
rect 5570 5097 5600 5183
rect 5670 5097 5700 5183
rect 2970 4727 3000 4813
rect 3070 4727 3100 4813
rect 3170 4727 3200 4813
rect 3270 4727 3300 4813
rect 3370 4727 3400 4813
rect 3470 4727 3500 4813
rect 3570 4727 3600 4813
rect 3670 4727 3700 4813
rect 3770 4727 3800 4813
rect 3870 4727 3900 4813
rect 3970 4727 4000 4813
rect 4070 4727 4100 4813
rect 4170 4727 4200 4813
rect 4270 4727 4300 4813
rect 4370 4727 4400 4813
rect 4470 4727 4500 4813
rect 4570 4727 4600 4813
rect 2170 4587 2200 4673
rect 2270 4587 2300 4673
rect 2370 4587 2400 4673
rect 2470 4587 2500 4673
rect 2570 4587 2600 4673
rect 2670 4587 2700 4673
rect 2770 4587 2800 4673
rect 2870 4587 2900 4673
rect 2970 4587 3000 4673
rect 3070 4587 3100 4673
rect 3170 4587 3200 4673
rect 1770 4447 1800 4533
rect 1870 4447 1900 4533
rect 1970 4447 2000 4533
rect 2070 4447 2100 4533
rect 2170 4447 2200 4533
rect 2270 4447 2300 4533
rect 2370 4447 2400 4533
rect 870 4307 900 4393
rect 970 4307 1000 4393
rect 1070 4307 1100 4393
rect 1170 4307 1200 4393
rect 1270 4307 1300 4393
rect 1370 4307 1400 4393
rect 1470 4307 1500 4393
rect 1570 4307 1600 4393
rect 1670 4307 1700 4393
rect 1770 4307 1800 4393
rect 1870 4307 1900 4393
rect 1970 4307 2000 4393
rect 2070 4307 2100 4393
rect 2170 4307 2200 4393
rect 2270 4307 2300 4393
rect 2370 4307 2400 4393
rect 470 4167 500 4253
rect 570 4167 600 4253
rect 670 4167 700 4253
rect 770 4167 800 4253
rect 870 4167 900 4253
rect 970 4167 1000 4253
rect 1070 4167 1100 4253
rect 1170 4167 1200 4253
rect 1270 4167 1300 4253
rect 1370 4167 1400 4253
rect 70 4027 100 4113
rect 170 4027 200 4113
rect 270 4027 300 4113
rect 370 4027 400 4113
rect 570 4027 600 4113
rect 70 3887 100 3973
rect 170 3887 200 3973
rect 270 3887 300 3973
rect 370 3887 400 3973
rect 470 3887 500 3973
rect 3370 4587 3400 4673
rect 3470 4587 3500 4673
rect 3570 4587 3600 4673
rect 3670 4587 3700 4673
rect 3770 4587 3800 4673
rect 3870 4587 3900 4673
rect 3970 4587 4000 4673
rect 4070 4587 4100 4673
rect 4170 4587 4200 4673
rect 4270 4587 4300 4673
rect 4370 4587 4400 4673
rect 4470 4587 4500 4673
rect 2570 4447 2600 4533
rect 2670 4447 2700 4533
rect 2770 4447 2800 4533
rect 2870 4447 2900 4533
rect 2970 4447 3000 4533
rect 3070 4447 3100 4533
rect 3170 4447 3200 4533
rect 3270 4447 3300 4533
rect 2570 4307 2600 4393
rect 2670 4307 2700 4393
rect 2770 4307 2800 4393
rect 2970 4307 3000 4393
rect 3070 4307 3100 4393
rect 3170 4307 3200 4393
rect 3470 4447 3500 4533
rect 3570 4447 3600 4533
rect 3670 4447 3700 4533
rect 3770 4447 3800 4533
rect 3870 4447 3900 4533
rect 3970 4447 4000 4533
rect 4070 4447 4100 4533
rect 4170 4447 4200 4533
rect 4270 4447 4300 4533
rect 4770 4727 4800 4813
rect 4870 4727 4900 4813
rect 4970 4727 5000 4813
rect 5070 4727 5100 4813
rect 5170 4727 5200 4813
rect 5270 4727 5300 4813
rect 5370 4727 5400 4813
rect 5870 5097 5900 5183
rect 5970 5097 6000 5183
rect 6070 5097 6100 5183
rect 6170 5097 6200 5183
rect 6270 5097 6300 5183
rect 6370 5097 6400 5183
rect 6570 5097 6600 5183
rect 6670 5097 6700 5183
rect 6880 5097 6910 5183
rect 6980 5097 7010 5183
rect 7080 5097 7110 5183
rect 7180 5097 7210 5183
rect 7280 5097 7310 5183
rect 7380 5097 7410 5183
rect 5570 4727 5600 4813
rect 5670 4727 5700 4813
rect 5770 4727 5800 4813
rect 5870 4727 5900 4813
rect 6070 4727 6100 4813
rect 4670 4587 4700 4673
rect 4770 4587 4800 4673
rect 4870 4587 4900 4673
rect 4970 4587 5000 4673
rect 5070 4587 5100 4673
rect 5170 4587 5200 4673
rect 5270 4587 5300 4673
rect 5370 4587 5400 4673
rect 5470 4587 5500 4673
rect 5570 4587 5600 4673
rect 5670 4587 5700 4673
rect 5770 4587 5800 4673
rect 5870 4587 5900 4673
rect 5970 4587 6000 4673
rect 4470 4447 4500 4533
rect 4570 4447 4600 4533
rect 4670 4447 4700 4533
rect 4770 4447 4800 4533
rect 4870 4447 4900 4533
rect 4970 4447 5000 4533
rect 5070 4447 5100 4533
rect 5170 4447 5200 4533
rect 3370 4307 3400 4393
rect 3470 4307 3500 4393
rect 3570 4307 3600 4393
rect 3670 4307 3700 4393
rect 3770 4307 3800 4393
rect 3870 4307 3900 4393
rect 3970 4307 4000 4393
rect 4070 4307 4100 4393
rect 4170 4307 4200 4393
rect 4270 4307 4300 4393
rect 4370 4307 4400 4393
rect 4470 4307 4500 4393
rect 4570 4307 4600 4393
rect 4670 4307 4700 4393
rect 4770 4307 4800 4393
rect 4870 4307 4900 4393
rect 4970 4307 5000 4393
rect 1570 4167 1600 4253
rect 1670 4167 1700 4253
rect 1770 4167 1800 4253
rect 1870 4167 1900 4253
rect 1970 4167 2000 4253
rect 2070 4167 2100 4253
rect 2170 4167 2200 4253
rect 2270 4167 2300 4253
rect 2370 4167 2400 4253
rect 2470 4167 2500 4253
rect 2570 4167 2600 4253
rect 2670 4167 2700 4253
rect 2770 4167 2800 4253
rect 2870 4167 2900 4253
rect 2970 4167 3000 4253
rect 3070 4167 3100 4253
rect 3170 4167 3200 4253
rect 3270 4167 3300 4253
rect 3370 4167 3400 4253
rect 770 4027 800 4113
rect 870 4027 900 4113
rect 970 4027 1000 4113
rect 1070 4027 1100 4113
rect 1170 4027 1200 4113
rect 1270 4027 1300 4113
rect 1370 4027 1400 4113
rect 1470 4027 1500 4113
rect 1670 4027 1700 4113
rect 1870 4027 1900 4113
rect 2070 4027 2100 4113
rect 2170 4027 2200 4113
rect 670 3887 700 3973
rect 770 3887 800 3973
rect 870 3887 900 3973
rect 970 3887 1000 3973
rect 1070 3887 1100 3973
rect 1170 3887 1200 3973
rect 1270 3887 1300 3973
rect 1370 3887 1400 3973
rect 1470 3887 1500 3973
rect 1570 3887 1600 3973
rect 1670 3887 1700 3973
rect 1770 3887 1800 3973
rect 1870 3887 1900 3973
rect 1970 3887 2000 3973
rect 2070 3887 2100 3973
rect 70 3747 100 3833
rect 170 3747 200 3833
rect 270 3747 300 3833
rect 370 3747 400 3833
rect 470 3747 500 3833
rect 570 3747 600 3833
rect 670 3747 700 3833
rect 770 3747 800 3833
rect 870 3747 900 3833
rect 970 3747 1000 3833
rect 1070 3747 1100 3833
rect 1170 3747 1200 3833
rect 70 3517 100 3603
rect 170 3517 200 3603
rect 1370 3747 1400 3833
rect 370 3517 400 3603
rect 470 3517 500 3603
rect 570 3517 600 3603
rect 670 3517 700 3603
rect 770 3517 800 3603
rect 870 3517 900 3603
rect 970 3517 1000 3603
rect 1070 3517 1100 3603
rect 1170 3517 1200 3603
rect 1270 3517 1300 3603
rect 70 3377 100 3463
rect 170 3377 200 3463
rect 270 3377 300 3463
rect 370 3377 400 3463
rect 470 3377 500 3463
rect 670 3377 700 3463
rect 1570 3747 1600 3833
rect 1670 3747 1700 3833
rect 1470 3517 1500 3603
rect 2370 4027 2400 4113
rect 2570 4027 2600 4113
rect 2670 4027 2700 4113
rect 2770 4027 2800 4113
rect 2870 4027 2900 4113
rect 2970 4027 3000 4113
rect 3070 4027 3100 4113
rect 3170 4027 3200 4113
rect 2270 3887 2300 3973
rect 2370 3887 2400 3973
rect 2470 3887 2500 3973
rect 2570 3887 2600 3973
rect 2670 3887 2700 3973
rect 2770 3887 2800 3973
rect 2870 3887 2900 3973
rect 2970 3887 3000 3973
rect 3070 3887 3100 3973
rect 3170 3887 3200 3973
rect 3370 4027 3400 4113
rect 3570 4167 3600 4253
rect 3770 4167 3800 4253
rect 3870 4167 3900 4253
rect 3970 4167 4000 4253
rect 4070 4167 4100 4253
rect 4170 4167 4200 4253
rect 4270 4167 4300 4253
rect 4370 4167 4400 4253
rect 4570 4167 4600 4253
rect 4670 4167 4700 4253
rect 4770 4167 4800 4253
rect 4870 4167 4900 4253
rect 4970 4167 5000 4253
rect 3570 4027 3600 4113
rect 3670 4027 3700 4113
rect 3770 4027 3800 4113
rect 3870 4027 3900 4113
rect 3970 4027 4000 4113
rect 4070 4027 4100 4113
rect 4170 4027 4200 4113
rect 4270 4027 4300 4113
rect 4370 4027 4400 4113
rect 4470 4027 4500 4113
rect 4570 4027 4600 4113
rect 4670 4027 4700 4113
rect 3370 3887 3400 3973
rect 3470 3887 3500 3973
rect 3570 3887 3600 3973
rect 3670 3887 3700 3973
rect 3770 3887 3800 3973
rect 3870 3887 3900 3973
rect 3970 3887 4000 3973
rect 4070 3887 4100 3973
rect 1870 3747 1900 3833
rect 1970 3747 2000 3833
rect 2070 3747 2100 3833
rect 2170 3747 2200 3833
rect 2270 3747 2300 3833
rect 2370 3747 2400 3833
rect 2470 3747 2500 3833
rect 2570 3747 2600 3833
rect 2670 3747 2700 3833
rect 2770 3747 2800 3833
rect 2870 3747 2900 3833
rect 2970 3747 3000 3833
rect 3070 3747 3100 3833
rect 3170 3747 3200 3833
rect 3270 3747 3300 3833
rect 3370 3747 3400 3833
rect 1670 3517 1700 3603
rect 1770 3517 1800 3603
rect 1870 3517 1900 3603
rect 1970 3517 2000 3603
rect 2070 3517 2100 3603
rect 2170 3517 2200 3603
rect 870 3377 900 3463
rect 970 3377 1000 3463
rect 1070 3377 1100 3463
rect 1170 3377 1200 3463
rect 1270 3377 1300 3463
rect 1370 3377 1400 3463
rect 1470 3377 1500 3463
rect 1570 3377 1600 3463
rect 1670 3377 1700 3463
rect 1770 3377 1800 3463
rect 1870 3377 1900 3463
rect 70 3237 100 3323
rect 170 3237 200 3323
rect 270 3237 300 3323
rect 370 3237 400 3323
rect 470 3237 500 3323
rect 570 3237 600 3323
rect 670 3237 700 3323
rect 770 3237 800 3323
rect 870 3237 900 3323
rect 970 3237 1000 3323
rect 1070 3237 1100 3323
rect 1170 3237 1200 3323
rect 70 3097 100 3183
rect 170 3097 200 3183
rect 270 3097 300 3183
rect 370 3097 400 3183
rect 570 3097 600 3183
rect 670 3097 700 3183
rect 770 3097 800 3183
rect 870 3097 900 3183
rect 970 3097 1000 3183
rect 1070 3097 1100 3183
rect 4270 3887 4300 3973
rect 4370 3887 4400 3973
rect 4470 3887 4500 3973
rect 5370 4447 5400 4533
rect 5470 4447 5500 4533
rect 5570 4447 5600 4533
rect 5670 4447 5700 4533
rect 5170 4307 5200 4393
rect 5270 4307 5300 4393
rect 5370 4307 5400 4393
rect 5170 4167 5200 4253
rect 5270 4167 5300 4253
rect 5370 4167 5400 4253
rect 6270 4727 6300 4813
rect 6370 4727 6400 4813
rect 6570 4727 6600 4813
rect 6670 4727 6700 4813
rect 6880 4727 6910 4813
rect 6980 4727 7010 4813
rect 7080 4727 7110 4813
rect 7180 4727 7210 4813
rect 7280 4727 7310 4813
rect 7380 4727 7410 4813
rect 6170 4587 6200 4673
rect 5870 4447 5900 4533
rect 5970 4447 6000 4533
rect 6070 4447 6100 4533
rect 6170 4447 6200 4533
rect 5570 4307 5600 4393
rect 5670 4307 5700 4393
rect 5770 4307 5800 4393
rect 5870 4307 5900 4393
rect 5970 4307 6000 4393
rect 5570 4167 5600 4253
rect 5670 4167 5700 4253
rect 5770 4167 5800 4253
rect 4870 4027 4900 4113
rect 4970 4027 5000 4113
rect 5070 4027 5100 4113
rect 5170 4027 5200 4113
rect 5270 4027 5300 4113
rect 5370 4027 5400 4113
rect 5470 4027 5500 4113
rect 5570 4027 5600 4113
rect 6170 4307 6200 4393
rect 6370 4587 6400 4673
rect 6570 4587 6600 4673
rect 6670 4587 6700 4673
rect 6880 4587 6910 4673
rect 6980 4587 7010 4673
rect 7080 4587 7110 4673
rect 7180 4587 7210 4673
rect 7280 4587 7310 4673
rect 7380 4587 7410 4673
rect 6370 4447 6400 4533
rect 6570 4447 6600 4533
rect 6670 4447 6700 4533
rect 6880 4447 6910 4533
rect 6980 4447 7010 4533
rect 7080 4447 7110 4533
rect 7180 4447 7210 4533
rect 7280 4447 7310 4533
rect 7380 4447 7410 4533
rect 6370 4307 6400 4393
rect 6570 4307 6600 4393
rect 6670 4307 6700 4393
rect 6880 4307 6910 4393
rect 6980 4307 7010 4393
rect 7080 4307 7110 4393
rect 7180 4307 7210 4393
rect 7280 4307 7310 4393
rect 7380 4307 7410 4393
rect 5970 4167 6000 4253
rect 6070 4167 6100 4253
rect 6170 4167 6200 4253
rect 6270 4167 6300 4253
rect 6370 4167 6400 4253
rect 6570 4167 6600 4253
rect 6670 4167 6700 4253
rect 6880 4167 6910 4253
rect 6980 4167 7010 4253
rect 7080 4167 7110 4253
rect 7180 4167 7210 4253
rect 7280 4167 7310 4253
rect 7380 4167 7410 4253
rect 5770 4027 5800 4113
rect 5870 4027 5900 4113
rect 5970 4027 6000 4113
rect 6070 4027 6100 4113
rect 6170 4027 6200 4113
rect 6270 4027 6300 4113
rect 6370 4027 6400 4113
rect 6570 4027 6600 4113
rect 6670 4027 6700 4113
rect 6880 4027 6910 4113
rect 6980 4027 7010 4113
rect 7080 4027 7110 4113
rect 7180 4027 7210 4113
rect 7280 4027 7310 4113
rect 7380 4027 7410 4113
rect 4670 3887 4700 3973
rect 4770 3887 4800 3973
rect 4870 3887 4900 3973
rect 4970 3887 5000 3973
rect 5070 3887 5100 3973
rect 5170 3887 5200 3973
rect 5270 3887 5300 3973
rect 5370 3887 5400 3973
rect 5470 3887 5500 3973
rect 5570 3887 5600 3973
rect 5670 3887 5700 3973
rect 5770 3887 5800 3973
rect 5870 3887 5900 3973
rect 5970 3887 6000 3973
rect 3570 3747 3600 3833
rect 3670 3747 3700 3833
rect 3770 3747 3800 3833
rect 3870 3747 3900 3833
rect 3970 3747 4000 3833
rect 4070 3747 4100 3833
rect 4170 3747 4200 3833
rect 4270 3747 4300 3833
rect 4370 3747 4400 3833
rect 4470 3747 4500 3833
rect 4570 3747 4600 3833
rect 4670 3747 4700 3833
rect 2370 3517 2400 3603
rect 2470 3517 2500 3603
rect 2570 3517 2600 3603
rect 2670 3517 2700 3603
rect 2770 3517 2800 3603
rect 2870 3517 2900 3603
rect 2970 3517 3000 3603
rect 3070 3517 3100 3603
rect 3170 3517 3200 3603
rect 3270 3517 3300 3603
rect 3370 3517 3400 3603
rect 3470 3517 3500 3603
rect 2070 3377 2100 3463
rect 2170 3377 2200 3463
rect 2270 3377 2300 3463
rect 2370 3377 2400 3463
rect 2470 3377 2500 3463
rect 2570 3377 2600 3463
rect 2670 3377 2700 3463
rect 2770 3377 2800 3463
rect 1370 3237 1400 3323
rect 1470 3237 1500 3323
rect 1570 3237 1600 3323
rect 1670 3237 1700 3323
rect 1770 3237 1800 3323
rect 1870 3237 1900 3323
rect 1970 3237 2000 3323
rect 2070 3237 2100 3323
rect 2170 3237 2200 3323
rect 2270 3237 2300 3323
rect 2370 3237 2400 3323
rect 2470 3237 2500 3323
rect 2570 3237 2600 3323
rect 2670 3237 2700 3323
rect 1270 3097 1300 3183
rect 1370 3097 1400 3183
rect 1470 3097 1500 3183
rect 1570 3097 1600 3183
rect 1670 3097 1700 3183
rect 1770 3097 1800 3183
rect 1870 3097 1900 3183
rect 1970 3097 2000 3183
rect 2070 3097 2100 3183
rect 2170 3097 2200 3183
rect 2270 3097 2300 3183
rect 2370 3097 2400 3183
rect 3670 3517 3700 3603
rect 3870 3517 3900 3603
rect 3970 3517 4000 3603
rect 4070 3517 4100 3603
rect 4170 3517 4200 3603
rect 4870 3747 4900 3833
rect 4970 3747 5000 3833
rect 5070 3747 5100 3833
rect 5170 3747 5200 3833
rect 5270 3747 5300 3833
rect 5370 3747 5400 3833
rect 5470 3747 5500 3833
rect 5570 3747 5600 3833
rect 4370 3517 4400 3603
rect 4470 3517 4500 3603
rect 4570 3517 4600 3603
rect 4670 3517 4700 3603
rect 4870 3517 4900 3603
rect 4970 3517 5000 3603
rect 5070 3517 5100 3603
rect 5170 3517 5200 3603
rect 6170 3887 6200 3973
rect 6270 3887 6300 3973
rect 6370 3887 6400 3973
rect 6570 3887 6600 3973
rect 6670 3887 6700 3973
rect 6880 3887 6910 3973
rect 6980 3887 7010 3973
rect 7080 3887 7110 3973
rect 7180 3887 7210 3973
rect 7280 3887 7310 3973
rect 7380 3887 7410 3973
rect 5770 3747 5800 3833
rect 5870 3747 5900 3833
rect 5970 3747 6000 3833
rect 6070 3747 6100 3833
rect 6170 3747 6200 3833
rect 6270 3747 6300 3833
rect 6370 3747 6400 3833
rect 6570 3747 6600 3833
rect 6670 3747 6700 3833
rect 6880 3747 6910 3833
rect 6980 3747 7010 3833
rect 7080 3747 7110 3833
rect 7180 3747 7210 3833
rect 7280 3747 7310 3833
rect 7380 3747 7410 3833
rect 5370 3517 5400 3603
rect 5470 3517 5500 3603
rect 5570 3517 5600 3603
rect 5670 3517 5700 3603
rect 5770 3517 5800 3603
rect 5870 3517 5900 3603
rect 5970 3517 6000 3603
rect 6070 3517 6100 3603
rect 6170 3517 6200 3603
rect 6270 3517 6300 3603
rect 6370 3517 6400 3603
rect 6570 3517 6600 3603
rect 6670 3517 6700 3603
rect 6880 3517 6910 3603
rect 6980 3517 7010 3603
rect 7080 3517 7110 3603
rect 7180 3517 7210 3603
rect 7280 3517 7310 3603
rect 7380 3517 7410 3603
rect 2970 3377 3000 3463
rect 3070 3377 3100 3463
rect 3170 3377 3200 3463
rect 3270 3377 3300 3463
rect 3370 3377 3400 3463
rect 3470 3377 3500 3463
rect 3570 3377 3600 3463
rect 3670 3377 3700 3463
rect 3770 3377 3800 3463
rect 3870 3377 3900 3463
rect 3970 3377 4000 3463
rect 4070 3377 4100 3463
rect 4170 3377 4200 3463
rect 4270 3377 4300 3463
rect 4370 3377 4400 3463
rect 4470 3377 4500 3463
rect 4570 3377 4600 3463
rect 4670 3377 4700 3463
rect 4770 3377 4800 3463
rect 4870 3377 4900 3463
rect 4970 3377 5000 3463
rect 5070 3377 5100 3463
rect 5170 3377 5200 3463
rect 5270 3377 5300 3463
rect 5370 3377 5400 3463
rect 5470 3377 5500 3463
rect 5570 3377 5600 3463
rect 5670 3377 5700 3463
rect 5770 3377 5800 3463
rect 5870 3377 5900 3463
rect 2870 3237 2900 3323
rect 3070 3237 3100 3323
rect 3170 3237 3200 3323
rect 3270 3237 3300 3323
rect 3370 3237 3400 3323
rect 3470 3237 3500 3323
rect 3570 3237 3600 3323
rect 3670 3237 3700 3323
rect 3770 3237 3800 3323
rect 3870 3237 3900 3323
rect 3970 3237 4000 3323
rect 4070 3237 4100 3323
rect 4170 3237 4200 3323
rect 4270 3237 4300 3323
rect 2570 3097 2600 3183
rect 2670 3097 2700 3183
rect 2770 3097 2800 3183
rect 2870 3097 2900 3183
rect 2970 3097 3000 3183
rect 3070 3097 3100 3183
rect 3170 3097 3200 3183
rect 3370 3097 3400 3183
rect 3470 3097 3500 3183
rect 3570 3097 3600 3183
rect 70 2957 100 3043
rect 170 2957 200 3043
rect 270 2957 300 3043
rect 370 2957 400 3043
rect 470 2957 500 3043
rect 570 2957 600 3043
rect 670 2957 700 3043
rect 770 2957 800 3043
rect 870 2957 900 3043
rect 970 2957 1000 3043
rect 1070 2957 1100 3043
rect 1170 2957 1200 3043
rect 1270 2957 1300 3043
rect 1370 2957 1400 3043
rect 1470 2957 1500 3043
rect 1570 2957 1600 3043
rect 1670 2957 1700 3043
rect 1770 2957 1800 3043
rect 1870 2957 1900 3043
rect 1970 2957 2000 3043
rect 2070 2957 2100 3043
rect 2170 2957 2200 3043
rect 2270 2957 2300 3043
rect 2370 2957 2400 3043
rect 2470 2957 2500 3043
rect 2570 2957 2600 3043
rect 2670 2957 2700 3043
rect 2770 2957 2800 3043
rect 2870 2957 2900 3043
rect 2970 2957 3000 3043
rect 3070 2957 3100 3043
rect 3170 2957 3200 3043
rect 3270 2957 3300 3043
rect 70 2817 100 2903
rect 170 2817 200 2903
rect 270 2817 300 2903
rect 470 2817 500 2903
rect 570 2817 600 2903
rect 670 2817 700 2903
rect 870 2817 900 2903
rect 970 2817 1000 2903
rect 1070 2817 1100 2903
rect 1170 2817 1200 2903
rect 1270 2817 1300 2903
rect 1370 2817 1400 2903
rect 70 2677 100 2763
rect 170 2677 200 2763
rect 270 2677 300 2763
rect 370 2677 400 2763
rect 470 2677 500 2763
rect 570 2677 600 2763
rect 670 2677 700 2763
rect 770 2677 800 2763
rect 870 2677 900 2763
rect 970 2677 1000 2763
rect 1070 2677 1100 2763
rect 1170 2677 1200 2763
rect 1270 2677 1300 2763
rect 1570 2817 1600 2903
rect 1670 2817 1700 2903
rect 1770 2817 1800 2903
rect 1870 2817 1900 2903
rect 1970 2817 2000 2903
rect 2070 2817 2100 2903
rect 1470 2677 1500 2763
rect 70 2537 100 2623
rect 170 2537 200 2623
rect 270 2537 300 2623
rect 370 2537 400 2623
rect 470 2537 500 2623
rect 570 2537 600 2623
rect 670 2537 700 2623
rect 770 2537 800 2623
rect 870 2537 900 2623
rect 970 2537 1000 2623
rect 1070 2537 1100 2623
rect 1170 2537 1200 2623
rect 1270 2537 1300 2623
rect 1370 2537 1400 2623
rect 1470 2537 1500 2623
rect 1670 2677 1700 2763
rect 1770 2677 1800 2763
rect 1870 2677 1900 2763
rect 1970 2677 2000 2763
rect 2270 2817 2300 2903
rect 2470 2817 2500 2903
rect 2670 2817 2700 2903
rect 2770 2817 2800 2903
rect 2870 2817 2900 2903
rect 2970 2817 3000 2903
rect 2170 2677 2200 2763
rect 2270 2677 2300 2763
rect 2370 2677 2400 2763
rect 2470 2677 2500 2763
rect 2570 2677 2600 2763
rect 2670 2677 2700 2763
rect 2770 2677 2800 2763
rect 1670 2537 1700 2623
rect 1770 2537 1800 2623
rect 1870 2537 1900 2623
rect 1970 2537 2000 2623
rect 2070 2537 2100 2623
rect 2270 2537 2300 2623
rect 2370 2537 2400 2623
rect 2570 2537 2600 2623
rect 3770 3097 3800 3183
rect 3870 3097 3900 3183
rect 3970 3097 4000 3183
rect 4070 3097 4100 3183
rect 4170 3097 4200 3183
rect 3470 2957 3500 3043
rect 3570 2957 3600 3043
rect 3670 2957 3700 3043
rect 3770 2957 3800 3043
rect 3970 2957 4000 3043
rect 4470 3237 4500 3323
rect 4570 3237 4600 3323
rect 4670 3237 4700 3323
rect 4770 3237 4800 3323
rect 4370 3097 4400 3183
rect 4470 3097 4500 3183
rect 4170 2957 4200 3043
rect 4270 2957 4300 3043
rect 4370 2957 4400 3043
rect 4470 2957 4500 3043
rect 4670 3097 4700 3183
rect 4970 3237 5000 3323
rect 5070 3237 5100 3323
rect 5170 3237 5200 3323
rect 5270 3237 5300 3323
rect 5370 3237 5400 3323
rect 5470 3237 5500 3323
rect 4870 3097 4900 3183
rect 4970 3097 5000 3183
rect 5170 3097 5200 3183
rect 5270 3097 5300 3183
rect 5370 3097 5400 3183
rect 5470 3097 5500 3183
rect 6070 3377 6100 3463
rect 6170 3377 6200 3463
rect 6270 3377 6300 3463
rect 6370 3377 6400 3463
rect 6570 3377 6600 3463
rect 6670 3377 6700 3463
rect 6880 3377 6910 3463
rect 6980 3377 7010 3463
rect 7080 3377 7110 3463
rect 7180 3377 7210 3463
rect 7280 3377 7310 3463
rect 7380 3377 7410 3463
rect 5670 3237 5700 3323
rect 5770 3237 5800 3323
rect 5870 3237 5900 3323
rect 5970 3237 6000 3323
rect 6070 3237 6100 3323
rect 6170 3237 6200 3323
rect 6270 3237 6300 3323
rect 6370 3237 6400 3323
rect 6570 3237 6600 3323
rect 6670 3237 6700 3323
rect 6880 3237 6910 3323
rect 6980 3237 7010 3323
rect 7080 3237 7110 3323
rect 7180 3237 7210 3323
rect 7280 3237 7310 3323
rect 7380 3237 7410 3323
rect 5670 3097 5700 3183
rect 5870 3097 5900 3183
rect 5970 3097 6000 3183
rect 6070 3097 6100 3183
rect 6170 3097 6200 3183
rect 6270 3097 6300 3183
rect 6370 3097 6400 3183
rect 6570 3097 6600 3183
rect 6670 3097 6700 3183
rect 6880 3097 6910 3183
rect 6980 3097 7010 3183
rect 7080 3097 7110 3183
rect 7180 3097 7210 3183
rect 7280 3097 7310 3183
rect 7380 3097 7410 3183
rect 4670 2957 4700 3043
rect 4770 2957 4800 3043
rect 4870 2957 4900 3043
rect 4970 2957 5000 3043
rect 5070 2957 5100 3043
rect 5170 2957 5200 3043
rect 5270 2957 5300 3043
rect 5370 2957 5400 3043
rect 5470 2957 5500 3043
rect 5570 2957 5600 3043
rect 5670 2957 5700 3043
rect 5770 2957 5800 3043
rect 5870 2957 5900 3043
rect 6070 2957 6100 3043
rect 6170 2957 6200 3043
rect 6270 2957 6300 3043
rect 6370 2957 6400 3043
rect 6570 2957 6600 3043
rect 6670 2957 6700 3043
rect 6880 2957 6910 3043
rect 6980 2957 7010 3043
rect 7080 2957 7110 3043
rect 7180 2957 7210 3043
rect 7280 2957 7310 3043
rect 7380 2957 7410 3043
rect 3170 2817 3200 2903
rect 3270 2817 3300 2903
rect 3370 2817 3400 2903
rect 3470 2817 3500 2903
rect 3570 2817 3600 2903
rect 3670 2817 3700 2903
rect 3770 2817 3800 2903
rect 3870 2817 3900 2903
rect 3970 2817 4000 2903
rect 4070 2817 4100 2903
rect 4170 2817 4200 2903
rect 4270 2817 4300 2903
rect 4370 2817 4400 2903
rect 4470 2817 4500 2903
rect 4570 2817 4600 2903
rect 4670 2817 4700 2903
rect 4770 2817 4800 2903
rect 4870 2817 4900 2903
rect 4970 2817 5000 2903
rect 5070 2817 5100 2903
rect 5170 2817 5200 2903
rect 5270 2817 5300 2903
rect 5370 2817 5400 2903
rect 5470 2817 5500 2903
rect 5570 2817 5600 2903
rect 5670 2817 5700 2903
rect 5770 2817 5800 2903
rect 5870 2817 5900 2903
rect 5970 2817 6000 2903
rect 2970 2677 3000 2763
rect 3070 2677 3100 2763
rect 3270 2677 3300 2763
rect 3370 2677 3400 2763
rect 3470 2677 3500 2763
rect 3570 2677 3600 2763
rect 3670 2677 3700 2763
rect 3770 2677 3800 2763
rect 3870 2677 3900 2763
rect 3970 2677 4000 2763
rect 4070 2677 4100 2763
rect 4170 2677 4200 2763
rect 4270 2677 4300 2763
rect 4370 2677 4400 2763
rect 2770 2537 2800 2623
rect 2870 2537 2900 2623
rect 2970 2537 3000 2623
rect 3070 2537 3100 2623
rect 3170 2537 3200 2623
rect 3370 2537 3400 2623
rect 4570 2677 4600 2763
rect 4770 2677 4800 2763
rect 4870 2677 4900 2763
rect 4970 2677 5000 2763
rect 5070 2677 5100 2763
rect 5170 2677 5200 2763
rect 5270 2677 5300 2763
rect 5370 2677 5400 2763
rect 6170 2817 6200 2903
rect 6270 2817 6300 2903
rect 6370 2817 6400 2903
rect 6570 2817 6600 2903
rect 6670 2817 6700 2903
rect 6880 2817 6910 2903
rect 6980 2817 7010 2903
rect 7080 2817 7110 2903
rect 7180 2817 7210 2903
rect 7280 2817 7310 2903
rect 7380 2817 7410 2903
rect 5570 2677 5600 2763
rect 5670 2677 5700 2763
rect 5770 2677 5800 2763
rect 5870 2677 5900 2763
rect 5970 2677 6000 2763
rect 6070 2677 6100 2763
rect 6170 2677 6200 2763
rect 6270 2677 6300 2763
rect 6370 2677 6400 2763
rect 6570 2677 6600 2763
rect 6670 2677 6700 2763
rect 6880 2677 6910 2763
rect 6980 2677 7010 2763
rect 7080 2677 7110 2763
rect 7180 2677 7210 2763
rect 7280 2677 7310 2763
rect 7380 2677 7410 2763
rect 3570 2537 3600 2623
rect 3670 2537 3700 2623
rect 3770 2537 3800 2623
rect 3870 2537 3900 2623
rect 3970 2537 4000 2623
rect 4070 2537 4100 2623
rect 4170 2537 4200 2623
rect 4270 2537 4300 2623
rect 4370 2537 4400 2623
rect 4470 2537 4500 2623
rect 4570 2537 4600 2623
rect 4670 2537 4700 2623
rect 4770 2537 4800 2623
rect 4870 2537 4900 2623
rect 4970 2537 5000 2623
rect 5070 2537 5100 2623
rect 5170 2537 5200 2623
rect 5270 2537 5300 2623
rect 5370 2537 5400 2623
rect 5470 2537 5500 2623
rect 5670 2537 5700 2623
rect 5770 2537 5800 2623
rect 5870 2537 5900 2623
rect 5970 2537 6000 2623
rect 6070 2537 6100 2623
rect 6170 2537 6200 2623
rect 6270 2537 6300 2623
rect 6370 2537 6400 2623
rect 6570 2537 6600 2623
rect 6670 2537 6700 2623
rect 6880 2537 6910 2623
rect 6980 2537 7010 2623
rect 7080 2537 7110 2623
rect 7180 2537 7210 2623
rect 7280 2537 7310 2623
rect 7380 2537 7410 2623
rect 70 2307 100 2393
rect 170 2307 200 2393
rect 270 2307 300 2393
rect 370 2307 400 2393
rect 470 2307 500 2393
rect 570 2307 600 2393
rect 670 2307 700 2393
rect 770 2307 800 2393
rect 870 2307 900 2393
rect 970 2307 1000 2393
rect 1070 2307 1100 2393
rect 1170 2307 1200 2393
rect 1270 2307 1300 2393
rect 1370 2307 1400 2393
rect 1470 2307 1500 2393
rect 1570 2307 1600 2393
rect 1670 2307 1700 2393
rect 1770 2307 1800 2393
rect 1870 2307 1900 2393
rect 1970 2307 2000 2393
rect 2070 2307 2100 2393
rect 2170 2307 2200 2393
rect 2270 2307 2300 2393
rect 2370 2307 2400 2393
rect 2470 2307 2500 2393
rect 2570 2307 2600 2393
rect 2670 2307 2700 2393
rect 2770 2307 2800 2393
rect 2870 2307 2900 2393
rect 2970 2307 3000 2393
rect 3070 2307 3100 2393
rect 3170 2307 3200 2393
rect 3270 2307 3300 2393
rect 3370 2307 3400 2393
rect 3470 2307 3500 2393
rect 3570 2307 3600 2393
rect 3670 2307 3700 2393
rect 3770 2307 3800 2393
rect 3870 2307 3900 2393
rect 3970 2307 4000 2393
rect 4070 2307 4100 2393
rect 4170 2307 4200 2393
rect 4270 2307 4300 2393
rect 4370 2307 4400 2393
rect 4470 2307 4500 2393
rect 4570 2307 4600 2393
rect 4670 2307 4700 2393
rect 4770 2307 4800 2393
rect 4870 2307 4900 2393
rect 4970 2307 5000 2393
rect 5070 2307 5100 2393
rect 5170 2307 5200 2393
rect 5270 2307 5300 2393
rect 5370 2307 5400 2393
rect 70 2167 100 2253
rect 170 2167 200 2253
rect 370 2167 400 2253
rect 470 2167 500 2253
rect 570 2167 600 2253
rect 670 2167 700 2253
rect 770 2167 800 2253
rect 870 2167 900 2253
rect 970 2167 1000 2253
rect 1070 2167 1100 2253
rect 1170 2167 1200 2253
rect 1270 2167 1300 2253
rect 70 2027 100 2113
rect 170 2027 200 2113
rect 270 2027 300 2113
rect 70 1887 100 1973
rect 170 1887 200 1973
rect 270 1887 300 1973
rect 470 2027 500 2113
rect 570 2027 600 2113
rect 670 2027 700 2113
rect 770 2027 800 2113
rect 870 2027 900 2113
rect 970 2027 1000 2113
rect 1070 2027 1100 2113
rect 1170 2027 1200 2113
rect 1270 2027 1300 2113
rect 1470 2167 1500 2253
rect 1470 2027 1500 2113
rect 470 1887 500 1973
rect 570 1887 600 1973
rect 670 1887 700 1973
rect 770 1887 800 1973
rect 870 1887 900 1973
rect 970 1887 1000 1973
rect 1070 1887 1100 1973
rect 1170 1887 1200 1973
rect 1270 1887 1300 1973
rect 1370 1887 1400 1973
rect 70 1747 100 1833
rect 170 1747 200 1833
rect 270 1747 300 1833
rect 370 1747 400 1833
rect 470 1747 500 1833
rect 570 1747 600 1833
rect 670 1747 700 1833
rect 770 1747 800 1833
rect 870 1747 900 1833
rect 70 1607 100 1693
rect 70 1467 100 1553
rect 270 1607 300 1693
rect 370 1607 400 1693
rect 470 1607 500 1693
rect 570 1607 600 1693
rect 670 1607 700 1693
rect 270 1467 300 1553
rect 370 1467 400 1553
rect 70 1327 100 1413
rect 170 1327 200 1413
rect 870 1607 900 1693
rect 1670 2167 1700 2253
rect 1770 2167 1800 2253
rect 1670 2027 1700 2113
rect 1770 2027 1800 2113
rect 1970 2167 2000 2253
rect 2070 2167 2100 2253
rect 2170 2167 2200 2253
rect 1970 2027 2000 2113
rect 2070 2027 2100 2113
rect 2170 2027 2200 2113
rect 2370 2167 2400 2253
rect 2470 2167 2500 2253
rect 2570 2167 2600 2253
rect 2670 2167 2700 2253
rect 2770 2167 2800 2253
rect 2370 2027 2400 2113
rect 1570 1887 1600 1973
rect 1670 1887 1700 1973
rect 1770 1887 1800 1973
rect 1870 1887 1900 1973
rect 1970 1887 2000 1973
rect 2070 1887 2100 1973
rect 2170 1887 2200 1973
rect 2270 1887 2300 1973
rect 2370 1887 2400 1973
rect 1070 1747 1100 1833
rect 1170 1747 1200 1833
rect 1270 1747 1300 1833
rect 1370 1747 1400 1833
rect 1470 1747 1500 1833
rect 1570 1747 1600 1833
rect 1670 1747 1700 1833
rect 1770 1747 1800 1833
rect 1070 1607 1100 1693
rect 1170 1607 1200 1693
rect 1270 1607 1300 1693
rect 1370 1607 1400 1693
rect 1470 1607 1500 1693
rect 1670 1607 1700 1693
rect 570 1467 600 1553
rect 670 1467 700 1553
rect 770 1467 800 1553
rect 870 1467 900 1553
rect 970 1467 1000 1553
rect 1070 1467 1100 1553
rect 1170 1467 1200 1553
rect 1270 1467 1300 1553
rect 1370 1467 1400 1553
rect 1470 1467 1500 1553
rect 1570 1467 1600 1553
rect 370 1327 400 1413
rect 470 1327 500 1413
rect 70 1097 100 1183
rect 170 1097 200 1183
rect 270 1097 300 1183
rect 670 1327 700 1413
rect 770 1327 800 1413
rect 870 1327 900 1413
rect 970 1327 1000 1413
rect 1070 1327 1100 1413
rect 1170 1327 1200 1413
rect 1270 1327 1300 1413
rect 1370 1327 1400 1413
rect 1470 1327 1500 1413
rect 470 1097 500 1183
rect 670 1097 700 1183
rect 870 1097 900 1183
rect 970 1097 1000 1183
rect 1070 1097 1100 1183
rect 1170 1097 1200 1183
rect 70 957 100 1043
rect 170 957 200 1043
rect 270 957 300 1043
rect 370 957 400 1043
rect 470 957 500 1043
rect 570 957 600 1043
rect 670 957 700 1043
rect 770 957 800 1043
rect 870 957 900 1043
rect 1070 957 1100 1043
rect 70 817 100 903
rect 170 817 200 903
rect 270 817 300 903
rect 370 817 400 903
rect 470 817 500 903
rect 570 817 600 903
rect 670 817 700 903
rect 770 817 800 903
rect 870 817 900 903
rect 970 817 1000 903
rect 70 677 100 763
rect 170 677 200 763
rect 270 677 300 763
rect 370 677 400 763
rect 470 677 500 763
rect 570 677 600 763
rect 670 677 700 763
rect 770 677 800 763
rect 870 677 900 763
rect 70 537 100 623
rect 170 537 200 623
rect 270 537 300 623
rect 370 537 400 623
rect 470 537 500 623
rect 70 397 100 483
rect 170 397 200 483
rect 370 397 400 483
rect 2970 2167 3000 2253
rect 3070 2167 3100 2253
rect 3170 2167 3200 2253
rect 3270 2167 3300 2253
rect 3370 2167 3400 2253
rect 3470 2167 3500 2253
rect 2570 2027 2600 2113
rect 2670 2027 2700 2113
rect 2770 2027 2800 2113
rect 2870 2027 2900 2113
rect 2970 2027 3000 2113
rect 3070 2027 3100 2113
rect 3170 2027 3200 2113
rect 3270 2027 3300 2113
rect 2570 1887 2600 1973
rect 2670 1887 2700 1973
rect 2770 1887 2800 1973
rect 2870 1887 2900 1973
rect 2970 1887 3000 1973
rect 3670 2167 3700 2253
rect 3770 2167 3800 2253
rect 3870 2167 3900 2253
rect 3970 2167 4000 2253
rect 4070 2167 4100 2253
rect 4170 2167 4200 2253
rect 3470 2027 3500 2113
rect 3570 2027 3600 2113
rect 3770 2027 3800 2113
rect 3870 2027 3900 2113
rect 3170 1887 3200 1973
rect 3270 1887 3300 1973
rect 3370 1887 3400 1973
rect 3470 1887 3500 1973
rect 3570 1887 3600 1973
rect 3670 1887 3700 1973
rect 3770 1887 3800 1973
rect 1970 1747 2000 1833
rect 2070 1747 2100 1833
rect 2170 1747 2200 1833
rect 2270 1747 2300 1833
rect 2370 1747 2400 1833
rect 2470 1747 2500 1833
rect 2570 1747 2600 1833
rect 2670 1747 2700 1833
rect 2770 1747 2800 1833
rect 2870 1747 2900 1833
rect 2970 1747 3000 1833
rect 3070 1747 3100 1833
rect 3170 1747 3200 1833
rect 3270 1747 3300 1833
rect 3370 1747 3400 1833
rect 1870 1607 1900 1693
rect 2070 1607 2100 1693
rect 2170 1607 2200 1693
rect 2270 1607 2300 1693
rect 2370 1607 2400 1693
rect 2470 1607 2500 1693
rect 2570 1607 2600 1693
rect 2770 1607 2800 1693
rect 2870 1607 2900 1693
rect 2970 1607 3000 1693
rect 3070 1607 3100 1693
rect 3170 1607 3200 1693
rect 3270 1607 3300 1693
rect 3370 1607 3400 1693
rect 3570 1747 3600 1833
rect 4370 2167 4400 2253
rect 4070 2027 4100 2113
rect 4170 2027 4200 2113
rect 4270 2027 4300 2113
rect 4370 2027 4400 2113
rect 3970 1887 4000 1973
rect 4070 1887 4100 1973
rect 4170 1887 4200 1973
rect 4270 1887 4300 1973
rect 4370 1887 4400 1973
rect 3770 1747 3800 1833
rect 3870 1747 3900 1833
rect 3570 1607 3600 1693
rect 3670 1607 3700 1693
rect 5570 2307 5600 2393
rect 5670 2307 5700 2393
rect 5770 2307 5800 2393
rect 5870 2307 5900 2393
rect 5970 2307 6000 2393
rect 6070 2307 6100 2393
rect 6170 2307 6200 2393
rect 6270 2307 6300 2393
rect 6370 2307 6400 2393
rect 6570 2307 6600 2393
rect 6670 2307 6700 2393
rect 6880 2307 6910 2393
rect 6980 2307 7010 2393
rect 7080 2307 7110 2393
rect 7180 2307 7210 2393
rect 7280 2307 7310 2393
rect 7380 2307 7410 2393
rect 4570 2167 4600 2253
rect 4670 2167 4700 2253
rect 4770 2167 4800 2253
rect 4870 2167 4900 2253
rect 4970 2167 5000 2253
rect 5070 2167 5100 2253
rect 5170 2167 5200 2253
rect 5270 2167 5300 2253
rect 5370 2167 5400 2253
rect 5470 2167 5500 2253
rect 5570 2167 5600 2253
rect 5670 2167 5700 2253
rect 5770 2167 5800 2253
rect 5870 2167 5900 2253
rect 5970 2167 6000 2253
rect 6070 2167 6100 2253
rect 6170 2167 6200 2253
rect 6270 2167 6300 2253
rect 6370 2167 6400 2253
rect 6570 2167 6600 2253
rect 6670 2167 6700 2253
rect 6880 2167 6910 2253
rect 6980 2167 7010 2253
rect 7080 2167 7110 2253
rect 7180 2167 7210 2253
rect 7280 2167 7310 2253
rect 7380 2167 7410 2253
rect 4570 2027 4600 2113
rect 4670 2027 4700 2113
rect 4770 2027 4800 2113
rect 4870 2027 4900 2113
rect 4970 2027 5000 2113
rect 5070 2027 5100 2113
rect 5170 2027 5200 2113
rect 5270 2027 5300 2113
rect 5370 2027 5400 2113
rect 5470 2027 5500 2113
rect 5570 2027 5600 2113
rect 5670 2027 5700 2113
rect 5770 2027 5800 2113
rect 5870 2027 5900 2113
rect 5970 2027 6000 2113
rect 6070 2027 6100 2113
rect 6170 2027 6200 2113
rect 6270 2027 6300 2113
rect 6370 2027 6400 2113
rect 6570 2027 6600 2113
rect 6670 2027 6700 2113
rect 6880 2027 6910 2113
rect 6980 2027 7010 2113
rect 7080 2027 7110 2113
rect 7180 2027 7210 2113
rect 7280 2027 7310 2113
rect 7380 2027 7410 2113
rect 4570 1887 4600 1973
rect 4670 1887 4700 1973
rect 4770 1887 4800 1973
rect 4870 1887 4900 1973
rect 4070 1747 4100 1833
rect 4170 1747 4200 1833
rect 4270 1747 4300 1833
rect 4370 1747 4400 1833
rect 4470 1747 4500 1833
rect 4570 1747 4600 1833
rect 4670 1747 4700 1833
rect 4770 1747 4800 1833
rect 3870 1607 3900 1693
rect 3970 1607 4000 1693
rect 4070 1607 4100 1693
rect 4170 1607 4200 1693
rect 4270 1607 4300 1693
rect 4370 1607 4400 1693
rect 1770 1467 1800 1553
rect 1870 1467 1900 1553
rect 1970 1467 2000 1553
rect 2070 1467 2100 1553
rect 2170 1467 2200 1553
rect 2270 1467 2300 1553
rect 2370 1467 2400 1553
rect 2470 1467 2500 1553
rect 2570 1467 2600 1553
rect 2670 1467 2700 1553
rect 2770 1467 2800 1553
rect 2870 1467 2900 1553
rect 2970 1467 3000 1553
rect 3070 1467 3100 1553
rect 3170 1467 3200 1553
rect 3270 1467 3300 1553
rect 3370 1467 3400 1553
rect 3470 1467 3500 1553
rect 3570 1467 3600 1553
rect 3670 1467 3700 1553
rect 3770 1467 3800 1553
rect 3870 1467 3900 1553
rect 3970 1467 4000 1553
rect 4070 1467 4100 1553
rect 1670 1327 1700 1413
rect 1870 1327 1900 1413
rect 1970 1327 2000 1413
rect 2070 1327 2100 1413
rect 2170 1327 2200 1413
rect 2270 1327 2300 1413
rect 2370 1327 2400 1413
rect 2470 1327 2500 1413
rect 2570 1327 2600 1413
rect 2670 1327 2700 1413
rect 2770 1327 2800 1413
rect 2870 1327 2900 1413
rect 1370 1097 1400 1183
rect 1470 1097 1500 1183
rect 1570 1097 1600 1183
rect 1670 1097 1700 1183
rect 1770 1097 1800 1183
rect 1870 1097 1900 1183
rect 1970 1097 2000 1183
rect 2070 1097 2100 1183
rect 2170 1097 2200 1183
rect 2270 1097 2300 1183
rect 2370 1097 2400 1183
rect 2470 1097 2500 1183
rect 1270 957 1300 1043
rect 1370 957 1400 1043
rect 1470 957 1500 1043
rect 1570 957 1600 1043
rect 1670 957 1700 1043
rect 1770 957 1800 1043
rect 1870 957 1900 1043
rect 1970 957 2000 1043
rect 2070 957 2100 1043
rect 1170 817 1200 903
rect 1270 817 1300 903
rect 1370 817 1400 903
rect 1470 817 1500 903
rect 1570 817 1600 903
rect 1670 817 1700 903
rect 2270 957 2300 1043
rect 2370 957 2400 1043
rect 2670 1097 2700 1183
rect 3070 1327 3100 1413
rect 3170 1327 3200 1413
rect 3270 1327 3300 1413
rect 3370 1327 3400 1413
rect 3470 1327 3500 1413
rect 3670 1327 3700 1413
rect 3770 1327 3800 1413
rect 4270 1467 4300 1553
rect 4370 1467 4400 1553
rect 5070 1887 5100 1973
rect 5270 1887 5300 1973
rect 5470 1887 5500 1973
rect 5570 1887 5600 1973
rect 5670 1887 5700 1973
rect 5870 1887 5900 1973
rect 5970 1887 6000 1973
rect 6170 1887 6200 1973
rect 6270 1887 6300 1973
rect 6370 1887 6400 1973
rect 6570 1887 6600 1973
rect 6670 1887 6700 1973
rect 6880 1887 6910 1973
rect 6980 1887 7010 1973
rect 7080 1887 7110 1973
rect 7180 1887 7210 1973
rect 7280 1887 7310 1973
rect 7380 1887 7410 1973
rect 4970 1747 5000 1833
rect 5070 1747 5100 1833
rect 5170 1747 5200 1833
rect 5270 1747 5300 1833
rect 5370 1747 5400 1833
rect 5470 1747 5500 1833
rect 5570 1747 5600 1833
rect 5670 1747 5700 1833
rect 5770 1747 5800 1833
rect 5870 1747 5900 1833
rect 5970 1747 6000 1833
rect 6070 1747 6100 1833
rect 6170 1747 6200 1833
rect 6270 1747 6300 1833
rect 6370 1747 6400 1833
rect 6570 1747 6600 1833
rect 6670 1747 6700 1833
rect 6880 1747 6910 1833
rect 6980 1747 7010 1833
rect 7080 1747 7110 1833
rect 7180 1747 7210 1833
rect 7280 1747 7310 1833
rect 7380 1747 7410 1833
rect 4570 1607 4600 1693
rect 4670 1607 4700 1693
rect 4770 1607 4800 1693
rect 4870 1607 4900 1693
rect 4970 1607 5000 1693
rect 5070 1607 5100 1693
rect 5170 1607 5200 1693
rect 5270 1607 5300 1693
rect 4570 1467 4600 1553
rect 4670 1467 4700 1553
rect 4770 1467 4800 1553
rect 4870 1467 4900 1553
rect 4970 1467 5000 1553
rect 3970 1327 4000 1413
rect 4070 1327 4100 1413
rect 4170 1327 4200 1413
rect 4270 1327 4300 1413
rect 4370 1327 4400 1413
rect 4470 1327 4500 1413
rect 4570 1327 4600 1413
rect 4670 1327 4700 1413
rect 4770 1327 4800 1413
rect 2870 1097 2900 1183
rect 2970 1097 3000 1183
rect 3070 1097 3100 1183
rect 3170 1097 3200 1183
rect 3270 1097 3300 1183
rect 3370 1097 3400 1183
rect 3470 1097 3500 1183
rect 3570 1097 3600 1183
rect 3670 1097 3700 1183
rect 3770 1097 3800 1183
rect 3870 1097 3900 1183
rect 3970 1097 4000 1183
rect 4070 1097 4100 1183
rect 4170 1097 4200 1183
rect 2570 957 2600 1043
rect 2670 957 2700 1043
rect 2770 957 2800 1043
rect 2870 957 2900 1043
rect 2970 957 3000 1043
rect 3070 957 3100 1043
rect 3170 957 3200 1043
rect 3270 957 3300 1043
rect 3370 957 3400 1043
rect 3470 957 3500 1043
rect 3570 957 3600 1043
rect 3670 957 3700 1043
rect 3770 957 3800 1043
rect 3870 957 3900 1043
rect 3970 957 4000 1043
rect 4070 957 4100 1043
rect 4170 957 4200 1043
rect 4970 1327 5000 1413
rect 5170 1467 5200 1553
rect 5470 1607 5500 1693
rect 5570 1607 5600 1693
rect 5670 1607 5700 1693
rect 5370 1467 5400 1553
rect 5570 1467 5600 1553
rect 5670 1467 5700 1553
rect 5870 1607 5900 1693
rect 5870 1467 5900 1553
rect 6070 1607 6100 1693
rect 6170 1607 6200 1693
rect 6270 1607 6300 1693
rect 6370 1607 6400 1693
rect 6570 1607 6600 1693
rect 6670 1607 6700 1693
rect 6880 1607 6910 1693
rect 6980 1607 7010 1693
rect 7080 1607 7110 1693
rect 7180 1607 7210 1693
rect 7280 1607 7310 1693
rect 7380 1607 7410 1693
rect 6070 1467 6100 1553
rect 6170 1467 6200 1553
rect 5170 1327 5200 1413
rect 5270 1327 5300 1413
rect 5370 1327 5400 1413
rect 5470 1327 5500 1413
rect 5570 1327 5600 1413
rect 5670 1327 5700 1413
rect 5770 1327 5800 1413
rect 5870 1327 5900 1413
rect 5970 1327 6000 1413
rect 6070 1327 6100 1413
rect 4370 1097 4400 1183
rect 4470 1097 4500 1183
rect 4570 1097 4600 1183
rect 4670 1097 4700 1183
rect 4770 1097 4800 1183
rect 4870 1097 4900 1183
rect 4970 1097 5000 1183
rect 5070 1097 5100 1183
rect 5170 1097 5200 1183
rect 5270 1097 5300 1183
rect 5370 1097 5400 1183
rect 4370 957 4400 1043
rect 4470 957 4500 1043
rect 4570 957 4600 1043
rect 4670 957 4700 1043
rect 4770 957 4800 1043
rect 1870 817 1900 903
rect 1970 817 2000 903
rect 2070 817 2100 903
rect 2170 817 2200 903
rect 2270 817 2300 903
rect 2370 817 2400 903
rect 2470 817 2500 903
rect 2570 817 2600 903
rect 2670 817 2700 903
rect 2770 817 2800 903
rect 2870 817 2900 903
rect 2970 817 3000 903
rect 3070 817 3100 903
rect 3170 817 3200 903
rect 3270 817 3300 903
rect 3370 817 3400 903
rect 3470 817 3500 903
rect 3570 817 3600 903
rect 3670 817 3700 903
rect 3770 817 3800 903
rect 3870 817 3900 903
rect 3970 817 4000 903
rect 4070 817 4100 903
rect 4170 817 4200 903
rect 4270 817 4300 903
rect 1070 677 1100 763
rect 1170 677 1200 763
rect 1270 677 1300 763
rect 1370 677 1400 763
rect 1470 677 1500 763
rect 1570 677 1600 763
rect 1670 677 1700 763
rect 1770 677 1800 763
rect 1870 677 1900 763
rect 1970 677 2000 763
rect 670 537 700 623
rect 770 537 800 623
rect 870 537 900 623
rect 970 537 1000 623
rect 2170 677 2200 763
rect 4470 817 4500 903
rect 2370 677 2400 763
rect 2470 677 2500 763
rect 2570 677 2600 763
rect 2670 677 2700 763
rect 2770 677 2800 763
rect 2870 677 2900 763
rect 2970 677 3000 763
rect 3070 677 3100 763
rect 3170 677 3200 763
rect 3270 677 3300 763
rect 3370 677 3400 763
rect 3470 677 3500 763
rect 3570 677 3600 763
rect 3670 677 3700 763
rect 3770 677 3800 763
rect 3870 677 3900 763
rect 3970 677 4000 763
rect 4070 677 4100 763
rect 4170 677 4200 763
rect 4270 677 4300 763
rect 4370 677 4400 763
rect 1170 537 1200 623
rect 1270 537 1300 623
rect 1370 537 1400 623
rect 1470 537 1500 623
rect 1570 537 1600 623
rect 1670 537 1700 623
rect 1770 537 1800 623
rect 1870 537 1900 623
rect 1970 537 2000 623
rect 2070 537 2100 623
rect 2170 537 2200 623
rect 2270 537 2300 623
rect 2370 537 2400 623
rect 2470 537 2500 623
rect 2570 537 2600 623
rect 2670 537 2700 623
rect 2770 537 2800 623
rect 2870 537 2900 623
rect 2970 537 3000 623
rect 3070 537 3100 623
rect 3170 537 3200 623
rect 3270 537 3300 623
rect 3370 537 3400 623
rect 3470 537 3500 623
rect 3570 537 3600 623
rect 3670 537 3700 623
rect 570 397 600 483
rect 670 397 700 483
rect 770 397 800 483
rect 870 397 900 483
rect 970 397 1000 483
rect 1070 397 1100 483
rect 1170 397 1200 483
rect 1270 397 1300 483
rect 1370 397 1400 483
rect 70 257 100 343
rect 170 257 200 343
rect 270 257 300 343
rect 370 257 400 343
rect 470 257 500 343
rect 570 257 600 343
rect 1570 397 1600 483
rect 1670 397 1700 483
rect 1770 397 1800 483
rect 1870 397 1900 483
rect 1970 397 2000 483
rect 2070 397 2100 483
rect 2170 397 2200 483
rect 2270 397 2300 483
rect 2370 397 2400 483
rect 2470 397 2500 483
rect 2570 397 2600 483
rect 2670 397 2700 483
rect 2770 397 2800 483
rect 2870 397 2900 483
rect 2970 397 3000 483
rect 770 257 800 343
rect 870 257 900 343
rect 970 257 1000 343
rect 1070 257 1100 343
rect 1170 257 1200 343
rect 1270 257 1300 343
rect 1370 257 1400 343
rect 1470 257 1500 343
rect 70 117 100 203
rect 170 117 200 203
rect 270 117 300 203
rect 370 117 400 203
rect 470 117 500 203
rect 570 117 600 203
rect 670 117 700 203
rect 770 117 800 203
rect 1670 257 1700 343
rect 1770 257 1800 343
rect 1870 257 1900 343
rect 1970 257 2000 343
rect 2070 257 2100 343
rect 2170 257 2200 343
rect 970 117 1000 203
rect 1070 117 1100 203
rect 1170 117 1200 203
rect 1270 117 1300 203
rect 1370 117 1400 203
rect 1470 117 1500 203
rect 1570 117 1600 203
rect 1670 117 1700 203
rect 1770 117 1800 203
rect 1870 117 1900 203
rect 2370 257 2400 343
rect 2570 257 2600 343
rect 2770 257 2800 343
rect 3170 397 3200 483
rect 3370 397 3400 483
rect 3470 397 3500 483
rect 2970 257 3000 343
rect 3070 257 3100 343
rect 3170 257 3200 343
rect 3270 257 3300 343
rect 3370 257 3400 343
rect 3470 257 3500 343
rect 2070 117 2100 203
rect 2170 117 2200 203
rect 2270 117 2300 203
rect 2370 117 2400 203
rect 2470 117 2500 203
rect 2570 117 2600 203
rect 2670 117 2700 203
rect 2770 117 2800 203
rect 2870 117 2900 203
rect 2970 117 3000 203
rect 3070 117 3100 203
rect 3170 117 3200 203
rect 3270 117 3300 203
rect 3370 117 3400 203
rect 3470 117 3500 203
rect 3670 397 3700 483
rect 3870 537 3900 623
rect 3970 537 4000 623
rect 4170 537 4200 623
rect 4970 957 5000 1043
rect 5570 1097 5600 1183
rect 5670 1097 5700 1183
rect 5770 1097 5800 1183
rect 5870 1097 5900 1183
rect 6370 1467 6400 1553
rect 6570 1467 6600 1553
rect 6670 1467 6700 1553
rect 6880 1467 6910 1553
rect 6980 1467 7010 1553
rect 7080 1467 7110 1553
rect 7180 1467 7210 1553
rect 7280 1467 7310 1553
rect 7380 1467 7410 1553
rect 6270 1327 6300 1413
rect 6370 1327 6400 1413
rect 6570 1327 6600 1413
rect 6670 1327 6700 1413
rect 6880 1327 6910 1413
rect 6980 1327 7010 1413
rect 7080 1327 7110 1413
rect 7180 1327 7210 1413
rect 7280 1327 7310 1413
rect 7380 1327 7410 1413
rect 6070 1097 6100 1183
rect 6170 1097 6200 1183
rect 6270 1097 6300 1183
rect 6370 1097 6400 1183
rect 6570 1097 6600 1183
rect 6670 1097 6700 1183
rect 6880 1097 6910 1183
rect 6980 1097 7010 1183
rect 7080 1097 7110 1183
rect 7180 1097 7210 1183
rect 7280 1097 7310 1183
rect 7380 1097 7410 1183
rect 5170 957 5200 1043
rect 5270 957 5300 1043
rect 5370 957 5400 1043
rect 5470 957 5500 1043
rect 5570 957 5600 1043
rect 5670 957 5700 1043
rect 5770 957 5800 1043
rect 5870 957 5900 1043
rect 5970 957 6000 1043
rect 6070 957 6100 1043
rect 6170 957 6200 1043
rect 6370 957 6400 1043
rect 6570 957 6600 1043
rect 6670 957 6700 1043
rect 6880 957 6910 1043
rect 6980 957 7010 1043
rect 7080 957 7110 1043
rect 7180 957 7210 1043
rect 7280 957 7310 1043
rect 7380 957 7410 1043
rect 4670 817 4700 903
rect 4770 817 4800 903
rect 4870 817 4900 903
rect 4970 817 5000 903
rect 5070 817 5100 903
rect 5170 817 5200 903
rect 5270 817 5300 903
rect 5370 817 5400 903
rect 5470 817 5500 903
rect 5570 817 5600 903
rect 5670 817 5700 903
rect 5770 817 5800 903
rect 5870 817 5900 903
rect 5970 817 6000 903
rect 6070 817 6100 903
rect 6170 817 6200 903
rect 6270 817 6300 903
rect 6370 817 6400 903
rect 6570 817 6600 903
rect 6670 817 6700 903
rect 6880 817 6910 903
rect 6980 817 7010 903
rect 7080 817 7110 903
rect 7180 817 7210 903
rect 7280 817 7310 903
rect 7380 817 7410 903
rect 4570 677 4600 763
rect 4670 677 4700 763
rect 4770 677 4800 763
rect 4870 677 4900 763
rect 4970 677 5000 763
rect 5070 677 5100 763
rect 5170 677 5200 763
rect 5270 677 5300 763
rect 5370 677 5400 763
rect 5470 677 5500 763
rect 4370 537 4400 623
rect 4470 537 4500 623
rect 4570 537 4600 623
rect 4770 537 4800 623
rect 4870 537 4900 623
rect 4970 537 5000 623
rect 5070 537 5100 623
rect 5170 537 5200 623
rect 5670 677 5700 763
rect 5870 677 5900 763
rect 5970 677 6000 763
rect 6070 677 6100 763
rect 6170 677 6200 763
rect 6270 677 6300 763
rect 6370 677 6400 763
rect 6570 677 6600 763
rect 6670 677 6700 763
rect 6880 677 6910 763
rect 6980 677 7010 763
rect 7080 677 7110 763
rect 7180 677 7210 763
rect 7280 677 7310 763
rect 7380 677 7410 763
rect 5370 537 5400 623
rect 5470 537 5500 623
rect 5570 537 5600 623
rect 5670 537 5700 623
rect 5770 537 5800 623
rect 5870 537 5900 623
rect 5970 537 6000 623
rect 3870 397 3900 483
rect 3970 397 4000 483
rect 4070 397 4100 483
rect 4170 397 4200 483
rect 4270 397 4300 483
rect 4370 397 4400 483
rect 4470 397 4500 483
rect 4570 397 4600 483
rect 4670 397 4700 483
rect 4770 397 4800 483
rect 4870 397 4900 483
rect 4970 397 5000 483
rect 5070 397 5100 483
rect 5170 397 5200 483
rect 5270 397 5300 483
rect 5370 397 5400 483
rect 5470 397 5500 483
rect 6170 537 6200 623
rect 6270 537 6300 623
rect 6370 537 6400 623
rect 6570 537 6600 623
rect 6670 537 6700 623
rect 6880 537 6910 623
rect 6980 537 7010 623
rect 7080 537 7110 623
rect 7180 537 7210 623
rect 7280 537 7310 623
rect 7380 537 7410 623
rect 5670 397 5700 483
rect 5770 397 5800 483
rect 5870 397 5900 483
rect 5970 397 6000 483
rect 6070 397 6100 483
rect 6170 397 6200 483
rect 3670 257 3700 343
rect 3770 257 3800 343
rect 3870 257 3900 343
rect 3970 257 4000 343
rect 4070 257 4100 343
rect 4170 257 4200 343
rect 4270 257 4300 343
rect 4370 257 4400 343
rect 4470 257 4500 343
rect 4570 257 4600 343
rect 4670 257 4700 343
rect 4770 257 4800 343
rect 4870 257 4900 343
rect 4970 257 5000 343
rect 5070 257 5100 343
rect 5170 257 5200 343
rect 5270 257 5300 343
rect 5370 257 5400 343
rect 5470 257 5500 343
rect 5570 257 5600 343
rect 3670 117 3700 203
rect 3770 117 3800 203
rect 3870 117 3900 203
rect 3970 117 4000 203
rect 4070 117 4100 203
rect 4170 117 4200 203
rect 4270 117 4300 203
rect 4370 117 4400 203
rect 4470 117 4500 203
rect 4570 117 4600 203
rect 4670 117 4700 203
rect 6370 397 6400 483
rect 6570 397 6600 483
rect 6670 397 6700 483
rect 6880 397 6910 483
rect 6980 397 7010 483
rect 7080 397 7110 483
rect 7180 397 7210 483
rect 7280 397 7310 483
rect 7380 397 7410 483
rect 5770 257 5800 343
rect 5870 257 5900 343
rect 5970 257 6000 343
rect 6070 257 6100 343
rect 6170 257 6200 343
rect 6270 257 6300 343
rect 6370 257 6400 343
rect 6570 257 6600 343
rect 6670 257 6700 343
rect 6880 257 6910 343
rect 6980 257 7010 343
rect 7080 257 7110 343
rect 7180 257 7210 343
rect 7280 257 7310 343
rect 7380 257 7410 343
rect 4870 117 4900 203
rect 4970 117 5000 203
rect 5070 117 5100 203
rect 5170 117 5200 203
rect 5270 117 5300 203
rect 5370 117 5400 203
rect 5470 117 5500 203
rect 5570 117 5600 203
rect 5670 117 5700 203
rect 5770 117 5800 203
rect 5870 117 5900 203
rect 5970 117 6000 203
rect 6070 117 6100 203
rect 6270 117 6300 203
rect 6370 117 6400 203
rect 6570 117 6600 203
rect 6670 117 6700 203
rect 6880 117 6910 203
rect 6980 117 7010 203
rect 7080 117 7110 203
rect 7180 117 7210 203
rect 7280 117 7310 203
rect 7380 117 7410 203
rect -10 -940 108 -910
rect 162 -940 280 -910
rect 390 -940 508 -910
rect 562 -940 680 -910
rect 790 -940 908 -910
rect 962 -940 1080 -910
rect 1190 -940 1308 -910
rect 1362 -940 1480 -910
rect -10 -1040 108 -1010
rect 162 -1040 280 -1010
rect 390 -1040 508 -1010
rect 562 -1040 680 -1010
rect 1590 -940 1708 -910
rect 1762 -940 1880 -910
rect 1990 -940 2108 -910
rect 2162 -940 2280 -910
rect 790 -1040 908 -1010
rect 962 -1040 1080 -1010
rect 1190 -1040 1308 -1010
rect 1362 -1040 1480 -1010
rect -10 -1140 108 -1110
rect 162 -1140 280 -1110
rect 390 -1140 508 -1110
rect 562 -1140 680 -1110
rect 2390 -940 2508 -910
rect 2562 -940 2680 -910
rect 2790 -940 2908 -910
rect 2962 -940 3080 -910
rect 1590 -1040 1708 -1010
rect 1762 -1040 1880 -1010
rect 1990 -1040 2108 -1010
rect 2162 -1040 2280 -1010
rect 790 -1140 908 -1110
rect 962 -1140 1080 -1110
rect 1190 -1140 1308 -1110
rect 1362 -1140 1480 -1110
rect -10 -1240 108 -1210
rect 162 -1240 280 -1210
rect 390 -1240 508 -1210
rect 562 -1240 680 -1210
rect 3190 -940 3308 -910
rect 3362 -940 3480 -910
rect 3590 -940 3708 -910
rect 3762 -940 3880 -910
rect 2390 -1040 2508 -1010
rect 2562 -1040 2680 -1010
rect 2790 -1040 2908 -1010
rect 2962 -1040 3080 -1010
rect 1590 -1140 1708 -1110
rect 1762 -1140 1880 -1110
rect 1990 -1140 2108 -1110
rect 2162 -1140 2280 -1110
rect 790 -1240 908 -1210
rect 962 -1240 1080 -1210
rect 1190 -1240 1308 -1210
rect 1362 -1240 1480 -1210
rect -10 -1340 108 -1310
rect 162 -1340 280 -1310
rect 390 -1340 508 -1310
rect 562 -1340 680 -1310
rect 3990 -940 4108 -910
rect 4162 -940 4280 -910
rect 4390 -940 4508 -910
rect 4562 -940 4680 -910
rect 3190 -1040 3308 -1010
rect 3362 -1040 3480 -1010
rect 3590 -1040 3708 -1010
rect 3762 -1040 3880 -1010
rect 2390 -1140 2508 -1110
rect 2562 -1140 2680 -1110
rect 2790 -1140 2908 -1110
rect 2962 -1140 3080 -1110
rect 1590 -1240 1708 -1210
rect 1762 -1240 1880 -1210
rect 1990 -1240 2108 -1210
rect 2162 -1240 2280 -1210
rect 790 -1340 908 -1310
rect 962 -1340 1080 -1310
rect 1190 -1340 1308 -1310
rect 1362 -1340 1480 -1310
rect -10 -1440 108 -1410
rect 162 -1440 280 -1410
rect 390 -1440 508 -1410
rect 562 -1440 680 -1410
rect 4790 -940 4908 -910
rect 4962 -940 5080 -910
rect 5190 -940 5308 -910
rect 5362 -940 5480 -910
rect 3990 -1040 4108 -1010
rect 4162 -1040 4280 -1010
rect 4390 -1040 4508 -1010
rect 4562 -1040 4680 -1010
rect 3190 -1140 3308 -1110
rect 3362 -1140 3480 -1110
rect 3590 -1140 3708 -1110
rect 3762 -1140 3880 -1110
rect 2390 -1240 2508 -1210
rect 2562 -1240 2680 -1210
rect 2790 -1240 2908 -1210
rect 2962 -1240 3080 -1210
rect 1590 -1340 1708 -1310
rect 1762 -1340 1880 -1310
rect 1990 -1340 2108 -1310
rect 2162 -1340 2280 -1310
rect 790 -1440 908 -1410
rect 962 -1440 1080 -1410
rect 1190 -1440 1308 -1410
rect 1362 -1440 1480 -1410
rect -10 -1540 108 -1510
rect 162 -1540 280 -1510
rect 390 -1540 508 -1510
rect 562 -1540 680 -1510
rect 5590 -940 5708 -910
rect 5762 -940 5880 -910
rect 5990 -940 6108 -910
rect 6162 -940 6280 -910
rect 4790 -1040 4908 -1010
rect 4962 -1040 5080 -1010
rect 5190 -1040 5308 -1010
rect 5362 -1040 5480 -1010
rect 3990 -1140 4108 -1110
rect 4162 -1140 4280 -1110
rect 4390 -1140 4508 -1110
rect 4562 -1140 4680 -1110
rect 3190 -1240 3308 -1210
rect 3362 -1240 3480 -1210
rect 3590 -1240 3708 -1210
rect 3762 -1240 3880 -1210
rect 2390 -1340 2508 -1310
rect 2562 -1340 2680 -1310
rect 2790 -1340 2908 -1310
rect 2962 -1340 3080 -1310
rect 1590 -1440 1708 -1410
rect 1762 -1440 1880 -1410
rect 1990 -1440 2108 -1410
rect 2162 -1440 2280 -1410
rect 790 -1540 908 -1510
rect 962 -1540 1080 -1510
rect 1190 -1540 1308 -1510
rect 1362 -1540 1480 -1510
rect -10 -1640 108 -1610
rect 162 -1640 280 -1610
rect 390 -1640 508 -1610
rect 562 -1640 680 -1610
rect 5590 -1040 5708 -1010
rect 5762 -1040 5880 -1010
rect 5990 -1040 6108 -1010
rect 6162 -1040 6280 -1010
rect 4790 -1140 4908 -1110
rect 4962 -1140 5080 -1110
rect 5190 -1140 5308 -1110
rect 5362 -1140 5480 -1110
rect 3990 -1240 4108 -1210
rect 4162 -1240 4280 -1210
rect 4390 -1240 4508 -1210
rect 4562 -1240 4680 -1210
rect 3190 -1340 3308 -1310
rect 3362 -1340 3480 -1310
rect 3590 -1340 3708 -1310
rect 3762 -1340 3880 -1310
rect 2390 -1440 2508 -1410
rect 2562 -1440 2680 -1410
rect 2790 -1440 2908 -1410
rect 2962 -1440 3080 -1410
rect 1590 -1540 1708 -1510
rect 1762 -1540 1880 -1510
rect 1990 -1540 2108 -1510
rect 2162 -1540 2280 -1510
rect 790 -1640 908 -1610
rect 962 -1640 1080 -1610
rect 1190 -1640 1308 -1610
rect 1362 -1640 1480 -1610
rect -10 -1740 108 -1710
rect 162 -1740 280 -1710
rect 390 -1740 508 -1710
rect 562 -1740 680 -1710
rect 5590 -1140 5708 -1110
rect 5762 -1140 5880 -1110
rect 5990 -1140 6108 -1110
rect 6162 -1140 6280 -1110
rect 4790 -1240 4908 -1210
rect 4962 -1240 5080 -1210
rect 5190 -1240 5308 -1210
rect 5362 -1240 5480 -1210
rect 3990 -1340 4108 -1310
rect 4162 -1340 4280 -1310
rect 4390 -1340 4508 -1310
rect 4562 -1340 4680 -1310
rect 3190 -1440 3308 -1410
rect 3362 -1440 3480 -1410
rect 3590 -1440 3708 -1410
rect 3762 -1440 3880 -1410
rect 2390 -1540 2508 -1510
rect 2562 -1540 2680 -1510
rect 2790 -1540 2908 -1510
rect 2962 -1540 3080 -1510
rect 1590 -1640 1708 -1610
rect 1762 -1640 1880 -1610
rect 1990 -1640 2108 -1610
rect 2162 -1640 2280 -1610
rect 790 -1740 908 -1710
rect 962 -1740 1080 -1710
rect 1190 -1740 1308 -1710
rect 1362 -1740 1480 -1710
rect -10 -1840 108 -1810
rect 162 -1840 280 -1810
rect 390 -1840 508 -1810
rect 562 -1840 680 -1810
rect 5590 -1240 5708 -1210
rect 5762 -1240 5880 -1210
rect 5990 -1240 6108 -1210
rect 6162 -1240 6280 -1210
rect 4790 -1340 4908 -1310
rect 4962 -1340 5080 -1310
rect 5190 -1340 5308 -1310
rect 5362 -1340 5480 -1310
rect 3990 -1440 4108 -1410
rect 4162 -1440 4280 -1410
rect 4390 -1440 4508 -1410
rect 4562 -1440 4680 -1410
rect 3190 -1540 3308 -1510
rect 3362 -1540 3480 -1510
rect 3590 -1540 3708 -1510
rect 3762 -1540 3880 -1510
rect 2390 -1640 2508 -1610
rect 2562 -1640 2680 -1610
rect 2790 -1640 2908 -1610
rect 2962 -1640 3080 -1610
rect 1590 -1740 1708 -1710
rect 1762 -1740 1880 -1710
rect 1990 -1740 2108 -1710
rect 2162 -1740 2280 -1710
rect 790 -1840 908 -1810
rect 962 -1840 1080 -1810
rect 1190 -1840 1308 -1810
rect 1362 -1840 1480 -1810
rect 5590 -1340 5708 -1310
rect 5762 -1340 5880 -1310
rect 5990 -1340 6108 -1310
rect 6162 -1340 6280 -1310
rect 4790 -1440 4908 -1410
rect 4962 -1440 5080 -1410
rect 5190 -1440 5308 -1410
rect 5362 -1440 5480 -1410
rect 3990 -1540 4108 -1510
rect 4162 -1540 4280 -1510
rect 4390 -1540 4508 -1510
rect 4562 -1540 4680 -1510
rect 3190 -1640 3308 -1610
rect 3362 -1640 3480 -1610
rect 3590 -1640 3708 -1610
rect 3762 -1640 3880 -1610
rect 2390 -1740 2508 -1710
rect 2562 -1740 2680 -1710
rect 2790 -1740 2908 -1710
rect 2962 -1740 3080 -1710
rect 1590 -1840 1708 -1810
rect 1762 -1840 1880 -1810
rect 1990 -1840 2108 -1810
rect 2162 -1840 2280 -1810
rect 5590 -1440 5708 -1410
rect 5762 -1440 5880 -1410
rect 5990 -1440 6108 -1410
rect 6162 -1440 6280 -1410
rect 4790 -1540 4908 -1510
rect 4962 -1540 5080 -1510
rect 5190 -1540 5308 -1510
rect 5362 -1540 5480 -1510
rect 3990 -1640 4108 -1610
rect 4162 -1640 4280 -1610
rect 4390 -1640 4508 -1610
rect 4562 -1640 4680 -1610
rect 3190 -1740 3308 -1710
rect 3362 -1740 3480 -1710
rect 3590 -1740 3708 -1710
rect 3762 -1740 3880 -1710
rect 2390 -1840 2508 -1810
rect 2562 -1840 2680 -1810
rect 2790 -1840 2908 -1810
rect 2962 -1840 3080 -1810
rect 5590 -1540 5708 -1510
rect 5762 -1540 5880 -1510
rect 5990 -1540 6108 -1510
rect 6162 -1540 6280 -1510
rect 4790 -1640 4908 -1610
rect 4962 -1640 5080 -1610
rect 5190 -1640 5308 -1610
rect 5362 -1640 5480 -1610
rect 3990 -1740 4108 -1710
rect 4162 -1740 4280 -1710
rect 4390 -1740 4508 -1710
rect 4562 -1740 4680 -1710
rect 3190 -1840 3308 -1810
rect 3362 -1840 3480 -1810
rect 3590 -1840 3708 -1810
rect 3762 -1840 3880 -1810
rect 5590 -1640 5708 -1610
rect 5762 -1640 5880 -1610
rect 5990 -1640 6108 -1610
rect 6162 -1640 6280 -1610
rect 4790 -1740 4908 -1710
rect 4962 -1740 5080 -1710
rect 5190 -1740 5308 -1710
rect 5362 -1740 5480 -1710
rect 3990 -1840 4108 -1810
rect 4162 -1840 4280 -1810
rect 4390 -1840 4508 -1810
rect 4562 -1840 4680 -1810
rect 5590 -1740 5708 -1710
rect 5762 -1740 5880 -1710
rect 5990 -1740 6108 -1710
rect 6162 -1740 6280 -1710
rect 4790 -1840 4908 -1810
rect 4962 -1840 5080 -1810
rect 5190 -1840 5308 -1810
rect 5362 -1840 5480 -1810
rect 5590 -1840 5708 -1810
rect 5762 -1840 5880 -1810
rect 5990 -1840 6108 -1810
rect 6162 -1840 6280 -1810
<< ndiff >>
rect 16 9707 70 9793
rect 100 9767 170 9793
rect 100 9733 118 9767
rect 152 9733 170 9767
rect 100 9707 170 9733
rect 200 9767 270 9793
rect 200 9733 218 9767
rect 252 9733 270 9767
rect 200 9707 270 9733
rect 300 9707 370 9793
rect 400 9707 470 9793
rect 500 9767 570 9793
rect 500 9733 518 9767
rect 552 9733 570 9767
rect 500 9707 570 9733
rect 600 9767 670 9793
rect 600 9733 618 9767
rect 652 9733 670 9767
rect 600 9707 670 9733
rect 700 9707 770 9793
rect 800 9707 870 9793
rect 900 9767 970 9793
rect 900 9733 918 9767
rect 952 9733 970 9767
rect 900 9707 970 9733
rect 1000 9767 1070 9793
rect 1000 9733 1018 9767
rect 1052 9733 1070 9767
rect 1000 9707 1070 9733
rect 1100 9767 1170 9793
rect 1100 9733 1118 9767
rect 1152 9733 1170 9767
rect 1100 9707 1170 9733
rect 1200 9707 1270 9793
rect 1300 9707 1370 9793
rect 1400 9767 1470 9793
rect 1400 9733 1418 9767
rect 1452 9733 1470 9767
rect 1400 9707 1470 9733
rect 1500 9767 1554 9793
rect 1500 9733 1512 9767
rect 1546 9733 1554 9767
rect 1500 9707 1554 9733
rect 16 9567 70 9653
rect 100 9567 170 9653
rect 200 9627 270 9653
rect 200 9593 218 9627
rect 252 9593 270 9627
rect 200 9567 270 9593
rect 300 9627 370 9653
rect 300 9593 318 9627
rect 352 9593 370 9627
rect 300 9567 370 9593
rect 400 9567 470 9653
rect 500 9627 570 9653
rect 500 9593 518 9627
rect 552 9593 570 9627
rect 500 9567 570 9593
rect 600 9627 654 9653
rect 600 9593 612 9627
rect 646 9593 654 9627
rect 600 9567 654 9593
rect 16 9427 70 9513
rect 100 9487 170 9513
rect 100 9453 118 9487
rect 152 9453 170 9487
rect 100 9427 170 9453
rect 200 9487 270 9513
rect 200 9453 218 9487
rect 252 9453 270 9487
rect 200 9427 270 9453
rect 300 9487 370 9513
rect 300 9453 318 9487
rect 352 9453 370 9487
rect 300 9427 370 9453
rect 400 9487 454 9513
rect 400 9453 412 9487
rect 446 9453 454 9487
rect 400 9427 454 9453
rect 1616 9767 1670 9793
rect 1616 9733 1624 9767
rect 1658 9733 1670 9767
rect 1616 9707 1670 9733
rect 1700 9767 1770 9793
rect 1700 9733 1718 9767
rect 1752 9733 1770 9767
rect 1700 9707 1770 9733
rect 1800 9707 1870 9793
rect 1900 9767 1970 9793
rect 1900 9733 1918 9767
rect 1952 9733 1970 9767
rect 1900 9707 1970 9733
rect 2000 9767 2070 9793
rect 2000 9733 2018 9767
rect 2052 9733 2070 9767
rect 2000 9707 2070 9733
rect 2100 9767 2154 9793
rect 2100 9733 2112 9767
rect 2146 9733 2154 9767
rect 2100 9707 2154 9733
rect 716 9627 770 9653
rect 716 9593 724 9627
rect 758 9593 770 9627
rect 716 9567 770 9593
rect 800 9627 870 9653
rect 800 9593 818 9627
rect 852 9593 870 9627
rect 800 9567 870 9593
rect 900 9567 970 9653
rect 1000 9567 1070 9653
rect 1100 9567 1170 9653
rect 1200 9627 1270 9653
rect 1200 9593 1218 9627
rect 1252 9593 1270 9627
rect 1200 9567 1270 9593
rect 1300 9627 1370 9653
rect 1300 9593 1318 9627
rect 1352 9593 1370 9627
rect 1300 9567 1370 9593
rect 1400 9627 1470 9653
rect 1400 9593 1418 9627
rect 1452 9593 1470 9627
rect 1400 9567 1470 9593
rect 1500 9627 1570 9653
rect 1500 9593 1518 9627
rect 1552 9593 1570 9627
rect 1500 9567 1570 9593
rect 1600 9627 1670 9653
rect 1600 9593 1618 9627
rect 1652 9593 1670 9627
rect 1600 9567 1670 9593
rect 1700 9627 1770 9653
rect 1700 9593 1718 9627
rect 1752 9593 1770 9627
rect 1700 9567 1770 9593
rect 1800 9567 1870 9653
rect 1900 9567 1970 9653
rect 2000 9627 2070 9653
rect 2000 9593 2018 9627
rect 2052 9593 2070 9627
rect 2000 9567 2070 9593
rect 2100 9627 2154 9653
rect 2100 9593 2112 9627
rect 2146 9593 2154 9627
rect 2100 9567 2154 9593
rect 516 9487 570 9513
rect 516 9453 524 9487
rect 558 9453 570 9487
rect 516 9427 570 9453
rect 600 9487 670 9513
rect 600 9453 618 9487
rect 652 9453 670 9487
rect 600 9427 670 9453
rect 700 9487 770 9513
rect 700 9453 718 9487
rect 752 9453 770 9487
rect 700 9427 770 9453
rect 800 9487 870 9513
rect 800 9453 818 9487
rect 852 9453 870 9487
rect 800 9427 870 9453
rect 900 9487 954 9513
rect 900 9453 912 9487
rect 946 9453 954 9487
rect 900 9427 954 9453
rect 1016 9487 1070 9513
rect 1016 9453 1024 9487
rect 1058 9453 1070 9487
rect 1016 9427 1070 9453
rect 1100 9487 1154 9513
rect 1100 9453 1112 9487
rect 1146 9453 1154 9487
rect 1100 9427 1154 9453
rect 1216 9487 1270 9513
rect 1216 9453 1224 9487
rect 1258 9453 1270 9487
rect 1216 9427 1270 9453
rect 1300 9487 1370 9513
rect 1300 9453 1318 9487
rect 1352 9453 1370 9487
rect 1300 9427 1370 9453
rect 1400 9427 1470 9513
rect 1500 9427 1570 9513
rect 1600 9487 1670 9513
rect 1600 9453 1618 9487
rect 1652 9453 1670 9487
rect 1600 9427 1670 9453
rect 1700 9487 1754 9513
rect 1700 9453 1712 9487
rect 1746 9453 1754 9487
rect 1700 9427 1754 9453
rect 16 9287 70 9373
rect 100 9287 170 9373
rect 200 9287 270 9373
rect 300 9287 370 9373
rect 400 9347 470 9373
rect 400 9313 418 9347
rect 452 9313 470 9347
rect 400 9287 470 9313
rect 500 9347 570 9373
rect 500 9313 518 9347
rect 552 9313 570 9347
rect 500 9287 570 9313
rect 600 9347 670 9373
rect 600 9313 618 9347
rect 652 9313 670 9347
rect 600 9287 670 9313
rect 700 9347 770 9373
rect 700 9313 718 9347
rect 752 9313 770 9347
rect 700 9287 770 9313
rect 800 9287 870 9373
rect 900 9347 970 9373
rect 900 9313 918 9347
rect 952 9313 970 9347
rect 900 9287 970 9313
rect 1000 9347 1070 9373
rect 1000 9313 1018 9347
rect 1052 9313 1070 9347
rect 1000 9287 1070 9313
rect 1100 9347 1170 9373
rect 1100 9313 1118 9347
rect 1152 9313 1170 9347
rect 1100 9287 1170 9313
rect 1200 9347 1270 9373
rect 1200 9313 1218 9347
rect 1252 9313 1270 9347
rect 1200 9287 1270 9313
rect 1300 9287 1370 9373
rect 1400 9287 1470 9373
rect 1500 9347 1570 9373
rect 1500 9313 1518 9347
rect 1552 9313 1570 9347
rect 1500 9287 1570 9313
rect 1600 9347 1670 9373
rect 1600 9313 1618 9347
rect 1652 9313 1670 9347
rect 1600 9287 1670 9313
rect 1700 9347 1754 9373
rect 1700 9313 1712 9347
rect 1746 9313 1754 9347
rect 1700 9287 1754 9313
rect 16 9207 70 9233
rect 16 9173 24 9207
rect 58 9173 70 9207
rect 16 9147 70 9173
rect 100 9207 170 9233
rect 100 9173 118 9207
rect 152 9173 170 9207
rect 100 9147 170 9173
rect 200 9207 270 9233
rect 200 9173 218 9207
rect 252 9173 270 9207
rect 200 9147 270 9173
rect 300 9207 370 9233
rect 300 9173 318 9207
rect 352 9173 370 9207
rect 300 9147 370 9173
rect 400 9207 470 9233
rect 400 9173 418 9207
rect 452 9173 470 9207
rect 400 9147 470 9173
rect 500 9147 570 9233
rect 600 9207 670 9233
rect 600 9173 618 9207
rect 652 9173 670 9207
rect 600 9147 670 9173
rect 700 9207 770 9233
rect 700 9173 718 9207
rect 752 9173 770 9207
rect 700 9147 770 9173
rect 800 9207 870 9233
rect 800 9173 818 9207
rect 852 9173 870 9207
rect 800 9147 870 9173
rect 900 9207 970 9233
rect 900 9173 918 9207
rect 952 9173 970 9207
rect 900 9147 970 9173
rect 1000 9207 1070 9233
rect 1000 9173 1018 9207
rect 1052 9173 1070 9207
rect 1000 9147 1070 9173
rect 1100 9147 1170 9233
rect 1200 9207 1270 9233
rect 1200 9173 1218 9207
rect 1252 9173 1270 9207
rect 1200 9147 1270 9173
rect 1300 9207 1370 9233
rect 1300 9173 1318 9207
rect 1352 9173 1370 9207
rect 1300 9147 1370 9173
rect 1400 9207 1470 9233
rect 1400 9173 1418 9207
rect 1452 9173 1470 9207
rect 1400 9147 1470 9173
rect 1500 9207 1554 9233
rect 1500 9173 1512 9207
rect 1546 9173 1554 9207
rect 1500 9147 1554 9173
rect 16 9007 70 9093
rect 100 9067 170 9093
rect 100 9033 118 9067
rect 152 9033 170 9067
rect 100 9007 170 9033
rect 200 9067 270 9093
rect 200 9033 218 9067
rect 252 9033 270 9067
rect 200 9007 270 9033
rect 300 9007 370 9093
rect 400 9007 470 9093
rect 500 9067 570 9093
rect 500 9033 518 9067
rect 552 9033 570 9067
rect 500 9007 570 9033
rect 600 9067 654 9093
rect 600 9033 612 9067
rect 646 9033 654 9067
rect 600 9007 654 9033
rect 1816 9487 1870 9513
rect 1816 9453 1824 9487
rect 1858 9453 1870 9487
rect 1816 9427 1870 9453
rect 1900 9487 1970 9513
rect 1900 9453 1918 9487
rect 1952 9453 1970 9487
rect 1900 9427 1970 9453
rect 2000 9487 2054 9513
rect 2000 9453 2012 9487
rect 2046 9453 2054 9487
rect 2000 9427 2054 9453
rect 2216 9767 2270 9793
rect 2216 9733 2224 9767
rect 2258 9733 2270 9767
rect 2216 9707 2270 9733
rect 2300 9767 2370 9793
rect 2300 9733 2318 9767
rect 2352 9733 2370 9767
rect 2300 9707 2370 9733
rect 2400 9707 2470 9793
rect 2500 9707 2570 9793
rect 2600 9767 2670 9793
rect 2600 9733 2618 9767
rect 2652 9733 2670 9767
rect 2600 9707 2670 9733
rect 2700 9767 2754 9793
rect 2700 9733 2712 9767
rect 2746 9733 2754 9767
rect 2700 9707 2754 9733
rect 2216 9627 2270 9653
rect 2216 9593 2224 9627
rect 2258 9593 2270 9627
rect 2216 9567 2270 9593
rect 2300 9627 2354 9653
rect 2300 9593 2312 9627
rect 2346 9593 2354 9627
rect 2300 9567 2354 9593
rect 2116 9487 2170 9513
rect 2116 9453 2124 9487
rect 2158 9453 2170 9487
rect 2116 9427 2170 9453
rect 2200 9487 2270 9513
rect 2200 9453 2218 9487
rect 2252 9453 2270 9487
rect 2200 9427 2270 9453
rect 2300 9487 2354 9513
rect 2300 9453 2312 9487
rect 2346 9453 2354 9487
rect 2300 9427 2354 9453
rect 2816 9767 2870 9793
rect 2816 9733 2824 9767
rect 2858 9733 2870 9767
rect 2816 9707 2870 9733
rect 2900 9767 2970 9793
rect 2900 9733 2918 9767
rect 2952 9733 2970 9767
rect 2900 9707 2970 9733
rect 3000 9707 3070 9793
rect 3100 9767 3170 9793
rect 3100 9733 3118 9767
rect 3152 9733 3170 9767
rect 3100 9707 3170 9733
rect 3200 9767 3254 9793
rect 3200 9733 3212 9767
rect 3246 9733 3254 9767
rect 3200 9707 3254 9733
rect 2416 9627 2470 9653
rect 2416 9593 2424 9627
rect 2458 9593 2470 9627
rect 2416 9567 2470 9593
rect 2500 9627 2570 9653
rect 2500 9593 2518 9627
rect 2552 9593 2570 9627
rect 2500 9567 2570 9593
rect 2600 9567 2670 9653
rect 2700 9567 2770 9653
rect 2800 9627 2870 9653
rect 2800 9593 2818 9627
rect 2852 9593 2870 9627
rect 2800 9567 2870 9593
rect 2900 9627 2954 9653
rect 2900 9593 2912 9627
rect 2946 9593 2954 9627
rect 2900 9567 2954 9593
rect 2416 9487 2470 9513
rect 2416 9453 2424 9487
rect 2458 9453 2470 9487
rect 2416 9427 2470 9453
rect 2500 9487 2554 9513
rect 2500 9453 2512 9487
rect 2546 9453 2554 9487
rect 2500 9427 2554 9453
rect 2616 9487 2670 9513
rect 2616 9453 2624 9487
rect 2658 9453 2670 9487
rect 2616 9427 2670 9453
rect 2700 9487 2754 9513
rect 2700 9453 2712 9487
rect 2746 9453 2754 9487
rect 2700 9427 2754 9453
rect 3316 9767 3370 9793
rect 3316 9733 3324 9767
rect 3358 9733 3370 9767
rect 3316 9707 3370 9733
rect 3400 9767 3470 9793
rect 3400 9733 3418 9767
rect 3452 9733 3470 9767
rect 3400 9707 3470 9733
rect 3500 9767 3554 9793
rect 3500 9733 3512 9767
rect 3546 9733 3554 9767
rect 3500 9707 3554 9733
rect 3616 9767 3670 9793
rect 3616 9733 3624 9767
rect 3658 9733 3670 9767
rect 3616 9707 3670 9733
rect 3700 9767 3770 9793
rect 3700 9733 3718 9767
rect 3752 9733 3770 9767
rect 3700 9707 3770 9733
rect 3800 9767 3870 9793
rect 3800 9733 3818 9767
rect 3852 9733 3870 9767
rect 3800 9707 3870 9733
rect 3900 9707 3970 9793
rect 4000 9767 4070 9793
rect 4000 9733 4018 9767
rect 4052 9733 4070 9767
rect 4000 9707 4070 9733
rect 4100 9767 4170 9793
rect 4100 9733 4118 9767
rect 4152 9733 4170 9767
rect 4100 9707 4170 9733
rect 4200 9767 4270 9793
rect 4200 9733 4218 9767
rect 4252 9733 4270 9767
rect 4200 9707 4270 9733
rect 4300 9707 4370 9793
rect 4400 9707 4470 9793
rect 4500 9707 4570 9793
rect 4600 9707 4670 9793
rect 4700 9707 4770 9793
rect 4800 9767 4870 9793
rect 4800 9733 4818 9767
rect 4852 9733 4870 9767
rect 4800 9707 4870 9733
rect 4900 9767 4970 9793
rect 4900 9733 4918 9767
rect 4952 9733 4970 9767
rect 4900 9707 4970 9733
rect 5000 9707 5070 9793
rect 5100 9707 5170 9793
rect 5200 9707 5270 9793
rect 5300 9767 5370 9793
rect 5300 9733 5318 9767
rect 5352 9733 5370 9767
rect 5300 9707 5370 9733
rect 5400 9767 5454 9793
rect 5400 9733 5412 9767
rect 5446 9733 5454 9767
rect 5400 9707 5454 9733
rect 3016 9627 3070 9653
rect 3016 9593 3024 9627
rect 3058 9593 3070 9627
rect 3016 9567 3070 9593
rect 3100 9627 3170 9653
rect 3100 9593 3118 9627
rect 3152 9593 3170 9627
rect 3100 9567 3170 9593
rect 3200 9627 3270 9653
rect 3200 9593 3218 9627
rect 3252 9593 3270 9627
rect 3200 9567 3270 9593
rect 3300 9627 3370 9653
rect 3300 9593 3318 9627
rect 3352 9593 3370 9627
rect 3300 9567 3370 9593
rect 3400 9627 3470 9653
rect 3400 9593 3418 9627
rect 3452 9593 3470 9627
rect 3400 9567 3470 9593
rect 3500 9627 3570 9653
rect 3500 9593 3518 9627
rect 3552 9593 3570 9627
rect 3500 9567 3570 9593
rect 3600 9627 3670 9653
rect 3600 9593 3618 9627
rect 3652 9593 3670 9627
rect 3600 9567 3670 9593
rect 3700 9567 3770 9653
rect 3800 9567 3870 9653
rect 3900 9627 3970 9653
rect 3900 9593 3918 9627
rect 3952 9593 3970 9627
rect 3900 9567 3970 9593
rect 4000 9627 4054 9653
rect 4000 9593 4012 9627
rect 4046 9593 4054 9627
rect 4000 9567 4054 9593
rect 2816 9487 2870 9513
rect 2816 9453 2824 9487
rect 2858 9453 2870 9487
rect 2816 9427 2870 9453
rect 2900 9487 2970 9513
rect 2900 9453 2918 9487
rect 2952 9453 2970 9487
rect 2900 9427 2970 9453
rect 3000 9427 3070 9513
rect 3100 9427 3170 9513
rect 3200 9427 3270 9513
rect 3300 9427 3370 9513
rect 3400 9487 3470 9513
rect 3400 9453 3418 9487
rect 3452 9453 3470 9487
rect 3400 9427 3470 9453
rect 3500 9487 3570 9513
rect 3500 9453 3518 9487
rect 3552 9453 3570 9487
rect 3500 9427 3570 9453
rect 3600 9487 3670 9513
rect 3600 9453 3618 9487
rect 3652 9453 3670 9487
rect 3600 9427 3670 9453
rect 3700 9427 3770 9513
rect 3800 9487 3870 9513
rect 3800 9453 3818 9487
rect 3852 9453 3870 9487
rect 3800 9427 3870 9453
rect 3900 9487 3970 9513
rect 3900 9453 3918 9487
rect 3952 9453 3970 9487
rect 3900 9427 3970 9453
rect 4000 9487 4054 9513
rect 4000 9453 4012 9487
rect 4046 9453 4054 9487
rect 4000 9427 4054 9453
rect 5516 9767 5570 9793
rect 5516 9733 5524 9767
rect 5558 9733 5570 9767
rect 5516 9707 5570 9733
rect 5600 9767 5670 9793
rect 5600 9733 5618 9767
rect 5652 9733 5670 9767
rect 5600 9707 5670 9733
rect 5700 9767 5754 9793
rect 5700 9733 5712 9767
rect 5746 9733 5754 9767
rect 5700 9707 5754 9733
rect 5816 9767 5870 9793
rect 5816 9733 5824 9767
rect 5858 9733 5870 9767
rect 5816 9707 5870 9733
rect 5900 9767 5954 9793
rect 5900 9733 5912 9767
rect 5946 9733 5954 9767
rect 5900 9707 5954 9733
rect 4116 9627 4170 9653
rect 4116 9593 4124 9627
rect 4158 9593 4170 9627
rect 4116 9567 4170 9593
rect 4200 9627 4270 9653
rect 4200 9593 4218 9627
rect 4252 9593 4270 9627
rect 4200 9567 4270 9593
rect 4300 9627 4370 9653
rect 4300 9593 4318 9627
rect 4352 9593 4370 9627
rect 4300 9567 4370 9593
rect 4400 9567 4470 9653
rect 4500 9567 4570 9653
rect 4600 9627 4670 9653
rect 4600 9593 4618 9627
rect 4652 9593 4670 9627
rect 4600 9567 4670 9593
rect 4700 9627 4770 9653
rect 4700 9593 4718 9627
rect 4752 9593 4770 9627
rect 4700 9567 4770 9593
rect 4800 9627 4870 9653
rect 4800 9593 4818 9627
rect 4852 9593 4870 9627
rect 4800 9567 4870 9593
rect 4900 9627 4970 9653
rect 4900 9593 4918 9627
rect 4952 9593 4970 9627
rect 4900 9567 4970 9593
rect 5000 9567 5070 9653
rect 5100 9567 5170 9653
rect 5200 9567 5270 9653
rect 5300 9567 5370 9653
rect 5400 9567 5470 9653
rect 5500 9627 5570 9653
rect 5500 9593 5518 9627
rect 5552 9593 5570 9627
rect 5500 9567 5570 9593
rect 5600 9627 5670 9653
rect 5600 9593 5618 9627
rect 5652 9593 5670 9627
rect 5600 9567 5670 9593
rect 5700 9627 5770 9653
rect 5700 9593 5718 9627
rect 5752 9593 5770 9627
rect 5700 9567 5770 9593
rect 5800 9627 5870 9653
rect 5800 9593 5818 9627
rect 5852 9593 5870 9627
rect 5800 9567 5870 9593
rect 5900 9627 5954 9653
rect 5900 9593 5912 9627
rect 5946 9593 5954 9627
rect 5900 9567 5954 9593
rect 4116 9487 4170 9513
rect 4116 9453 4124 9487
rect 4158 9453 4170 9487
rect 4116 9427 4170 9453
rect 4200 9487 4270 9513
rect 4200 9453 4218 9487
rect 4252 9453 4270 9487
rect 4200 9427 4270 9453
rect 4300 9487 4370 9513
rect 4300 9453 4318 9487
rect 4352 9453 4370 9487
rect 4300 9427 4370 9453
rect 4400 9487 4470 9513
rect 4400 9453 4418 9487
rect 4452 9453 4470 9487
rect 4400 9427 4470 9453
rect 4500 9487 4554 9513
rect 4500 9453 4512 9487
rect 4546 9453 4554 9487
rect 4500 9427 4554 9453
rect 1816 9347 1870 9373
rect 1816 9313 1824 9347
rect 1858 9313 1870 9347
rect 1816 9287 1870 9313
rect 1900 9347 1970 9373
rect 1900 9313 1918 9347
rect 1952 9313 1970 9347
rect 1900 9287 1970 9313
rect 2000 9347 2070 9373
rect 2000 9313 2018 9347
rect 2052 9313 2070 9347
rect 2000 9287 2070 9313
rect 2100 9287 2170 9373
rect 2200 9287 2270 9373
rect 2300 9287 2370 9373
rect 2400 9287 2470 9373
rect 2500 9287 2570 9373
rect 2600 9287 2670 9373
rect 2700 9347 2770 9373
rect 2700 9313 2718 9347
rect 2752 9313 2770 9347
rect 2700 9287 2770 9313
rect 2800 9347 2870 9373
rect 2800 9313 2818 9347
rect 2852 9313 2870 9347
rect 2800 9287 2870 9313
rect 2900 9347 2970 9373
rect 2900 9313 2918 9347
rect 2952 9313 2970 9347
rect 2900 9287 2970 9313
rect 3000 9287 3070 9373
rect 3100 9287 3170 9373
rect 3200 9347 3270 9373
rect 3200 9313 3218 9347
rect 3252 9313 3270 9347
rect 3200 9287 3270 9313
rect 3300 9347 3370 9373
rect 3300 9313 3318 9347
rect 3352 9313 3370 9347
rect 3300 9287 3370 9313
rect 3400 9287 3470 9373
rect 3500 9347 3570 9373
rect 3500 9313 3518 9347
rect 3552 9313 3570 9347
rect 3500 9287 3570 9313
rect 3600 9347 3670 9373
rect 3600 9313 3618 9347
rect 3652 9313 3670 9347
rect 3600 9287 3670 9313
rect 3700 9347 3770 9373
rect 3700 9313 3718 9347
rect 3752 9313 3770 9347
rect 3700 9287 3770 9313
rect 3800 9347 3870 9373
rect 3800 9313 3818 9347
rect 3852 9313 3870 9347
rect 3800 9287 3870 9313
rect 3900 9287 3970 9373
rect 4000 9347 4070 9373
rect 4000 9313 4018 9347
rect 4052 9313 4070 9347
rect 4000 9287 4070 9313
rect 4100 9347 4154 9373
rect 4100 9313 4112 9347
rect 4146 9313 4154 9347
rect 4100 9287 4154 9313
rect 1616 9207 1670 9233
rect 1616 9173 1624 9207
rect 1658 9173 1670 9207
rect 1616 9147 1670 9173
rect 1700 9207 1770 9233
rect 1700 9173 1718 9207
rect 1752 9173 1770 9207
rect 1700 9147 1770 9173
rect 1800 9207 1870 9233
rect 1800 9173 1818 9207
rect 1852 9173 1870 9207
rect 1800 9147 1870 9173
rect 1900 9147 1970 9233
rect 2000 9207 2070 9233
rect 2000 9173 2018 9207
rect 2052 9173 2070 9207
rect 2000 9147 2070 9173
rect 2100 9207 2170 9233
rect 2100 9173 2118 9207
rect 2152 9173 2170 9207
rect 2100 9147 2170 9173
rect 2200 9207 2270 9233
rect 2200 9173 2218 9207
rect 2252 9173 2270 9207
rect 2200 9147 2270 9173
rect 2300 9207 2370 9233
rect 2300 9173 2318 9207
rect 2352 9173 2370 9207
rect 2300 9147 2370 9173
rect 2400 9207 2454 9233
rect 2400 9173 2412 9207
rect 2446 9173 2454 9207
rect 2400 9147 2454 9173
rect 716 9067 770 9093
rect 716 9033 724 9067
rect 758 9033 770 9067
rect 716 9007 770 9033
rect 800 9067 870 9093
rect 800 9033 818 9067
rect 852 9033 870 9067
rect 800 9007 870 9033
rect 900 9067 970 9093
rect 900 9033 918 9067
rect 952 9033 970 9067
rect 900 9007 970 9033
rect 1000 9007 1070 9093
rect 1100 9067 1170 9093
rect 1100 9033 1118 9067
rect 1152 9033 1170 9067
rect 1100 9007 1170 9033
rect 1200 9067 1270 9093
rect 1200 9033 1218 9067
rect 1252 9033 1270 9067
rect 1200 9007 1270 9033
rect 1300 9007 1370 9093
rect 1400 9007 1470 9093
rect 1500 9067 1570 9093
rect 1500 9033 1518 9067
rect 1552 9033 1570 9067
rect 1500 9007 1570 9033
rect 1600 9067 1670 9093
rect 1600 9033 1618 9067
rect 1652 9033 1670 9067
rect 1600 9007 1670 9033
rect 1700 9067 1754 9093
rect 1700 9033 1712 9067
rect 1746 9033 1754 9067
rect 1700 9007 1754 9033
rect 1816 9067 1870 9093
rect 1816 9033 1824 9067
rect 1858 9033 1870 9067
rect 1816 9007 1870 9033
rect 1900 9067 1954 9093
rect 1900 9033 1912 9067
rect 1946 9033 1954 9067
rect 1900 9007 1954 9033
rect 2516 9207 2570 9233
rect 2516 9173 2524 9207
rect 2558 9173 2570 9207
rect 2516 9147 2570 9173
rect 2600 9207 2670 9233
rect 2600 9173 2618 9207
rect 2652 9173 2670 9207
rect 2600 9147 2670 9173
rect 2700 9207 2770 9233
rect 2700 9173 2718 9207
rect 2752 9173 2770 9207
rect 2700 9147 2770 9173
rect 2800 9147 2870 9233
rect 2900 9147 2970 9233
rect 3000 9147 3070 9233
rect 3100 9147 3170 9233
rect 3200 9147 3270 9233
rect 3300 9207 3370 9233
rect 3300 9173 3318 9207
rect 3352 9173 3370 9207
rect 3300 9147 3370 9173
rect 3400 9207 3470 9233
rect 3400 9173 3418 9207
rect 3452 9173 3470 9207
rect 3400 9147 3470 9173
rect 3500 9147 3570 9233
rect 3600 9147 3670 9233
rect 3700 9207 3770 9233
rect 3700 9173 3718 9207
rect 3752 9173 3770 9207
rect 3700 9147 3770 9173
rect 3800 9207 3870 9233
rect 3800 9173 3818 9207
rect 3852 9173 3870 9207
rect 3800 9147 3870 9173
rect 3900 9207 3970 9233
rect 3900 9173 3918 9207
rect 3952 9173 3970 9207
rect 3900 9147 3970 9173
rect 4000 9207 4054 9233
rect 4000 9173 4012 9207
rect 4046 9173 4054 9207
rect 4000 9147 4054 9173
rect 2016 9067 2070 9093
rect 2016 9033 2024 9067
rect 2058 9033 2070 9067
rect 2016 9007 2070 9033
rect 2100 9067 2170 9093
rect 2100 9033 2118 9067
rect 2152 9033 2170 9067
rect 2100 9007 2170 9033
rect 2200 9007 2270 9093
rect 2300 9007 2370 9093
rect 2400 9067 2470 9093
rect 2400 9033 2418 9067
rect 2452 9033 2470 9067
rect 2400 9007 2470 9033
rect 2500 9067 2570 9093
rect 2500 9033 2518 9067
rect 2552 9033 2570 9067
rect 2500 9007 2570 9033
rect 2600 9067 2654 9093
rect 2600 9033 2612 9067
rect 2646 9033 2654 9067
rect 2600 9007 2654 9033
rect 16 8867 70 8953
rect 100 8867 170 8953
rect 200 8927 270 8953
rect 200 8893 218 8927
rect 252 8893 270 8927
rect 200 8867 270 8893
rect 300 8927 370 8953
rect 300 8893 318 8927
rect 352 8893 370 8927
rect 300 8867 370 8893
rect 400 8927 470 8953
rect 400 8893 418 8927
rect 452 8893 470 8927
rect 400 8867 470 8893
rect 500 8867 570 8953
rect 600 8867 670 8953
rect 700 8867 770 8953
rect 800 8867 870 8953
rect 900 8927 970 8953
rect 900 8893 918 8927
rect 952 8893 970 8927
rect 900 8867 970 8893
rect 1000 8927 1070 8953
rect 1000 8893 1018 8927
rect 1052 8893 1070 8927
rect 1000 8867 1070 8893
rect 1100 8927 1170 8953
rect 1100 8893 1118 8927
rect 1152 8893 1170 8927
rect 1100 8867 1170 8893
rect 1200 8927 1270 8953
rect 1200 8893 1218 8927
rect 1252 8893 1270 8927
rect 1200 8867 1270 8893
rect 1300 8927 1370 8953
rect 1300 8893 1318 8927
rect 1352 8893 1370 8927
rect 1300 8867 1370 8893
rect 1400 8927 1470 8953
rect 1400 8893 1418 8927
rect 1452 8893 1470 8927
rect 1400 8867 1470 8893
rect 1500 8927 1570 8953
rect 1500 8893 1518 8927
rect 1552 8893 1570 8927
rect 1500 8867 1570 8893
rect 1600 8867 1670 8953
rect 1700 8867 1770 8953
rect 1800 8867 1870 8953
rect 1900 8927 1970 8953
rect 1900 8893 1918 8927
rect 1952 8893 1970 8927
rect 1900 8867 1970 8893
rect 2000 8927 2070 8953
rect 2000 8893 2018 8927
rect 2052 8893 2070 8927
rect 2000 8867 2070 8893
rect 2100 8927 2170 8953
rect 2100 8893 2118 8927
rect 2152 8893 2170 8927
rect 2100 8867 2170 8893
rect 2200 8927 2270 8953
rect 2200 8893 2218 8927
rect 2252 8893 2270 8927
rect 2200 8867 2270 8893
rect 2300 8867 2370 8953
rect 2400 8867 2470 8953
rect 2500 8927 2570 8953
rect 2500 8893 2518 8927
rect 2552 8893 2570 8927
rect 2500 8867 2570 8893
rect 2600 8927 2654 8953
rect 2600 8893 2612 8927
rect 2646 8893 2654 8927
rect 2600 8867 2654 8893
rect 16 8787 70 8813
rect 16 8753 24 8787
rect 58 8753 70 8787
rect 16 8727 70 8753
rect 100 8787 170 8813
rect 100 8753 118 8787
rect 152 8753 170 8787
rect 100 8727 170 8753
rect 200 8787 254 8813
rect 200 8753 212 8787
rect 246 8753 254 8787
rect 200 8727 254 8753
rect 316 8787 370 8813
rect 316 8753 324 8787
rect 358 8753 370 8787
rect 316 8727 370 8753
rect 400 8787 470 8813
rect 400 8753 418 8787
rect 452 8753 470 8787
rect 400 8727 470 8753
rect 500 8727 570 8813
rect 600 8787 670 8813
rect 600 8753 618 8787
rect 652 8753 670 8787
rect 600 8727 670 8753
rect 700 8787 770 8813
rect 700 8753 718 8787
rect 752 8753 770 8787
rect 700 8727 770 8753
rect 800 8727 870 8813
rect 900 8787 970 8813
rect 900 8753 918 8787
rect 952 8753 970 8787
rect 900 8727 970 8753
rect 1000 8787 1070 8813
rect 1000 8753 1018 8787
rect 1052 8753 1070 8787
rect 1000 8727 1070 8753
rect 1100 8787 1170 8813
rect 1100 8753 1118 8787
rect 1152 8753 1170 8787
rect 1100 8727 1170 8753
rect 1200 8787 1270 8813
rect 1200 8753 1218 8787
rect 1252 8753 1270 8787
rect 1200 8727 1270 8753
rect 1300 8787 1370 8813
rect 1300 8753 1318 8787
rect 1352 8753 1370 8787
rect 1300 8727 1370 8753
rect 1400 8727 1470 8813
rect 1500 8787 1570 8813
rect 1500 8753 1518 8787
rect 1552 8753 1570 8787
rect 1500 8727 1570 8753
rect 1600 8787 1670 8813
rect 1600 8753 1618 8787
rect 1652 8753 1670 8787
rect 1600 8727 1670 8753
rect 1700 8787 1770 8813
rect 1700 8753 1718 8787
rect 1752 8753 1770 8787
rect 1700 8727 1770 8753
rect 1800 8727 1870 8813
rect 1900 8787 1970 8813
rect 1900 8753 1918 8787
rect 1952 8753 1970 8787
rect 1900 8727 1970 8753
rect 2000 8787 2070 8813
rect 2000 8753 2018 8787
rect 2052 8753 2070 8787
rect 2000 8727 2070 8753
rect 2100 8787 2170 8813
rect 2100 8753 2118 8787
rect 2152 8753 2170 8787
rect 2100 8727 2170 8753
rect 2200 8787 2270 8813
rect 2200 8753 2218 8787
rect 2252 8753 2270 8787
rect 2200 8727 2270 8753
rect 2300 8787 2370 8813
rect 2300 8753 2318 8787
rect 2352 8753 2370 8787
rect 2300 8727 2370 8753
rect 2400 8787 2470 8813
rect 2400 8753 2418 8787
rect 2452 8753 2470 8787
rect 2400 8727 2470 8753
rect 2500 8787 2570 8813
rect 2500 8753 2518 8787
rect 2552 8753 2570 8787
rect 2500 8727 2570 8753
rect 2600 8787 2654 8813
rect 2600 8753 2612 8787
rect 2646 8753 2654 8787
rect 2600 8727 2654 8753
rect 16 8497 70 8583
rect 100 8497 170 8583
rect 200 8557 270 8583
rect 200 8523 218 8557
rect 252 8523 270 8557
rect 200 8497 270 8523
rect 300 8557 370 8583
rect 300 8523 318 8557
rect 352 8523 370 8557
rect 300 8497 370 8523
rect 400 8497 470 8583
rect 500 8557 570 8583
rect 500 8523 518 8557
rect 552 8523 570 8557
rect 500 8497 570 8523
rect 600 8557 670 8583
rect 600 8523 618 8557
rect 652 8523 670 8557
rect 600 8497 670 8523
rect 700 8557 770 8583
rect 700 8523 718 8557
rect 752 8523 770 8557
rect 700 8497 770 8523
rect 800 8557 854 8583
rect 800 8523 812 8557
rect 846 8523 854 8557
rect 800 8497 854 8523
rect 916 8557 970 8583
rect 916 8523 924 8557
rect 958 8523 970 8557
rect 916 8497 970 8523
rect 1000 8557 1054 8583
rect 1000 8523 1012 8557
rect 1046 8523 1054 8557
rect 1000 8497 1054 8523
rect 2716 9067 2770 9093
rect 2716 9033 2724 9067
rect 2758 9033 2770 9067
rect 2716 9007 2770 9033
rect 2800 9067 2854 9093
rect 2800 9033 2812 9067
rect 2846 9033 2854 9067
rect 2800 9007 2854 9033
rect 2916 9067 2970 9093
rect 2916 9033 2924 9067
rect 2958 9033 2970 9067
rect 2916 9007 2970 9033
rect 3000 9067 3070 9093
rect 3000 9033 3018 9067
rect 3052 9033 3070 9067
rect 3000 9007 3070 9033
rect 3100 9067 3170 9093
rect 3100 9033 3118 9067
rect 3152 9033 3170 9067
rect 3100 9007 3170 9033
rect 3200 9067 3254 9093
rect 3200 9033 3212 9067
rect 3246 9033 3254 9067
rect 3200 9007 3254 9033
rect 4616 9487 4670 9513
rect 4616 9453 4624 9487
rect 4658 9453 4670 9487
rect 4616 9427 4670 9453
rect 4700 9487 4770 9513
rect 4700 9453 4718 9487
rect 4752 9453 4770 9487
rect 4700 9427 4770 9453
rect 4800 9487 4854 9513
rect 4800 9453 4812 9487
rect 4846 9453 4854 9487
rect 4800 9427 4854 9453
rect 4916 9487 4970 9513
rect 4916 9453 4924 9487
rect 4958 9453 4970 9487
rect 4916 9427 4970 9453
rect 5000 9487 5054 9513
rect 5000 9453 5012 9487
rect 5046 9453 5054 9487
rect 5000 9427 5054 9453
rect 5116 9487 5170 9513
rect 5116 9453 5124 9487
rect 5158 9453 5170 9487
rect 5116 9427 5170 9453
rect 5200 9487 5254 9513
rect 5200 9453 5212 9487
rect 5246 9453 5254 9487
rect 5200 9427 5254 9453
rect 5316 9487 5370 9513
rect 5316 9453 5324 9487
rect 5358 9453 5370 9487
rect 5316 9427 5370 9453
rect 5400 9487 5470 9513
rect 5400 9453 5418 9487
rect 5452 9453 5470 9487
rect 5400 9427 5470 9453
rect 5500 9487 5570 9513
rect 5500 9453 5518 9487
rect 5552 9453 5570 9487
rect 5500 9427 5570 9453
rect 5600 9487 5654 9513
rect 5600 9453 5612 9487
rect 5646 9453 5654 9487
rect 5600 9427 5654 9453
rect 5716 9487 5770 9513
rect 5716 9453 5724 9487
rect 5758 9453 5770 9487
rect 5716 9427 5770 9453
rect 5800 9487 5854 9513
rect 5800 9453 5812 9487
rect 5846 9453 5854 9487
rect 5800 9427 5854 9453
rect 6016 9767 6070 9793
rect 6016 9733 6024 9767
rect 6058 9733 6070 9767
rect 6016 9707 6070 9733
rect 6100 9767 6170 9793
rect 6100 9733 6118 9767
rect 6152 9733 6170 9767
rect 6100 9707 6170 9733
rect 6200 9767 6270 9793
rect 6200 9733 6218 9767
rect 6252 9733 6270 9767
rect 6200 9707 6270 9733
rect 6300 9767 6370 9793
rect 6300 9733 6318 9767
rect 6352 9733 6370 9767
rect 6300 9707 6370 9733
rect 6400 9767 6454 9793
rect 6400 9733 6412 9767
rect 6446 9733 6454 9767
rect 6400 9707 6454 9733
rect 6512 9782 6570 9793
rect 6512 9748 6524 9782
rect 6558 9748 6570 9782
rect 6512 9707 6570 9748
rect 6600 9767 6670 9793
rect 6600 9733 6618 9767
rect 6652 9733 6670 9767
rect 6600 9707 6670 9733
rect 6700 9752 6758 9793
rect 6700 9718 6712 9752
rect 6746 9718 6758 9752
rect 6700 9707 6758 9718
rect 6820 9767 6880 9793
rect 6820 9733 6828 9767
rect 6862 9733 6880 9767
rect 6820 9707 6880 9733
rect 6910 9767 6980 9793
rect 6910 9733 6928 9767
rect 6962 9733 6980 9767
rect 6910 9707 6980 9733
rect 7010 9767 7080 9793
rect 7010 9733 7028 9767
rect 7062 9733 7080 9767
rect 7010 9707 7080 9733
rect 7110 9767 7180 9793
rect 7110 9733 7128 9767
rect 7162 9733 7180 9767
rect 7110 9707 7180 9733
rect 7210 9767 7280 9793
rect 7210 9733 7228 9767
rect 7262 9733 7280 9767
rect 7210 9707 7280 9733
rect 7310 9767 7380 9793
rect 7310 9733 7328 9767
rect 7362 9733 7380 9767
rect 7310 9707 7380 9733
rect 7410 9767 7470 9793
rect 7410 9733 7428 9767
rect 7462 9733 7470 9767
rect 7410 9707 7470 9733
rect 6016 9627 6070 9653
rect 6016 9593 6024 9627
rect 6058 9593 6070 9627
rect 6016 9567 6070 9593
rect 6100 9627 6170 9653
rect 6100 9593 6118 9627
rect 6152 9593 6170 9627
rect 6100 9567 6170 9593
rect 6200 9567 6270 9653
rect 6300 9627 6370 9653
rect 6300 9593 6318 9627
rect 6352 9593 6370 9627
rect 6300 9567 6370 9593
rect 6400 9627 6454 9653
rect 6400 9593 6412 9627
rect 6446 9593 6454 9627
rect 6400 9567 6454 9593
rect 6512 9642 6570 9653
rect 6512 9608 6524 9642
rect 6558 9608 6570 9642
rect 6512 9567 6570 9608
rect 6600 9627 6670 9653
rect 6600 9593 6618 9627
rect 6652 9593 6670 9627
rect 6600 9567 6670 9593
rect 6700 9612 6758 9653
rect 6700 9578 6712 9612
rect 6746 9578 6758 9612
rect 6700 9567 6758 9578
rect 6820 9627 6880 9653
rect 6820 9593 6828 9627
rect 6862 9593 6880 9627
rect 6820 9567 6880 9593
rect 6910 9627 6980 9653
rect 6910 9593 6928 9627
rect 6962 9593 6980 9627
rect 6910 9567 6980 9593
rect 7010 9627 7080 9653
rect 7010 9593 7028 9627
rect 7062 9593 7080 9627
rect 7010 9567 7080 9593
rect 7110 9627 7180 9653
rect 7110 9593 7128 9627
rect 7162 9593 7180 9627
rect 7110 9567 7180 9593
rect 7210 9627 7280 9653
rect 7210 9593 7228 9627
rect 7262 9593 7280 9627
rect 7210 9567 7280 9593
rect 7310 9627 7380 9653
rect 7310 9593 7328 9627
rect 7362 9593 7380 9627
rect 7310 9567 7380 9593
rect 7410 9627 7470 9653
rect 7410 9593 7428 9627
rect 7462 9593 7470 9627
rect 7410 9567 7470 9593
rect 5916 9487 5970 9513
rect 5916 9453 5924 9487
rect 5958 9453 5970 9487
rect 5916 9427 5970 9453
rect 6000 9487 6070 9513
rect 6000 9453 6018 9487
rect 6052 9453 6070 9487
rect 6000 9427 6070 9453
rect 6100 9487 6154 9513
rect 6100 9453 6112 9487
rect 6146 9453 6154 9487
rect 6100 9427 6154 9453
rect 6216 9487 6270 9513
rect 6216 9453 6224 9487
rect 6258 9453 6270 9487
rect 6216 9427 6270 9453
rect 6300 9487 6370 9513
rect 6300 9453 6318 9487
rect 6352 9453 6370 9487
rect 6300 9427 6370 9453
rect 6400 9487 6454 9513
rect 6400 9453 6412 9487
rect 6446 9453 6454 9487
rect 6400 9427 6454 9453
rect 6512 9502 6570 9513
rect 6512 9468 6524 9502
rect 6558 9468 6570 9502
rect 6512 9427 6570 9468
rect 6600 9487 6670 9513
rect 6600 9453 6618 9487
rect 6652 9453 6670 9487
rect 6600 9427 6670 9453
rect 6700 9472 6758 9513
rect 6700 9438 6712 9472
rect 6746 9438 6758 9472
rect 6700 9427 6758 9438
rect 6820 9487 6880 9513
rect 6820 9453 6828 9487
rect 6862 9453 6880 9487
rect 6820 9427 6880 9453
rect 6910 9487 6980 9513
rect 6910 9453 6928 9487
rect 6962 9453 6980 9487
rect 6910 9427 6980 9453
rect 7010 9487 7080 9513
rect 7010 9453 7028 9487
rect 7062 9453 7080 9487
rect 7010 9427 7080 9453
rect 7110 9487 7180 9513
rect 7110 9453 7128 9487
rect 7162 9453 7180 9487
rect 7110 9427 7180 9453
rect 7210 9487 7280 9513
rect 7210 9453 7228 9487
rect 7262 9453 7280 9487
rect 7210 9427 7280 9453
rect 7310 9487 7380 9513
rect 7310 9453 7328 9487
rect 7362 9453 7380 9487
rect 7310 9427 7380 9453
rect 7410 9487 7470 9513
rect 7410 9453 7428 9487
rect 7462 9453 7470 9487
rect 7410 9427 7470 9453
rect 4216 9347 4270 9373
rect 4216 9313 4224 9347
rect 4258 9313 4270 9347
rect 4216 9287 4270 9313
rect 4300 9347 4370 9373
rect 4300 9313 4318 9347
rect 4352 9313 4370 9347
rect 4300 9287 4370 9313
rect 4400 9287 4470 9373
rect 4500 9347 4570 9373
rect 4500 9313 4518 9347
rect 4552 9313 4570 9347
rect 4500 9287 4570 9313
rect 4600 9347 4670 9373
rect 4600 9313 4618 9347
rect 4652 9313 4670 9347
rect 4600 9287 4670 9313
rect 4700 9287 4770 9373
rect 4800 9347 4870 9373
rect 4800 9313 4818 9347
rect 4852 9313 4870 9347
rect 4800 9287 4870 9313
rect 4900 9347 4970 9373
rect 4900 9313 4918 9347
rect 4952 9313 4970 9347
rect 4900 9287 4970 9313
rect 5000 9287 5070 9373
rect 5100 9347 5170 9373
rect 5100 9313 5118 9347
rect 5152 9313 5170 9347
rect 5100 9287 5170 9313
rect 5200 9347 5270 9373
rect 5200 9313 5218 9347
rect 5252 9313 5270 9347
rect 5200 9287 5270 9313
rect 5300 9347 5370 9373
rect 5300 9313 5318 9347
rect 5352 9313 5370 9347
rect 5300 9287 5370 9313
rect 5400 9347 5470 9373
rect 5400 9313 5418 9347
rect 5452 9313 5470 9347
rect 5400 9287 5470 9313
rect 5500 9347 5570 9373
rect 5500 9313 5518 9347
rect 5552 9313 5570 9347
rect 5500 9287 5570 9313
rect 5600 9287 5670 9373
rect 5700 9287 5770 9373
rect 5800 9347 5870 9373
rect 5800 9313 5818 9347
rect 5852 9313 5870 9347
rect 5800 9287 5870 9313
rect 5900 9347 5970 9373
rect 5900 9313 5918 9347
rect 5952 9313 5970 9347
rect 5900 9287 5970 9313
rect 6000 9287 6070 9373
rect 6100 9347 6170 9373
rect 6100 9313 6118 9347
rect 6152 9313 6170 9347
rect 6100 9287 6170 9313
rect 6200 9347 6270 9373
rect 6200 9313 6218 9347
rect 6252 9313 6270 9347
rect 6200 9287 6270 9313
rect 6300 9347 6370 9373
rect 6300 9313 6318 9347
rect 6352 9313 6370 9347
rect 6300 9287 6370 9313
rect 6400 9347 6454 9373
rect 6400 9313 6412 9347
rect 6446 9313 6454 9347
rect 6400 9287 6454 9313
rect 6512 9362 6570 9373
rect 6512 9328 6524 9362
rect 6558 9328 6570 9362
rect 6512 9287 6570 9328
rect 6600 9347 6670 9373
rect 6600 9313 6618 9347
rect 6652 9313 6670 9347
rect 6600 9287 6670 9313
rect 6700 9332 6758 9373
rect 6700 9298 6712 9332
rect 6746 9298 6758 9332
rect 6700 9287 6758 9298
rect 6820 9347 6880 9373
rect 6820 9313 6828 9347
rect 6862 9313 6880 9347
rect 6820 9287 6880 9313
rect 6910 9347 6980 9373
rect 6910 9313 6928 9347
rect 6962 9313 6980 9347
rect 6910 9287 6980 9313
rect 7010 9347 7080 9373
rect 7010 9313 7028 9347
rect 7062 9313 7080 9347
rect 7010 9287 7080 9313
rect 7110 9347 7180 9373
rect 7110 9313 7128 9347
rect 7162 9313 7180 9347
rect 7110 9287 7180 9313
rect 7210 9347 7280 9373
rect 7210 9313 7228 9347
rect 7262 9313 7280 9347
rect 7210 9287 7280 9313
rect 7310 9347 7380 9373
rect 7310 9313 7328 9347
rect 7362 9313 7380 9347
rect 7310 9287 7380 9313
rect 7410 9347 7470 9373
rect 7410 9313 7428 9347
rect 7462 9313 7470 9347
rect 7410 9287 7470 9313
rect 4116 9207 4170 9233
rect 4116 9173 4124 9207
rect 4158 9173 4170 9207
rect 4116 9147 4170 9173
rect 4200 9207 4270 9233
rect 4200 9173 4218 9207
rect 4252 9173 4270 9207
rect 4200 9147 4270 9173
rect 4300 9147 4370 9233
rect 4400 9207 4470 9233
rect 4400 9173 4418 9207
rect 4452 9173 4470 9207
rect 4400 9147 4470 9173
rect 4500 9207 4570 9233
rect 4500 9173 4518 9207
rect 4552 9173 4570 9207
rect 4500 9147 4570 9173
rect 4600 9147 4670 9233
rect 4700 9147 4770 9233
rect 4800 9147 4870 9233
rect 4900 9207 4970 9233
rect 4900 9173 4918 9207
rect 4952 9173 4970 9207
rect 4900 9147 4970 9173
rect 5000 9207 5054 9233
rect 5000 9173 5012 9207
rect 5046 9173 5054 9207
rect 5000 9147 5054 9173
rect 3316 9067 3370 9093
rect 3316 9033 3324 9067
rect 3358 9033 3370 9067
rect 3316 9007 3370 9033
rect 3400 9067 3470 9093
rect 3400 9033 3418 9067
rect 3452 9033 3470 9067
rect 3400 9007 3470 9033
rect 3500 9067 3570 9093
rect 3500 9033 3518 9067
rect 3552 9033 3570 9067
rect 3500 9007 3570 9033
rect 3600 9067 3670 9093
rect 3600 9033 3618 9067
rect 3652 9033 3670 9067
rect 3600 9007 3670 9033
rect 3700 9007 3770 9093
rect 3800 9007 3870 9093
rect 3900 9007 3970 9093
rect 4000 9067 4070 9093
rect 4000 9033 4018 9067
rect 4052 9033 4070 9067
rect 4000 9007 4070 9033
rect 4100 9067 4170 9093
rect 4100 9033 4118 9067
rect 4152 9033 4170 9067
rect 4100 9007 4170 9033
rect 4200 9067 4270 9093
rect 4200 9033 4218 9067
rect 4252 9033 4270 9067
rect 4200 9007 4270 9033
rect 4300 9007 4370 9093
rect 4400 9067 4470 9093
rect 4400 9033 4418 9067
rect 4452 9033 4470 9067
rect 4400 9007 4470 9033
rect 4500 9067 4554 9093
rect 4500 9033 4512 9067
rect 4546 9033 4554 9067
rect 4500 9007 4554 9033
rect 2716 8927 2770 8953
rect 2716 8893 2724 8927
rect 2758 8893 2770 8927
rect 2716 8867 2770 8893
rect 2800 8927 2870 8953
rect 2800 8893 2818 8927
rect 2852 8893 2870 8927
rect 2800 8867 2870 8893
rect 2900 8867 2970 8953
rect 3000 8927 3070 8953
rect 3000 8893 3018 8927
rect 3052 8893 3070 8927
rect 3000 8867 3070 8893
rect 3100 8927 3170 8953
rect 3100 8893 3118 8927
rect 3152 8893 3170 8927
rect 3100 8867 3170 8893
rect 3200 8867 3270 8953
rect 3300 8867 3370 8953
rect 3400 8867 3470 8953
rect 3500 8867 3570 8953
rect 3600 8867 3670 8953
rect 3700 8867 3770 8953
rect 3800 8927 3870 8953
rect 3800 8893 3818 8927
rect 3852 8893 3870 8927
rect 3800 8867 3870 8893
rect 3900 8927 3970 8953
rect 3900 8893 3918 8927
rect 3952 8893 3970 8927
rect 3900 8867 3970 8893
rect 4000 8867 4070 8953
rect 4100 8927 4170 8953
rect 4100 8893 4118 8927
rect 4152 8893 4170 8927
rect 4100 8867 4170 8893
rect 4200 8927 4270 8953
rect 4200 8893 4218 8927
rect 4252 8893 4270 8927
rect 4200 8867 4270 8893
rect 4300 8927 4370 8953
rect 4300 8893 4318 8927
rect 4352 8893 4370 8927
rect 4300 8867 4370 8893
rect 4400 8927 4454 8953
rect 4400 8893 4412 8927
rect 4446 8893 4454 8927
rect 4400 8867 4454 8893
rect 2716 8787 2770 8813
rect 2716 8753 2724 8787
rect 2758 8753 2770 8787
rect 2716 8727 2770 8753
rect 2800 8787 2870 8813
rect 2800 8753 2818 8787
rect 2852 8753 2870 8787
rect 2800 8727 2870 8753
rect 2900 8727 2970 8813
rect 3000 8787 3070 8813
rect 3000 8753 3018 8787
rect 3052 8753 3070 8787
rect 3000 8727 3070 8753
rect 3100 8787 3154 8813
rect 3100 8753 3112 8787
rect 3146 8753 3154 8787
rect 3100 8727 3154 8753
rect 1116 8557 1170 8583
rect 1116 8523 1124 8557
rect 1158 8523 1170 8557
rect 1116 8497 1170 8523
rect 1200 8557 1270 8583
rect 1200 8523 1218 8557
rect 1252 8523 1270 8557
rect 1200 8497 1270 8523
rect 1300 8497 1370 8583
rect 1400 8497 1470 8583
rect 1500 8497 1570 8583
rect 1600 8497 1670 8583
rect 1700 8497 1770 8583
rect 1800 8557 1870 8583
rect 1800 8523 1818 8557
rect 1852 8523 1870 8557
rect 1800 8497 1870 8523
rect 1900 8557 1970 8583
rect 1900 8523 1918 8557
rect 1952 8523 1970 8557
rect 1900 8497 1970 8523
rect 2000 8557 2070 8583
rect 2000 8523 2018 8557
rect 2052 8523 2070 8557
rect 2000 8497 2070 8523
rect 2100 8557 2170 8583
rect 2100 8523 2118 8557
rect 2152 8523 2170 8557
rect 2100 8497 2170 8523
rect 2200 8497 2270 8583
rect 2300 8557 2370 8583
rect 2300 8523 2318 8557
rect 2352 8523 2370 8557
rect 2300 8497 2370 8523
rect 2400 8557 2470 8583
rect 2400 8523 2418 8557
rect 2452 8523 2470 8557
rect 2400 8497 2470 8523
rect 2500 8497 2570 8583
rect 2600 8557 2670 8583
rect 2600 8523 2618 8557
rect 2652 8523 2670 8557
rect 2600 8497 2670 8523
rect 2700 8557 2754 8583
rect 2700 8523 2712 8557
rect 2746 8523 2754 8557
rect 2700 8497 2754 8523
rect 16 8417 70 8443
rect 16 8383 24 8417
rect 58 8383 70 8417
rect 16 8357 70 8383
rect 100 8417 170 8443
rect 100 8383 118 8417
rect 152 8383 170 8417
rect 100 8357 170 8383
rect 200 8357 270 8443
rect 300 8357 370 8443
rect 400 8417 470 8443
rect 400 8383 418 8417
rect 452 8383 470 8417
rect 400 8357 470 8383
rect 500 8417 570 8443
rect 500 8383 518 8417
rect 552 8383 570 8417
rect 500 8357 570 8383
rect 600 8417 670 8443
rect 600 8383 618 8417
rect 652 8383 670 8417
rect 600 8357 670 8383
rect 700 8417 770 8443
rect 700 8383 718 8417
rect 752 8383 770 8417
rect 700 8357 770 8383
rect 800 8417 870 8443
rect 800 8383 818 8417
rect 852 8383 870 8417
rect 800 8357 870 8383
rect 900 8357 970 8443
rect 1000 8357 1070 8443
rect 1100 8417 1170 8443
rect 1100 8383 1118 8417
rect 1152 8383 1170 8417
rect 1100 8357 1170 8383
rect 1200 8417 1270 8443
rect 1200 8383 1218 8417
rect 1252 8383 1270 8417
rect 1200 8357 1270 8383
rect 1300 8417 1354 8443
rect 1300 8383 1312 8417
rect 1346 8383 1354 8417
rect 1300 8357 1354 8383
rect 16 8217 70 8303
rect 100 8277 170 8303
rect 100 8243 118 8277
rect 152 8243 170 8277
rect 100 8217 170 8243
rect 200 8277 270 8303
rect 200 8243 218 8277
rect 252 8243 270 8277
rect 200 8217 270 8243
rect 300 8277 370 8303
rect 300 8243 318 8277
rect 352 8243 370 8277
rect 300 8217 370 8243
rect 400 8217 470 8303
rect 500 8277 570 8303
rect 500 8243 518 8277
rect 552 8243 570 8277
rect 500 8217 570 8243
rect 600 8277 654 8303
rect 600 8243 612 8277
rect 646 8243 654 8277
rect 600 8217 654 8243
rect 716 8277 770 8303
rect 716 8243 724 8277
rect 758 8243 770 8277
rect 716 8217 770 8243
rect 800 8277 854 8303
rect 800 8243 812 8277
rect 846 8243 854 8277
rect 800 8217 854 8243
rect 1416 8417 1470 8443
rect 1416 8383 1424 8417
rect 1458 8383 1470 8417
rect 1416 8357 1470 8383
rect 1500 8417 1570 8443
rect 1500 8383 1518 8417
rect 1552 8383 1570 8417
rect 1500 8357 1570 8383
rect 1600 8417 1670 8443
rect 1600 8383 1618 8417
rect 1652 8383 1670 8417
rect 1600 8357 1670 8383
rect 1700 8417 1770 8443
rect 1700 8383 1718 8417
rect 1752 8383 1770 8417
rect 1700 8357 1770 8383
rect 1800 8417 1854 8443
rect 1800 8383 1812 8417
rect 1846 8383 1854 8417
rect 1800 8357 1854 8383
rect 1916 8417 1970 8443
rect 1916 8383 1924 8417
rect 1958 8383 1970 8417
rect 1916 8357 1970 8383
rect 2000 8417 2054 8443
rect 2000 8383 2012 8417
rect 2046 8383 2054 8417
rect 2000 8357 2054 8383
rect 916 8277 970 8303
rect 916 8243 924 8277
rect 958 8243 970 8277
rect 916 8217 970 8243
rect 1000 8277 1070 8303
rect 1000 8243 1018 8277
rect 1052 8243 1070 8277
rect 1000 8217 1070 8243
rect 1100 8217 1170 8303
rect 1200 8217 1270 8303
rect 1300 8217 1370 8303
rect 1400 8277 1470 8303
rect 1400 8243 1418 8277
rect 1452 8243 1470 8277
rect 1400 8217 1470 8243
rect 1500 8277 1570 8303
rect 1500 8243 1518 8277
rect 1552 8243 1570 8277
rect 1500 8217 1570 8243
rect 1600 8277 1670 8303
rect 1600 8243 1618 8277
rect 1652 8243 1670 8277
rect 1600 8217 1670 8243
rect 1700 8217 1770 8303
rect 1800 8277 1870 8303
rect 1800 8243 1818 8277
rect 1852 8243 1870 8277
rect 1800 8217 1870 8243
rect 1900 8277 1954 8303
rect 1900 8243 1912 8277
rect 1946 8243 1954 8277
rect 1900 8217 1954 8243
rect 16 8077 70 8163
rect 100 8077 170 8163
rect 200 8137 270 8163
rect 200 8103 218 8137
rect 252 8103 270 8137
rect 200 8077 270 8103
rect 300 8137 370 8163
rect 300 8103 318 8137
rect 352 8103 370 8137
rect 300 8077 370 8103
rect 400 8077 470 8163
rect 500 8137 570 8163
rect 500 8103 518 8137
rect 552 8103 570 8137
rect 500 8077 570 8103
rect 600 8137 670 8163
rect 600 8103 618 8137
rect 652 8103 670 8137
rect 600 8077 670 8103
rect 700 8077 770 8163
rect 800 8077 870 8163
rect 900 8077 970 8163
rect 1000 8137 1070 8163
rect 1000 8103 1018 8137
rect 1052 8103 1070 8137
rect 1000 8077 1070 8103
rect 1100 8137 1170 8163
rect 1100 8103 1118 8137
rect 1152 8103 1170 8137
rect 1100 8077 1170 8103
rect 1200 8137 1254 8163
rect 1200 8103 1212 8137
rect 1246 8103 1254 8137
rect 1200 8077 1254 8103
rect 16 7937 70 8023
rect 100 7997 170 8023
rect 100 7963 118 7997
rect 152 7963 170 7997
rect 100 7937 170 7963
rect 200 7997 254 8023
rect 200 7963 212 7997
rect 246 7963 254 7997
rect 200 7937 254 7963
rect 316 7997 370 8023
rect 316 7963 324 7997
rect 358 7963 370 7997
rect 316 7937 370 7963
rect 400 7997 470 8023
rect 400 7963 418 7997
rect 452 7963 470 7997
rect 400 7937 470 7963
rect 500 7937 570 8023
rect 600 7997 670 8023
rect 600 7963 618 7997
rect 652 7963 670 7997
rect 600 7937 670 7963
rect 700 7997 770 8023
rect 700 7963 718 7997
rect 752 7963 770 7997
rect 700 7937 770 7963
rect 800 7997 870 8023
rect 800 7963 818 7997
rect 852 7963 870 7997
rect 800 7937 870 7963
rect 900 7997 970 8023
rect 900 7963 918 7997
rect 952 7963 970 7997
rect 900 7937 970 7963
rect 1000 7997 1054 8023
rect 1000 7963 1012 7997
rect 1046 7963 1054 7997
rect 1000 7937 1054 7963
rect 16 7857 70 7883
rect 16 7823 24 7857
rect 58 7823 70 7857
rect 16 7797 70 7823
rect 100 7857 170 7883
rect 100 7823 118 7857
rect 152 7823 170 7857
rect 100 7797 170 7823
rect 200 7857 270 7883
rect 200 7823 218 7857
rect 252 7823 270 7857
rect 200 7797 270 7823
rect 300 7857 370 7883
rect 300 7823 318 7857
rect 352 7823 370 7857
rect 300 7797 370 7823
rect 400 7797 470 7883
rect 500 7857 570 7883
rect 500 7823 518 7857
rect 552 7823 570 7857
rect 500 7797 570 7823
rect 600 7857 654 7883
rect 600 7823 612 7857
rect 646 7823 654 7857
rect 600 7797 654 7823
rect 716 7857 770 7883
rect 716 7823 724 7857
rect 758 7823 770 7857
rect 716 7797 770 7823
rect 800 7857 854 7883
rect 800 7823 812 7857
rect 846 7823 854 7857
rect 800 7797 854 7823
rect 2116 8417 2170 8443
rect 2116 8383 2124 8417
rect 2158 8383 2170 8417
rect 2116 8357 2170 8383
rect 2200 8417 2270 8443
rect 2200 8383 2218 8417
rect 2252 8383 2270 8417
rect 2200 8357 2270 8383
rect 2300 8417 2354 8443
rect 2300 8383 2312 8417
rect 2346 8383 2354 8417
rect 2300 8357 2354 8383
rect 2016 8277 2070 8303
rect 2016 8243 2024 8277
rect 2058 8243 2070 8277
rect 2016 8217 2070 8243
rect 2100 8277 2170 8303
rect 2100 8243 2118 8277
rect 2152 8243 2170 8277
rect 2100 8217 2170 8243
rect 2200 8277 2270 8303
rect 2200 8243 2218 8277
rect 2252 8243 2270 8277
rect 2200 8217 2270 8243
rect 2300 8277 2354 8303
rect 2300 8243 2312 8277
rect 2346 8243 2354 8277
rect 2300 8217 2354 8243
rect 4616 9067 4670 9093
rect 4616 9033 4624 9067
rect 4658 9033 4670 9067
rect 4616 9007 4670 9033
rect 4700 9067 4754 9093
rect 4700 9033 4712 9067
rect 4746 9033 4754 9067
rect 4700 9007 4754 9033
rect 4516 8927 4570 8953
rect 4516 8893 4524 8927
rect 4558 8893 4570 8927
rect 4516 8867 4570 8893
rect 4600 8927 4654 8953
rect 4600 8893 4612 8927
rect 4646 8893 4654 8927
rect 4600 8867 4654 8893
rect 5116 9207 5170 9233
rect 5116 9173 5124 9207
rect 5158 9173 5170 9207
rect 5116 9147 5170 9173
rect 5200 9207 5270 9233
rect 5200 9173 5218 9207
rect 5252 9173 5270 9207
rect 5200 9147 5270 9173
rect 5300 9207 5370 9233
rect 5300 9173 5318 9207
rect 5352 9173 5370 9207
rect 5300 9147 5370 9173
rect 5400 9207 5454 9233
rect 5400 9173 5412 9207
rect 5446 9173 5454 9207
rect 5400 9147 5454 9173
rect 4816 9067 4870 9093
rect 4816 9033 4824 9067
rect 4858 9033 4870 9067
rect 4816 9007 4870 9033
rect 4900 9067 4970 9093
rect 4900 9033 4918 9067
rect 4952 9033 4970 9067
rect 4900 9007 4970 9033
rect 5000 9007 5070 9093
rect 5100 9067 5170 9093
rect 5100 9033 5118 9067
rect 5152 9033 5170 9067
rect 5100 9007 5170 9033
rect 5200 9067 5254 9093
rect 5200 9033 5212 9067
rect 5246 9033 5254 9067
rect 5200 9007 5254 9033
rect 4716 8927 4770 8953
rect 4716 8893 4724 8927
rect 4758 8893 4770 8927
rect 4716 8867 4770 8893
rect 4800 8927 4854 8953
rect 4800 8893 4812 8927
rect 4846 8893 4854 8927
rect 4800 8867 4854 8893
rect 5516 9207 5570 9233
rect 5516 9173 5524 9207
rect 5558 9173 5570 9207
rect 5516 9147 5570 9173
rect 5600 9207 5670 9233
rect 5600 9173 5618 9207
rect 5652 9173 5670 9207
rect 5600 9147 5670 9173
rect 5700 9207 5754 9233
rect 5700 9173 5712 9207
rect 5746 9173 5754 9207
rect 5700 9147 5754 9173
rect 5816 9207 5870 9233
rect 5816 9173 5824 9207
rect 5858 9173 5870 9207
rect 5816 9147 5870 9173
rect 5900 9207 5970 9233
rect 5900 9173 5918 9207
rect 5952 9173 5970 9207
rect 5900 9147 5970 9173
rect 6000 9147 6070 9233
rect 6100 9207 6170 9233
rect 6100 9173 6118 9207
rect 6152 9173 6170 9207
rect 6100 9147 6170 9173
rect 6200 9207 6270 9233
rect 6200 9173 6218 9207
rect 6252 9173 6270 9207
rect 6200 9147 6270 9173
rect 6300 9207 6370 9233
rect 6300 9173 6318 9207
rect 6352 9173 6370 9207
rect 6300 9147 6370 9173
rect 6400 9147 6454 9233
rect 6512 9222 6570 9233
rect 6512 9188 6524 9222
rect 6558 9188 6570 9222
rect 6512 9147 6570 9188
rect 6600 9207 6670 9233
rect 6600 9173 6618 9207
rect 6652 9173 6670 9207
rect 6600 9147 6670 9173
rect 6700 9192 6758 9233
rect 6700 9158 6712 9192
rect 6746 9158 6758 9192
rect 6700 9147 6758 9158
rect 6820 9207 6880 9233
rect 6820 9173 6828 9207
rect 6862 9173 6880 9207
rect 6820 9147 6880 9173
rect 6910 9207 6980 9233
rect 6910 9173 6928 9207
rect 6962 9173 6980 9207
rect 6910 9147 6980 9173
rect 7010 9207 7080 9233
rect 7010 9173 7028 9207
rect 7062 9173 7080 9207
rect 7010 9147 7080 9173
rect 7110 9207 7180 9233
rect 7110 9173 7128 9207
rect 7162 9173 7180 9207
rect 7110 9147 7180 9173
rect 7210 9207 7280 9233
rect 7210 9173 7228 9207
rect 7262 9173 7280 9207
rect 7210 9147 7280 9173
rect 7310 9207 7380 9233
rect 7310 9173 7328 9207
rect 7362 9173 7380 9207
rect 7310 9147 7380 9173
rect 7410 9207 7470 9233
rect 7410 9173 7428 9207
rect 7462 9173 7470 9207
rect 7410 9147 7470 9173
rect 5316 9067 5370 9093
rect 5316 9033 5324 9067
rect 5358 9033 5370 9067
rect 5316 9007 5370 9033
rect 5400 9067 5470 9093
rect 5400 9033 5418 9067
rect 5452 9033 5470 9067
rect 5400 9007 5470 9033
rect 5500 9007 5570 9093
rect 5600 9007 5670 9093
rect 5700 9007 5770 9093
rect 5800 9067 5870 9093
rect 5800 9033 5818 9067
rect 5852 9033 5870 9067
rect 5800 9007 5870 9033
rect 5900 9067 5970 9093
rect 5900 9033 5918 9067
rect 5952 9033 5970 9067
rect 5900 9007 5970 9033
rect 6000 9067 6070 9093
rect 6000 9033 6018 9067
rect 6052 9033 6070 9067
rect 6000 9007 6070 9033
rect 6100 9007 6170 9093
rect 6200 9067 6270 9093
rect 6200 9033 6218 9067
rect 6252 9033 6270 9067
rect 6200 9007 6270 9033
rect 6300 9067 6370 9093
rect 6300 9033 6318 9067
rect 6352 9033 6370 9067
rect 6300 9007 6370 9033
rect 6400 9067 6454 9093
rect 6400 9033 6412 9067
rect 6446 9033 6454 9067
rect 6400 9007 6454 9033
rect 6512 9082 6570 9093
rect 6512 9048 6524 9082
rect 6558 9048 6570 9082
rect 6512 9007 6570 9048
rect 6600 9067 6670 9093
rect 6600 9033 6618 9067
rect 6652 9033 6670 9067
rect 6600 9007 6670 9033
rect 6700 9052 6758 9093
rect 6700 9018 6712 9052
rect 6746 9018 6758 9052
rect 6700 9007 6758 9018
rect 6820 9067 6880 9093
rect 6820 9033 6828 9067
rect 6862 9033 6880 9067
rect 6820 9007 6880 9033
rect 6910 9067 6980 9093
rect 6910 9033 6928 9067
rect 6962 9033 6980 9067
rect 6910 9007 6980 9033
rect 7010 9067 7080 9093
rect 7010 9033 7028 9067
rect 7062 9033 7080 9067
rect 7010 9007 7080 9033
rect 7110 9067 7180 9093
rect 7110 9033 7128 9067
rect 7162 9033 7180 9067
rect 7110 9007 7180 9033
rect 7210 9067 7280 9093
rect 7210 9033 7228 9067
rect 7262 9033 7280 9067
rect 7210 9007 7280 9033
rect 7310 9067 7380 9093
rect 7310 9033 7328 9067
rect 7362 9033 7380 9067
rect 7310 9007 7380 9033
rect 7410 9067 7470 9093
rect 7410 9033 7428 9067
rect 7462 9033 7470 9067
rect 7410 9007 7470 9033
rect 4916 8927 4970 8953
rect 4916 8893 4924 8927
rect 4958 8893 4970 8927
rect 4916 8867 4970 8893
rect 5000 8927 5070 8953
rect 5000 8893 5018 8927
rect 5052 8893 5070 8927
rect 5000 8867 5070 8893
rect 5100 8927 5170 8953
rect 5100 8893 5118 8927
rect 5152 8893 5170 8927
rect 5100 8867 5170 8893
rect 5200 8927 5270 8953
rect 5200 8893 5218 8927
rect 5252 8893 5270 8927
rect 5200 8867 5270 8893
rect 5300 8927 5370 8953
rect 5300 8893 5318 8927
rect 5352 8893 5370 8927
rect 5300 8867 5370 8893
rect 5400 8867 5470 8953
rect 5500 8927 5570 8953
rect 5500 8893 5518 8927
rect 5552 8893 5570 8927
rect 5500 8867 5570 8893
rect 5600 8927 5654 8953
rect 5600 8893 5612 8927
rect 5646 8893 5654 8927
rect 5600 8867 5654 8893
rect 3216 8787 3270 8813
rect 3216 8753 3224 8787
rect 3258 8753 3270 8787
rect 3216 8727 3270 8753
rect 3300 8787 3370 8813
rect 3300 8753 3318 8787
rect 3352 8753 3370 8787
rect 3300 8727 3370 8753
rect 3400 8787 3470 8813
rect 3400 8753 3418 8787
rect 3452 8753 3470 8787
rect 3400 8727 3470 8753
rect 3500 8727 3570 8813
rect 3600 8787 3670 8813
rect 3600 8753 3618 8787
rect 3652 8753 3670 8787
rect 3600 8727 3670 8753
rect 3700 8787 3770 8813
rect 3700 8753 3718 8787
rect 3752 8753 3770 8787
rect 3700 8727 3770 8753
rect 3800 8727 3870 8813
rect 3900 8787 3970 8813
rect 3900 8753 3918 8787
rect 3952 8753 3970 8787
rect 3900 8727 3970 8753
rect 4000 8787 4070 8813
rect 4000 8753 4018 8787
rect 4052 8753 4070 8787
rect 4000 8727 4070 8753
rect 4100 8787 4170 8813
rect 4100 8753 4118 8787
rect 4152 8753 4170 8787
rect 4100 8727 4170 8753
rect 4200 8727 4270 8813
rect 4300 8727 4370 8813
rect 4400 8727 4470 8813
rect 4500 8787 4570 8813
rect 4500 8753 4518 8787
rect 4552 8753 4570 8787
rect 4500 8727 4570 8753
rect 4600 8787 4670 8813
rect 4600 8753 4618 8787
rect 4652 8753 4670 8787
rect 4600 8727 4670 8753
rect 4700 8787 4770 8813
rect 4700 8753 4718 8787
rect 4752 8753 4770 8787
rect 4700 8727 4770 8753
rect 4800 8727 4870 8813
rect 4900 8727 4970 8813
rect 5000 8727 5070 8813
rect 5100 8787 5170 8813
rect 5100 8753 5118 8787
rect 5152 8753 5170 8787
rect 5100 8727 5170 8753
rect 5200 8787 5270 8813
rect 5200 8753 5218 8787
rect 5252 8753 5270 8787
rect 5200 8727 5270 8753
rect 5300 8727 5370 8813
rect 5400 8787 5470 8813
rect 5400 8753 5418 8787
rect 5452 8753 5470 8787
rect 5400 8727 5470 8753
rect 5500 8787 5554 8813
rect 5500 8753 5512 8787
rect 5546 8753 5554 8787
rect 5500 8727 5554 8753
rect 2816 8557 2870 8583
rect 2816 8523 2824 8557
rect 2858 8523 2870 8557
rect 2816 8497 2870 8523
rect 2900 8557 2970 8583
rect 2900 8523 2918 8557
rect 2952 8523 2970 8557
rect 2900 8497 2970 8523
rect 3000 8497 3070 8583
rect 3100 8557 3170 8583
rect 3100 8523 3118 8557
rect 3152 8523 3170 8557
rect 3100 8497 3170 8523
rect 3200 8557 3270 8583
rect 3200 8523 3218 8557
rect 3252 8523 3270 8557
rect 3200 8497 3270 8523
rect 3300 8557 3354 8583
rect 3300 8523 3312 8557
rect 3346 8523 3354 8557
rect 3300 8497 3354 8523
rect 3416 8557 3470 8583
rect 3416 8523 3424 8557
rect 3458 8523 3470 8557
rect 3416 8497 3470 8523
rect 3500 8557 3554 8583
rect 3500 8523 3512 8557
rect 3546 8523 3554 8557
rect 3500 8497 3554 8523
rect 3616 8557 3670 8583
rect 3616 8523 3624 8557
rect 3658 8523 3670 8557
rect 3616 8497 3670 8523
rect 3700 8557 3770 8583
rect 3700 8523 3718 8557
rect 3752 8523 3770 8557
rect 3700 8497 3770 8523
rect 3800 8497 3870 8583
rect 3900 8557 3970 8583
rect 3900 8523 3918 8557
rect 3952 8523 3970 8557
rect 3900 8497 3970 8523
rect 4000 8557 4054 8583
rect 4000 8523 4012 8557
rect 4046 8523 4054 8557
rect 4000 8497 4054 8523
rect 2416 8417 2470 8443
rect 2416 8383 2424 8417
rect 2458 8383 2470 8417
rect 2416 8357 2470 8383
rect 2500 8417 2570 8443
rect 2500 8383 2518 8417
rect 2552 8383 2570 8417
rect 2500 8357 2570 8383
rect 2600 8417 2670 8443
rect 2600 8383 2618 8417
rect 2652 8383 2670 8417
rect 2600 8357 2670 8383
rect 2700 8417 2770 8443
rect 2700 8383 2718 8417
rect 2752 8383 2770 8417
rect 2700 8357 2770 8383
rect 2800 8417 2870 8443
rect 2800 8383 2818 8417
rect 2852 8383 2870 8417
rect 2800 8357 2870 8383
rect 2900 8357 2970 8443
rect 3000 8417 3070 8443
rect 3000 8383 3018 8417
rect 3052 8383 3070 8417
rect 3000 8357 3070 8383
rect 3100 8417 3170 8443
rect 3100 8383 3118 8417
rect 3152 8383 3170 8417
rect 3100 8357 3170 8383
rect 3200 8417 3270 8443
rect 3200 8383 3218 8417
rect 3252 8383 3270 8417
rect 3200 8357 3270 8383
rect 3300 8357 3370 8443
rect 3400 8417 3470 8443
rect 3400 8383 3418 8417
rect 3452 8383 3470 8417
rect 3400 8357 3470 8383
rect 3500 8417 3570 8443
rect 3500 8383 3518 8417
rect 3552 8383 3570 8417
rect 3500 8357 3570 8383
rect 3600 8417 3670 8443
rect 3600 8383 3618 8417
rect 3652 8383 3670 8417
rect 3600 8357 3670 8383
rect 3700 8417 3770 8443
rect 3700 8383 3718 8417
rect 3752 8383 3770 8417
rect 3700 8357 3770 8383
rect 3800 8417 3854 8443
rect 3800 8383 3812 8417
rect 3846 8383 3854 8417
rect 3800 8357 3854 8383
rect 2416 8277 2470 8303
rect 2416 8243 2424 8277
rect 2458 8243 2470 8277
rect 2416 8217 2470 8243
rect 2500 8277 2554 8303
rect 2500 8243 2512 8277
rect 2546 8243 2554 8277
rect 2500 8217 2554 8243
rect 2616 8277 2670 8303
rect 2616 8243 2624 8277
rect 2658 8243 2670 8277
rect 2616 8217 2670 8243
rect 2700 8277 2770 8303
rect 2700 8243 2718 8277
rect 2752 8243 2770 8277
rect 2700 8217 2770 8243
rect 2800 8217 2870 8303
rect 2900 8277 2970 8303
rect 2900 8243 2918 8277
rect 2952 8243 2970 8277
rect 2900 8217 2970 8243
rect 3000 8277 3070 8303
rect 3000 8243 3018 8277
rect 3052 8243 3070 8277
rect 3000 8217 3070 8243
rect 3100 8277 3154 8303
rect 3100 8243 3112 8277
rect 3146 8243 3154 8277
rect 3100 8217 3154 8243
rect 1316 8137 1370 8163
rect 1316 8103 1324 8137
rect 1358 8103 1370 8137
rect 1316 8077 1370 8103
rect 1400 8137 1470 8163
rect 1400 8103 1418 8137
rect 1452 8103 1470 8137
rect 1400 8077 1470 8103
rect 1500 8137 1570 8163
rect 1500 8103 1518 8137
rect 1552 8103 1570 8137
rect 1500 8077 1570 8103
rect 1600 8077 1670 8163
rect 1700 8077 1770 8163
rect 1800 8077 1870 8163
rect 1900 8137 1970 8163
rect 1900 8103 1918 8137
rect 1952 8103 1970 8137
rect 1900 8077 1970 8103
rect 2000 8137 2070 8163
rect 2000 8103 2018 8137
rect 2052 8103 2070 8137
rect 2000 8077 2070 8103
rect 2100 8137 2170 8163
rect 2100 8103 2118 8137
rect 2152 8103 2170 8137
rect 2100 8077 2170 8103
rect 2200 8137 2270 8163
rect 2200 8103 2218 8137
rect 2252 8103 2270 8137
rect 2200 8077 2270 8103
rect 2300 8137 2370 8163
rect 2300 8103 2318 8137
rect 2352 8103 2370 8137
rect 2300 8077 2370 8103
rect 2400 8077 2470 8163
rect 2500 8137 2570 8163
rect 2500 8103 2518 8137
rect 2552 8103 2570 8137
rect 2500 8077 2570 8103
rect 2600 8137 2654 8163
rect 2600 8103 2612 8137
rect 2646 8103 2654 8137
rect 2600 8077 2654 8103
rect 1116 7997 1170 8023
rect 1116 7963 1124 7997
rect 1158 7963 1170 7997
rect 1116 7937 1170 7963
rect 1200 7997 1270 8023
rect 1200 7963 1218 7997
rect 1252 7963 1270 7997
rect 1200 7937 1270 7963
rect 1300 7997 1354 8023
rect 1300 7963 1312 7997
rect 1346 7963 1354 7997
rect 1300 7937 1354 7963
rect 1416 7997 1470 8023
rect 1416 7963 1424 7997
rect 1458 7963 1470 7997
rect 1416 7937 1470 7963
rect 1500 7997 1570 8023
rect 1500 7963 1518 7997
rect 1552 7963 1570 7997
rect 1500 7937 1570 7963
rect 1600 7997 1670 8023
rect 1600 7963 1618 7997
rect 1652 7963 1670 7997
rect 1600 7937 1670 7963
rect 1700 7997 1754 8023
rect 1700 7963 1712 7997
rect 1746 7963 1754 7997
rect 1700 7937 1754 7963
rect 916 7857 970 7883
rect 916 7823 924 7857
rect 958 7823 970 7857
rect 916 7797 970 7823
rect 1000 7857 1070 7883
rect 1000 7823 1018 7857
rect 1052 7823 1070 7857
rect 1000 7797 1070 7823
rect 1100 7857 1170 7883
rect 1100 7823 1118 7857
rect 1152 7823 1170 7857
rect 1100 7797 1170 7823
rect 1200 7857 1270 7883
rect 1200 7823 1218 7857
rect 1252 7823 1270 7857
rect 1200 7797 1270 7823
rect 1300 7857 1370 7883
rect 1300 7823 1318 7857
rect 1352 7823 1370 7857
rect 1300 7797 1370 7823
rect 1400 7857 1454 7883
rect 1400 7823 1412 7857
rect 1446 7823 1454 7857
rect 1400 7797 1454 7823
rect 1516 7857 1570 7883
rect 1516 7823 1524 7857
rect 1558 7823 1570 7857
rect 1516 7797 1570 7823
rect 1600 7857 1654 7883
rect 1600 7823 1612 7857
rect 1646 7823 1654 7857
rect 1600 7797 1654 7823
rect 16 7717 70 7743
rect 16 7683 24 7717
rect 58 7683 70 7717
rect 16 7657 70 7683
rect 100 7717 170 7743
rect 100 7683 118 7717
rect 152 7683 170 7717
rect 100 7657 170 7683
rect 200 7717 270 7743
rect 200 7683 218 7717
rect 252 7683 270 7717
rect 200 7657 270 7683
rect 300 7657 370 7743
rect 400 7657 470 7743
rect 500 7717 570 7743
rect 500 7683 518 7717
rect 552 7683 570 7717
rect 500 7657 570 7683
rect 600 7717 670 7743
rect 600 7683 618 7717
rect 652 7683 670 7717
rect 600 7657 670 7683
rect 700 7657 770 7743
rect 800 7657 870 7743
rect 900 7657 970 7743
rect 1000 7657 1070 7743
rect 1100 7717 1170 7743
rect 1100 7683 1118 7717
rect 1152 7683 1170 7717
rect 1100 7657 1170 7683
rect 1200 7717 1270 7743
rect 1200 7683 1218 7717
rect 1252 7683 1270 7717
rect 1200 7657 1270 7683
rect 1300 7657 1370 7743
rect 1400 7717 1470 7743
rect 1400 7683 1418 7717
rect 1452 7683 1470 7717
rect 1400 7657 1470 7683
rect 1500 7717 1554 7743
rect 1500 7683 1512 7717
rect 1546 7683 1554 7717
rect 1500 7657 1554 7683
rect 16 7577 70 7603
rect 16 7543 24 7577
rect 58 7543 70 7577
rect 16 7517 70 7543
rect 100 7577 170 7603
rect 100 7543 118 7577
rect 152 7543 170 7577
rect 100 7517 170 7543
rect 200 7577 270 7603
rect 200 7543 218 7577
rect 252 7543 270 7577
rect 200 7517 270 7543
rect 300 7517 370 7603
rect 400 7517 470 7603
rect 500 7517 570 7603
rect 600 7517 670 7603
rect 700 7517 770 7603
rect 800 7517 870 7603
rect 900 7577 970 7603
rect 900 7543 918 7577
rect 952 7543 970 7577
rect 900 7517 970 7543
rect 1000 7577 1054 7603
rect 1000 7543 1012 7577
rect 1046 7543 1054 7577
rect 1000 7517 1054 7543
rect 1116 7577 1170 7603
rect 1116 7543 1124 7577
rect 1158 7543 1170 7577
rect 1116 7517 1170 7543
rect 1200 7577 1270 7603
rect 1200 7543 1218 7577
rect 1252 7543 1270 7577
rect 1200 7517 1270 7543
rect 1300 7577 1354 7603
rect 1300 7543 1312 7577
rect 1346 7543 1354 7577
rect 1300 7517 1354 7543
rect 1816 7997 1870 8023
rect 1816 7963 1824 7997
rect 1858 7963 1870 7997
rect 1816 7937 1870 7963
rect 1900 7997 1970 8023
rect 1900 7963 1918 7997
rect 1952 7963 1970 7997
rect 1900 7937 1970 7963
rect 2000 7997 2054 8023
rect 2000 7963 2012 7997
rect 2046 7963 2054 7997
rect 2000 7937 2054 7963
rect 2716 8137 2770 8163
rect 2716 8103 2724 8137
rect 2758 8103 2770 8137
rect 2716 8077 2770 8103
rect 2800 8137 2854 8163
rect 2800 8103 2812 8137
rect 2846 8103 2854 8137
rect 2800 8077 2854 8103
rect 2116 7997 2170 8023
rect 2116 7963 2124 7997
rect 2158 7963 2170 7997
rect 2116 7937 2170 7963
rect 2200 7997 2270 8023
rect 2200 7963 2218 7997
rect 2252 7963 2270 7997
rect 2200 7937 2270 7963
rect 2300 7997 2370 8023
rect 2300 7963 2318 7997
rect 2352 7963 2370 7997
rect 2300 7937 2370 7963
rect 2400 7937 2470 8023
rect 2500 7997 2570 8023
rect 2500 7963 2518 7997
rect 2552 7963 2570 7997
rect 2500 7937 2570 7963
rect 2600 7997 2670 8023
rect 2600 7963 2618 7997
rect 2652 7963 2670 7997
rect 2600 7937 2670 7963
rect 2700 7997 2754 8023
rect 2700 7963 2712 7997
rect 2746 7963 2754 7997
rect 2700 7937 2754 7963
rect 1716 7857 1770 7883
rect 1716 7823 1724 7857
rect 1758 7823 1770 7857
rect 1716 7797 1770 7823
rect 1800 7857 1870 7883
rect 1800 7823 1818 7857
rect 1852 7823 1870 7857
rect 1800 7797 1870 7823
rect 1900 7797 1970 7883
rect 2000 7857 2070 7883
rect 2000 7823 2018 7857
rect 2052 7823 2070 7857
rect 2000 7797 2070 7823
rect 2100 7857 2170 7883
rect 2100 7823 2118 7857
rect 2152 7823 2170 7857
rect 2100 7797 2170 7823
rect 2200 7797 2270 7883
rect 2300 7857 2370 7883
rect 2300 7823 2318 7857
rect 2352 7823 2370 7857
rect 2300 7797 2370 7823
rect 2400 7857 2470 7883
rect 2400 7823 2418 7857
rect 2452 7823 2470 7857
rect 2400 7797 2470 7823
rect 2500 7857 2554 7883
rect 2500 7823 2512 7857
rect 2546 7823 2554 7857
rect 2500 7797 2554 7823
rect 1616 7717 1670 7743
rect 1616 7683 1624 7717
rect 1658 7683 1670 7717
rect 1616 7657 1670 7683
rect 1700 7717 1754 7743
rect 1700 7683 1712 7717
rect 1746 7683 1754 7717
rect 1700 7657 1754 7683
rect 3216 8277 3270 8303
rect 3216 8243 3224 8277
rect 3258 8243 3270 8277
rect 3216 8217 3270 8243
rect 3300 8277 3370 8303
rect 3300 8243 3318 8277
rect 3352 8243 3370 8277
rect 3300 8217 3370 8243
rect 3400 8277 3470 8303
rect 3400 8243 3418 8277
rect 3452 8243 3470 8277
rect 3400 8217 3470 8243
rect 3500 8277 3554 8303
rect 3500 8243 3512 8277
rect 3546 8243 3554 8277
rect 3500 8217 3554 8243
rect 4116 8557 4170 8583
rect 4116 8523 4124 8557
rect 4158 8523 4170 8557
rect 4116 8497 4170 8523
rect 4200 8557 4270 8583
rect 4200 8523 4218 8557
rect 4252 8523 4270 8557
rect 4200 8497 4270 8523
rect 4300 8557 4354 8583
rect 4300 8523 4312 8557
rect 4346 8523 4354 8557
rect 4300 8497 4354 8523
rect 4416 8557 4470 8583
rect 4416 8523 4424 8557
rect 4458 8523 4470 8557
rect 4416 8497 4470 8523
rect 4500 8557 4570 8583
rect 4500 8523 4518 8557
rect 4552 8523 4570 8557
rect 4500 8497 4570 8523
rect 4600 8557 4670 8583
rect 4600 8523 4618 8557
rect 4652 8523 4670 8557
rect 4600 8497 4670 8523
rect 4700 8557 4754 8583
rect 4700 8523 4712 8557
rect 4746 8523 4754 8557
rect 4700 8497 4754 8523
rect 3916 8417 3970 8443
rect 3916 8383 3924 8417
rect 3958 8383 3970 8417
rect 3916 8357 3970 8383
rect 4000 8417 4070 8443
rect 4000 8383 4018 8417
rect 4052 8383 4070 8417
rect 4000 8357 4070 8383
rect 4100 8357 4170 8443
rect 4200 8417 4270 8443
rect 4200 8383 4218 8417
rect 4252 8383 4270 8417
rect 4200 8357 4270 8383
rect 4300 8417 4370 8443
rect 4300 8383 4318 8417
rect 4352 8383 4370 8417
rect 4300 8357 4370 8383
rect 4400 8357 4470 8443
rect 4500 8417 4570 8443
rect 4500 8383 4518 8417
rect 4552 8383 4570 8417
rect 4500 8357 4570 8383
rect 4600 8417 4670 8443
rect 4600 8383 4618 8417
rect 4652 8383 4670 8417
rect 4600 8357 4670 8383
rect 4700 8417 4754 8443
rect 4700 8383 4712 8417
rect 4746 8383 4754 8417
rect 4700 8357 4754 8383
rect 5716 8927 5770 8953
rect 5716 8893 5724 8927
rect 5758 8893 5770 8927
rect 5716 8867 5770 8893
rect 5800 8927 5870 8953
rect 5800 8893 5818 8927
rect 5852 8893 5870 8927
rect 5800 8867 5870 8893
rect 5900 8867 5970 8953
rect 6000 8927 6070 8953
rect 6000 8893 6018 8927
rect 6052 8893 6070 8927
rect 6000 8867 6070 8893
rect 6100 8927 6154 8953
rect 6100 8893 6112 8927
rect 6146 8893 6154 8927
rect 6100 8867 6154 8893
rect 5616 8787 5670 8813
rect 5616 8753 5624 8787
rect 5658 8753 5670 8787
rect 5616 8727 5670 8753
rect 5700 8787 5770 8813
rect 5700 8753 5718 8787
rect 5752 8753 5770 8787
rect 5700 8727 5770 8753
rect 5800 8787 5870 8813
rect 5800 8753 5818 8787
rect 5852 8753 5870 8787
rect 5800 8727 5870 8753
rect 5900 8787 5954 8813
rect 5900 8753 5912 8787
rect 5946 8753 5954 8787
rect 5900 8727 5954 8753
rect 4816 8557 4870 8583
rect 4816 8523 4824 8557
rect 4858 8523 4870 8557
rect 4816 8497 4870 8523
rect 4900 8557 4970 8583
rect 4900 8523 4918 8557
rect 4952 8523 4970 8557
rect 4900 8497 4970 8523
rect 5000 8557 5070 8583
rect 5000 8523 5018 8557
rect 5052 8523 5070 8557
rect 5000 8497 5070 8523
rect 5100 8497 5170 8583
rect 5200 8557 5270 8583
rect 5200 8523 5218 8557
rect 5252 8523 5270 8557
rect 5200 8497 5270 8523
rect 5300 8557 5370 8583
rect 5300 8523 5318 8557
rect 5352 8523 5370 8557
rect 5300 8497 5370 8523
rect 5400 8557 5470 8583
rect 5400 8523 5418 8557
rect 5452 8523 5470 8557
rect 5400 8497 5470 8523
rect 5500 8557 5570 8583
rect 5500 8523 5518 8557
rect 5552 8523 5570 8557
rect 5500 8497 5570 8523
rect 5600 8557 5654 8583
rect 5600 8523 5612 8557
rect 5646 8523 5654 8557
rect 5600 8497 5654 8523
rect 4816 8417 4870 8443
rect 4816 8383 4824 8417
rect 4858 8383 4870 8417
rect 4816 8357 4870 8383
rect 4900 8417 4954 8443
rect 4900 8383 4912 8417
rect 4946 8383 4954 8417
rect 4900 8357 4954 8383
rect 6216 8927 6270 8953
rect 6216 8893 6224 8927
rect 6258 8893 6270 8927
rect 6216 8867 6270 8893
rect 6300 8927 6370 8953
rect 6300 8893 6318 8927
rect 6352 8893 6370 8927
rect 6300 8867 6370 8893
rect 6400 8867 6454 8953
rect 6512 8942 6570 8953
rect 6512 8908 6524 8942
rect 6558 8908 6570 8942
rect 6512 8867 6570 8908
rect 6600 8927 6670 8953
rect 6600 8893 6618 8927
rect 6652 8893 6670 8927
rect 6600 8867 6670 8893
rect 6700 8912 6758 8953
rect 6700 8878 6712 8912
rect 6746 8878 6758 8912
rect 6700 8867 6758 8878
rect 6820 8927 6880 8953
rect 6820 8893 6828 8927
rect 6862 8893 6880 8927
rect 6820 8867 6880 8893
rect 6910 8927 6980 8953
rect 6910 8893 6928 8927
rect 6962 8893 6980 8927
rect 6910 8867 6980 8893
rect 7010 8927 7080 8953
rect 7010 8893 7028 8927
rect 7062 8893 7080 8927
rect 7010 8867 7080 8893
rect 7110 8927 7180 8953
rect 7110 8893 7128 8927
rect 7162 8893 7180 8927
rect 7110 8867 7180 8893
rect 7210 8927 7280 8953
rect 7210 8893 7228 8927
rect 7262 8893 7280 8927
rect 7210 8867 7280 8893
rect 7310 8927 7380 8953
rect 7310 8893 7328 8927
rect 7362 8893 7380 8927
rect 7310 8867 7380 8893
rect 7410 8927 7470 8953
rect 7410 8893 7428 8927
rect 7462 8893 7470 8927
rect 7410 8867 7470 8893
rect 6016 8787 6070 8813
rect 6016 8753 6024 8787
rect 6058 8753 6070 8787
rect 6016 8727 6070 8753
rect 6100 8787 6170 8813
rect 6100 8753 6118 8787
rect 6152 8753 6170 8787
rect 6100 8727 6170 8753
rect 6200 8787 6270 8813
rect 6200 8753 6218 8787
rect 6252 8753 6270 8787
rect 6200 8727 6270 8753
rect 6300 8787 6370 8813
rect 6300 8753 6318 8787
rect 6352 8753 6370 8787
rect 6300 8727 6370 8753
rect 6400 8727 6454 8813
rect 6512 8802 6570 8813
rect 6512 8768 6524 8802
rect 6558 8768 6570 8802
rect 6512 8727 6570 8768
rect 6600 8787 6670 8813
rect 6600 8753 6618 8787
rect 6652 8753 6670 8787
rect 6600 8727 6670 8753
rect 6700 8772 6758 8813
rect 6700 8738 6712 8772
rect 6746 8738 6758 8772
rect 6700 8727 6758 8738
rect 6820 8787 6880 8813
rect 6820 8753 6828 8787
rect 6862 8753 6880 8787
rect 6820 8727 6880 8753
rect 6910 8787 6980 8813
rect 6910 8753 6928 8787
rect 6962 8753 6980 8787
rect 6910 8727 6980 8753
rect 7010 8787 7080 8813
rect 7010 8753 7028 8787
rect 7062 8753 7080 8787
rect 7010 8727 7080 8753
rect 7110 8787 7180 8813
rect 7110 8753 7128 8787
rect 7162 8753 7180 8787
rect 7110 8727 7180 8753
rect 7210 8787 7280 8813
rect 7210 8753 7228 8787
rect 7262 8753 7280 8787
rect 7210 8727 7280 8753
rect 7310 8787 7380 8813
rect 7310 8753 7328 8787
rect 7362 8753 7380 8787
rect 7310 8727 7380 8753
rect 7410 8787 7470 8813
rect 7410 8753 7428 8787
rect 7462 8753 7470 8787
rect 7410 8727 7470 8753
rect 5716 8557 5770 8583
rect 5716 8523 5724 8557
rect 5758 8523 5770 8557
rect 5716 8497 5770 8523
rect 5800 8557 5870 8583
rect 5800 8523 5818 8557
rect 5852 8523 5870 8557
rect 5800 8497 5870 8523
rect 5900 8497 5970 8583
rect 6000 8497 6070 8583
rect 6100 8497 6170 8583
rect 6200 8557 6270 8583
rect 6200 8523 6218 8557
rect 6252 8523 6270 8557
rect 6200 8497 6270 8523
rect 6300 8557 6370 8583
rect 6300 8523 6318 8557
rect 6352 8523 6370 8557
rect 6300 8497 6370 8523
rect 6400 8497 6454 8583
rect 6512 8572 6570 8583
rect 6512 8538 6524 8572
rect 6558 8538 6570 8572
rect 6512 8497 6570 8538
rect 6600 8557 6670 8583
rect 6600 8523 6618 8557
rect 6652 8523 6670 8557
rect 6600 8497 6670 8523
rect 6700 8542 6758 8583
rect 6700 8508 6712 8542
rect 6746 8508 6758 8542
rect 6700 8497 6758 8508
rect 6820 8557 6880 8583
rect 6820 8523 6828 8557
rect 6862 8523 6880 8557
rect 6820 8497 6880 8523
rect 6910 8557 6980 8583
rect 6910 8523 6928 8557
rect 6962 8523 6980 8557
rect 6910 8497 6980 8523
rect 7010 8557 7080 8583
rect 7010 8523 7028 8557
rect 7062 8523 7080 8557
rect 7010 8497 7080 8523
rect 7110 8557 7180 8583
rect 7110 8523 7128 8557
rect 7162 8523 7180 8557
rect 7110 8497 7180 8523
rect 7210 8557 7280 8583
rect 7210 8523 7228 8557
rect 7262 8523 7280 8557
rect 7210 8497 7280 8523
rect 7310 8557 7380 8583
rect 7310 8523 7328 8557
rect 7362 8523 7380 8557
rect 7310 8497 7380 8523
rect 7410 8557 7470 8583
rect 7410 8523 7428 8557
rect 7462 8523 7470 8557
rect 7410 8497 7470 8523
rect 5016 8417 5070 8443
rect 5016 8383 5024 8417
rect 5058 8383 5070 8417
rect 5016 8357 5070 8383
rect 5100 8417 5170 8443
rect 5100 8383 5118 8417
rect 5152 8383 5170 8417
rect 5100 8357 5170 8383
rect 5200 8417 5270 8443
rect 5200 8383 5218 8417
rect 5252 8383 5270 8417
rect 5200 8357 5270 8383
rect 5300 8417 5370 8443
rect 5300 8383 5318 8417
rect 5352 8383 5370 8417
rect 5300 8357 5370 8383
rect 5400 8357 5470 8443
rect 5500 8357 5570 8443
rect 5600 8357 5670 8443
rect 5700 8417 5770 8443
rect 5700 8383 5718 8417
rect 5752 8383 5770 8417
rect 5700 8357 5770 8383
rect 5800 8417 5854 8443
rect 5800 8383 5812 8417
rect 5846 8383 5854 8417
rect 5800 8357 5854 8383
rect 5916 8417 5970 8443
rect 5916 8383 5924 8417
rect 5958 8383 5970 8417
rect 5916 8357 5970 8383
rect 6000 8417 6070 8443
rect 6000 8383 6018 8417
rect 6052 8383 6070 8417
rect 6000 8357 6070 8383
rect 6100 8417 6170 8443
rect 6100 8383 6118 8417
rect 6152 8383 6170 8417
rect 6100 8357 6170 8383
rect 6200 8357 6270 8443
rect 6300 8417 6370 8443
rect 6300 8383 6318 8417
rect 6352 8383 6370 8417
rect 6300 8357 6370 8383
rect 6400 8417 6454 8443
rect 6400 8383 6412 8417
rect 6446 8383 6454 8417
rect 6400 8357 6454 8383
rect 6512 8432 6570 8443
rect 6512 8398 6524 8432
rect 6558 8398 6570 8432
rect 6512 8357 6570 8398
rect 6600 8417 6670 8443
rect 6600 8383 6618 8417
rect 6652 8383 6670 8417
rect 6600 8357 6670 8383
rect 6700 8402 6758 8443
rect 6700 8368 6712 8402
rect 6746 8368 6758 8402
rect 6700 8357 6758 8368
rect 6820 8417 6880 8443
rect 6820 8383 6828 8417
rect 6862 8383 6880 8417
rect 6820 8357 6880 8383
rect 6910 8417 6980 8443
rect 6910 8383 6928 8417
rect 6962 8383 6980 8417
rect 6910 8357 6980 8383
rect 7010 8417 7080 8443
rect 7010 8383 7028 8417
rect 7062 8383 7080 8417
rect 7010 8357 7080 8383
rect 7110 8417 7180 8443
rect 7110 8383 7128 8417
rect 7162 8383 7180 8417
rect 7110 8357 7180 8383
rect 7210 8417 7280 8443
rect 7210 8383 7228 8417
rect 7262 8383 7280 8417
rect 7210 8357 7280 8383
rect 7310 8417 7380 8443
rect 7310 8383 7328 8417
rect 7362 8383 7380 8417
rect 7310 8357 7380 8383
rect 7410 8417 7470 8443
rect 7410 8383 7428 8417
rect 7462 8383 7470 8417
rect 7410 8357 7470 8383
rect 3616 8277 3670 8303
rect 3616 8243 3624 8277
rect 3658 8243 3670 8277
rect 3616 8217 3670 8243
rect 3700 8277 3770 8303
rect 3700 8243 3718 8277
rect 3752 8243 3770 8277
rect 3700 8217 3770 8243
rect 3800 8277 3870 8303
rect 3800 8243 3818 8277
rect 3852 8243 3870 8277
rect 3800 8217 3870 8243
rect 3900 8217 3970 8303
rect 4000 8217 4070 8303
rect 4100 8217 4170 8303
rect 4200 8277 4270 8303
rect 4200 8243 4218 8277
rect 4252 8243 4270 8277
rect 4200 8217 4270 8243
rect 4300 8277 4370 8303
rect 4300 8243 4318 8277
rect 4352 8243 4370 8277
rect 4300 8217 4370 8243
rect 4400 8217 4470 8303
rect 4500 8217 4570 8303
rect 4600 8277 4670 8303
rect 4600 8243 4618 8277
rect 4652 8243 4670 8277
rect 4600 8217 4670 8243
rect 4700 8277 4770 8303
rect 4700 8243 4718 8277
rect 4752 8243 4770 8277
rect 4700 8217 4770 8243
rect 4800 8217 4870 8303
rect 4900 8217 4970 8303
rect 5000 8277 5070 8303
rect 5000 8243 5018 8277
rect 5052 8243 5070 8277
rect 5000 8217 5070 8243
rect 5100 8277 5170 8303
rect 5100 8243 5118 8277
rect 5152 8243 5170 8277
rect 5100 8217 5170 8243
rect 5200 8277 5270 8303
rect 5200 8243 5218 8277
rect 5252 8243 5270 8277
rect 5200 8217 5270 8243
rect 5300 8217 5370 8303
rect 5400 8217 5470 8303
rect 5500 8277 5570 8303
rect 5500 8243 5518 8277
rect 5552 8243 5570 8277
rect 5500 8217 5570 8243
rect 5600 8277 5670 8303
rect 5600 8243 5618 8277
rect 5652 8243 5670 8277
rect 5600 8217 5670 8243
rect 5700 8217 5770 8303
rect 5800 8217 5870 8303
rect 5900 8217 5970 8303
rect 6000 8217 6070 8303
rect 6100 8277 6170 8303
rect 6100 8243 6118 8277
rect 6152 8243 6170 8277
rect 6100 8217 6170 8243
rect 6200 8277 6270 8303
rect 6200 8243 6218 8277
rect 6252 8243 6270 8277
rect 6200 8217 6270 8243
rect 6300 8277 6370 8303
rect 6300 8243 6318 8277
rect 6352 8243 6370 8277
rect 6300 8217 6370 8243
rect 6400 8277 6454 8303
rect 6400 8243 6412 8277
rect 6446 8243 6454 8277
rect 6400 8217 6454 8243
rect 6512 8292 6570 8303
rect 6512 8258 6524 8292
rect 6558 8258 6570 8292
rect 6512 8217 6570 8258
rect 6600 8277 6670 8303
rect 6600 8243 6618 8277
rect 6652 8243 6670 8277
rect 6600 8217 6670 8243
rect 6700 8262 6758 8303
rect 6700 8228 6712 8262
rect 6746 8228 6758 8262
rect 6700 8217 6758 8228
rect 6820 8277 6880 8303
rect 6820 8243 6828 8277
rect 6862 8243 6880 8277
rect 6820 8217 6880 8243
rect 6910 8277 6980 8303
rect 6910 8243 6928 8277
rect 6962 8243 6980 8277
rect 6910 8217 6980 8243
rect 7010 8277 7080 8303
rect 7010 8243 7028 8277
rect 7062 8243 7080 8277
rect 7010 8217 7080 8243
rect 7110 8277 7180 8303
rect 7110 8243 7128 8277
rect 7162 8243 7180 8277
rect 7110 8217 7180 8243
rect 7210 8277 7280 8303
rect 7210 8243 7228 8277
rect 7262 8243 7280 8277
rect 7210 8217 7280 8243
rect 7310 8277 7380 8303
rect 7310 8243 7328 8277
rect 7362 8243 7380 8277
rect 7310 8217 7380 8243
rect 7410 8277 7470 8303
rect 7410 8243 7428 8277
rect 7462 8243 7470 8277
rect 7410 8217 7470 8243
rect 2916 8137 2970 8163
rect 2916 8103 2924 8137
rect 2958 8103 2970 8137
rect 2916 8077 2970 8103
rect 3000 8137 3070 8163
rect 3000 8103 3018 8137
rect 3052 8103 3070 8137
rect 3000 8077 3070 8103
rect 3100 8077 3170 8163
rect 3200 8077 3270 8163
rect 3300 8077 3370 8163
rect 3400 8077 3470 8163
rect 3500 8137 3570 8163
rect 3500 8103 3518 8137
rect 3552 8103 3570 8137
rect 3500 8077 3570 8103
rect 3600 8137 3670 8163
rect 3600 8103 3618 8137
rect 3652 8103 3670 8137
rect 3600 8077 3670 8103
rect 3700 8137 3754 8163
rect 3700 8103 3712 8137
rect 3746 8103 3754 8137
rect 3700 8077 3754 8103
rect 2816 7997 2870 8023
rect 2816 7963 2824 7997
rect 2858 7963 2870 7997
rect 2816 7937 2870 7963
rect 2900 7997 2954 8023
rect 2900 7963 2912 7997
rect 2946 7963 2954 7997
rect 2900 7937 2954 7963
rect 3816 8137 3870 8163
rect 3816 8103 3824 8137
rect 3858 8103 3870 8137
rect 3816 8077 3870 8103
rect 3900 8137 3970 8163
rect 3900 8103 3918 8137
rect 3952 8103 3970 8137
rect 3900 8077 3970 8103
rect 4000 8137 4070 8163
rect 4000 8103 4018 8137
rect 4052 8103 4070 8137
rect 4000 8077 4070 8103
rect 4100 8137 4170 8163
rect 4100 8103 4118 8137
rect 4152 8103 4170 8137
rect 4100 8077 4170 8103
rect 4200 8137 4270 8163
rect 4200 8103 4218 8137
rect 4252 8103 4270 8137
rect 4200 8077 4270 8103
rect 4300 8137 4370 8163
rect 4300 8103 4318 8137
rect 4352 8103 4370 8137
rect 4300 8077 4370 8103
rect 4400 8137 4470 8163
rect 4400 8103 4418 8137
rect 4452 8103 4470 8137
rect 4400 8077 4470 8103
rect 4500 8077 4570 8163
rect 4600 8077 4670 8163
rect 4700 8137 4770 8163
rect 4700 8103 4718 8137
rect 4752 8103 4770 8137
rect 4700 8077 4770 8103
rect 4800 8137 4870 8163
rect 4800 8103 4818 8137
rect 4852 8103 4870 8137
rect 4800 8077 4870 8103
rect 4900 8137 4970 8163
rect 4900 8103 4918 8137
rect 4952 8103 4970 8137
rect 4900 8077 4970 8103
rect 5000 8077 5070 8163
rect 5100 8077 5170 8163
rect 5200 8137 5270 8163
rect 5200 8103 5218 8137
rect 5252 8103 5270 8137
rect 5200 8077 5270 8103
rect 5300 8137 5370 8163
rect 5300 8103 5318 8137
rect 5352 8103 5370 8137
rect 5300 8077 5370 8103
rect 5400 8137 5470 8163
rect 5400 8103 5418 8137
rect 5452 8103 5470 8137
rect 5400 8077 5470 8103
rect 5500 8137 5570 8163
rect 5500 8103 5518 8137
rect 5552 8103 5570 8137
rect 5500 8077 5570 8103
rect 5600 8077 5670 8163
rect 5700 8137 5770 8163
rect 5700 8103 5718 8137
rect 5752 8103 5770 8137
rect 5700 8077 5770 8103
rect 5800 8137 5870 8163
rect 5800 8103 5818 8137
rect 5852 8103 5870 8137
rect 5800 8077 5870 8103
rect 5900 8137 5970 8163
rect 5900 8103 5918 8137
rect 5952 8103 5970 8137
rect 5900 8077 5970 8103
rect 6000 8137 6070 8163
rect 6000 8103 6018 8137
rect 6052 8103 6070 8137
rect 6000 8077 6070 8103
rect 6100 8137 6170 8163
rect 6100 8103 6118 8137
rect 6152 8103 6170 8137
rect 6100 8077 6170 8103
rect 6200 8137 6270 8163
rect 6200 8103 6218 8137
rect 6252 8103 6270 8137
rect 6200 8077 6270 8103
rect 6300 8077 6370 8163
rect 6400 8077 6454 8163
rect 6512 8152 6570 8163
rect 6512 8118 6524 8152
rect 6558 8118 6570 8152
rect 6512 8077 6570 8118
rect 6600 8137 6670 8163
rect 6600 8103 6618 8137
rect 6652 8103 6670 8137
rect 6600 8077 6670 8103
rect 6700 8122 6758 8163
rect 6700 8088 6712 8122
rect 6746 8088 6758 8122
rect 6700 8077 6758 8088
rect 6820 8137 6880 8163
rect 6820 8103 6828 8137
rect 6862 8103 6880 8137
rect 6820 8077 6880 8103
rect 6910 8137 6980 8163
rect 6910 8103 6928 8137
rect 6962 8103 6980 8137
rect 6910 8077 6980 8103
rect 7010 8137 7080 8163
rect 7010 8103 7028 8137
rect 7062 8103 7080 8137
rect 7010 8077 7080 8103
rect 7110 8137 7180 8163
rect 7110 8103 7128 8137
rect 7162 8103 7180 8137
rect 7110 8077 7180 8103
rect 7210 8137 7280 8163
rect 7210 8103 7228 8137
rect 7262 8103 7280 8137
rect 7210 8077 7280 8103
rect 7310 8137 7380 8163
rect 7310 8103 7328 8137
rect 7362 8103 7380 8137
rect 7310 8077 7380 8103
rect 7410 8137 7470 8163
rect 7410 8103 7428 8137
rect 7462 8103 7470 8137
rect 7410 8077 7470 8103
rect 3016 7997 3070 8023
rect 3016 7963 3024 7997
rect 3058 7963 3070 7997
rect 3016 7937 3070 7963
rect 3100 7997 3170 8023
rect 3100 7963 3118 7997
rect 3152 7963 3170 7997
rect 3100 7937 3170 7963
rect 3200 7937 3270 8023
rect 3300 7997 3370 8023
rect 3300 7963 3318 7997
rect 3352 7963 3370 7997
rect 3300 7937 3370 7963
rect 3400 7997 3470 8023
rect 3400 7963 3418 7997
rect 3452 7963 3470 7997
rect 3400 7937 3470 7963
rect 3500 7937 3570 8023
rect 3600 7997 3670 8023
rect 3600 7963 3618 7997
rect 3652 7963 3670 7997
rect 3600 7937 3670 7963
rect 3700 7997 3770 8023
rect 3700 7963 3718 7997
rect 3752 7963 3770 7997
rect 3700 7937 3770 7963
rect 3800 7937 3870 8023
rect 3900 7997 3970 8023
rect 3900 7963 3918 7997
rect 3952 7963 3970 7997
rect 3900 7937 3970 7963
rect 4000 7997 4070 8023
rect 4000 7963 4018 7997
rect 4052 7963 4070 7997
rect 4000 7937 4070 7963
rect 4100 7997 4170 8023
rect 4100 7963 4118 7997
rect 4152 7963 4170 7997
rect 4100 7937 4170 7963
rect 4200 7937 4270 8023
rect 4300 7997 4370 8023
rect 4300 7963 4318 7997
rect 4352 7963 4370 7997
rect 4300 7937 4370 7963
rect 4400 7997 4470 8023
rect 4400 7963 4418 7997
rect 4452 7963 4470 7997
rect 4400 7937 4470 7963
rect 4500 7997 4570 8023
rect 4500 7963 4518 7997
rect 4552 7963 4570 7997
rect 4500 7937 4570 7963
rect 4600 7937 4670 8023
rect 4700 7997 4770 8023
rect 4700 7963 4718 7997
rect 4752 7963 4770 7997
rect 4700 7937 4770 7963
rect 4800 7997 4870 8023
rect 4800 7963 4818 7997
rect 4852 7963 4870 7997
rect 4800 7937 4870 7963
rect 4900 7997 4954 8023
rect 4900 7963 4912 7997
rect 4946 7963 4954 7997
rect 4900 7937 4954 7963
rect 2616 7857 2670 7883
rect 2616 7823 2624 7857
rect 2658 7823 2670 7857
rect 2616 7797 2670 7823
rect 2700 7857 2770 7883
rect 2700 7823 2718 7857
rect 2752 7823 2770 7857
rect 2700 7797 2770 7823
rect 2800 7797 2870 7883
rect 2900 7857 2970 7883
rect 2900 7823 2918 7857
rect 2952 7823 2970 7857
rect 2900 7797 2970 7823
rect 3000 7857 3070 7883
rect 3000 7823 3018 7857
rect 3052 7823 3070 7857
rect 3000 7797 3070 7823
rect 3100 7797 3170 7883
rect 3200 7857 3270 7883
rect 3200 7823 3218 7857
rect 3252 7823 3270 7857
rect 3200 7797 3270 7823
rect 3300 7857 3354 7883
rect 3300 7823 3312 7857
rect 3346 7823 3354 7857
rect 3300 7797 3354 7823
rect 1816 7717 1870 7743
rect 1816 7683 1824 7717
rect 1858 7683 1870 7717
rect 1816 7657 1870 7683
rect 1900 7717 1970 7743
rect 1900 7683 1918 7717
rect 1952 7683 1970 7717
rect 1900 7657 1970 7683
rect 2000 7717 2070 7743
rect 2000 7683 2018 7717
rect 2052 7683 2070 7717
rect 2000 7657 2070 7683
rect 2100 7717 2170 7743
rect 2100 7683 2118 7717
rect 2152 7683 2170 7717
rect 2100 7657 2170 7683
rect 2200 7657 2270 7743
rect 2300 7657 2370 7743
rect 2400 7657 2470 7743
rect 2500 7717 2570 7743
rect 2500 7683 2518 7717
rect 2552 7683 2570 7717
rect 2500 7657 2570 7683
rect 2600 7717 2670 7743
rect 2600 7683 2618 7717
rect 2652 7683 2670 7717
rect 2600 7657 2670 7683
rect 2700 7717 2754 7743
rect 2700 7683 2712 7717
rect 2746 7683 2754 7717
rect 2700 7657 2754 7683
rect 1416 7577 1470 7603
rect 1416 7543 1424 7577
rect 1458 7543 1470 7577
rect 1416 7517 1470 7543
rect 1500 7577 1570 7603
rect 1500 7543 1518 7577
rect 1552 7543 1570 7577
rect 1500 7517 1570 7543
rect 1600 7577 1670 7603
rect 1600 7543 1618 7577
rect 1652 7543 1670 7577
rect 1600 7517 1670 7543
rect 1700 7577 1770 7603
rect 1700 7543 1718 7577
rect 1752 7543 1770 7577
rect 1700 7517 1770 7543
rect 1800 7517 1870 7603
rect 1900 7577 1970 7603
rect 1900 7543 1918 7577
rect 1952 7543 1970 7577
rect 1900 7517 1970 7543
rect 2000 7577 2070 7603
rect 2000 7543 2018 7577
rect 2052 7543 2070 7577
rect 2000 7517 2070 7543
rect 2100 7517 2170 7603
rect 2200 7517 2270 7603
rect 2300 7577 2370 7603
rect 2300 7543 2318 7577
rect 2352 7543 2370 7577
rect 2300 7517 2370 7543
rect 2400 7577 2470 7603
rect 2400 7543 2418 7577
rect 2452 7543 2470 7577
rect 2400 7517 2470 7543
rect 2500 7517 2570 7603
rect 2600 7577 2670 7603
rect 2600 7543 2618 7577
rect 2652 7543 2670 7577
rect 2600 7517 2670 7543
rect 2700 7577 2754 7603
rect 2700 7543 2712 7577
rect 2746 7543 2754 7577
rect 2700 7517 2754 7543
rect 16 7287 70 7373
rect 100 7287 170 7373
rect 200 7347 270 7373
rect 200 7313 218 7347
rect 252 7313 270 7347
rect 200 7287 270 7313
rect 300 7347 370 7373
rect 300 7313 318 7347
rect 352 7313 370 7347
rect 300 7287 370 7313
rect 400 7347 470 7373
rect 400 7313 418 7347
rect 452 7313 470 7347
rect 400 7287 470 7313
rect 500 7347 570 7373
rect 500 7313 518 7347
rect 552 7313 570 7347
rect 500 7287 570 7313
rect 600 7287 670 7373
rect 700 7287 770 7373
rect 800 7347 870 7373
rect 800 7313 818 7347
rect 852 7313 870 7347
rect 800 7287 870 7313
rect 900 7347 970 7373
rect 900 7313 918 7347
rect 952 7313 970 7347
rect 900 7287 970 7313
rect 1000 7347 1070 7373
rect 1000 7313 1018 7347
rect 1052 7313 1070 7347
rect 1000 7287 1070 7313
rect 1100 7347 1170 7373
rect 1100 7313 1118 7347
rect 1152 7313 1170 7347
rect 1100 7287 1170 7313
rect 1200 7347 1254 7373
rect 1200 7313 1212 7347
rect 1246 7313 1254 7347
rect 1200 7287 1254 7313
rect 16 7147 70 7233
rect 100 7207 170 7233
rect 100 7173 118 7207
rect 152 7173 170 7207
rect 100 7147 170 7173
rect 200 7207 270 7233
rect 200 7173 218 7207
rect 252 7173 270 7207
rect 200 7147 270 7173
rect 300 7207 354 7233
rect 300 7173 312 7207
rect 346 7173 354 7207
rect 300 7147 354 7173
rect 16 7067 70 7093
rect 16 7033 24 7067
rect 58 7033 70 7067
rect 16 7007 70 7033
rect 100 7067 170 7093
rect 100 7033 118 7067
rect 152 7033 170 7067
rect 100 7007 170 7033
rect 200 7067 270 7093
rect 200 7033 218 7067
rect 252 7033 270 7067
rect 200 7007 270 7033
rect 300 7067 354 7093
rect 300 7033 312 7067
rect 346 7033 354 7067
rect 300 7007 354 7033
rect 1316 7347 1370 7373
rect 1316 7313 1324 7347
rect 1358 7313 1370 7347
rect 1316 7287 1370 7313
rect 1400 7347 1470 7373
rect 1400 7313 1418 7347
rect 1452 7313 1470 7347
rect 1400 7287 1470 7313
rect 1500 7347 1554 7373
rect 1500 7313 1512 7347
rect 1546 7313 1554 7347
rect 1500 7287 1554 7313
rect 1616 7347 1670 7373
rect 1616 7313 1624 7347
rect 1658 7313 1670 7347
rect 1616 7287 1670 7313
rect 1700 7347 1770 7373
rect 1700 7313 1718 7347
rect 1752 7313 1770 7347
rect 1700 7287 1770 7313
rect 1800 7287 1870 7373
rect 1900 7287 1970 7373
rect 2000 7347 2070 7373
rect 2000 7313 2018 7347
rect 2052 7313 2070 7347
rect 2000 7287 2070 7313
rect 2100 7347 2154 7373
rect 2100 7313 2112 7347
rect 2146 7313 2154 7347
rect 2100 7287 2154 7313
rect 2216 7347 2270 7373
rect 2216 7313 2224 7347
rect 2258 7313 2270 7347
rect 2216 7287 2270 7313
rect 2300 7347 2354 7373
rect 2300 7313 2312 7347
rect 2346 7313 2354 7347
rect 2300 7287 2354 7313
rect 2416 7347 2470 7373
rect 2416 7313 2424 7347
rect 2458 7313 2470 7347
rect 2416 7287 2470 7313
rect 2500 7347 2554 7373
rect 2500 7313 2512 7347
rect 2546 7313 2554 7347
rect 2500 7287 2554 7313
rect 416 7207 470 7233
rect 416 7173 424 7207
rect 458 7173 470 7207
rect 416 7147 470 7173
rect 500 7207 570 7233
rect 500 7173 518 7207
rect 552 7173 570 7207
rect 500 7147 570 7173
rect 600 7207 670 7233
rect 600 7173 618 7207
rect 652 7173 670 7207
rect 600 7147 670 7173
rect 700 7207 770 7233
rect 700 7173 718 7207
rect 752 7173 770 7207
rect 700 7147 770 7173
rect 800 7207 870 7233
rect 800 7173 818 7207
rect 852 7173 870 7207
rect 800 7147 870 7173
rect 900 7207 970 7233
rect 900 7173 918 7207
rect 952 7173 970 7207
rect 900 7147 970 7173
rect 1000 7207 1070 7233
rect 1000 7173 1018 7207
rect 1052 7173 1070 7207
rect 1000 7147 1070 7173
rect 1100 7147 1170 7233
rect 1200 7147 1270 7233
rect 1300 7207 1370 7233
rect 1300 7173 1318 7207
rect 1352 7173 1370 7207
rect 1300 7147 1370 7173
rect 1400 7207 1470 7233
rect 1400 7173 1418 7207
rect 1452 7173 1470 7207
rect 1400 7147 1470 7173
rect 1500 7207 1570 7233
rect 1500 7173 1518 7207
rect 1552 7173 1570 7207
rect 1500 7147 1570 7173
rect 1600 7147 1670 7233
rect 1700 7147 1770 7233
rect 1800 7147 1870 7233
rect 1900 7207 1970 7233
rect 1900 7173 1918 7207
rect 1952 7173 1970 7207
rect 1900 7147 1970 7173
rect 2000 7207 2070 7233
rect 2000 7173 2018 7207
rect 2052 7173 2070 7207
rect 2000 7147 2070 7173
rect 2100 7207 2170 7233
rect 2100 7173 2118 7207
rect 2152 7173 2170 7207
rect 2100 7147 2170 7173
rect 2200 7207 2270 7233
rect 2200 7173 2218 7207
rect 2252 7173 2270 7207
rect 2200 7147 2270 7173
rect 2300 7207 2370 7233
rect 2300 7173 2318 7207
rect 2352 7173 2370 7207
rect 2300 7147 2370 7173
rect 2400 7207 2470 7233
rect 2400 7173 2418 7207
rect 2452 7173 2470 7207
rect 2400 7147 2470 7173
rect 2500 7207 2554 7233
rect 2500 7173 2512 7207
rect 2546 7173 2554 7207
rect 2500 7147 2554 7173
rect 416 7067 470 7093
rect 416 7033 424 7067
rect 458 7033 470 7067
rect 416 7007 470 7033
rect 500 7067 570 7093
rect 500 7033 518 7067
rect 552 7033 570 7067
rect 500 7007 570 7033
rect 600 7067 670 7093
rect 600 7033 618 7067
rect 652 7033 670 7067
rect 600 7007 670 7033
rect 700 7067 770 7093
rect 700 7033 718 7067
rect 752 7033 770 7067
rect 700 7007 770 7033
rect 800 7067 870 7093
rect 800 7033 818 7067
rect 852 7033 870 7067
rect 800 7007 870 7033
rect 900 7067 970 7093
rect 900 7033 918 7067
rect 952 7033 970 7067
rect 900 7007 970 7033
rect 1000 7067 1070 7093
rect 1000 7033 1018 7067
rect 1052 7033 1070 7067
rect 1000 7007 1070 7033
rect 1100 7067 1170 7093
rect 1100 7033 1118 7067
rect 1152 7033 1170 7067
rect 1100 7007 1170 7033
rect 1200 7067 1254 7093
rect 1200 7033 1212 7067
rect 1246 7033 1254 7067
rect 1200 7007 1254 7033
rect 1316 7067 1370 7093
rect 1316 7033 1324 7067
rect 1358 7033 1370 7067
rect 1316 7007 1370 7033
rect 1400 7067 1470 7093
rect 1400 7033 1418 7067
rect 1452 7033 1470 7067
rect 1400 7007 1470 7033
rect 1500 7067 1570 7093
rect 1500 7033 1518 7067
rect 1552 7033 1570 7067
rect 1500 7007 1570 7033
rect 1600 7067 1670 7093
rect 1600 7033 1618 7067
rect 1652 7033 1670 7067
rect 1600 7007 1670 7033
rect 1700 7067 1770 7093
rect 1700 7033 1718 7067
rect 1752 7033 1770 7067
rect 1700 7007 1770 7033
rect 1800 7007 1870 7093
rect 1900 7007 1970 7093
rect 2000 7067 2070 7093
rect 2000 7033 2018 7067
rect 2052 7033 2070 7067
rect 2000 7007 2070 7033
rect 2100 7067 2170 7093
rect 2100 7033 2118 7067
rect 2152 7033 2170 7067
rect 2100 7007 2170 7033
rect 2200 7067 2254 7093
rect 2200 7033 2212 7067
rect 2246 7033 2254 7067
rect 2200 7007 2254 7033
rect 16 6927 70 6953
rect 16 6893 24 6927
rect 58 6893 70 6927
rect 16 6867 70 6893
rect 100 6927 170 6953
rect 100 6893 118 6927
rect 152 6893 170 6927
rect 100 6867 170 6893
rect 200 6927 270 6953
rect 200 6893 218 6927
rect 252 6893 270 6927
rect 200 6867 270 6893
rect 300 6867 370 6953
rect 400 6867 470 6953
rect 500 6867 570 6953
rect 600 6927 670 6953
rect 600 6893 618 6927
rect 652 6893 670 6927
rect 600 6867 670 6893
rect 700 6927 770 6953
rect 700 6893 718 6927
rect 752 6893 770 6927
rect 700 6867 770 6893
rect 800 6867 870 6953
rect 900 6867 970 6953
rect 1000 6867 1070 6953
rect 1100 6927 1170 6953
rect 1100 6893 1118 6927
rect 1152 6893 1170 6927
rect 1100 6867 1170 6893
rect 1200 6927 1270 6953
rect 1200 6893 1218 6927
rect 1252 6893 1270 6927
rect 1200 6867 1270 6893
rect 1300 6927 1370 6953
rect 1300 6893 1318 6927
rect 1352 6893 1370 6927
rect 1300 6867 1370 6893
rect 1400 6927 1454 6953
rect 1400 6893 1412 6927
rect 1446 6893 1454 6927
rect 1400 6867 1454 6893
rect 16 6727 70 6813
rect 100 6727 170 6813
rect 200 6787 270 6813
rect 200 6753 218 6787
rect 252 6753 270 6787
rect 200 6727 270 6753
rect 300 6787 370 6813
rect 300 6753 318 6787
rect 352 6753 370 6787
rect 300 6727 370 6753
rect 400 6727 470 6813
rect 500 6787 570 6813
rect 500 6753 518 6787
rect 552 6753 570 6787
rect 500 6727 570 6753
rect 600 6787 670 6813
rect 600 6753 618 6787
rect 652 6753 670 6787
rect 600 6727 670 6753
rect 700 6787 770 6813
rect 700 6753 718 6787
rect 752 6753 770 6787
rect 700 6727 770 6753
rect 800 6787 870 6813
rect 800 6753 818 6787
rect 852 6753 870 6787
rect 800 6727 870 6753
rect 900 6787 970 6813
rect 900 6753 918 6787
rect 952 6753 970 6787
rect 900 6727 970 6753
rect 1000 6787 1070 6813
rect 1000 6753 1018 6787
rect 1052 6753 1070 6787
rect 1000 6727 1070 6753
rect 1100 6787 1170 6813
rect 1100 6753 1118 6787
rect 1152 6753 1170 6787
rect 1100 6727 1170 6753
rect 1200 6787 1270 6813
rect 1200 6753 1218 6787
rect 1252 6753 1270 6787
rect 1200 6727 1270 6753
rect 1300 6787 1354 6813
rect 1300 6753 1312 6787
rect 1346 6753 1354 6787
rect 1300 6727 1354 6753
rect 16 6647 70 6673
rect 16 6613 24 6647
rect 58 6613 70 6647
rect 16 6587 70 6613
rect 100 6647 170 6673
rect 100 6613 118 6647
rect 152 6613 170 6647
rect 100 6587 170 6613
rect 200 6647 254 6673
rect 200 6613 212 6647
rect 246 6613 254 6647
rect 200 6587 254 6613
rect 316 6647 370 6673
rect 316 6613 324 6647
rect 358 6613 370 6647
rect 316 6587 370 6613
rect 400 6647 470 6673
rect 400 6613 418 6647
rect 452 6613 470 6647
rect 400 6587 470 6613
rect 500 6647 570 6673
rect 500 6613 518 6647
rect 552 6613 570 6647
rect 500 6587 570 6613
rect 600 6587 670 6673
rect 700 6587 770 6673
rect 800 6647 870 6673
rect 800 6613 818 6647
rect 852 6613 870 6647
rect 800 6587 870 6613
rect 900 6647 970 6673
rect 900 6613 918 6647
rect 952 6613 970 6647
rect 900 6587 970 6613
rect 1000 6647 1054 6673
rect 1000 6613 1012 6647
rect 1046 6613 1054 6647
rect 1000 6587 1054 6613
rect 16 6447 70 6533
rect 100 6507 170 6533
rect 100 6473 118 6507
rect 152 6473 170 6507
rect 100 6447 170 6473
rect 200 6507 270 6533
rect 200 6473 218 6507
rect 252 6473 270 6507
rect 200 6447 270 6473
rect 300 6507 370 6533
rect 300 6473 318 6507
rect 352 6473 370 6507
rect 300 6447 370 6473
rect 400 6507 470 6533
rect 400 6473 418 6507
rect 452 6473 470 6507
rect 400 6447 470 6473
rect 500 6507 554 6533
rect 500 6473 512 6507
rect 546 6473 554 6507
rect 500 6447 554 6473
rect 16 6367 70 6393
rect 16 6333 24 6367
rect 58 6333 70 6367
rect 16 6307 70 6333
rect 100 6367 154 6393
rect 100 6333 112 6367
rect 146 6333 154 6367
rect 100 6307 154 6333
rect 1116 6647 1170 6673
rect 1116 6613 1124 6647
rect 1158 6613 1170 6647
rect 1116 6587 1170 6613
rect 1200 6647 1254 6673
rect 1200 6613 1212 6647
rect 1246 6613 1254 6647
rect 1200 6587 1254 6613
rect 1516 6927 1570 6953
rect 1516 6893 1524 6927
rect 1558 6893 1570 6927
rect 1516 6867 1570 6893
rect 1600 6927 1670 6953
rect 1600 6893 1618 6927
rect 1652 6893 1670 6927
rect 1600 6867 1670 6893
rect 1700 6927 1770 6953
rect 1700 6893 1718 6927
rect 1752 6893 1770 6927
rect 1700 6867 1770 6893
rect 1800 6927 1870 6953
rect 1800 6893 1818 6927
rect 1852 6893 1870 6927
rect 1800 6867 1870 6893
rect 1900 6927 1970 6953
rect 1900 6893 1918 6927
rect 1952 6893 1970 6927
rect 1900 6867 1970 6893
rect 2000 6927 2054 6953
rect 2000 6893 2012 6927
rect 2046 6893 2054 6927
rect 2000 6867 2054 6893
rect 1416 6787 1470 6813
rect 1416 6753 1424 6787
rect 1458 6753 1470 6787
rect 1416 6727 1470 6753
rect 1500 6787 1554 6813
rect 1500 6753 1512 6787
rect 1546 6753 1554 6787
rect 1500 6727 1554 6753
rect 3416 7857 3470 7883
rect 3416 7823 3424 7857
rect 3458 7823 3470 7857
rect 3416 7797 3470 7823
rect 3500 7857 3570 7883
rect 3500 7823 3518 7857
rect 3552 7823 3570 7857
rect 3500 7797 3570 7823
rect 3600 7857 3670 7883
rect 3600 7823 3618 7857
rect 3652 7823 3670 7857
rect 3600 7797 3670 7823
rect 3700 7857 3754 7883
rect 3700 7823 3712 7857
rect 3746 7823 3754 7857
rect 3700 7797 3754 7823
rect 3816 7857 3870 7883
rect 3816 7823 3824 7857
rect 3858 7823 3870 7857
rect 3816 7797 3870 7823
rect 3900 7857 3954 7883
rect 3900 7823 3912 7857
rect 3946 7823 3954 7857
rect 3900 7797 3954 7823
rect 4016 7857 4070 7883
rect 4016 7823 4024 7857
rect 4058 7823 4070 7857
rect 4016 7797 4070 7823
rect 4100 7857 4154 7883
rect 4100 7823 4112 7857
rect 4146 7823 4154 7857
rect 4100 7797 4154 7823
rect 2816 7717 2870 7743
rect 2816 7683 2824 7717
rect 2858 7683 2870 7717
rect 2816 7657 2870 7683
rect 2900 7717 2970 7743
rect 2900 7683 2918 7717
rect 2952 7683 2970 7717
rect 2900 7657 2970 7683
rect 3000 7717 3070 7743
rect 3000 7683 3018 7717
rect 3052 7683 3070 7717
rect 3000 7657 3070 7683
rect 3100 7717 3170 7743
rect 3100 7683 3118 7717
rect 3152 7683 3170 7717
rect 3100 7657 3170 7683
rect 3200 7717 3270 7743
rect 3200 7683 3218 7717
rect 3252 7683 3270 7717
rect 3200 7657 3270 7683
rect 3300 7657 3370 7743
rect 3400 7657 3470 7743
rect 3500 7717 3570 7743
rect 3500 7683 3518 7717
rect 3552 7683 3570 7717
rect 3500 7657 3570 7683
rect 3600 7717 3670 7743
rect 3600 7683 3618 7717
rect 3652 7683 3670 7717
rect 3600 7657 3670 7683
rect 3700 7717 3770 7743
rect 3700 7683 3718 7717
rect 3752 7683 3770 7717
rect 3700 7657 3770 7683
rect 3800 7717 3870 7743
rect 3800 7683 3818 7717
rect 3852 7683 3870 7717
rect 3800 7657 3870 7683
rect 3900 7657 3970 7743
rect 4000 7717 4070 7743
rect 4000 7683 4018 7717
rect 4052 7683 4070 7717
rect 4000 7657 4070 7683
rect 4100 7717 4154 7743
rect 4100 7683 4112 7717
rect 4146 7683 4154 7717
rect 4100 7657 4154 7683
rect 2816 7577 2870 7603
rect 2816 7543 2824 7577
rect 2858 7543 2870 7577
rect 2816 7517 2870 7543
rect 2900 7577 2970 7603
rect 2900 7543 2918 7577
rect 2952 7543 2970 7577
rect 2900 7517 2970 7543
rect 3000 7577 3054 7603
rect 3000 7543 3012 7577
rect 3046 7543 3054 7577
rect 3000 7517 3054 7543
rect 3116 7577 3170 7603
rect 3116 7543 3124 7577
rect 3158 7543 3170 7577
rect 3116 7517 3170 7543
rect 3200 7577 3254 7603
rect 3200 7543 3212 7577
rect 3246 7543 3254 7577
rect 3200 7517 3254 7543
rect 3316 7577 3370 7603
rect 3316 7543 3324 7577
rect 3358 7543 3370 7577
rect 3316 7517 3370 7543
rect 3400 7577 3470 7603
rect 3400 7543 3418 7577
rect 3452 7543 3470 7577
rect 3400 7517 3470 7543
rect 3500 7517 3570 7603
rect 3600 7517 3670 7603
rect 3700 7517 3770 7603
rect 3800 7577 3870 7603
rect 3800 7543 3818 7577
rect 3852 7543 3870 7577
rect 3800 7517 3870 7543
rect 3900 7577 3954 7603
rect 3900 7543 3912 7577
rect 3946 7543 3954 7577
rect 3900 7517 3954 7543
rect 4216 7857 4270 7883
rect 4216 7823 4224 7857
rect 4258 7823 4270 7857
rect 4216 7797 4270 7823
rect 4300 7857 4370 7883
rect 4300 7823 4318 7857
rect 4352 7823 4370 7857
rect 4300 7797 4370 7823
rect 4400 7857 4470 7883
rect 4400 7823 4418 7857
rect 4452 7823 4470 7857
rect 4400 7797 4470 7823
rect 4500 7857 4554 7883
rect 4500 7823 4512 7857
rect 4546 7823 4554 7857
rect 4500 7797 4554 7823
rect 4216 7717 4270 7743
rect 4216 7683 4224 7717
rect 4258 7683 4270 7717
rect 4216 7657 4270 7683
rect 4300 7717 4354 7743
rect 4300 7683 4312 7717
rect 4346 7683 4354 7717
rect 4300 7657 4354 7683
rect 4616 7857 4670 7883
rect 4616 7823 4624 7857
rect 4658 7823 4670 7857
rect 4616 7797 4670 7823
rect 4700 7857 4754 7883
rect 4700 7823 4712 7857
rect 4746 7823 4754 7857
rect 4700 7797 4754 7823
rect 4816 7857 4870 7883
rect 4816 7823 4824 7857
rect 4858 7823 4870 7857
rect 4816 7797 4870 7823
rect 4900 7857 4954 7883
rect 4900 7823 4912 7857
rect 4946 7823 4954 7857
rect 4900 7797 4954 7823
rect 5016 7997 5070 8023
rect 5016 7963 5024 7997
rect 5058 7963 5070 7997
rect 5016 7937 5070 7963
rect 5100 7997 5170 8023
rect 5100 7963 5118 7997
rect 5152 7963 5170 7997
rect 5100 7937 5170 7963
rect 5200 7937 5270 8023
rect 5300 7937 5370 8023
rect 5400 7937 5470 8023
rect 5500 7997 5570 8023
rect 5500 7963 5518 7997
rect 5552 7963 5570 7997
rect 5500 7937 5570 7963
rect 5600 7997 5670 8023
rect 5600 7963 5618 7997
rect 5652 7963 5670 7997
rect 5600 7937 5670 7963
rect 5700 7997 5770 8023
rect 5700 7963 5718 7997
rect 5752 7963 5770 7997
rect 5700 7937 5770 7963
rect 5800 7937 5870 8023
rect 5900 7997 5970 8023
rect 5900 7963 5918 7997
rect 5952 7963 5970 7997
rect 5900 7937 5970 7963
rect 6000 7997 6070 8023
rect 6000 7963 6018 7997
rect 6052 7963 6070 7997
rect 6000 7937 6070 7963
rect 6100 7937 6170 8023
rect 6200 7937 6270 8023
rect 6300 7937 6370 8023
rect 6400 7937 6454 8023
rect 6512 8012 6570 8023
rect 6512 7978 6524 8012
rect 6558 7978 6570 8012
rect 6512 7937 6570 7978
rect 6600 7997 6670 8023
rect 6600 7963 6618 7997
rect 6652 7963 6670 7997
rect 6600 7937 6670 7963
rect 6700 7982 6758 8023
rect 6700 7948 6712 7982
rect 6746 7948 6758 7982
rect 6700 7937 6758 7948
rect 6820 7997 6880 8023
rect 6820 7963 6828 7997
rect 6862 7963 6880 7997
rect 6820 7937 6880 7963
rect 6910 7997 6980 8023
rect 6910 7963 6928 7997
rect 6962 7963 6980 7997
rect 6910 7937 6980 7963
rect 7010 7997 7080 8023
rect 7010 7963 7028 7997
rect 7062 7963 7080 7997
rect 7010 7937 7080 7963
rect 7110 7997 7180 8023
rect 7110 7963 7128 7997
rect 7162 7963 7180 7997
rect 7110 7937 7180 7963
rect 7210 7997 7280 8023
rect 7210 7963 7228 7997
rect 7262 7963 7280 7997
rect 7210 7937 7280 7963
rect 7310 7997 7380 8023
rect 7310 7963 7328 7997
rect 7362 7963 7380 7997
rect 7310 7937 7380 7963
rect 7410 7997 7470 8023
rect 7410 7963 7428 7997
rect 7462 7963 7470 7997
rect 7410 7937 7470 7963
rect 5016 7857 5070 7883
rect 5016 7823 5024 7857
rect 5058 7823 5070 7857
rect 5016 7797 5070 7823
rect 5100 7857 5170 7883
rect 5100 7823 5118 7857
rect 5152 7823 5170 7857
rect 5100 7797 5170 7823
rect 5200 7857 5270 7883
rect 5200 7823 5218 7857
rect 5252 7823 5270 7857
rect 5200 7797 5270 7823
rect 5300 7857 5370 7883
rect 5300 7823 5318 7857
rect 5352 7823 5370 7857
rect 5300 7797 5370 7823
rect 5400 7857 5470 7883
rect 5400 7823 5418 7857
rect 5452 7823 5470 7857
rect 5400 7797 5470 7823
rect 5500 7857 5554 7883
rect 5500 7823 5512 7857
rect 5546 7823 5554 7857
rect 5500 7797 5554 7823
rect 4416 7717 4470 7743
rect 4416 7683 4424 7717
rect 4458 7683 4470 7717
rect 4416 7657 4470 7683
rect 4500 7717 4570 7743
rect 4500 7683 4518 7717
rect 4552 7683 4570 7717
rect 4500 7657 4570 7683
rect 4600 7657 4670 7743
rect 4700 7657 4770 7743
rect 4800 7717 4870 7743
rect 4800 7683 4818 7717
rect 4852 7683 4870 7717
rect 4800 7657 4870 7683
rect 4900 7717 4970 7743
rect 4900 7683 4918 7717
rect 4952 7683 4970 7717
rect 4900 7657 4970 7683
rect 5000 7717 5070 7743
rect 5000 7683 5018 7717
rect 5052 7683 5070 7717
rect 5000 7657 5070 7683
rect 5100 7717 5170 7743
rect 5100 7683 5118 7717
rect 5152 7683 5170 7717
rect 5100 7657 5170 7683
rect 5200 7657 5270 7743
rect 5300 7657 5370 7743
rect 5400 7717 5470 7743
rect 5400 7683 5418 7717
rect 5452 7683 5470 7717
rect 5400 7657 5470 7683
rect 5500 7717 5554 7743
rect 5500 7683 5512 7717
rect 5546 7683 5554 7717
rect 5500 7657 5554 7683
rect 4016 7577 4070 7603
rect 4016 7543 4024 7577
rect 4058 7543 4070 7577
rect 4016 7517 4070 7543
rect 4100 7577 4170 7603
rect 4100 7543 4118 7577
rect 4152 7543 4170 7577
rect 4100 7517 4170 7543
rect 4200 7577 4270 7603
rect 4200 7543 4218 7577
rect 4252 7543 4270 7577
rect 4200 7517 4270 7543
rect 4300 7517 4370 7603
rect 4400 7517 4470 7603
rect 4500 7517 4570 7603
rect 4600 7577 4670 7603
rect 4600 7543 4618 7577
rect 4652 7543 4670 7577
rect 4600 7517 4670 7543
rect 4700 7577 4770 7603
rect 4700 7543 4718 7577
rect 4752 7543 4770 7577
rect 4700 7517 4770 7543
rect 4800 7577 4870 7603
rect 4800 7543 4818 7577
rect 4852 7543 4870 7577
rect 4800 7517 4870 7543
rect 4900 7577 4954 7603
rect 4900 7543 4912 7577
rect 4946 7543 4954 7577
rect 4900 7517 4954 7543
rect 5016 7577 5070 7603
rect 5016 7543 5024 7577
rect 5058 7543 5070 7577
rect 5016 7517 5070 7543
rect 5100 7577 5154 7603
rect 5100 7543 5112 7577
rect 5146 7543 5154 7577
rect 5100 7517 5154 7543
rect 5616 7857 5670 7883
rect 5616 7823 5624 7857
rect 5658 7823 5670 7857
rect 5616 7797 5670 7823
rect 5700 7857 5754 7883
rect 5700 7823 5712 7857
rect 5746 7823 5754 7857
rect 5700 7797 5754 7823
rect 5616 7717 5670 7743
rect 5616 7683 5624 7717
rect 5658 7683 5670 7717
rect 5616 7657 5670 7683
rect 5700 7717 5754 7743
rect 5700 7683 5712 7717
rect 5746 7683 5754 7717
rect 5700 7657 5754 7683
rect 5816 7857 5870 7883
rect 5816 7823 5824 7857
rect 5858 7823 5870 7857
rect 5816 7797 5870 7823
rect 5900 7857 5970 7883
rect 5900 7823 5918 7857
rect 5952 7823 5970 7857
rect 5900 7797 5970 7823
rect 6000 7857 6070 7883
rect 6000 7823 6018 7857
rect 6052 7823 6070 7857
rect 6000 7797 6070 7823
rect 6100 7797 6170 7883
rect 6200 7857 6270 7883
rect 6200 7823 6218 7857
rect 6252 7823 6270 7857
rect 6200 7797 6270 7823
rect 6300 7857 6370 7883
rect 6300 7823 6318 7857
rect 6352 7823 6370 7857
rect 6300 7797 6370 7823
rect 6400 7857 6454 7883
rect 6400 7823 6412 7857
rect 6446 7823 6454 7857
rect 6400 7797 6454 7823
rect 6512 7872 6570 7883
rect 6512 7838 6524 7872
rect 6558 7838 6570 7872
rect 6512 7797 6570 7838
rect 6600 7857 6670 7883
rect 6600 7823 6618 7857
rect 6652 7823 6670 7857
rect 6600 7797 6670 7823
rect 6700 7842 6758 7883
rect 6700 7808 6712 7842
rect 6746 7808 6758 7842
rect 6700 7797 6758 7808
rect 6820 7857 6880 7883
rect 6820 7823 6828 7857
rect 6862 7823 6880 7857
rect 6820 7797 6880 7823
rect 6910 7857 6980 7883
rect 6910 7823 6928 7857
rect 6962 7823 6980 7857
rect 6910 7797 6980 7823
rect 7010 7857 7080 7883
rect 7010 7823 7028 7857
rect 7062 7823 7080 7857
rect 7010 7797 7080 7823
rect 7110 7857 7180 7883
rect 7110 7823 7128 7857
rect 7162 7823 7180 7857
rect 7110 7797 7180 7823
rect 7210 7857 7280 7883
rect 7210 7823 7228 7857
rect 7262 7823 7280 7857
rect 7210 7797 7280 7823
rect 7310 7857 7380 7883
rect 7310 7823 7328 7857
rect 7362 7823 7380 7857
rect 7310 7797 7380 7823
rect 7410 7857 7470 7883
rect 7410 7823 7428 7857
rect 7462 7823 7470 7857
rect 7410 7797 7470 7823
rect 5816 7717 5870 7743
rect 5816 7683 5824 7717
rect 5858 7683 5870 7717
rect 5816 7657 5870 7683
rect 5900 7717 5970 7743
rect 5900 7683 5918 7717
rect 5952 7683 5970 7717
rect 5900 7657 5970 7683
rect 6000 7657 6070 7743
rect 6100 7717 6170 7743
rect 6100 7683 6118 7717
rect 6152 7683 6170 7717
rect 6100 7657 6170 7683
rect 6200 7717 6270 7743
rect 6200 7683 6218 7717
rect 6252 7683 6270 7717
rect 6200 7657 6270 7683
rect 6300 7717 6370 7743
rect 6300 7683 6318 7717
rect 6352 7683 6370 7717
rect 6300 7657 6370 7683
rect 6400 7657 6454 7743
rect 6512 7732 6570 7743
rect 6512 7698 6524 7732
rect 6558 7698 6570 7732
rect 6512 7657 6570 7698
rect 6600 7717 6670 7743
rect 6600 7683 6618 7717
rect 6652 7683 6670 7717
rect 6600 7657 6670 7683
rect 6700 7702 6758 7743
rect 6700 7668 6712 7702
rect 6746 7668 6758 7702
rect 6700 7657 6758 7668
rect 6820 7717 6880 7743
rect 6820 7683 6828 7717
rect 6862 7683 6880 7717
rect 6820 7657 6880 7683
rect 6910 7717 6980 7743
rect 6910 7683 6928 7717
rect 6962 7683 6980 7717
rect 6910 7657 6980 7683
rect 7010 7717 7080 7743
rect 7010 7683 7028 7717
rect 7062 7683 7080 7717
rect 7010 7657 7080 7683
rect 7110 7717 7180 7743
rect 7110 7683 7128 7717
rect 7162 7683 7180 7717
rect 7110 7657 7180 7683
rect 7210 7717 7280 7743
rect 7210 7683 7228 7717
rect 7262 7683 7280 7717
rect 7210 7657 7280 7683
rect 7310 7717 7380 7743
rect 7310 7683 7328 7717
rect 7362 7683 7380 7717
rect 7310 7657 7380 7683
rect 7410 7717 7470 7743
rect 7410 7683 7428 7717
rect 7462 7683 7470 7717
rect 7410 7657 7470 7683
rect 5216 7577 5270 7603
rect 5216 7543 5224 7577
rect 5258 7543 5270 7577
rect 5216 7517 5270 7543
rect 5300 7577 5370 7603
rect 5300 7543 5318 7577
rect 5352 7543 5370 7577
rect 5300 7517 5370 7543
rect 5400 7577 5470 7603
rect 5400 7543 5418 7577
rect 5452 7543 5470 7577
rect 5400 7517 5470 7543
rect 5500 7577 5570 7603
rect 5500 7543 5518 7577
rect 5552 7543 5570 7577
rect 5500 7517 5570 7543
rect 5600 7577 5670 7603
rect 5600 7543 5618 7577
rect 5652 7543 5670 7577
rect 5600 7517 5670 7543
rect 5700 7577 5770 7603
rect 5700 7543 5718 7577
rect 5752 7543 5770 7577
rect 5700 7517 5770 7543
rect 5800 7577 5870 7603
rect 5800 7543 5818 7577
rect 5852 7543 5870 7577
rect 5800 7517 5870 7543
rect 5900 7577 5970 7603
rect 5900 7543 5918 7577
rect 5952 7543 5970 7577
rect 5900 7517 5970 7543
rect 6000 7577 6070 7603
rect 6000 7543 6018 7577
rect 6052 7543 6070 7577
rect 6000 7517 6070 7543
rect 6100 7577 6170 7603
rect 6100 7543 6118 7577
rect 6152 7543 6170 7577
rect 6100 7517 6170 7543
rect 6200 7517 6270 7603
rect 6300 7577 6370 7603
rect 6300 7543 6318 7577
rect 6352 7543 6370 7577
rect 6300 7517 6370 7543
rect 6400 7577 6454 7603
rect 6400 7543 6412 7577
rect 6446 7543 6454 7577
rect 6400 7517 6454 7543
rect 6512 7592 6570 7603
rect 6512 7558 6524 7592
rect 6558 7558 6570 7592
rect 6512 7517 6570 7558
rect 6600 7577 6670 7603
rect 6600 7543 6618 7577
rect 6652 7543 6670 7577
rect 6600 7517 6670 7543
rect 6700 7562 6758 7603
rect 6700 7528 6712 7562
rect 6746 7528 6758 7562
rect 6700 7517 6758 7528
rect 6820 7577 6880 7603
rect 6820 7543 6828 7577
rect 6862 7543 6880 7577
rect 6820 7517 6880 7543
rect 6910 7577 6980 7603
rect 6910 7543 6928 7577
rect 6962 7543 6980 7577
rect 6910 7517 6980 7543
rect 7010 7577 7080 7603
rect 7010 7543 7028 7577
rect 7062 7543 7080 7577
rect 7010 7517 7080 7543
rect 7110 7577 7180 7603
rect 7110 7543 7128 7577
rect 7162 7543 7180 7577
rect 7110 7517 7180 7543
rect 7210 7577 7280 7603
rect 7210 7543 7228 7577
rect 7262 7543 7280 7577
rect 7210 7517 7280 7543
rect 7310 7577 7380 7603
rect 7310 7543 7328 7577
rect 7362 7543 7380 7577
rect 7310 7517 7380 7543
rect 7410 7577 7470 7603
rect 7410 7543 7428 7577
rect 7462 7543 7470 7577
rect 7410 7517 7470 7543
rect 2616 7347 2670 7373
rect 2616 7313 2624 7347
rect 2658 7313 2670 7347
rect 2616 7287 2670 7313
rect 2700 7347 2770 7373
rect 2700 7313 2718 7347
rect 2752 7313 2770 7347
rect 2700 7287 2770 7313
rect 2800 7347 2870 7373
rect 2800 7313 2818 7347
rect 2852 7313 2870 7347
rect 2800 7287 2870 7313
rect 2900 7347 2970 7373
rect 2900 7313 2918 7347
rect 2952 7313 2970 7347
rect 2900 7287 2970 7313
rect 3000 7347 3070 7373
rect 3000 7313 3018 7347
rect 3052 7313 3070 7347
rect 3000 7287 3070 7313
rect 3100 7287 3170 7373
rect 3200 7347 3270 7373
rect 3200 7313 3218 7347
rect 3252 7313 3270 7347
rect 3200 7287 3270 7313
rect 3300 7347 3370 7373
rect 3300 7313 3318 7347
rect 3352 7313 3370 7347
rect 3300 7287 3370 7313
rect 3400 7347 3470 7373
rect 3400 7313 3418 7347
rect 3452 7313 3470 7347
rect 3400 7287 3470 7313
rect 3500 7287 3570 7373
rect 3600 7347 3670 7373
rect 3600 7313 3618 7347
rect 3652 7313 3670 7347
rect 3600 7287 3670 7313
rect 3700 7347 3770 7373
rect 3700 7313 3718 7347
rect 3752 7313 3770 7347
rect 3700 7287 3770 7313
rect 3800 7347 3870 7373
rect 3800 7313 3818 7347
rect 3852 7313 3870 7347
rect 3800 7287 3870 7313
rect 3900 7287 3970 7373
rect 4000 7347 4070 7373
rect 4000 7313 4018 7347
rect 4052 7313 4070 7347
rect 4000 7287 4070 7313
rect 4100 7347 4170 7373
rect 4100 7313 4118 7347
rect 4152 7313 4170 7347
rect 4100 7287 4170 7313
rect 4200 7287 4270 7373
rect 4300 7287 4370 7373
rect 4400 7287 4470 7373
rect 4500 7347 4570 7373
rect 4500 7313 4518 7347
rect 4552 7313 4570 7347
rect 4500 7287 4570 7313
rect 4600 7347 4670 7373
rect 4600 7313 4618 7347
rect 4652 7313 4670 7347
rect 4600 7287 4670 7313
rect 4700 7347 4770 7373
rect 4700 7313 4718 7347
rect 4752 7313 4770 7347
rect 4700 7287 4770 7313
rect 4800 7347 4870 7373
rect 4800 7313 4818 7347
rect 4852 7313 4870 7347
rect 4800 7287 4870 7313
rect 4900 7347 4970 7373
rect 4900 7313 4918 7347
rect 4952 7313 4970 7347
rect 4900 7287 4970 7313
rect 5000 7347 5070 7373
rect 5000 7313 5018 7347
rect 5052 7313 5070 7347
rect 5000 7287 5070 7313
rect 5100 7287 5170 7373
rect 5200 7347 5270 7373
rect 5200 7313 5218 7347
rect 5252 7313 5270 7347
rect 5200 7287 5270 7313
rect 5300 7347 5370 7373
rect 5300 7313 5318 7347
rect 5352 7313 5370 7347
rect 5300 7287 5370 7313
rect 5400 7287 5470 7373
rect 5500 7287 5570 7373
rect 5600 7347 5670 7373
rect 5600 7313 5618 7347
rect 5652 7313 5670 7347
rect 5600 7287 5670 7313
rect 5700 7347 5770 7373
rect 5700 7313 5718 7347
rect 5752 7313 5770 7347
rect 5700 7287 5770 7313
rect 5800 7287 5870 7373
rect 5900 7287 5970 7373
rect 6000 7287 6070 7373
rect 6100 7287 6170 7373
rect 6200 7287 6270 7373
rect 6300 7287 6370 7373
rect 6400 7287 6454 7373
rect 6512 7362 6570 7373
rect 6512 7328 6524 7362
rect 6558 7328 6570 7362
rect 6512 7287 6570 7328
rect 6600 7347 6670 7373
rect 6600 7313 6618 7347
rect 6652 7313 6670 7347
rect 6600 7287 6670 7313
rect 6700 7332 6758 7373
rect 6700 7298 6712 7332
rect 6746 7298 6758 7332
rect 6700 7287 6758 7298
rect 6820 7347 6880 7373
rect 6820 7313 6828 7347
rect 6862 7313 6880 7347
rect 6820 7287 6880 7313
rect 6910 7347 6980 7373
rect 6910 7313 6928 7347
rect 6962 7313 6980 7347
rect 6910 7287 6980 7313
rect 7010 7347 7080 7373
rect 7010 7313 7028 7347
rect 7062 7313 7080 7347
rect 7010 7287 7080 7313
rect 7110 7347 7180 7373
rect 7110 7313 7128 7347
rect 7162 7313 7180 7347
rect 7110 7287 7180 7313
rect 7210 7347 7280 7373
rect 7210 7313 7228 7347
rect 7262 7313 7280 7347
rect 7210 7287 7280 7313
rect 7310 7347 7380 7373
rect 7310 7313 7328 7347
rect 7362 7313 7380 7347
rect 7310 7287 7380 7313
rect 7410 7347 7470 7373
rect 7410 7313 7428 7347
rect 7462 7313 7470 7347
rect 7410 7287 7470 7313
rect 2616 7207 2670 7233
rect 2616 7173 2624 7207
rect 2658 7173 2670 7207
rect 2616 7147 2670 7173
rect 2700 7207 2770 7233
rect 2700 7173 2718 7207
rect 2752 7173 2770 7207
rect 2700 7147 2770 7173
rect 2800 7207 2870 7233
rect 2800 7173 2818 7207
rect 2852 7173 2870 7207
rect 2800 7147 2870 7173
rect 2900 7207 2954 7233
rect 2900 7173 2912 7207
rect 2946 7173 2954 7207
rect 2900 7147 2954 7173
rect 3016 7207 3070 7233
rect 3016 7173 3024 7207
rect 3058 7173 3070 7207
rect 3016 7147 3070 7173
rect 3100 7207 3170 7233
rect 3100 7173 3118 7207
rect 3152 7173 3170 7207
rect 3100 7147 3170 7173
rect 3200 7207 3254 7233
rect 3200 7173 3212 7207
rect 3246 7173 3254 7207
rect 3200 7147 3254 7173
rect 2316 7067 2370 7093
rect 2316 7033 2324 7067
rect 2358 7033 2370 7067
rect 2316 7007 2370 7033
rect 2400 7067 2470 7093
rect 2400 7033 2418 7067
rect 2452 7033 2470 7067
rect 2400 7007 2470 7033
rect 2500 7067 2570 7093
rect 2500 7033 2518 7067
rect 2552 7033 2570 7067
rect 2500 7007 2570 7033
rect 2600 7067 2670 7093
rect 2600 7033 2618 7067
rect 2652 7033 2670 7067
rect 2600 7007 2670 7033
rect 2700 7067 2770 7093
rect 2700 7033 2718 7067
rect 2752 7033 2770 7067
rect 2700 7007 2770 7033
rect 2800 7067 2870 7093
rect 2800 7033 2818 7067
rect 2852 7033 2870 7067
rect 2800 7007 2870 7033
rect 2900 7067 2970 7093
rect 2900 7033 2918 7067
rect 2952 7033 2970 7067
rect 2900 7007 2970 7033
rect 3000 7067 3054 7093
rect 3000 7033 3012 7067
rect 3046 7033 3054 7067
rect 3000 7007 3054 7033
rect 2116 6927 2170 6953
rect 2116 6893 2124 6927
rect 2158 6893 2170 6927
rect 2116 6867 2170 6893
rect 2200 6927 2270 6953
rect 2200 6893 2218 6927
rect 2252 6893 2270 6927
rect 2200 6867 2270 6893
rect 2300 6927 2370 6953
rect 2300 6893 2318 6927
rect 2352 6893 2370 6927
rect 2300 6867 2370 6893
rect 2400 6867 2470 6953
rect 2500 6867 2570 6953
rect 2600 6867 2670 6953
rect 2700 6927 2770 6953
rect 2700 6893 2718 6927
rect 2752 6893 2770 6927
rect 2700 6867 2770 6893
rect 2800 6927 2870 6953
rect 2800 6893 2818 6927
rect 2852 6893 2870 6927
rect 2800 6867 2870 6893
rect 2900 6927 2954 6953
rect 2900 6893 2912 6927
rect 2946 6893 2954 6927
rect 2900 6867 2954 6893
rect 1616 6787 1670 6813
rect 1616 6753 1624 6787
rect 1658 6753 1670 6787
rect 1616 6727 1670 6753
rect 1700 6787 1770 6813
rect 1700 6753 1718 6787
rect 1752 6753 1770 6787
rect 1700 6727 1770 6753
rect 1800 6727 1870 6813
rect 1900 6787 1970 6813
rect 1900 6753 1918 6787
rect 1952 6753 1970 6787
rect 1900 6727 1970 6753
rect 2000 6787 2070 6813
rect 2000 6753 2018 6787
rect 2052 6753 2070 6787
rect 2000 6727 2070 6753
rect 2100 6787 2154 6813
rect 2100 6753 2112 6787
rect 2146 6753 2154 6787
rect 2100 6727 2154 6753
rect 3316 7207 3370 7233
rect 3316 7173 3324 7207
rect 3358 7173 3370 7207
rect 3316 7147 3370 7173
rect 3400 7207 3470 7233
rect 3400 7173 3418 7207
rect 3452 7173 3470 7207
rect 3400 7147 3470 7173
rect 3500 7147 3570 7233
rect 3600 7147 3670 7233
rect 3700 7147 3770 7233
rect 3800 7207 3870 7233
rect 3800 7173 3818 7207
rect 3852 7173 3870 7207
rect 3800 7147 3870 7173
rect 3900 7207 3970 7233
rect 3900 7173 3918 7207
rect 3952 7173 3970 7207
rect 3900 7147 3970 7173
rect 4000 7207 4070 7233
rect 4000 7173 4018 7207
rect 4052 7173 4070 7207
rect 4000 7147 4070 7173
rect 4100 7147 4170 7233
rect 4200 7207 4270 7233
rect 4200 7173 4218 7207
rect 4252 7173 4270 7207
rect 4200 7147 4270 7173
rect 4300 7207 4354 7233
rect 4300 7173 4312 7207
rect 4346 7173 4354 7207
rect 4300 7147 4354 7173
rect 3116 7067 3170 7093
rect 3116 7033 3124 7067
rect 3158 7033 3170 7067
rect 3116 7007 3170 7033
rect 3200 7067 3270 7093
rect 3200 7033 3218 7067
rect 3252 7033 3270 7067
rect 3200 7007 3270 7033
rect 3300 7067 3370 7093
rect 3300 7033 3318 7067
rect 3352 7033 3370 7067
rect 3300 7007 3370 7033
rect 3400 7067 3454 7093
rect 3400 7033 3412 7067
rect 3446 7033 3454 7067
rect 3400 7007 3454 7033
rect 3016 6927 3070 6953
rect 3016 6893 3024 6927
rect 3058 6893 3070 6927
rect 3016 6867 3070 6893
rect 3100 6927 3154 6953
rect 3100 6893 3112 6927
rect 3146 6893 3154 6927
rect 3100 6867 3154 6893
rect 3216 6927 3270 6953
rect 3216 6893 3224 6927
rect 3258 6893 3270 6927
rect 3216 6867 3270 6893
rect 3300 6927 3370 6953
rect 3300 6893 3318 6927
rect 3352 6893 3370 6927
rect 3300 6867 3370 6893
rect 3400 6927 3454 6953
rect 3400 6893 3412 6927
rect 3446 6893 3454 6927
rect 3400 6867 3454 6893
rect 3516 7067 3570 7093
rect 3516 7033 3524 7067
rect 3558 7033 3570 7067
rect 3516 7007 3570 7033
rect 3600 7067 3670 7093
rect 3600 7033 3618 7067
rect 3652 7033 3670 7067
rect 3600 7007 3670 7033
rect 3700 7067 3770 7093
rect 3700 7033 3718 7067
rect 3752 7033 3770 7067
rect 3700 7007 3770 7033
rect 3800 7067 3870 7093
rect 3800 7033 3818 7067
rect 3852 7033 3870 7067
rect 3800 7007 3870 7033
rect 3900 7067 3970 7093
rect 3900 7033 3918 7067
rect 3952 7033 3970 7067
rect 3900 7007 3970 7033
rect 4000 7067 4054 7093
rect 4000 7033 4012 7067
rect 4046 7033 4054 7067
rect 4000 7007 4054 7033
rect 4416 7207 4470 7233
rect 4416 7173 4424 7207
rect 4458 7173 4470 7207
rect 4416 7147 4470 7173
rect 4500 7207 4570 7233
rect 4500 7173 4518 7207
rect 4552 7173 4570 7207
rect 4500 7147 4570 7173
rect 4600 7207 4654 7233
rect 4600 7173 4612 7207
rect 4646 7173 4654 7207
rect 4600 7147 4654 7173
rect 4716 7207 4770 7233
rect 4716 7173 4724 7207
rect 4758 7173 4770 7207
rect 4716 7147 4770 7173
rect 4800 7207 4870 7233
rect 4800 7173 4818 7207
rect 4852 7173 4870 7207
rect 4800 7147 4870 7173
rect 4900 7207 4970 7233
rect 4900 7173 4918 7207
rect 4952 7173 4970 7207
rect 4900 7147 4970 7173
rect 5000 7207 5054 7233
rect 5000 7173 5012 7207
rect 5046 7173 5054 7207
rect 5000 7147 5054 7173
rect 5116 7207 5170 7233
rect 5116 7173 5124 7207
rect 5158 7173 5170 7207
rect 5116 7147 5170 7173
rect 5200 7207 5270 7233
rect 5200 7173 5218 7207
rect 5252 7173 5270 7207
rect 5200 7147 5270 7173
rect 5300 7147 5370 7233
rect 5400 7147 5470 7233
rect 5500 7147 5570 7233
rect 5600 7207 5670 7233
rect 5600 7173 5618 7207
rect 5652 7173 5670 7207
rect 5600 7147 5670 7173
rect 5700 7207 5770 7233
rect 5700 7173 5718 7207
rect 5752 7173 5770 7207
rect 5700 7147 5770 7173
rect 5800 7147 5870 7233
rect 5900 7207 5970 7233
rect 5900 7173 5918 7207
rect 5952 7173 5970 7207
rect 5900 7147 5970 7173
rect 6000 7207 6054 7233
rect 6000 7173 6012 7207
rect 6046 7173 6054 7207
rect 6000 7147 6054 7173
rect 4116 7067 4170 7093
rect 4116 7033 4124 7067
rect 4158 7033 4170 7067
rect 4116 7007 4170 7033
rect 4200 7067 4270 7093
rect 4200 7033 4218 7067
rect 4252 7033 4270 7067
rect 4200 7007 4270 7033
rect 4300 7067 4370 7093
rect 4300 7033 4318 7067
rect 4352 7033 4370 7067
rect 4300 7007 4370 7033
rect 4400 7007 4470 7093
rect 4500 7007 4570 7093
rect 4600 7067 4670 7093
rect 4600 7033 4618 7067
rect 4652 7033 4670 7067
rect 4600 7007 4670 7033
rect 4700 7067 4770 7093
rect 4700 7033 4718 7067
rect 4752 7033 4770 7067
rect 4700 7007 4770 7033
rect 4800 7007 4870 7093
rect 4900 7007 4970 7093
rect 5000 7067 5070 7093
rect 5000 7033 5018 7067
rect 5052 7033 5070 7067
rect 5000 7007 5070 7033
rect 5100 7067 5154 7093
rect 5100 7033 5112 7067
rect 5146 7033 5154 7067
rect 5100 7007 5154 7033
rect 3516 6927 3570 6953
rect 3516 6893 3524 6927
rect 3558 6893 3570 6927
rect 3516 6867 3570 6893
rect 3600 6927 3670 6953
rect 3600 6893 3618 6927
rect 3652 6893 3670 6927
rect 3600 6867 3670 6893
rect 3700 6867 3770 6953
rect 3800 6867 3870 6953
rect 3900 6927 3970 6953
rect 3900 6893 3918 6927
rect 3952 6893 3970 6927
rect 3900 6867 3970 6893
rect 4000 6927 4070 6953
rect 4000 6893 4018 6927
rect 4052 6893 4070 6927
rect 4000 6867 4070 6893
rect 4100 6927 4170 6953
rect 4100 6893 4118 6927
rect 4152 6893 4170 6927
rect 4100 6867 4170 6893
rect 4200 6927 4254 6953
rect 4200 6893 4212 6927
rect 4246 6893 4254 6927
rect 4200 6867 4254 6893
rect 4316 6927 4370 6953
rect 4316 6893 4324 6927
rect 4358 6893 4370 6927
rect 4316 6867 4370 6893
rect 4400 6927 4470 6953
rect 4400 6893 4418 6927
rect 4452 6893 4470 6927
rect 4400 6867 4470 6893
rect 4500 6927 4570 6953
rect 4500 6893 4518 6927
rect 4552 6893 4570 6927
rect 4500 6867 4570 6893
rect 4600 6927 4670 6953
rect 4600 6893 4618 6927
rect 4652 6893 4670 6927
rect 4600 6867 4670 6893
rect 4700 6927 4770 6953
rect 4700 6893 4718 6927
rect 4752 6893 4770 6927
rect 4700 6867 4770 6893
rect 4800 6927 4854 6953
rect 4800 6893 4812 6927
rect 4846 6893 4854 6927
rect 4800 6867 4854 6893
rect 4916 6927 4970 6953
rect 4916 6893 4924 6927
rect 4958 6893 4970 6927
rect 4916 6867 4970 6893
rect 5000 6927 5070 6953
rect 5000 6893 5018 6927
rect 5052 6893 5070 6927
rect 5000 6867 5070 6893
rect 5100 6927 5154 6953
rect 5100 6893 5112 6927
rect 5146 6893 5154 6927
rect 5100 6867 5154 6893
rect 6116 7207 6170 7233
rect 6116 7173 6124 7207
rect 6158 7173 6170 7207
rect 6116 7147 6170 7173
rect 6200 7207 6270 7233
rect 6200 7173 6218 7207
rect 6252 7173 6270 7207
rect 6200 7147 6270 7173
rect 6300 7207 6370 7233
rect 6300 7173 6318 7207
rect 6352 7173 6370 7207
rect 6300 7147 6370 7173
rect 6400 7207 6454 7233
rect 6400 7173 6412 7207
rect 6446 7173 6454 7207
rect 6400 7147 6454 7173
rect 6512 7222 6570 7233
rect 6512 7188 6524 7222
rect 6558 7188 6570 7222
rect 6512 7147 6570 7188
rect 6600 7207 6670 7233
rect 6600 7173 6618 7207
rect 6652 7173 6670 7207
rect 6600 7147 6670 7173
rect 6700 7192 6758 7233
rect 6700 7158 6712 7192
rect 6746 7158 6758 7192
rect 6700 7147 6758 7158
rect 6820 7207 6880 7233
rect 6820 7173 6828 7207
rect 6862 7173 6880 7207
rect 6820 7147 6880 7173
rect 6910 7207 6980 7233
rect 6910 7173 6928 7207
rect 6962 7173 6980 7207
rect 6910 7147 6980 7173
rect 7010 7207 7080 7233
rect 7010 7173 7028 7207
rect 7062 7173 7080 7207
rect 7010 7147 7080 7173
rect 7110 7207 7180 7233
rect 7110 7173 7128 7207
rect 7162 7173 7180 7207
rect 7110 7147 7180 7173
rect 7210 7207 7280 7233
rect 7210 7173 7228 7207
rect 7262 7173 7280 7207
rect 7210 7147 7280 7173
rect 7310 7207 7380 7233
rect 7310 7173 7328 7207
rect 7362 7173 7380 7207
rect 7310 7147 7380 7173
rect 7410 7207 7470 7233
rect 7410 7173 7428 7207
rect 7462 7173 7470 7207
rect 7410 7147 7470 7173
rect 5216 7067 5270 7093
rect 5216 7033 5224 7067
rect 5258 7033 5270 7067
rect 5216 7007 5270 7033
rect 5300 7067 5370 7093
rect 5300 7033 5318 7067
rect 5352 7033 5370 7067
rect 5300 7007 5370 7033
rect 5400 7067 5470 7093
rect 5400 7033 5418 7067
rect 5452 7033 5470 7067
rect 5400 7007 5470 7033
rect 5500 7067 5570 7093
rect 5500 7033 5518 7067
rect 5552 7033 5570 7067
rect 5500 7007 5570 7033
rect 5600 7067 5670 7093
rect 5600 7033 5618 7067
rect 5652 7033 5670 7067
rect 5600 7007 5670 7033
rect 5700 7067 5770 7093
rect 5700 7033 5718 7067
rect 5752 7033 5770 7067
rect 5700 7007 5770 7033
rect 5800 7067 5870 7093
rect 5800 7033 5818 7067
rect 5852 7033 5870 7067
rect 5800 7007 5870 7033
rect 5900 7007 5970 7093
rect 6000 7067 6070 7093
rect 6000 7033 6018 7067
rect 6052 7033 6070 7067
rect 6000 7007 6070 7033
rect 6100 7067 6154 7093
rect 6100 7033 6112 7067
rect 6146 7033 6154 7067
rect 6100 7007 6154 7033
rect 5216 6927 5270 6953
rect 5216 6893 5224 6927
rect 5258 6893 5270 6927
rect 5216 6867 5270 6893
rect 5300 6927 5354 6953
rect 5300 6893 5312 6927
rect 5346 6893 5354 6927
rect 5300 6867 5354 6893
rect 5416 6927 5470 6953
rect 5416 6893 5424 6927
rect 5458 6893 5470 6927
rect 5416 6867 5470 6893
rect 5500 6927 5570 6953
rect 5500 6893 5518 6927
rect 5552 6893 5570 6927
rect 5500 6867 5570 6893
rect 5600 6867 5670 6953
rect 5700 6927 5770 6953
rect 5700 6893 5718 6927
rect 5752 6893 5770 6927
rect 5700 6867 5770 6893
rect 5800 6927 5870 6953
rect 5800 6893 5818 6927
rect 5852 6893 5870 6927
rect 5800 6867 5870 6893
rect 5900 6867 5970 6953
rect 6000 6927 6070 6953
rect 6000 6893 6018 6927
rect 6052 6893 6070 6927
rect 6000 6867 6070 6893
rect 6100 6927 6154 6953
rect 6100 6893 6112 6927
rect 6146 6893 6154 6927
rect 6100 6867 6154 6893
rect 2216 6787 2270 6813
rect 2216 6753 2224 6787
rect 2258 6753 2270 6787
rect 2216 6727 2270 6753
rect 2300 6787 2370 6813
rect 2300 6753 2318 6787
rect 2352 6753 2370 6787
rect 2300 6727 2370 6753
rect 2400 6727 2470 6813
rect 2500 6727 2570 6813
rect 2600 6727 2670 6813
rect 2700 6727 2770 6813
rect 2800 6787 2870 6813
rect 2800 6753 2818 6787
rect 2852 6753 2870 6787
rect 2800 6727 2870 6753
rect 2900 6787 2970 6813
rect 2900 6753 2918 6787
rect 2952 6753 2970 6787
rect 2900 6727 2970 6753
rect 3000 6727 3070 6813
rect 3100 6727 3170 6813
rect 3200 6727 3270 6813
rect 3300 6727 3370 6813
rect 3400 6727 3470 6813
rect 3500 6727 3570 6813
rect 3600 6727 3670 6813
rect 3700 6727 3770 6813
rect 3800 6727 3870 6813
rect 3900 6727 3970 6813
rect 4000 6787 4070 6813
rect 4000 6753 4018 6787
rect 4052 6753 4070 6787
rect 4000 6727 4070 6753
rect 4100 6787 4170 6813
rect 4100 6753 4118 6787
rect 4152 6753 4170 6787
rect 4100 6727 4170 6753
rect 4200 6727 4270 6813
rect 4300 6787 4370 6813
rect 4300 6753 4318 6787
rect 4352 6753 4370 6787
rect 4300 6727 4370 6753
rect 4400 6787 4470 6813
rect 4400 6753 4418 6787
rect 4452 6753 4470 6787
rect 4400 6727 4470 6753
rect 4500 6787 4570 6813
rect 4500 6753 4518 6787
rect 4552 6753 4570 6787
rect 4500 6727 4570 6753
rect 4600 6727 4670 6813
rect 4700 6787 4770 6813
rect 4700 6753 4718 6787
rect 4752 6753 4770 6787
rect 4700 6727 4770 6753
rect 4800 6787 4870 6813
rect 4800 6753 4818 6787
rect 4852 6753 4870 6787
rect 4800 6727 4870 6753
rect 4900 6787 4970 6813
rect 4900 6753 4918 6787
rect 4952 6753 4970 6787
rect 4900 6727 4970 6753
rect 5000 6787 5070 6813
rect 5000 6753 5018 6787
rect 5052 6753 5070 6787
rect 5000 6727 5070 6753
rect 5100 6787 5170 6813
rect 5100 6753 5118 6787
rect 5152 6753 5170 6787
rect 5100 6727 5170 6753
rect 5200 6727 5270 6813
rect 5300 6787 5370 6813
rect 5300 6753 5318 6787
rect 5352 6753 5370 6787
rect 5300 6727 5370 6753
rect 5400 6787 5454 6813
rect 5400 6753 5412 6787
rect 5446 6753 5454 6787
rect 5400 6727 5454 6753
rect 1316 6647 1370 6673
rect 1316 6613 1324 6647
rect 1358 6613 1370 6647
rect 1316 6587 1370 6613
rect 1400 6647 1470 6673
rect 1400 6613 1418 6647
rect 1452 6613 1470 6647
rect 1400 6587 1470 6613
rect 1500 6587 1570 6673
rect 1600 6587 1670 6673
rect 1700 6587 1770 6673
rect 1800 6647 1870 6673
rect 1800 6613 1818 6647
rect 1852 6613 1870 6647
rect 1800 6587 1870 6613
rect 1900 6647 1970 6673
rect 1900 6613 1918 6647
rect 1952 6613 1970 6647
rect 1900 6587 1970 6613
rect 2000 6647 2070 6673
rect 2000 6613 2018 6647
rect 2052 6613 2070 6647
rect 2000 6587 2070 6613
rect 2100 6647 2170 6673
rect 2100 6613 2118 6647
rect 2152 6613 2170 6647
rect 2100 6587 2170 6613
rect 2200 6647 2270 6673
rect 2200 6613 2218 6647
rect 2252 6613 2270 6647
rect 2200 6587 2270 6613
rect 2300 6647 2370 6673
rect 2300 6613 2318 6647
rect 2352 6613 2370 6647
rect 2300 6587 2370 6613
rect 2400 6587 2470 6673
rect 2500 6647 2570 6673
rect 2500 6613 2518 6647
rect 2552 6613 2570 6647
rect 2500 6587 2570 6613
rect 2600 6647 2670 6673
rect 2600 6613 2618 6647
rect 2652 6613 2670 6647
rect 2600 6587 2670 6613
rect 2700 6587 2770 6673
rect 2800 6587 2870 6673
rect 2900 6587 2970 6673
rect 3000 6647 3070 6673
rect 3000 6613 3018 6647
rect 3052 6613 3070 6647
rect 3000 6587 3070 6613
rect 3100 6647 3170 6673
rect 3100 6613 3118 6647
rect 3152 6613 3170 6647
rect 3100 6587 3170 6613
rect 3200 6587 3270 6673
rect 3300 6647 3370 6673
rect 3300 6613 3318 6647
rect 3352 6613 3370 6647
rect 3300 6587 3370 6613
rect 3400 6647 3454 6673
rect 3400 6613 3412 6647
rect 3446 6613 3454 6647
rect 3400 6587 3454 6613
rect 616 6507 670 6533
rect 616 6473 624 6507
rect 658 6473 670 6507
rect 616 6447 670 6473
rect 700 6507 770 6533
rect 700 6473 718 6507
rect 752 6473 770 6507
rect 700 6447 770 6473
rect 800 6507 870 6533
rect 800 6473 818 6507
rect 852 6473 870 6507
rect 800 6447 870 6473
rect 900 6507 970 6533
rect 900 6473 918 6507
rect 952 6473 970 6507
rect 900 6447 970 6473
rect 1000 6507 1070 6533
rect 1000 6473 1018 6507
rect 1052 6473 1070 6507
rect 1000 6447 1070 6473
rect 1100 6507 1170 6533
rect 1100 6473 1118 6507
rect 1152 6473 1170 6507
rect 1100 6447 1170 6473
rect 1200 6507 1270 6533
rect 1200 6473 1218 6507
rect 1252 6473 1270 6507
rect 1200 6447 1270 6473
rect 1300 6447 1370 6533
rect 1400 6507 1470 6533
rect 1400 6473 1418 6507
rect 1452 6473 1470 6507
rect 1400 6447 1470 6473
rect 1500 6507 1570 6533
rect 1500 6473 1518 6507
rect 1552 6473 1570 6507
rect 1500 6447 1570 6473
rect 1600 6507 1654 6533
rect 1600 6473 1612 6507
rect 1646 6473 1654 6507
rect 1600 6447 1654 6473
rect 216 6367 270 6393
rect 216 6333 224 6367
rect 258 6333 270 6367
rect 216 6307 270 6333
rect 300 6367 370 6393
rect 300 6333 318 6367
rect 352 6333 370 6367
rect 300 6307 370 6333
rect 400 6367 470 6393
rect 400 6333 418 6367
rect 452 6333 470 6367
rect 400 6307 470 6333
rect 500 6367 570 6393
rect 500 6333 518 6367
rect 552 6333 570 6367
rect 500 6307 570 6333
rect 600 6307 670 6393
rect 700 6367 770 6393
rect 700 6333 718 6367
rect 752 6333 770 6367
rect 700 6307 770 6333
rect 800 6367 854 6393
rect 800 6333 812 6367
rect 846 6333 854 6367
rect 800 6307 854 6333
rect 916 6367 970 6393
rect 916 6333 924 6367
rect 958 6333 970 6367
rect 916 6307 970 6333
rect 1000 6367 1054 6393
rect 1000 6333 1012 6367
rect 1046 6333 1054 6367
rect 1000 6307 1054 6333
rect 1116 6367 1170 6393
rect 1116 6333 1124 6367
rect 1158 6333 1170 6367
rect 1116 6307 1170 6333
rect 1200 6367 1270 6393
rect 1200 6333 1218 6367
rect 1252 6333 1270 6367
rect 1200 6307 1270 6333
rect 1300 6367 1370 6393
rect 1300 6333 1318 6367
rect 1352 6333 1370 6367
rect 1300 6307 1370 6333
rect 1400 6307 1470 6393
rect 1500 6367 1570 6393
rect 1500 6333 1518 6367
rect 1552 6333 1570 6367
rect 1500 6307 1570 6333
rect 1600 6367 1654 6393
rect 1600 6333 1612 6367
rect 1646 6333 1654 6367
rect 1600 6307 1654 6333
rect 3516 6647 3570 6673
rect 3516 6613 3524 6647
rect 3558 6613 3570 6647
rect 3516 6587 3570 6613
rect 3600 6647 3654 6673
rect 3600 6613 3612 6647
rect 3646 6613 3654 6647
rect 3600 6587 3654 6613
rect 3716 6647 3770 6673
rect 3716 6613 3724 6647
rect 3758 6613 3770 6647
rect 3716 6587 3770 6613
rect 3800 6647 3870 6673
rect 3800 6613 3818 6647
rect 3852 6613 3870 6647
rect 3800 6587 3870 6613
rect 3900 6647 3970 6673
rect 3900 6613 3918 6647
rect 3952 6613 3970 6647
rect 3900 6587 3970 6613
rect 4000 6587 4070 6673
rect 4100 6587 4170 6673
rect 4200 6647 4270 6673
rect 4200 6613 4218 6647
rect 4252 6613 4270 6647
rect 4200 6587 4270 6613
rect 4300 6647 4370 6673
rect 4300 6613 4318 6647
rect 4352 6613 4370 6647
rect 4300 6587 4370 6613
rect 4400 6647 4454 6673
rect 4400 6613 4412 6647
rect 4446 6613 4454 6647
rect 4400 6587 4454 6613
rect 1716 6507 1770 6533
rect 1716 6473 1724 6507
rect 1758 6473 1770 6507
rect 1716 6447 1770 6473
rect 1800 6507 1870 6533
rect 1800 6473 1818 6507
rect 1852 6473 1870 6507
rect 1800 6447 1870 6473
rect 1900 6447 1970 6533
rect 2000 6447 2070 6533
rect 2100 6507 2170 6533
rect 2100 6473 2118 6507
rect 2152 6473 2170 6507
rect 2100 6447 2170 6473
rect 2200 6507 2270 6533
rect 2200 6473 2218 6507
rect 2252 6473 2270 6507
rect 2200 6447 2270 6473
rect 2300 6447 2370 6533
rect 2400 6447 2470 6533
rect 2500 6447 2570 6533
rect 2600 6447 2670 6533
rect 2700 6447 2770 6533
rect 2800 6447 2870 6533
rect 2900 6447 2970 6533
rect 3000 6447 3070 6533
rect 3100 6447 3170 6533
rect 3200 6507 3270 6533
rect 3200 6473 3218 6507
rect 3252 6473 3270 6507
rect 3200 6447 3270 6473
rect 3300 6507 3370 6533
rect 3300 6473 3318 6507
rect 3352 6473 3370 6507
rect 3300 6447 3370 6473
rect 3400 6507 3470 6533
rect 3400 6473 3418 6507
rect 3452 6473 3470 6507
rect 3400 6447 3470 6473
rect 3500 6447 3570 6533
rect 3600 6507 3670 6533
rect 3600 6473 3618 6507
rect 3652 6473 3670 6507
rect 3600 6447 3670 6473
rect 3700 6507 3754 6533
rect 3700 6473 3712 6507
rect 3746 6473 3754 6507
rect 3700 6447 3754 6473
rect 1716 6367 1770 6393
rect 1716 6333 1724 6367
rect 1758 6333 1770 6367
rect 1716 6307 1770 6333
rect 1800 6367 1870 6393
rect 1800 6333 1818 6367
rect 1852 6333 1870 6367
rect 1800 6307 1870 6333
rect 1900 6367 1954 6393
rect 1900 6333 1912 6367
rect 1946 6333 1954 6367
rect 1900 6307 1954 6333
rect 2016 6367 2070 6393
rect 2016 6333 2024 6367
rect 2058 6333 2070 6367
rect 2016 6307 2070 6333
rect 2100 6367 2170 6393
rect 2100 6333 2118 6367
rect 2152 6333 2170 6367
rect 2100 6307 2170 6333
rect 2200 6367 2270 6393
rect 2200 6333 2218 6367
rect 2252 6333 2270 6367
rect 2200 6307 2270 6333
rect 2300 6367 2370 6393
rect 2300 6333 2318 6367
rect 2352 6333 2370 6367
rect 2300 6307 2370 6333
rect 2400 6307 2470 6393
rect 2500 6307 2570 6393
rect 2600 6367 2670 6393
rect 2600 6333 2618 6367
rect 2652 6333 2670 6367
rect 2600 6307 2670 6333
rect 2700 6367 2770 6393
rect 2700 6333 2718 6367
rect 2752 6333 2770 6367
rect 2700 6307 2770 6333
rect 2800 6367 2854 6393
rect 2800 6333 2812 6367
rect 2846 6333 2854 6367
rect 2800 6307 2854 6333
rect 16 6077 70 6163
rect 100 6077 170 6163
rect 200 6077 270 6163
rect 300 6137 370 6163
rect 300 6103 318 6137
rect 352 6103 370 6137
rect 300 6077 370 6103
rect 400 6137 470 6163
rect 400 6103 418 6137
rect 452 6103 470 6137
rect 400 6077 470 6103
rect 500 6077 570 6163
rect 600 6077 670 6163
rect 700 6077 770 6163
rect 800 6137 870 6163
rect 800 6103 818 6137
rect 852 6103 870 6137
rect 800 6077 870 6103
rect 900 6137 970 6163
rect 900 6103 918 6137
rect 952 6103 970 6137
rect 900 6077 970 6103
rect 1000 6137 1070 6163
rect 1000 6103 1018 6137
rect 1052 6103 1070 6137
rect 1000 6077 1070 6103
rect 1100 6077 1170 6163
rect 1200 6137 1270 6163
rect 1200 6103 1218 6137
rect 1252 6103 1270 6137
rect 1200 6077 1270 6103
rect 1300 6137 1370 6163
rect 1300 6103 1318 6137
rect 1352 6103 1370 6137
rect 1300 6077 1370 6103
rect 1400 6077 1470 6163
rect 1500 6137 1570 6163
rect 1500 6103 1518 6137
rect 1552 6103 1570 6137
rect 1500 6077 1570 6103
rect 1600 6137 1670 6163
rect 1600 6103 1618 6137
rect 1652 6103 1670 6137
rect 1600 6077 1670 6103
rect 1700 6077 1770 6163
rect 1800 6077 1870 6163
rect 1900 6137 1970 6163
rect 1900 6103 1918 6137
rect 1952 6103 1970 6137
rect 1900 6077 1970 6103
rect 2000 6137 2070 6163
rect 2000 6103 2018 6137
rect 2052 6103 2070 6137
rect 2000 6077 2070 6103
rect 2100 6077 2170 6163
rect 2200 6137 2270 6163
rect 2200 6103 2218 6137
rect 2252 6103 2270 6137
rect 2200 6077 2270 6103
rect 2300 6137 2370 6163
rect 2300 6103 2318 6137
rect 2352 6103 2370 6137
rect 2300 6077 2370 6103
rect 2400 6137 2454 6163
rect 2400 6103 2412 6137
rect 2446 6103 2454 6137
rect 2400 6077 2454 6103
rect 16 5937 70 6023
rect 100 5937 170 6023
rect 200 5997 270 6023
rect 200 5963 218 5997
rect 252 5963 270 5997
rect 200 5937 270 5963
rect 300 5997 370 6023
rect 300 5963 318 5997
rect 352 5963 370 5997
rect 300 5937 370 5963
rect 400 5997 454 6023
rect 400 5963 412 5997
rect 446 5963 454 5997
rect 400 5937 454 5963
rect 516 5997 570 6023
rect 516 5963 524 5997
rect 558 5963 570 5997
rect 516 5937 570 5963
rect 600 5997 670 6023
rect 600 5963 618 5997
rect 652 5963 670 5997
rect 600 5937 670 5963
rect 700 5937 770 6023
rect 800 5997 870 6023
rect 800 5963 818 5997
rect 852 5963 870 5997
rect 800 5937 870 5963
rect 900 5997 970 6023
rect 900 5963 918 5997
rect 952 5963 970 5997
rect 900 5937 970 5963
rect 1000 5997 1070 6023
rect 1000 5963 1018 5997
rect 1052 5963 1070 5997
rect 1000 5937 1070 5963
rect 1100 5937 1170 6023
rect 1200 5997 1270 6023
rect 1200 5963 1218 5997
rect 1252 5963 1270 5997
rect 1200 5937 1270 5963
rect 1300 5997 1354 6023
rect 1300 5963 1312 5997
rect 1346 5963 1354 5997
rect 1300 5937 1354 5963
rect 2916 6367 2970 6393
rect 2916 6333 2924 6367
rect 2958 6333 2970 6367
rect 2916 6307 2970 6333
rect 3000 6367 3070 6393
rect 3000 6333 3018 6367
rect 3052 6333 3070 6367
rect 3000 6307 3070 6333
rect 3100 6307 3170 6393
rect 3200 6367 3270 6393
rect 3200 6333 3218 6367
rect 3252 6333 3270 6367
rect 3200 6307 3270 6333
rect 3300 6367 3354 6393
rect 3300 6333 3312 6367
rect 3346 6333 3354 6367
rect 3300 6307 3354 6333
rect 5516 6787 5570 6813
rect 5516 6753 5524 6787
rect 5558 6753 5570 6787
rect 5516 6727 5570 6753
rect 5600 6787 5654 6813
rect 5600 6753 5612 6787
rect 5646 6753 5654 6787
rect 5600 6727 5654 6753
rect 5716 6787 5770 6813
rect 5716 6753 5724 6787
rect 5758 6753 5770 6787
rect 5716 6727 5770 6753
rect 5800 6787 5854 6813
rect 5800 6753 5812 6787
rect 5846 6753 5854 6787
rect 5800 6727 5854 6753
rect 4516 6647 4570 6673
rect 4516 6613 4524 6647
rect 4558 6613 4570 6647
rect 4516 6587 4570 6613
rect 4600 6647 4670 6673
rect 4600 6613 4618 6647
rect 4652 6613 4670 6647
rect 4600 6587 4670 6613
rect 4700 6647 4770 6673
rect 4700 6613 4718 6647
rect 4752 6613 4770 6647
rect 4700 6587 4770 6613
rect 4800 6647 4870 6673
rect 4800 6613 4818 6647
rect 4852 6613 4870 6647
rect 4800 6587 4870 6613
rect 4900 6647 4970 6673
rect 4900 6613 4918 6647
rect 4952 6613 4970 6647
rect 4900 6587 4970 6613
rect 5000 6587 5070 6673
rect 5100 6587 5170 6673
rect 5200 6587 5270 6673
rect 5300 6587 5370 6673
rect 5400 6647 5470 6673
rect 5400 6613 5418 6647
rect 5452 6613 5470 6647
rect 5400 6587 5470 6613
rect 5500 6647 5570 6673
rect 5500 6613 5518 6647
rect 5552 6613 5570 6647
rect 5500 6587 5570 6613
rect 5600 6587 5670 6673
rect 5700 6647 5770 6673
rect 5700 6613 5718 6647
rect 5752 6613 5770 6647
rect 5700 6587 5770 6613
rect 5800 6647 5854 6673
rect 5800 6613 5812 6647
rect 5846 6613 5854 6647
rect 5800 6587 5854 6613
rect 3816 6507 3870 6533
rect 3816 6473 3824 6507
rect 3858 6473 3870 6507
rect 3816 6447 3870 6473
rect 3900 6507 3970 6533
rect 3900 6473 3918 6507
rect 3952 6473 3970 6507
rect 3900 6447 3970 6473
rect 4000 6507 4070 6533
rect 4000 6473 4018 6507
rect 4052 6473 4070 6507
rect 4000 6447 4070 6473
rect 4100 6507 4170 6533
rect 4100 6473 4118 6507
rect 4152 6473 4170 6507
rect 4100 6447 4170 6473
rect 4200 6507 4270 6533
rect 4200 6473 4218 6507
rect 4252 6473 4270 6507
rect 4200 6447 4270 6473
rect 4300 6447 4370 6533
rect 4400 6447 4470 6533
rect 4500 6447 4570 6533
rect 4600 6507 4670 6533
rect 4600 6473 4618 6507
rect 4652 6473 4670 6507
rect 4600 6447 4670 6473
rect 4700 6507 4770 6533
rect 4700 6473 4718 6507
rect 4752 6473 4770 6507
rect 4700 6447 4770 6473
rect 4800 6507 4870 6533
rect 4800 6473 4818 6507
rect 4852 6473 4870 6507
rect 4800 6447 4870 6473
rect 4900 6507 4970 6533
rect 4900 6473 4918 6507
rect 4952 6473 4970 6507
rect 4900 6447 4970 6473
rect 5000 6507 5070 6533
rect 5000 6473 5018 6507
rect 5052 6473 5070 6507
rect 5000 6447 5070 6473
rect 5100 6507 5154 6533
rect 5100 6473 5112 6507
rect 5146 6473 5154 6507
rect 5100 6447 5154 6473
rect 3416 6367 3470 6393
rect 3416 6333 3424 6367
rect 3458 6333 3470 6367
rect 3416 6307 3470 6333
rect 3500 6367 3570 6393
rect 3500 6333 3518 6367
rect 3552 6333 3570 6367
rect 3500 6307 3570 6333
rect 3600 6367 3670 6393
rect 3600 6333 3618 6367
rect 3652 6333 3670 6367
rect 3600 6307 3670 6333
rect 3700 6307 3770 6393
rect 3800 6307 3870 6393
rect 3900 6367 3970 6393
rect 3900 6333 3918 6367
rect 3952 6333 3970 6367
rect 3900 6307 3970 6333
rect 4000 6367 4070 6393
rect 4000 6333 4018 6367
rect 4052 6333 4070 6367
rect 4000 6307 4070 6333
rect 4100 6367 4170 6393
rect 4100 6333 4118 6367
rect 4152 6333 4170 6367
rect 4100 6307 4170 6333
rect 4200 6307 4270 6393
rect 4300 6307 4370 6393
rect 4400 6307 4470 6393
rect 4500 6367 4570 6393
rect 4500 6333 4518 6367
rect 4552 6333 4570 6367
rect 4500 6307 4570 6333
rect 4600 6367 4670 6393
rect 4600 6333 4618 6367
rect 4652 6333 4670 6367
rect 4600 6307 4670 6333
rect 4700 6307 4770 6393
rect 4800 6367 4870 6393
rect 4800 6333 4818 6367
rect 4852 6333 4870 6367
rect 4800 6307 4870 6333
rect 4900 6367 4970 6393
rect 4900 6333 4918 6367
rect 4952 6333 4970 6367
rect 4900 6307 4970 6333
rect 5000 6367 5054 6393
rect 5000 6333 5012 6367
rect 5046 6333 5054 6367
rect 5000 6307 5054 6333
rect 2516 6137 2570 6163
rect 2516 6103 2524 6137
rect 2558 6103 2570 6137
rect 2516 6077 2570 6103
rect 2600 6137 2670 6163
rect 2600 6103 2618 6137
rect 2652 6103 2670 6137
rect 2600 6077 2670 6103
rect 2700 6137 2770 6163
rect 2700 6103 2718 6137
rect 2752 6103 2770 6137
rect 2700 6077 2770 6103
rect 2800 6077 2870 6163
rect 2900 6137 2970 6163
rect 2900 6103 2918 6137
rect 2952 6103 2970 6137
rect 2900 6077 2970 6103
rect 3000 6137 3070 6163
rect 3000 6103 3018 6137
rect 3052 6103 3070 6137
rect 3000 6077 3070 6103
rect 3100 6077 3170 6163
rect 3200 6137 3270 6163
rect 3200 6103 3218 6137
rect 3252 6103 3270 6137
rect 3200 6077 3270 6103
rect 3300 6137 3370 6163
rect 3300 6103 3318 6137
rect 3352 6103 3370 6137
rect 3300 6077 3370 6103
rect 3400 6137 3470 6163
rect 3400 6103 3418 6137
rect 3452 6103 3470 6137
rect 3400 6077 3470 6103
rect 3500 6077 3570 6163
rect 3600 6137 3670 6163
rect 3600 6103 3618 6137
rect 3652 6103 3670 6137
rect 3600 6077 3670 6103
rect 3700 6137 3754 6163
rect 3700 6103 3712 6137
rect 3746 6103 3754 6137
rect 3700 6077 3754 6103
rect 1416 5997 1470 6023
rect 1416 5963 1424 5997
rect 1458 5963 1470 5997
rect 1416 5937 1470 5963
rect 1500 5997 1570 6023
rect 1500 5963 1518 5997
rect 1552 5963 1570 5997
rect 1500 5937 1570 5963
rect 1600 5997 1670 6023
rect 1600 5963 1618 5997
rect 1652 5963 1670 5997
rect 1600 5937 1670 5963
rect 1700 5997 1770 6023
rect 1700 5963 1718 5997
rect 1752 5963 1770 5997
rect 1700 5937 1770 5963
rect 1800 5997 1870 6023
rect 1800 5963 1818 5997
rect 1852 5963 1870 5997
rect 1800 5937 1870 5963
rect 1900 5997 1970 6023
rect 1900 5963 1918 5997
rect 1952 5963 1970 5997
rect 1900 5937 1970 5963
rect 2000 5937 2070 6023
rect 2100 5937 2170 6023
rect 2200 5937 2270 6023
rect 2300 5937 2370 6023
rect 2400 5937 2470 6023
rect 2500 5937 2570 6023
rect 2600 5997 2670 6023
rect 2600 5963 2618 5997
rect 2652 5963 2670 5997
rect 2600 5937 2670 5963
rect 2700 5997 2770 6023
rect 2700 5963 2718 5997
rect 2752 5963 2770 5997
rect 2700 5937 2770 5963
rect 2800 5997 2870 6023
rect 2800 5963 2818 5997
rect 2852 5963 2870 5997
rect 2800 5937 2870 5963
rect 2900 5997 2970 6023
rect 2900 5963 2918 5997
rect 2952 5963 2970 5997
rect 2900 5937 2970 5963
rect 3000 5937 3070 6023
rect 3100 5937 3170 6023
rect 3200 5997 3270 6023
rect 3200 5963 3218 5997
rect 3252 5963 3270 5997
rect 3200 5937 3270 5963
rect 3300 5997 3354 6023
rect 3300 5963 3312 5997
rect 3346 5963 3354 5997
rect 3300 5937 3354 5963
rect 16 5857 70 5883
rect 16 5823 24 5857
rect 58 5823 70 5857
rect 16 5797 70 5823
rect 100 5857 170 5883
rect 100 5823 118 5857
rect 152 5823 170 5857
rect 100 5797 170 5823
rect 200 5857 270 5883
rect 200 5823 218 5857
rect 252 5823 270 5857
rect 200 5797 270 5823
rect 300 5797 370 5883
rect 400 5797 470 5883
rect 500 5857 570 5883
rect 500 5823 518 5857
rect 552 5823 570 5857
rect 500 5797 570 5823
rect 600 5857 670 5883
rect 600 5823 618 5857
rect 652 5823 670 5857
rect 600 5797 670 5823
rect 700 5797 770 5883
rect 800 5797 870 5883
rect 900 5857 970 5883
rect 900 5823 918 5857
rect 952 5823 970 5857
rect 900 5797 970 5823
rect 1000 5857 1070 5883
rect 1000 5823 1018 5857
rect 1052 5823 1070 5857
rect 1000 5797 1070 5823
rect 1100 5857 1170 5883
rect 1100 5823 1118 5857
rect 1152 5823 1170 5857
rect 1100 5797 1170 5823
rect 1200 5797 1270 5883
rect 1300 5857 1370 5883
rect 1300 5823 1318 5857
rect 1352 5823 1370 5857
rect 1300 5797 1370 5823
rect 1400 5857 1470 5883
rect 1400 5823 1418 5857
rect 1452 5823 1470 5857
rect 1400 5797 1470 5823
rect 1500 5857 1570 5883
rect 1500 5823 1518 5857
rect 1552 5823 1570 5857
rect 1500 5797 1570 5823
rect 1600 5857 1670 5883
rect 1600 5823 1618 5857
rect 1652 5823 1670 5857
rect 1600 5797 1670 5823
rect 1700 5857 1770 5883
rect 1700 5823 1718 5857
rect 1752 5823 1770 5857
rect 1700 5797 1770 5823
rect 1800 5797 1870 5883
rect 1900 5857 1970 5883
rect 1900 5823 1918 5857
rect 1952 5823 1970 5857
rect 1900 5797 1970 5823
rect 2000 5857 2054 5883
rect 2000 5823 2012 5857
rect 2046 5823 2054 5857
rect 2000 5797 2054 5823
rect 16 5657 70 5743
rect 100 5657 170 5743
rect 200 5717 270 5743
rect 200 5683 218 5717
rect 252 5683 270 5717
rect 200 5657 270 5683
rect 300 5717 354 5743
rect 300 5683 312 5717
rect 346 5683 354 5717
rect 300 5657 354 5683
rect 416 5717 470 5743
rect 416 5683 424 5717
rect 458 5683 470 5717
rect 416 5657 470 5683
rect 500 5717 570 5743
rect 500 5683 518 5717
rect 552 5683 570 5717
rect 500 5657 570 5683
rect 600 5717 670 5743
rect 600 5683 618 5717
rect 652 5683 670 5717
rect 600 5657 670 5683
rect 700 5717 770 5743
rect 700 5683 718 5717
rect 752 5683 770 5717
rect 700 5657 770 5683
rect 800 5717 870 5743
rect 800 5683 818 5717
rect 852 5683 870 5717
rect 800 5657 870 5683
rect 900 5717 970 5743
rect 900 5683 918 5717
rect 952 5683 970 5717
rect 900 5657 970 5683
rect 1000 5717 1054 5743
rect 1000 5683 1012 5717
rect 1046 5683 1054 5717
rect 1000 5657 1054 5683
rect 3816 6137 3870 6163
rect 3816 6103 3824 6137
rect 3858 6103 3870 6137
rect 3816 6077 3870 6103
rect 3900 6137 3970 6163
rect 3900 6103 3918 6137
rect 3952 6103 3970 6137
rect 3900 6077 3970 6103
rect 4000 6137 4054 6163
rect 4000 6103 4012 6137
rect 4046 6103 4054 6137
rect 4000 6077 4054 6103
rect 4116 6137 4170 6163
rect 4116 6103 4124 6137
rect 4158 6103 4170 6137
rect 4116 6077 4170 6103
rect 4200 6137 4270 6163
rect 4200 6103 4218 6137
rect 4252 6103 4270 6137
rect 4200 6077 4270 6103
rect 4300 6137 4370 6163
rect 4300 6103 4318 6137
rect 4352 6103 4370 6137
rect 4300 6077 4370 6103
rect 4400 6137 4454 6163
rect 4400 6103 4412 6137
rect 4446 6103 4454 6137
rect 4400 6077 4454 6103
rect 4516 6137 4570 6163
rect 4516 6103 4524 6137
rect 4558 6103 4570 6137
rect 4516 6077 4570 6103
rect 4600 6137 4654 6163
rect 4600 6103 4612 6137
rect 4646 6103 4654 6137
rect 4600 6077 4654 6103
rect 5216 6507 5270 6533
rect 5216 6473 5224 6507
rect 5258 6473 5270 6507
rect 5216 6447 5270 6473
rect 5300 6507 5354 6533
rect 5300 6473 5312 6507
rect 5346 6473 5354 6507
rect 5300 6447 5354 6473
rect 5116 6367 5170 6393
rect 5116 6333 5124 6367
rect 5158 6333 5170 6367
rect 5116 6307 5170 6333
rect 5200 6367 5270 6393
rect 5200 6333 5218 6367
rect 5252 6333 5270 6367
rect 5200 6307 5270 6333
rect 5300 6367 5354 6393
rect 5300 6333 5312 6367
rect 5346 6333 5354 6367
rect 5300 6307 5354 6333
rect 6216 7067 6270 7093
rect 6216 7033 6224 7067
rect 6258 7033 6270 7067
rect 6216 7007 6270 7033
rect 6300 7067 6370 7093
rect 6300 7033 6318 7067
rect 6352 7033 6370 7067
rect 6300 7007 6370 7033
rect 6400 7007 6454 7093
rect 6512 7082 6570 7093
rect 6512 7048 6524 7082
rect 6558 7048 6570 7082
rect 6512 7007 6570 7048
rect 6600 7067 6670 7093
rect 6600 7033 6618 7067
rect 6652 7033 6670 7067
rect 6600 7007 6670 7033
rect 6700 7052 6758 7093
rect 6700 7018 6712 7052
rect 6746 7018 6758 7052
rect 6700 7007 6758 7018
rect 6820 7067 6880 7093
rect 6820 7033 6828 7067
rect 6862 7033 6880 7067
rect 6820 7007 6880 7033
rect 6910 7067 6980 7093
rect 6910 7033 6928 7067
rect 6962 7033 6980 7067
rect 6910 7007 6980 7033
rect 7010 7067 7080 7093
rect 7010 7033 7028 7067
rect 7062 7033 7080 7067
rect 7010 7007 7080 7033
rect 7110 7067 7180 7093
rect 7110 7033 7128 7067
rect 7162 7033 7180 7067
rect 7110 7007 7180 7033
rect 7210 7067 7280 7093
rect 7210 7033 7228 7067
rect 7262 7033 7280 7067
rect 7210 7007 7280 7033
rect 7310 7067 7380 7093
rect 7310 7033 7328 7067
rect 7362 7033 7380 7067
rect 7310 7007 7380 7033
rect 7410 7067 7470 7093
rect 7410 7033 7428 7067
rect 7462 7033 7470 7067
rect 7410 7007 7470 7033
rect 6216 6927 6270 6953
rect 6216 6893 6224 6927
rect 6258 6893 6270 6927
rect 6216 6867 6270 6893
rect 6300 6927 6370 6953
rect 6300 6893 6318 6927
rect 6352 6893 6370 6927
rect 6300 6867 6370 6893
rect 6400 6867 6454 6953
rect 6512 6942 6570 6953
rect 6512 6908 6524 6942
rect 6558 6908 6570 6942
rect 6512 6867 6570 6908
rect 6600 6927 6670 6953
rect 6600 6893 6618 6927
rect 6652 6893 6670 6927
rect 6600 6867 6670 6893
rect 6700 6912 6758 6953
rect 6700 6878 6712 6912
rect 6746 6878 6758 6912
rect 6700 6867 6758 6878
rect 6820 6927 6880 6953
rect 6820 6893 6828 6927
rect 6862 6893 6880 6927
rect 6820 6867 6880 6893
rect 6910 6927 6980 6953
rect 6910 6893 6928 6927
rect 6962 6893 6980 6927
rect 6910 6867 6980 6893
rect 7010 6927 7080 6953
rect 7010 6893 7028 6927
rect 7062 6893 7080 6927
rect 7010 6867 7080 6893
rect 7110 6927 7180 6953
rect 7110 6893 7128 6927
rect 7162 6893 7180 6927
rect 7110 6867 7180 6893
rect 7210 6927 7280 6953
rect 7210 6893 7228 6927
rect 7262 6893 7280 6927
rect 7210 6867 7280 6893
rect 7310 6927 7380 6953
rect 7310 6893 7328 6927
rect 7362 6893 7380 6927
rect 7310 6867 7380 6893
rect 7410 6927 7470 6953
rect 7410 6893 7428 6927
rect 7462 6893 7470 6927
rect 7410 6867 7470 6893
rect 5916 6787 5970 6813
rect 5916 6753 5924 6787
rect 5958 6753 5970 6787
rect 5916 6727 5970 6753
rect 6000 6787 6070 6813
rect 6000 6753 6018 6787
rect 6052 6753 6070 6787
rect 6000 6727 6070 6753
rect 6100 6787 6170 6813
rect 6100 6753 6118 6787
rect 6152 6753 6170 6787
rect 6100 6727 6170 6753
rect 6200 6787 6270 6813
rect 6200 6753 6218 6787
rect 6252 6753 6270 6787
rect 6200 6727 6270 6753
rect 6300 6787 6370 6813
rect 6300 6753 6318 6787
rect 6352 6753 6370 6787
rect 6300 6727 6370 6753
rect 6400 6727 6454 6813
rect 6512 6802 6570 6813
rect 6512 6768 6524 6802
rect 6558 6768 6570 6802
rect 6512 6727 6570 6768
rect 6600 6787 6670 6813
rect 6600 6753 6618 6787
rect 6652 6753 6670 6787
rect 6600 6727 6670 6753
rect 6700 6772 6758 6813
rect 6700 6738 6712 6772
rect 6746 6738 6758 6772
rect 6700 6727 6758 6738
rect 6820 6787 6880 6813
rect 6820 6753 6828 6787
rect 6862 6753 6880 6787
rect 6820 6727 6880 6753
rect 6910 6787 6980 6813
rect 6910 6753 6928 6787
rect 6962 6753 6980 6787
rect 6910 6727 6980 6753
rect 7010 6787 7080 6813
rect 7010 6753 7028 6787
rect 7062 6753 7080 6787
rect 7010 6727 7080 6753
rect 7110 6787 7180 6813
rect 7110 6753 7128 6787
rect 7162 6753 7180 6787
rect 7110 6727 7180 6753
rect 7210 6787 7280 6813
rect 7210 6753 7228 6787
rect 7262 6753 7280 6787
rect 7210 6727 7280 6753
rect 7310 6787 7380 6813
rect 7310 6753 7328 6787
rect 7362 6753 7380 6787
rect 7310 6727 7380 6753
rect 7410 6787 7470 6813
rect 7410 6753 7428 6787
rect 7462 6753 7470 6787
rect 7410 6727 7470 6753
rect 5916 6647 5970 6673
rect 5916 6613 5924 6647
rect 5958 6613 5970 6647
rect 5916 6587 5970 6613
rect 6000 6647 6070 6673
rect 6000 6613 6018 6647
rect 6052 6613 6070 6647
rect 6000 6587 6070 6613
rect 6100 6647 6170 6673
rect 6100 6613 6118 6647
rect 6152 6613 6170 6647
rect 6100 6587 6170 6613
rect 6200 6587 6270 6673
rect 6300 6587 6370 6673
rect 6400 6587 6454 6673
rect 6512 6662 6570 6673
rect 6512 6628 6524 6662
rect 6558 6628 6570 6662
rect 6512 6587 6570 6628
rect 6600 6647 6670 6673
rect 6600 6613 6618 6647
rect 6652 6613 6670 6647
rect 6600 6587 6670 6613
rect 6700 6632 6758 6673
rect 6700 6598 6712 6632
rect 6746 6598 6758 6632
rect 6700 6587 6758 6598
rect 6820 6647 6880 6673
rect 6820 6613 6828 6647
rect 6862 6613 6880 6647
rect 6820 6587 6880 6613
rect 6910 6647 6980 6673
rect 6910 6613 6928 6647
rect 6962 6613 6980 6647
rect 6910 6587 6980 6613
rect 7010 6647 7080 6673
rect 7010 6613 7028 6647
rect 7062 6613 7080 6647
rect 7010 6587 7080 6613
rect 7110 6647 7180 6673
rect 7110 6613 7128 6647
rect 7162 6613 7180 6647
rect 7110 6587 7180 6613
rect 7210 6647 7280 6673
rect 7210 6613 7228 6647
rect 7262 6613 7280 6647
rect 7210 6587 7280 6613
rect 7310 6647 7380 6673
rect 7310 6613 7328 6647
rect 7362 6613 7380 6647
rect 7310 6587 7380 6613
rect 7410 6647 7470 6673
rect 7410 6613 7428 6647
rect 7462 6613 7470 6647
rect 7410 6587 7470 6613
rect 5416 6507 5470 6533
rect 5416 6473 5424 6507
rect 5458 6473 5470 6507
rect 5416 6447 5470 6473
rect 5500 6507 5570 6533
rect 5500 6473 5518 6507
rect 5552 6473 5570 6507
rect 5500 6447 5570 6473
rect 5600 6507 5670 6533
rect 5600 6473 5618 6507
rect 5652 6473 5670 6507
rect 5600 6447 5670 6473
rect 5700 6507 5770 6533
rect 5700 6473 5718 6507
rect 5752 6473 5770 6507
rect 5700 6447 5770 6473
rect 5800 6507 5870 6533
rect 5800 6473 5818 6507
rect 5852 6473 5870 6507
rect 5800 6447 5870 6473
rect 5900 6507 5970 6533
rect 5900 6473 5918 6507
rect 5952 6473 5970 6507
rect 5900 6447 5970 6473
rect 6000 6507 6070 6533
rect 6000 6473 6018 6507
rect 6052 6473 6070 6507
rect 6000 6447 6070 6473
rect 6100 6447 6170 6533
rect 6200 6507 6270 6533
rect 6200 6473 6218 6507
rect 6252 6473 6270 6507
rect 6200 6447 6270 6473
rect 6300 6507 6370 6533
rect 6300 6473 6318 6507
rect 6352 6473 6370 6507
rect 6300 6447 6370 6473
rect 6400 6447 6454 6533
rect 6512 6522 6570 6533
rect 6512 6488 6524 6522
rect 6558 6488 6570 6522
rect 6512 6447 6570 6488
rect 6600 6507 6670 6533
rect 6600 6473 6618 6507
rect 6652 6473 6670 6507
rect 6600 6447 6670 6473
rect 6700 6492 6758 6533
rect 6700 6458 6712 6492
rect 6746 6458 6758 6492
rect 6700 6447 6758 6458
rect 6820 6507 6880 6533
rect 6820 6473 6828 6507
rect 6862 6473 6880 6507
rect 6820 6447 6880 6473
rect 6910 6507 6980 6533
rect 6910 6473 6928 6507
rect 6962 6473 6980 6507
rect 6910 6447 6980 6473
rect 7010 6507 7080 6533
rect 7010 6473 7028 6507
rect 7062 6473 7080 6507
rect 7010 6447 7080 6473
rect 7110 6507 7180 6533
rect 7110 6473 7128 6507
rect 7162 6473 7180 6507
rect 7110 6447 7180 6473
rect 7210 6507 7280 6533
rect 7210 6473 7228 6507
rect 7262 6473 7280 6507
rect 7210 6447 7280 6473
rect 7310 6507 7380 6533
rect 7310 6473 7328 6507
rect 7362 6473 7380 6507
rect 7310 6447 7380 6473
rect 7410 6507 7470 6533
rect 7410 6473 7428 6507
rect 7462 6473 7470 6507
rect 7410 6447 7470 6473
rect 5416 6367 5470 6393
rect 5416 6333 5424 6367
rect 5458 6333 5470 6367
rect 5416 6307 5470 6333
rect 5500 6367 5570 6393
rect 5500 6333 5518 6367
rect 5552 6333 5570 6367
rect 5500 6307 5570 6333
rect 5600 6307 5670 6393
rect 5700 6307 5770 6393
rect 5800 6367 5870 6393
rect 5800 6333 5818 6367
rect 5852 6333 5870 6367
rect 5800 6307 5870 6333
rect 5900 6367 5970 6393
rect 5900 6333 5918 6367
rect 5952 6333 5970 6367
rect 5900 6307 5970 6333
rect 6000 6367 6070 6393
rect 6000 6333 6018 6367
rect 6052 6333 6070 6367
rect 6000 6307 6070 6333
rect 6100 6367 6154 6393
rect 6100 6333 6112 6367
rect 6146 6333 6154 6367
rect 6100 6307 6154 6333
rect 6216 6367 6270 6393
rect 6216 6333 6224 6367
rect 6258 6333 6270 6367
rect 6216 6307 6270 6333
rect 6300 6367 6370 6393
rect 6300 6333 6318 6367
rect 6352 6333 6370 6367
rect 6300 6307 6370 6333
rect 6400 6367 6454 6393
rect 6400 6333 6412 6367
rect 6446 6333 6454 6367
rect 6400 6307 6454 6333
rect 6512 6382 6570 6393
rect 6512 6348 6524 6382
rect 6558 6348 6570 6382
rect 6512 6307 6570 6348
rect 6600 6367 6670 6393
rect 6600 6333 6618 6367
rect 6652 6333 6670 6367
rect 6600 6307 6670 6333
rect 6700 6352 6758 6393
rect 6700 6318 6712 6352
rect 6746 6318 6758 6352
rect 6700 6307 6758 6318
rect 6820 6367 6880 6393
rect 6820 6333 6828 6367
rect 6862 6333 6880 6367
rect 6820 6307 6880 6333
rect 6910 6367 6980 6393
rect 6910 6333 6928 6367
rect 6962 6333 6980 6367
rect 6910 6307 6980 6333
rect 7010 6367 7080 6393
rect 7010 6333 7028 6367
rect 7062 6333 7080 6367
rect 7010 6307 7080 6333
rect 7110 6367 7180 6393
rect 7110 6333 7128 6367
rect 7162 6333 7180 6367
rect 7110 6307 7180 6333
rect 7210 6367 7280 6393
rect 7210 6333 7228 6367
rect 7262 6333 7280 6367
rect 7210 6307 7280 6333
rect 7310 6367 7380 6393
rect 7310 6333 7328 6367
rect 7362 6333 7380 6367
rect 7310 6307 7380 6333
rect 7410 6367 7470 6393
rect 7410 6333 7428 6367
rect 7462 6333 7470 6367
rect 7410 6307 7470 6333
rect 4716 6137 4770 6163
rect 4716 6103 4724 6137
rect 4758 6103 4770 6137
rect 4716 6077 4770 6103
rect 4800 6137 4870 6163
rect 4800 6103 4818 6137
rect 4852 6103 4870 6137
rect 4800 6077 4870 6103
rect 4900 6137 4970 6163
rect 4900 6103 4918 6137
rect 4952 6103 4970 6137
rect 4900 6077 4970 6103
rect 5000 6077 5070 6163
rect 5100 6077 5170 6163
rect 5200 6077 5270 6163
rect 5300 6077 5370 6163
rect 5400 6137 5470 6163
rect 5400 6103 5418 6137
rect 5452 6103 5470 6137
rect 5400 6077 5470 6103
rect 5500 6137 5570 6163
rect 5500 6103 5518 6137
rect 5552 6103 5570 6137
rect 5500 6077 5570 6103
rect 5600 6077 5670 6163
rect 5700 6137 5770 6163
rect 5700 6103 5718 6137
rect 5752 6103 5770 6137
rect 5700 6077 5770 6103
rect 5800 6137 5870 6163
rect 5800 6103 5818 6137
rect 5852 6103 5870 6137
rect 5800 6077 5870 6103
rect 5900 6137 5970 6163
rect 5900 6103 5918 6137
rect 5952 6103 5970 6137
rect 5900 6077 5970 6103
rect 6000 6137 6054 6163
rect 6000 6103 6012 6137
rect 6046 6103 6054 6137
rect 6000 6077 6054 6103
rect 3416 5997 3470 6023
rect 3416 5963 3424 5997
rect 3458 5963 3470 5997
rect 3416 5937 3470 5963
rect 3500 5997 3570 6023
rect 3500 5963 3518 5997
rect 3552 5963 3570 5997
rect 3500 5937 3570 5963
rect 3600 5997 3670 6023
rect 3600 5963 3618 5997
rect 3652 5963 3670 5997
rect 3600 5937 3670 5963
rect 3700 5997 3770 6023
rect 3700 5963 3718 5997
rect 3752 5963 3770 5997
rect 3700 5937 3770 5963
rect 3800 5997 3870 6023
rect 3800 5963 3818 5997
rect 3852 5963 3870 5997
rect 3800 5937 3870 5963
rect 3900 5997 3970 6023
rect 3900 5963 3918 5997
rect 3952 5963 3970 5997
rect 3900 5937 3970 5963
rect 4000 5937 4070 6023
rect 4100 5937 4170 6023
rect 4200 5997 4270 6023
rect 4200 5963 4218 5997
rect 4252 5963 4270 5997
rect 4200 5937 4270 5963
rect 4300 5997 4370 6023
rect 4300 5963 4318 5997
rect 4352 5963 4370 5997
rect 4300 5937 4370 5963
rect 4400 5937 4470 6023
rect 4500 5997 4570 6023
rect 4500 5963 4518 5997
rect 4552 5963 4570 5997
rect 4500 5937 4570 5963
rect 4600 5997 4670 6023
rect 4600 5963 4618 5997
rect 4652 5963 4670 5997
rect 4600 5937 4670 5963
rect 4700 5937 4770 6023
rect 4800 5937 4870 6023
rect 4900 5997 4970 6023
rect 4900 5963 4918 5997
rect 4952 5963 4970 5997
rect 4900 5937 4970 5963
rect 5000 5997 5070 6023
rect 5000 5963 5018 5997
rect 5052 5963 5070 5997
rect 5000 5937 5070 5963
rect 5100 5997 5170 6023
rect 5100 5963 5118 5997
rect 5152 5963 5170 5997
rect 5100 5937 5170 5963
rect 5200 5997 5254 6023
rect 5200 5963 5212 5997
rect 5246 5963 5254 5997
rect 5200 5937 5254 5963
rect 2116 5857 2170 5883
rect 2116 5823 2124 5857
rect 2158 5823 2170 5857
rect 2116 5797 2170 5823
rect 2200 5857 2270 5883
rect 2200 5823 2218 5857
rect 2252 5823 2270 5857
rect 2200 5797 2270 5823
rect 2300 5857 2370 5883
rect 2300 5823 2318 5857
rect 2352 5823 2370 5857
rect 2300 5797 2370 5823
rect 2400 5797 2470 5883
rect 2500 5857 2570 5883
rect 2500 5823 2518 5857
rect 2552 5823 2570 5857
rect 2500 5797 2570 5823
rect 2600 5857 2670 5883
rect 2600 5823 2618 5857
rect 2652 5823 2670 5857
rect 2600 5797 2670 5823
rect 2700 5857 2770 5883
rect 2700 5823 2718 5857
rect 2752 5823 2770 5857
rect 2700 5797 2770 5823
rect 2800 5857 2870 5883
rect 2800 5823 2818 5857
rect 2852 5823 2870 5857
rect 2800 5797 2870 5823
rect 2900 5857 2970 5883
rect 2900 5823 2918 5857
rect 2952 5823 2970 5857
rect 2900 5797 2970 5823
rect 3000 5797 3070 5883
rect 3100 5857 3170 5883
rect 3100 5823 3118 5857
rect 3152 5823 3170 5857
rect 3100 5797 3170 5823
rect 3200 5857 3270 5883
rect 3200 5823 3218 5857
rect 3252 5823 3270 5857
rect 3200 5797 3270 5823
rect 3300 5857 3370 5883
rect 3300 5823 3318 5857
rect 3352 5823 3370 5857
rect 3300 5797 3370 5823
rect 3400 5857 3454 5883
rect 3400 5823 3412 5857
rect 3446 5823 3454 5857
rect 3400 5797 3454 5823
rect 1116 5717 1170 5743
rect 1116 5683 1124 5717
rect 1158 5683 1170 5717
rect 1116 5657 1170 5683
rect 1200 5717 1270 5743
rect 1200 5683 1218 5717
rect 1252 5683 1270 5717
rect 1200 5657 1270 5683
rect 1300 5717 1370 5743
rect 1300 5683 1318 5717
rect 1352 5683 1370 5717
rect 1300 5657 1370 5683
rect 1400 5717 1470 5743
rect 1400 5683 1418 5717
rect 1452 5683 1470 5717
rect 1400 5657 1470 5683
rect 1500 5717 1570 5743
rect 1500 5683 1518 5717
rect 1552 5683 1570 5717
rect 1500 5657 1570 5683
rect 1600 5717 1670 5743
rect 1600 5683 1618 5717
rect 1652 5683 1670 5717
rect 1600 5657 1670 5683
rect 1700 5717 1770 5743
rect 1700 5683 1718 5717
rect 1752 5683 1770 5717
rect 1700 5657 1770 5683
rect 1800 5717 1870 5743
rect 1800 5683 1818 5717
rect 1852 5683 1870 5717
rect 1800 5657 1870 5683
rect 1900 5717 1970 5743
rect 1900 5683 1918 5717
rect 1952 5683 1970 5717
rect 1900 5657 1970 5683
rect 2000 5657 2070 5743
rect 2100 5717 2170 5743
rect 2100 5683 2118 5717
rect 2152 5683 2170 5717
rect 2100 5657 2170 5683
rect 2200 5717 2270 5743
rect 2200 5683 2218 5717
rect 2252 5683 2270 5717
rect 2200 5657 2270 5683
rect 2300 5717 2370 5743
rect 2300 5683 2318 5717
rect 2352 5683 2370 5717
rect 2300 5657 2370 5683
rect 2400 5657 2470 5743
rect 2500 5657 2570 5743
rect 2600 5657 2670 5743
rect 2700 5717 2770 5743
rect 2700 5683 2718 5717
rect 2752 5683 2770 5717
rect 2700 5657 2770 5683
rect 2800 5717 2854 5743
rect 2800 5683 2812 5717
rect 2846 5683 2854 5717
rect 2800 5657 2854 5683
rect 16 5517 70 5603
rect 100 5577 170 5603
rect 100 5543 118 5577
rect 152 5543 170 5577
rect 100 5517 170 5543
rect 200 5577 270 5603
rect 200 5543 218 5577
rect 252 5543 270 5577
rect 200 5517 270 5543
rect 300 5577 370 5603
rect 300 5543 318 5577
rect 352 5543 370 5577
rect 300 5517 370 5543
rect 400 5577 470 5603
rect 400 5543 418 5577
rect 452 5543 470 5577
rect 400 5517 470 5543
rect 500 5577 570 5603
rect 500 5543 518 5577
rect 552 5543 570 5577
rect 500 5517 570 5543
rect 600 5517 670 5603
rect 700 5577 770 5603
rect 700 5543 718 5577
rect 752 5543 770 5577
rect 700 5517 770 5543
rect 800 5577 870 5603
rect 800 5543 818 5577
rect 852 5543 870 5577
rect 800 5517 870 5543
rect 900 5517 970 5603
rect 1000 5577 1070 5603
rect 1000 5543 1018 5577
rect 1052 5543 1070 5577
rect 1000 5517 1070 5543
rect 1100 5577 1154 5603
rect 1100 5543 1112 5577
rect 1146 5543 1154 5577
rect 1100 5517 1154 5543
rect 16 5437 70 5463
rect 16 5403 24 5437
rect 58 5403 70 5437
rect 16 5377 70 5403
rect 100 5437 170 5463
rect 100 5403 118 5437
rect 152 5403 170 5437
rect 100 5377 170 5403
rect 200 5437 270 5463
rect 200 5403 218 5437
rect 252 5403 270 5437
rect 200 5377 270 5403
rect 300 5437 370 5463
rect 300 5403 318 5437
rect 352 5403 370 5437
rect 300 5377 370 5403
rect 400 5437 454 5463
rect 400 5403 412 5437
rect 446 5403 454 5437
rect 400 5377 454 5403
rect 1216 5577 1270 5603
rect 1216 5543 1224 5577
rect 1258 5543 1270 5577
rect 1216 5517 1270 5543
rect 1300 5577 1354 5603
rect 1300 5543 1312 5577
rect 1346 5543 1354 5577
rect 1300 5517 1354 5543
rect 1416 5577 1470 5603
rect 1416 5543 1424 5577
rect 1458 5543 1470 5577
rect 1416 5517 1470 5543
rect 1500 5577 1570 5603
rect 1500 5543 1518 5577
rect 1552 5543 1570 5577
rect 1500 5517 1570 5543
rect 1600 5577 1670 5603
rect 1600 5543 1618 5577
rect 1652 5543 1670 5577
rect 1600 5517 1670 5543
rect 1700 5577 1770 5603
rect 1700 5543 1718 5577
rect 1752 5543 1770 5577
rect 1700 5517 1770 5543
rect 1800 5577 1870 5603
rect 1800 5543 1818 5577
rect 1852 5543 1870 5577
rect 1800 5517 1870 5543
rect 1900 5577 1954 5603
rect 1900 5543 1912 5577
rect 1946 5543 1954 5577
rect 1900 5517 1954 5543
rect 516 5437 570 5463
rect 516 5403 524 5437
rect 558 5403 570 5437
rect 516 5377 570 5403
rect 600 5437 670 5463
rect 600 5403 618 5437
rect 652 5403 670 5437
rect 600 5377 670 5403
rect 700 5437 770 5463
rect 700 5403 718 5437
rect 752 5403 770 5437
rect 700 5377 770 5403
rect 800 5377 870 5463
rect 900 5377 970 5463
rect 1000 5377 1070 5463
rect 1100 5377 1170 5463
rect 1200 5377 1270 5463
rect 1300 5437 1370 5463
rect 1300 5403 1318 5437
rect 1352 5403 1370 5437
rect 1300 5377 1370 5403
rect 1400 5437 1454 5463
rect 1400 5403 1412 5437
rect 1446 5403 1454 5437
rect 1400 5377 1454 5403
rect 1516 5437 1570 5463
rect 1516 5403 1524 5437
rect 1558 5403 1570 5437
rect 1516 5377 1570 5403
rect 1600 5437 1670 5463
rect 1600 5403 1618 5437
rect 1652 5403 1670 5437
rect 1600 5377 1670 5403
rect 1700 5437 1754 5463
rect 1700 5403 1712 5437
rect 1746 5403 1754 5437
rect 1700 5377 1754 5403
rect 2016 5577 2070 5603
rect 2016 5543 2024 5577
rect 2058 5543 2070 5577
rect 2016 5517 2070 5543
rect 2100 5577 2170 5603
rect 2100 5543 2118 5577
rect 2152 5543 2170 5577
rect 2100 5517 2170 5543
rect 2200 5577 2254 5603
rect 2200 5543 2212 5577
rect 2246 5543 2254 5577
rect 2200 5517 2254 5543
rect 1816 5437 1870 5463
rect 1816 5403 1824 5437
rect 1858 5403 1870 5437
rect 1816 5377 1870 5403
rect 1900 5437 1970 5463
rect 1900 5403 1918 5437
rect 1952 5403 1970 5437
rect 1900 5377 1970 5403
rect 2000 5437 2070 5463
rect 2000 5403 2018 5437
rect 2052 5403 2070 5437
rect 2000 5377 2070 5403
rect 2100 5437 2170 5463
rect 2100 5403 2118 5437
rect 2152 5403 2170 5437
rect 2100 5377 2170 5403
rect 2200 5437 2254 5463
rect 2200 5403 2212 5437
rect 2246 5403 2254 5437
rect 2200 5377 2254 5403
rect 16 5237 70 5323
rect 100 5237 170 5323
rect 200 5237 270 5323
rect 300 5297 370 5323
rect 300 5263 318 5297
rect 352 5263 370 5297
rect 300 5237 370 5263
rect 400 5297 470 5323
rect 400 5263 418 5297
rect 452 5263 470 5297
rect 400 5237 470 5263
rect 500 5237 570 5323
rect 600 5237 670 5323
rect 700 5297 770 5323
rect 700 5263 718 5297
rect 752 5263 770 5297
rect 700 5237 770 5263
rect 800 5297 870 5323
rect 800 5263 818 5297
rect 852 5263 870 5297
rect 800 5237 870 5263
rect 900 5237 970 5323
rect 1000 5237 1070 5323
rect 1100 5237 1170 5323
rect 1200 5297 1270 5323
rect 1200 5263 1218 5297
rect 1252 5263 1270 5297
rect 1200 5237 1270 5263
rect 1300 5297 1370 5323
rect 1300 5263 1318 5297
rect 1352 5263 1370 5297
rect 1300 5237 1370 5263
rect 1400 5297 1470 5323
rect 1400 5263 1418 5297
rect 1452 5263 1470 5297
rect 1400 5237 1470 5263
rect 1500 5237 1570 5323
rect 1600 5297 1670 5323
rect 1600 5263 1618 5297
rect 1652 5263 1670 5297
rect 1600 5237 1670 5263
rect 1700 5297 1770 5323
rect 1700 5263 1718 5297
rect 1752 5263 1770 5297
rect 1700 5237 1770 5263
rect 1800 5237 1870 5323
rect 1900 5237 1970 5323
rect 2000 5297 2070 5323
rect 2000 5263 2018 5297
rect 2052 5263 2070 5297
rect 2000 5237 2070 5263
rect 2100 5297 2154 5323
rect 2100 5263 2112 5297
rect 2146 5263 2154 5297
rect 2100 5237 2154 5263
rect 16 5097 70 5183
rect 100 5157 170 5183
rect 100 5123 118 5157
rect 152 5123 170 5157
rect 100 5097 170 5123
rect 200 5157 270 5183
rect 200 5123 218 5157
rect 252 5123 270 5157
rect 200 5097 270 5123
rect 300 5157 370 5183
rect 300 5123 318 5157
rect 352 5123 370 5157
rect 300 5097 370 5123
rect 400 5157 470 5183
rect 400 5123 418 5157
rect 452 5123 470 5157
rect 400 5097 470 5123
rect 500 5097 570 5183
rect 600 5157 670 5183
rect 600 5123 618 5157
rect 652 5123 670 5157
rect 600 5097 670 5123
rect 700 5157 770 5183
rect 700 5123 718 5157
rect 752 5123 770 5157
rect 700 5097 770 5123
rect 800 5157 870 5183
rect 800 5123 818 5157
rect 852 5123 870 5157
rect 800 5097 870 5123
rect 900 5097 970 5183
rect 1000 5097 1070 5183
rect 1100 5097 1170 5183
rect 1200 5157 1270 5183
rect 1200 5123 1218 5157
rect 1252 5123 1270 5157
rect 1200 5097 1270 5123
rect 1300 5157 1354 5183
rect 1300 5123 1312 5157
rect 1346 5123 1354 5157
rect 1300 5097 1354 5123
rect 16 4787 70 4813
rect 16 4753 24 4787
rect 58 4753 70 4787
rect 16 4727 70 4753
rect 100 4787 170 4813
rect 100 4753 118 4787
rect 152 4753 170 4787
rect 100 4727 170 4753
rect 200 4787 254 4813
rect 200 4753 212 4787
rect 246 4753 254 4787
rect 200 4727 254 4753
rect 316 4787 370 4813
rect 316 4753 324 4787
rect 358 4753 370 4787
rect 316 4727 370 4753
rect 400 4787 470 4813
rect 400 4753 418 4787
rect 452 4753 470 4787
rect 400 4727 470 4753
rect 500 4727 570 4813
rect 600 4787 670 4813
rect 600 4753 618 4787
rect 652 4753 670 4787
rect 600 4727 670 4753
rect 700 4787 770 4813
rect 700 4753 718 4787
rect 752 4753 770 4787
rect 700 4727 770 4753
rect 800 4727 870 4813
rect 900 4727 970 4813
rect 1000 4787 1070 4813
rect 1000 4753 1018 4787
rect 1052 4753 1070 4787
rect 1000 4727 1070 4753
rect 1100 4787 1154 4813
rect 1100 4753 1112 4787
rect 1146 4753 1154 4787
rect 1100 4727 1154 4753
rect 1416 5157 1470 5183
rect 1416 5123 1424 5157
rect 1458 5123 1470 5157
rect 1416 5097 1470 5123
rect 1500 5157 1570 5183
rect 1500 5123 1518 5157
rect 1552 5123 1570 5157
rect 1500 5097 1570 5123
rect 1600 5157 1670 5183
rect 1600 5123 1618 5157
rect 1652 5123 1670 5157
rect 1600 5097 1670 5123
rect 1700 5157 1770 5183
rect 1700 5123 1718 5157
rect 1752 5123 1770 5157
rect 1700 5097 1770 5123
rect 1800 5097 1870 5183
rect 1900 5097 1970 5183
rect 2000 5157 2070 5183
rect 2000 5123 2018 5157
rect 2052 5123 2070 5157
rect 2000 5097 2070 5123
rect 2100 5157 2154 5183
rect 2100 5123 2112 5157
rect 2146 5123 2154 5157
rect 2100 5097 2154 5123
rect 2916 5717 2970 5743
rect 2916 5683 2924 5717
rect 2958 5683 2970 5717
rect 2916 5657 2970 5683
rect 3000 5717 3054 5743
rect 3000 5683 3012 5717
rect 3046 5683 3054 5717
rect 3000 5657 3054 5683
rect 3116 5717 3170 5743
rect 3116 5683 3124 5717
rect 3158 5683 3170 5717
rect 3116 5657 3170 5683
rect 3200 5717 3254 5743
rect 3200 5683 3212 5717
rect 3246 5683 3254 5717
rect 3200 5657 3254 5683
rect 3316 5717 3370 5743
rect 3316 5683 3324 5717
rect 3358 5683 3370 5717
rect 3316 5657 3370 5683
rect 3400 5717 3454 5743
rect 3400 5683 3412 5717
rect 3446 5683 3454 5717
rect 3400 5657 3454 5683
rect 3516 5857 3570 5883
rect 3516 5823 3524 5857
rect 3558 5823 3570 5857
rect 3516 5797 3570 5823
rect 3600 5857 3670 5883
rect 3600 5823 3618 5857
rect 3652 5823 3670 5857
rect 3600 5797 3670 5823
rect 3700 5857 3770 5883
rect 3700 5823 3718 5857
rect 3752 5823 3770 5857
rect 3700 5797 3770 5823
rect 3800 5797 3870 5883
rect 3900 5797 3970 5883
rect 4000 5857 4070 5883
rect 4000 5823 4018 5857
rect 4052 5823 4070 5857
rect 4000 5797 4070 5823
rect 4100 5857 4154 5883
rect 4100 5823 4112 5857
rect 4146 5823 4154 5857
rect 4100 5797 4154 5823
rect 3516 5717 3570 5743
rect 3516 5683 3524 5717
rect 3558 5683 3570 5717
rect 3516 5657 3570 5683
rect 3600 5717 3654 5743
rect 3600 5683 3612 5717
rect 3646 5683 3654 5717
rect 3600 5657 3654 5683
rect 3716 5717 3770 5743
rect 3716 5683 3724 5717
rect 3758 5683 3770 5717
rect 3716 5657 3770 5683
rect 3800 5717 3870 5743
rect 3800 5683 3818 5717
rect 3852 5683 3870 5717
rect 3800 5657 3870 5683
rect 3900 5657 3970 5743
rect 4000 5717 4070 5743
rect 4000 5683 4018 5717
rect 4052 5683 4070 5717
rect 4000 5657 4070 5683
rect 4100 5717 4154 5743
rect 4100 5683 4112 5717
rect 4146 5683 4154 5717
rect 4100 5657 4154 5683
rect 2316 5577 2370 5603
rect 2316 5543 2324 5577
rect 2358 5543 2370 5577
rect 2316 5517 2370 5543
rect 2400 5577 2470 5603
rect 2400 5543 2418 5577
rect 2452 5543 2470 5577
rect 2400 5517 2470 5543
rect 2500 5577 2570 5603
rect 2500 5543 2518 5577
rect 2552 5543 2570 5577
rect 2500 5517 2570 5543
rect 2600 5517 2670 5603
rect 2700 5517 2770 5603
rect 2800 5517 2870 5603
rect 2900 5517 2970 5603
rect 3000 5577 3070 5603
rect 3000 5543 3018 5577
rect 3052 5543 3070 5577
rect 3000 5517 3070 5543
rect 3100 5577 3170 5603
rect 3100 5543 3118 5577
rect 3152 5543 3170 5577
rect 3100 5517 3170 5543
rect 3200 5577 3270 5603
rect 3200 5543 3218 5577
rect 3252 5543 3270 5577
rect 3200 5517 3270 5543
rect 3300 5577 3370 5603
rect 3300 5543 3318 5577
rect 3352 5543 3370 5577
rect 3300 5517 3370 5543
rect 3400 5577 3470 5603
rect 3400 5543 3418 5577
rect 3452 5543 3470 5577
rect 3400 5517 3470 5543
rect 3500 5577 3570 5603
rect 3500 5543 3518 5577
rect 3552 5543 3570 5577
rect 3500 5517 3570 5543
rect 3600 5577 3670 5603
rect 3600 5543 3618 5577
rect 3652 5543 3670 5577
rect 3600 5517 3670 5543
rect 3700 5517 3770 5603
rect 3800 5577 3870 5603
rect 3800 5543 3818 5577
rect 3852 5543 3870 5577
rect 3800 5517 3870 5543
rect 3900 5577 3970 5603
rect 3900 5543 3918 5577
rect 3952 5543 3970 5577
rect 3900 5517 3970 5543
rect 4000 5577 4054 5603
rect 4000 5543 4012 5577
rect 4046 5543 4054 5577
rect 4000 5517 4054 5543
rect 2316 5437 2370 5463
rect 2316 5403 2324 5437
rect 2358 5403 2370 5437
rect 2316 5377 2370 5403
rect 2400 5437 2470 5463
rect 2400 5403 2418 5437
rect 2452 5403 2470 5437
rect 2400 5377 2470 5403
rect 2500 5377 2570 5463
rect 2600 5377 2670 5463
rect 2700 5437 2770 5463
rect 2700 5403 2718 5437
rect 2752 5403 2770 5437
rect 2700 5377 2770 5403
rect 2800 5437 2870 5463
rect 2800 5403 2818 5437
rect 2852 5403 2870 5437
rect 2800 5377 2870 5403
rect 2900 5377 2970 5463
rect 3000 5437 3070 5463
rect 3000 5403 3018 5437
rect 3052 5403 3070 5437
rect 3000 5377 3070 5403
rect 3100 5437 3170 5463
rect 3100 5403 3118 5437
rect 3152 5403 3170 5437
rect 3100 5377 3170 5403
rect 3200 5377 3270 5463
rect 3300 5377 3370 5463
rect 3400 5377 3470 5463
rect 3500 5437 3570 5463
rect 3500 5403 3518 5437
rect 3552 5403 3570 5437
rect 3500 5377 3570 5403
rect 3600 5437 3670 5463
rect 3600 5403 3618 5437
rect 3652 5403 3670 5437
rect 3600 5377 3670 5403
rect 3700 5437 3754 5463
rect 3700 5403 3712 5437
rect 3746 5403 3754 5437
rect 3700 5377 3754 5403
rect 2216 5297 2270 5323
rect 2216 5263 2224 5297
rect 2258 5263 2270 5297
rect 2216 5237 2270 5263
rect 2300 5297 2354 5323
rect 2300 5263 2312 5297
rect 2346 5263 2354 5297
rect 2300 5237 2354 5263
rect 2416 5297 2470 5323
rect 2416 5263 2424 5297
rect 2458 5263 2470 5297
rect 2416 5237 2470 5263
rect 2500 5297 2570 5323
rect 2500 5263 2518 5297
rect 2552 5263 2570 5297
rect 2500 5237 2570 5263
rect 2600 5297 2654 5323
rect 2600 5263 2612 5297
rect 2646 5263 2654 5297
rect 2600 5237 2654 5263
rect 2716 5297 2770 5323
rect 2716 5263 2724 5297
rect 2758 5263 2770 5297
rect 2716 5237 2770 5263
rect 2800 5297 2870 5323
rect 2800 5263 2818 5297
rect 2852 5263 2870 5297
rect 2800 5237 2870 5263
rect 2900 5297 2954 5323
rect 2900 5263 2912 5297
rect 2946 5263 2954 5297
rect 2900 5237 2954 5263
rect 3016 5297 3070 5323
rect 3016 5263 3024 5297
rect 3058 5263 3070 5297
rect 3016 5237 3070 5263
rect 3100 5297 3154 5323
rect 3100 5263 3112 5297
rect 3146 5263 3154 5297
rect 3100 5237 3154 5263
rect 5316 5997 5370 6023
rect 5316 5963 5324 5997
rect 5358 5963 5370 5997
rect 5316 5937 5370 5963
rect 5400 5997 5470 6023
rect 5400 5963 5418 5997
rect 5452 5963 5470 5997
rect 5400 5937 5470 5963
rect 5500 5997 5570 6023
rect 5500 5963 5518 5997
rect 5552 5963 5570 5997
rect 5500 5937 5570 5963
rect 5600 5997 5670 6023
rect 5600 5963 5618 5997
rect 5652 5963 5670 5997
rect 5600 5937 5670 5963
rect 5700 5997 5770 6023
rect 5700 5963 5718 5997
rect 5752 5963 5770 5997
rect 5700 5937 5770 5963
rect 5800 5997 5854 6023
rect 5800 5963 5812 5997
rect 5846 5963 5854 5997
rect 5800 5937 5854 5963
rect 4216 5857 4270 5883
rect 4216 5823 4224 5857
rect 4258 5823 4270 5857
rect 4216 5797 4270 5823
rect 4300 5857 4370 5883
rect 4300 5823 4318 5857
rect 4352 5823 4370 5857
rect 4300 5797 4370 5823
rect 4400 5797 4470 5883
rect 4500 5857 4570 5883
rect 4500 5823 4518 5857
rect 4552 5823 4570 5857
rect 4500 5797 4570 5823
rect 4600 5857 4670 5883
rect 4600 5823 4618 5857
rect 4652 5823 4670 5857
rect 4600 5797 4670 5823
rect 4700 5857 4770 5883
rect 4700 5823 4718 5857
rect 4752 5823 4770 5857
rect 4700 5797 4770 5823
rect 4800 5797 4870 5883
rect 4900 5857 4970 5883
rect 4900 5823 4918 5857
rect 4952 5823 4970 5857
rect 4900 5797 4970 5823
rect 5000 5857 5070 5883
rect 5000 5823 5018 5857
rect 5052 5823 5070 5857
rect 5000 5797 5070 5823
rect 5100 5857 5170 5883
rect 5100 5823 5118 5857
rect 5152 5823 5170 5857
rect 5100 5797 5170 5823
rect 5200 5857 5270 5883
rect 5200 5823 5218 5857
rect 5252 5823 5270 5857
rect 5200 5797 5270 5823
rect 5300 5857 5370 5883
rect 5300 5823 5318 5857
rect 5352 5823 5370 5857
rect 5300 5797 5370 5823
rect 5400 5797 5470 5883
rect 5500 5797 5570 5883
rect 5600 5857 5670 5883
rect 5600 5823 5618 5857
rect 5652 5823 5670 5857
rect 5600 5797 5670 5823
rect 5700 5857 5754 5883
rect 5700 5823 5712 5857
rect 5746 5823 5754 5857
rect 5700 5797 5754 5823
rect 4216 5717 4270 5743
rect 4216 5683 4224 5717
rect 4258 5683 4270 5717
rect 4216 5657 4270 5683
rect 4300 5717 4354 5743
rect 4300 5683 4312 5717
rect 4346 5683 4354 5717
rect 4300 5657 4354 5683
rect 4416 5717 4470 5743
rect 4416 5683 4424 5717
rect 4458 5683 4470 5717
rect 4416 5657 4470 5683
rect 4500 5717 4554 5743
rect 4500 5683 4512 5717
rect 4546 5683 4554 5717
rect 4500 5657 4554 5683
rect 4616 5717 4670 5743
rect 4616 5683 4624 5717
rect 4658 5683 4670 5717
rect 4616 5657 4670 5683
rect 4700 5717 4770 5743
rect 4700 5683 4718 5717
rect 4752 5683 4770 5717
rect 4700 5657 4770 5683
rect 4800 5657 4870 5743
rect 4900 5717 4970 5743
rect 4900 5683 4918 5717
rect 4952 5683 4970 5717
rect 4900 5657 4970 5683
rect 5000 5717 5070 5743
rect 5000 5683 5018 5717
rect 5052 5683 5070 5717
rect 5000 5657 5070 5683
rect 5100 5657 5170 5743
rect 5200 5717 5270 5743
rect 5200 5683 5218 5717
rect 5252 5683 5270 5717
rect 5200 5657 5270 5683
rect 5300 5717 5370 5743
rect 5300 5683 5318 5717
rect 5352 5683 5370 5717
rect 5300 5657 5370 5683
rect 5400 5717 5470 5743
rect 5400 5683 5418 5717
rect 5452 5683 5470 5717
rect 5400 5657 5470 5683
rect 5500 5717 5554 5743
rect 5500 5683 5512 5717
rect 5546 5683 5554 5717
rect 5500 5657 5554 5683
rect 6116 6137 6170 6163
rect 6116 6103 6124 6137
rect 6158 6103 6170 6137
rect 6116 6077 6170 6103
rect 6200 6137 6254 6163
rect 6200 6103 6212 6137
rect 6246 6103 6254 6137
rect 6200 6077 6254 6103
rect 6316 6137 6370 6163
rect 6316 6103 6324 6137
rect 6358 6103 6370 6137
rect 6316 6077 6370 6103
rect 6400 6137 6454 6163
rect 6400 6103 6412 6137
rect 6446 6103 6454 6137
rect 6400 6077 6454 6103
rect 6512 6152 6570 6163
rect 6512 6118 6524 6152
rect 6558 6118 6570 6152
rect 6512 6077 6570 6118
rect 6600 6137 6670 6163
rect 6600 6103 6618 6137
rect 6652 6103 6670 6137
rect 6600 6077 6670 6103
rect 6700 6122 6758 6163
rect 6700 6088 6712 6122
rect 6746 6088 6758 6122
rect 6700 6077 6758 6088
rect 6820 6137 6880 6163
rect 6820 6103 6828 6137
rect 6862 6103 6880 6137
rect 6820 6077 6880 6103
rect 6910 6137 6980 6163
rect 6910 6103 6928 6137
rect 6962 6103 6980 6137
rect 6910 6077 6980 6103
rect 7010 6137 7080 6163
rect 7010 6103 7028 6137
rect 7062 6103 7080 6137
rect 7010 6077 7080 6103
rect 7110 6137 7180 6163
rect 7110 6103 7128 6137
rect 7162 6103 7180 6137
rect 7110 6077 7180 6103
rect 7210 6137 7280 6163
rect 7210 6103 7228 6137
rect 7262 6103 7280 6137
rect 7210 6077 7280 6103
rect 7310 6137 7380 6163
rect 7310 6103 7328 6137
rect 7362 6103 7380 6137
rect 7310 6077 7380 6103
rect 7410 6137 7470 6163
rect 7410 6103 7428 6137
rect 7462 6103 7470 6137
rect 7410 6077 7470 6103
rect 5916 5997 5970 6023
rect 5916 5963 5924 5997
rect 5958 5963 5970 5997
rect 5916 5937 5970 5963
rect 6000 5997 6070 6023
rect 6000 5963 6018 5997
rect 6052 5963 6070 5997
rect 6000 5937 6070 5963
rect 6100 5937 6170 6023
rect 6200 5937 6270 6023
rect 6300 5997 6370 6023
rect 6300 5963 6318 5997
rect 6352 5963 6370 5997
rect 6300 5937 6370 5963
rect 6400 5997 6454 6023
rect 6400 5963 6412 5997
rect 6446 5963 6454 5997
rect 6400 5937 6454 5963
rect 6512 6012 6570 6023
rect 6512 5978 6524 6012
rect 6558 5978 6570 6012
rect 6512 5937 6570 5978
rect 6600 5997 6670 6023
rect 6600 5963 6618 5997
rect 6652 5963 6670 5997
rect 6600 5937 6670 5963
rect 6700 5982 6758 6023
rect 6700 5948 6712 5982
rect 6746 5948 6758 5982
rect 6700 5937 6758 5948
rect 6820 5997 6880 6023
rect 6820 5963 6828 5997
rect 6862 5963 6880 5997
rect 6820 5937 6880 5963
rect 6910 5997 6980 6023
rect 6910 5963 6928 5997
rect 6962 5963 6980 5997
rect 6910 5937 6980 5963
rect 7010 5997 7080 6023
rect 7010 5963 7028 5997
rect 7062 5963 7080 5997
rect 7010 5937 7080 5963
rect 7110 5997 7180 6023
rect 7110 5963 7128 5997
rect 7162 5963 7180 5997
rect 7110 5937 7180 5963
rect 7210 5997 7280 6023
rect 7210 5963 7228 5997
rect 7262 5963 7280 5997
rect 7210 5937 7280 5963
rect 7310 5997 7380 6023
rect 7310 5963 7328 5997
rect 7362 5963 7380 5997
rect 7310 5937 7380 5963
rect 7410 5997 7470 6023
rect 7410 5963 7428 5997
rect 7462 5963 7470 5997
rect 7410 5937 7470 5963
rect 5816 5857 5870 5883
rect 5816 5823 5824 5857
rect 5858 5823 5870 5857
rect 5816 5797 5870 5823
rect 5900 5857 5954 5883
rect 5900 5823 5912 5857
rect 5946 5823 5954 5857
rect 5900 5797 5954 5823
rect 6016 5857 6070 5883
rect 6016 5823 6024 5857
rect 6058 5823 6070 5857
rect 6016 5797 6070 5823
rect 6100 5857 6170 5883
rect 6100 5823 6118 5857
rect 6152 5823 6170 5857
rect 6100 5797 6170 5823
rect 6200 5857 6270 5883
rect 6200 5823 6218 5857
rect 6252 5823 6270 5857
rect 6200 5797 6270 5823
rect 6300 5857 6370 5883
rect 6300 5823 6318 5857
rect 6352 5823 6370 5857
rect 6300 5797 6370 5823
rect 6400 5797 6454 5883
rect 6512 5872 6570 5883
rect 6512 5838 6524 5872
rect 6558 5838 6570 5872
rect 6512 5797 6570 5838
rect 6600 5857 6670 5883
rect 6600 5823 6618 5857
rect 6652 5823 6670 5857
rect 6600 5797 6670 5823
rect 6700 5842 6758 5883
rect 6700 5808 6712 5842
rect 6746 5808 6758 5842
rect 6700 5797 6758 5808
rect 6820 5857 6880 5883
rect 6820 5823 6828 5857
rect 6862 5823 6880 5857
rect 6820 5797 6880 5823
rect 6910 5857 6980 5883
rect 6910 5823 6928 5857
rect 6962 5823 6980 5857
rect 6910 5797 6980 5823
rect 7010 5857 7080 5883
rect 7010 5823 7028 5857
rect 7062 5823 7080 5857
rect 7010 5797 7080 5823
rect 7110 5857 7180 5883
rect 7110 5823 7128 5857
rect 7162 5823 7180 5857
rect 7110 5797 7180 5823
rect 7210 5857 7280 5883
rect 7210 5823 7228 5857
rect 7262 5823 7280 5857
rect 7210 5797 7280 5823
rect 7310 5857 7380 5883
rect 7310 5823 7328 5857
rect 7362 5823 7380 5857
rect 7310 5797 7380 5823
rect 7410 5857 7470 5883
rect 7410 5823 7428 5857
rect 7462 5823 7470 5857
rect 7410 5797 7470 5823
rect 5616 5717 5670 5743
rect 5616 5683 5624 5717
rect 5658 5683 5670 5717
rect 5616 5657 5670 5683
rect 5700 5717 5770 5743
rect 5700 5683 5718 5717
rect 5752 5683 5770 5717
rect 5700 5657 5770 5683
rect 5800 5717 5870 5743
rect 5800 5683 5818 5717
rect 5852 5683 5870 5717
rect 5800 5657 5870 5683
rect 5900 5657 5970 5743
rect 6000 5717 6070 5743
rect 6000 5683 6018 5717
rect 6052 5683 6070 5717
rect 6000 5657 6070 5683
rect 6100 5717 6170 5743
rect 6100 5683 6118 5717
rect 6152 5683 6170 5717
rect 6100 5657 6170 5683
rect 6200 5717 6270 5743
rect 6200 5683 6218 5717
rect 6252 5683 6270 5717
rect 6200 5657 6270 5683
rect 6300 5717 6370 5743
rect 6300 5683 6318 5717
rect 6352 5683 6370 5717
rect 6300 5657 6370 5683
rect 6400 5657 6454 5743
rect 6512 5732 6570 5743
rect 6512 5698 6524 5732
rect 6558 5698 6570 5732
rect 6512 5657 6570 5698
rect 6600 5717 6670 5743
rect 6600 5683 6618 5717
rect 6652 5683 6670 5717
rect 6600 5657 6670 5683
rect 6700 5702 6758 5743
rect 6700 5668 6712 5702
rect 6746 5668 6758 5702
rect 6700 5657 6758 5668
rect 6820 5717 6880 5743
rect 6820 5683 6828 5717
rect 6862 5683 6880 5717
rect 6820 5657 6880 5683
rect 6910 5717 6980 5743
rect 6910 5683 6928 5717
rect 6962 5683 6980 5717
rect 6910 5657 6980 5683
rect 7010 5717 7080 5743
rect 7010 5683 7028 5717
rect 7062 5683 7080 5717
rect 7010 5657 7080 5683
rect 7110 5717 7180 5743
rect 7110 5683 7128 5717
rect 7162 5683 7180 5717
rect 7110 5657 7180 5683
rect 7210 5717 7280 5743
rect 7210 5683 7228 5717
rect 7262 5683 7280 5717
rect 7210 5657 7280 5683
rect 7310 5717 7380 5743
rect 7310 5683 7328 5717
rect 7362 5683 7380 5717
rect 7310 5657 7380 5683
rect 7410 5717 7470 5743
rect 7410 5683 7428 5717
rect 7462 5683 7470 5717
rect 7410 5657 7470 5683
rect 4116 5577 4170 5603
rect 4116 5543 4124 5577
rect 4158 5543 4170 5577
rect 4116 5517 4170 5543
rect 4200 5577 4270 5603
rect 4200 5543 4218 5577
rect 4252 5543 4270 5577
rect 4200 5517 4270 5543
rect 4300 5517 4370 5603
rect 4400 5517 4470 5603
rect 4500 5577 4570 5603
rect 4500 5543 4518 5577
rect 4552 5543 4570 5577
rect 4500 5517 4570 5543
rect 4600 5577 4670 5603
rect 4600 5543 4618 5577
rect 4652 5543 4670 5577
rect 4600 5517 4670 5543
rect 4700 5577 4770 5603
rect 4700 5543 4718 5577
rect 4752 5543 4770 5577
rect 4700 5517 4770 5543
rect 4800 5577 4870 5603
rect 4800 5543 4818 5577
rect 4852 5543 4870 5577
rect 4800 5517 4870 5543
rect 4900 5517 4970 5603
rect 5000 5517 5070 5603
rect 5100 5577 5170 5603
rect 5100 5543 5118 5577
rect 5152 5543 5170 5577
rect 5100 5517 5170 5543
rect 5200 5577 5270 5603
rect 5200 5543 5218 5577
rect 5252 5543 5270 5577
rect 5200 5517 5270 5543
rect 5300 5577 5370 5603
rect 5300 5543 5318 5577
rect 5352 5543 5370 5577
rect 5300 5517 5370 5543
rect 5400 5577 5470 5603
rect 5400 5543 5418 5577
rect 5452 5543 5470 5577
rect 5400 5517 5470 5543
rect 5500 5517 5570 5603
rect 5600 5517 5670 5603
rect 5700 5577 5770 5603
rect 5700 5543 5718 5577
rect 5752 5543 5770 5577
rect 5700 5517 5770 5543
rect 5800 5577 5870 5603
rect 5800 5543 5818 5577
rect 5852 5543 5870 5577
rect 5800 5517 5870 5543
rect 5900 5577 5970 5603
rect 5900 5543 5918 5577
rect 5952 5543 5970 5577
rect 5900 5517 5970 5543
rect 6000 5577 6070 5603
rect 6000 5543 6018 5577
rect 6052 5543 6070 5577
rect 6000 5517 6070 5543
rect 6100 5517 6170 5603
rect 6200 5517 6270 5603
rect 6300 5517 6370 5603
rect 6400 5517 6454 5603
rect 6512 5592 6570 5603
rect 6512 5558 6524 5592
rect 6558 5558 6570 5592
rect 6512 5517 6570 5558
rect 6600 5577 6670 5603
rect 6600 5543 6618 5577
rect 6652 5543 6670 5577
rect 6600 5517 6670 5543
rect 6700 5562 6758 5603
rect 6700 5528 6712 5562
rect 6746 5528 6758 5562
rect 6700 5517 6758 5528
rect 6820 5577 6880 5603
rect 6820 5543 6828 5577
rect 6862 5543 6880 5577
rect 6820 5517 6880 5543
rect 6910 5577 6980 5603
rect 6910 5543 6928 5577
rect 6962 5543 6980 5577
rect 6910 5517 6980 5543
rect 7010 5577 7080 5603
rect 7010 5543 7028 5577
rect 7062 5543 7080 5577
rect 7010 5517 7080 5543
rect 7110 5577 7180 5603
rect 7110 5543 7128 5577
rect 7162 5543 7180 5577
rect 7110 5517 7180 5543
rect 7210 5577 7280 5603
rect 7210 5543 7228 5577
rect 7262 5543 7280 5577
rect 7210 5517 7280 5543
rect 7310 5577 7380 5603
rect 7310 5543 7328 5577
rect 7362 5543 7380 5577
rect 7310 5517 7380 5543
rect 7410 5577 7470 5603
rect 7410 5543 7428 5577
rect 7462 5543 7470 5577
rect 7410 5517 7470 5543
rect 3816 5437 3870 5463
rect 3816 5403 3824 5437
rect 3858 5403 3870 5437
rect 3816 5377 3870 5403
rect 3900 5437 3970 5463
rect 3900 5403 3918 5437
rect 3952 5403 3970 5437
rect 3900 5377 3970 5403
rect 4000 5437 4070 5463
rect 4000 5403 4018 5437
rect 4052 5403 4070 5437
rect 4000 5377 4070 5403
rect 4100 5437 4170 5463
rect 4100 5403 4118 5437
rect 4152 5403 4170 5437
rect 4100 5377 4170 5403
rect 4200 5437 4270 5463
rect 4200 5403 4218 5437
rect 4252 5403 4270 5437
rect 4200 5377 4270 5403
rect 4300 5377 4370 5463
rect 4400 5437 4470 5463
rect 4400 5403 4418 5437
rect 4452 5403 4470 5437
rect 4400 5377 4470 5403
rect 4500 5437 4570 5463
rect 4500 5403 4518 5437
rect 4552 5403 4570 5437
rect 4500 5377 4570 5403
rect 4600 5437 4670 5463
rect 4600 5403 4618 5437
rect 4652 5403 4670 5437
rect 4600 5377 4670 5403
rect 4700 5437 4770 5463
rect 4700 5403 4718 5437
rect 4752 5403 4770 5437
rect 4700 5377 4770 5403
rect 4800 5377 4870 5463
rect 4900 5377 4970 5463
rect 5000 5437 5070 5463
rect 5000 5403 5018 5437
rect 5052 5403 5070 5437
rect 5000 5377 5070 5403
rect 5100 5437 5154 5463
rect 5100 5403 5112 5437
rect 5146 5403 5154 5437
rect 5100 5377 5154 5403
rect 5216 5437 5270 5463
rect 5216 5403 5224 5437
rect 5258 5403 5270 5437
rect 5216 5377 5270 5403
rect 5300 5437 5354 5463
rect 5300 5403 5312 5437
rect 5346 5403 5354 5437
rect 5300 5377 5354 5403
rect 3216 5297 3270 5323
rect 3216 5263 3224 5297
rect 3258 5263 3270 5297
rect 3216 5237 3270 5263
rect 3300 5297 3370 5323
rect 3300 5263 3318 5297
rect 3352 5263 3370 5297
rect 3300 5237 3370 5263
rect 3400 5237 3470 5323
rect 3500 5297 3570 5323
rect 3500 5263 3518 5297
rect 3552 5263 3570 5297
rect 3500 5237 3570 5263
rect 3600 5297 3670 5323
rect 3600 5263 3618 5297
rect 3652 5263 3670 5297
rect 3600 5237 3670 5263
rect 3700 5237 3770 5323
rect 3800 5237 3870 5323
rect 3900 5237 3970 5323
rect 4000 5297 4070 5323
rect 4000 5263 4018 5297
rect 4052 5263 4070 5297
rect 4000 5237 4070 5263
rect 4100 5297 4170 5323
rect 4100 5263 4118 5297
rect 4152 5263 4170 5297
rect 4100 5237 4170 5263
rect 4200 5297 4270 5323
rect 4200 5263 4218 5297
rect 4252 5263 4270 5297
rect 4200 5237 4270 5263
rect 4300 5297 4370 5323
rect 4300 5263 4318 5297
rect 4352 5263 4370 5297
rect 4300 5237 4370 5263
rect 4400 5297 4470 5323
rect 4400 5263 4418 5297
rect 4452 5263 4470 5297
rect 4400 5237 4470 5263
rect 4500 5297 4570 5323
rect 4500 5263 4518 5297
rect 4552 5263 4570 5297
rect 4500 5237 4570 5263
rect 4600 5237 4670 5323
rect 4700 5297 4770 5323
rect 4700 5263 4718 5297
rect 4752 5263 4770 5297
rect 4700 5237 4770 5263
rect 4800 5297 4870 5323
rect 4800 5263 4818 5297
rect 4852 5263 4870 5297
rect 4800 5237 4870 5263
rect 4900 5297 4970 5323
rect 4900 5263 4918 5297
rect 4952 5263 4970 5297
rect 4900 5237 4970 5263
rect 5000 5297 5070 5323
rect 5000 5263 5018 5297
rect 5052 5263 5070 5297
rect 5000 5237 5070 5263
rect 5100 5297 5170 5323
rect 5100 5263 5118 5297
rect 5152 5263 5170 5297
rect 5100 5237 5170 5263
rect 5200 5297 5254 5323
rect 5200 5263 5212 5297
rect 5246 5263 5254 5297
rect 5200 5237 5254 5263
rect 2216 5157 2270 5183
rect 2216 5123 2224 5157
rect 2258 5123 2270 5157
rect 2216 5097 2270 5123
rect 2300 5157 2370 5183
rect 2300 5123 2318 5157
rect 2352 5123 2370 5157
rect 2300 5097 2370 5123
rect 2400 5157 2470 5183
rect 2400 5123 2418 5157
rect 2452 5123 2470 5157
rect 2400 5097 2470 5123
rect 2500 5157 2570 5183
rect 2500 5123 2518 5157
rect 2552 5123 2570 5157
rect 2500 5097 2570 5123
rect 2600 5097 2670 5183
rect 2700 5097 2770 5183
rect 2800 5157 2870 5183
rect 2800 5123 2818 5157
rect 2852 5123 2870 5157
rect 2800 5097 2870 5123
rect 2900 5157 2970 5183
rect 2900 5123 2918 5157
rect 2952 5123 2970 5157
rect 2900 5097 2970 5123
rect 3000 5157 3070 5183
rect 3000 5123 3018 5157
rect 3052 5123 3070 5157
rect 3000 5097 3070 5123
rect 3100 5157 3170 5183
rect 3100 5123 3118 5157
rect 3152 5123 3170 5157
rect 3100 5097 3170 5123
rect 3200 5097 3270 5183
rect 3300 5097 3370 5183
rect 3400 5097 3470 5183
rect 3500 5157 3570 5183
rect 3500 5123 3518 5157
rect 3552 5123 3570 5157
rect 3500 5097 3570 5123
rect 3600 5157 3670 5183
rect 3600 5123 3618 5157
rect 3652 5123 3670 5157
rect 3600 5097 3670 5123
rect 3700 5097 3770 5183
rect 3800 5097 3870 5183
rect 3900 5097 3970 5183
rect 4000 5157 4070 5183
rect 4000 5123 4018 5157
rect 4052 5123 4070 5157
rect 4000 5097 4070 5123
rect 4100 5157 4170 5183
rect 4100 5123 4118 5157
rect 4152 5123 4170 5157
rect 4100 5097 4170 5123
rect 4200 5157 4270 5183
rect 4200 5123 4218 5157
rect 4252 5123 4270 5157
rect 4200 5097 4270 5123
rect 4300 5157 4354 5183
rect 4300 5123 4312 5157
rect 4346 5123 4354 5157
rect 4300 5097 4354 5123
rect 1216 4787 1270 4813
rect 1216 4753 1224 4787
rect 1258 4753 1270 4787
rect 1216 4727 1270 4753
rect 1300 4787 1370 4813
rect 1300 4753 1318 4787
rect 1352 4753 1370 4787
rect 1300 4727 1370 4753
rect 1400 4727 1470 4813
rect 1500 4787 1570 4813
rect 1500 4753 1518 4787
rect 1552 4753 1570 4787
rect 1500 4727 1570 4753
rect 1600 4787 1670 4813
rect 1600 4753 1618 4787
rect 1652 4753 1670 4787
rect 1600 4727 1670 4753
rect 1700 4727 1770 4813
rect 1800 4727 1870 4813
rect 1900 4727 1970 4813
rect 2000 4787 2070 4813
rect 2000 4753 2018 4787
rect 2052 4753 2070 4787
rect 2000 4727 2070 4753
rect 2100 4787 2170 4813
rect 2100 4753 2118 4787
rect 2152 4753 2170 4787
rect 2100 4727 2170 4753
rect 2200 4787 2270 4813
rect 2200 4753 2218 4787
rect 2252 4753 2270 4787
rect 2200 4727 2270 4753
rect 2300 4727 2370 4813
rect 2400 4727 2470 4813
rect 2500 4727 2570 4813
rect 2600 4727 2670 4813
rect 2700 4787 2770 4813
rect 2700 4753 2718 4787
rect 2752 4753 2770 4787
rect 2700 4727 2770 4753
rect 2800 4787 2854 4813
rect 2800 4753 2812 4787
rect 2846 4753 2854 4787
rect 2800 4727 2854 4753
rect 16 4647 70 4673
rect 16 4613 24 4647
rect 58 4613 70 4647
rect 16 4587 70 4613
rect 100 4647 170 4673
rect 100 4613 118 4647
rect 152 4613 170 4647
rect 100 4587 170 4613
rect 200 4587 270 4673
rect 300 4647 370 4673
rect 300 4613 318 4647
rect 352 4613 370 4647
rect 300 4587 370 4613
rect 400 4647 470 4673
rect 400 4613 418 4647
rect 452 4613 470 4647
rect 400 4587 470 4613
rect 500 4647 570 4673
rect 500 4613 518 4647
rect 552 4613 570 4647
rect 500 4587 570 4613
rect 600 4587 670 4673
rect 700 4587 770 4673
rect 800 4647 870 4673
rect 800 4613 818 4647
rect 852 4613 870 4647
rect 800 4587 870 4613
rect 900 4647 970 4673
rect 900 4613 918 4647
rect 952 4613 970 4647
rect 900 4587 970 4613
rect 1000 4587 1070 4673
rect 1100 4587 1170 4673
rect 1200 4647 1270 4673
rect 1200 4613 1218 4647
rect 1252 4613 1270 4647
rect 1200 4587 1270 4613
rect 1300 4647 1370 4673
rect 1300 4613 1318 4647
rect 1352 4613 1370 4647
rect 1300 4587 1370 4613
rect 1400 4587 1470 4673
rect 1500 4647 1570 4673
rect 1500 4613 1518 4647
rect 1552 4613 1570 4647
rect 1500 4587 1570 4613
rect 1600 4647 1670 4673
rect 1600 4613 1618 4647
rect 1652 4613 1670 4647
rect 1600 4587 1670 4613
rect 1700 4647 1770 4673
rect 1700 4613 1718 4647
rect 1752 4613 1770 4647
rect 1700 4587 1770 4613
rect 1800 4647 1854 4673
rect 1800 4613 1812 4647
rect 1846 4613 1854 4647
rect 1800 4587 1854 4613
rect 16 4507 70 4533
rect 16 4473 24 4507
rect 58 4473 70 4507
rect 16 4447 70 4473
rect 100 4507 154 4533
rect 100 4473 112 4507
rect 146 4473 154 4507
rect 100 4447 154 4473
rect 216 4507 270 4533
rect 216 4473 224 4507
rect 258 4473 270 4507
rect 216 4447 270 4473
rect 300 4507 370 4533
rect 300 4473 318 4507
rect 352 4473 370 4507
rect 300 4447 370 4473
rect 400 4447 470 4533
rect 500 4447 570 4533
rect 600 4447 670 4533
rect 700 4507 770 4533
rect 700 4473 718 4507
rect 752 4473 770 4507
rect 700 4447 770 4473
rect 800 4507 870 4533
rect 800 4473 818 4507
rect 852 4473 870 4507
rect 800 4447 870 4473
rect 900 4507 970 4533
rect 900 4473 918 4507
rect 952 4473 970 4507
rect 900 4447 970 4473
rect 1000 4447 1070 4533
rect 1100 4447 1170 4533
rect 1200 4447 1270 4533
rect 1300 4507 1370 4533
rect 1300 4473 1318 4507
rect 1352 4473 1370 4507
rect 1300 4447 1370 4473
rect 1400 4507 1470 4533
rect 1400 4473 1418 4507
rect 1452 4473 1470 4507
rect 1400 4447 1470 4473
rect 1500 4507 1570 4533
rect 1500 4473 1518 4507
rect 1552 4473 1570 4507
rect 1500 4447 1570 4473
rect 1600 4507 1654 4533
rect 1600 4473 1612 4507
rect 1646 4473 1654 4507
rect 1600 4447 1654 4473
rect 16 4367 70 4393
rect 16 4333 24 4367
rect 58 4333 70 4367
rect 16 4307 70 4333
rect 100 4367 170 4393
rect 100 4333 118 4367
rect 152 4333 170 4367
rect 100 4307 170 4333
rect 200 4367 270 4393
rect 200 4333 218 4367
rect 252 4333 270 4367
rect 200 4307 270 4333
rect 300 4367 370 4393
rect 300 4333 318 4367
rect 352 4333 370 4367
rect 300 4307 370 4333
rect 400 4367 454 4393
rect 400 4333 412 4367
rect 446 4333 454 4367
rect 400 4307 454 4333
rect 16 4227 70 4253
rect 16 4193 24 4227
rect 58 4193 70 4227
rect 16 4167 70 4193
rect 100 4227 154 4253
rect 100 4193 112 4227
rect 146 4193 154 4227
rect 100 4167 154 4193
rect 216 4227 270 4253
rect 216 4193 224 4227
rect 258 4193 270 4227
rect 216 4167 270 4193
rect 300 4227 354 4253
rect 300 4193 312 4227
rect 346 4193 354 4227
rect 300 4167 354 4193
rect 516 4367 570 4393
rect 516 4333 524 4367
rect 558 4333 570 4367
rect 516 4307 570 4333
rect 600 4367 670 4393
rect 600 4333 618 4367
rect 652 4333 670 4367
rect 600 4307 670 4333
rect 700 4367 754 4393
rect 700 4333 712 4367
rect 746 4333 754 4367
rect 700 4307 754 4333
rect 1916 4647 1970 4673
rect 1916 4613 1924 4647
rect 1958 4613 1970 4647
rect 1916 4587 1970 4613
rect 2000 4647 2054 4673
rect 2000 4613 2012 4647
rect 2046 4613 2054 4647
rect 2000 4587 2054 4613
rect 4416 5157 4470 5183
rect 4416 5123 4424 5157
rect 4458 5123 4470 5157
rect 4416 5097 4470 5123
rect 4500 5157 4570 5183
rect 4500 5123 4518 5157
rect 4552 5123 4570 5157
rect 4500 5097 4570 5123
rect 4600 5157 4670 5183
rect 4600 5123 4618 5157
rect 4652 5123 4670 5157
rect 4600 5097 4670 5123
rect 4700 5157 4754 5183
rect 4700 5123 4712 5157
rect 4746 5123 4754 5157
rect 4700 5097 4754 5123
rect 5416 5437 5470 5463
rect 5416 5403 5424 5437
rect 5458 5403 5470 5437
rect 5416 5377 5470 5403
rect 5500 5437 5554 5463
rect 5500 5403 5512 5437
rect 5546 5403 5554 5437
rect 5500 5377 5554 5403
rect 5316 5297 5370 5323
rect 5316 5263 5324 5297
rect 5358 5263 5370 5297
rect 5316 5237 5370 5263
rect 5400 5297 5454 5323
rect 5400 5263 5412 5297
rect 5446 5263 5454 5297
rect 5400 5237 5454 5263
rect 5616 5437 5670 5463
rect 5616 5403 5624 5437
rect 5658 5403 5670 5437
rect 5616 5377 5670 5403
rect 5700 5437 5754 5463
rect 5700 5403 5712 5437
rect 5746 5403 5754 5437
rect 5700 5377 5754 5403
rect 5816 5437 5870 5463
rect 5816 5403 5824 5437
rect 5858 5403 5870 5437
rect 5816 5377 5870 5403
rect 5900 5437 5970 5463
rect 5900 5403 5918 5437
rect 5952 5403 5970 5437
rect 5900 5377 5970 5403
rect 6000 5437 6070 5463
rect 6000 5403 6018 5437
rect 6052 5403 6070 5437
rect 6000 5377 6070 5403
rect 6100 5377 6170 5463
rect 6200 5377 6270 5463
rect 6300 5377 6370 5463
rect 6400 5377 6454 5463
rect 6512 5452 6570 5463
rect 6512 5418 6524 5452
rect 6558 5418 6570 5452
rect 6512 5377 6570 5418
rect 6600 5437 6670 5463
rect 6600 5403 6618 5437
rect 6652 5403 6670 5437
rect 6600 5377 6670 5403
rect 6700 5422 6758 5463
rect 6700 5388 6712 5422
rect 6746 5388 6758 5422
rect 6700 5377 6758 5388
rect 6820 5437 6880 5463
rect 6820 5403 6828 5437
rect 6862 5403 6880 5437
rect 6820 5377 6880 5403
rect 6910 5437 6980 5463
rect 6910 5403 6928 5437
rect 6962 5403 6980 5437
rect 6910 5377 6980 5403
rect 7010 5437 7080 5463
rect 7010 5403 7028 5437
rect 7062 5403 7080 5437
rect 7010 5377 7080 5403
rect 7110 5437 7180 5463
rect 7110 5403 7128 5437
rect 7162 5403 7180 5437
rect 7110 5377 7180 5403
rect 7210 5437 7280 5463
rect 7210 5403 7228 5437
rect 7262 5403 7280 5437
rect 7210 5377 7280 5403
rect 7310 5437 7380 5463
rect 7310 5403 7328 5437
rect 7362 5403 7380 5437
rect 7310 5377 7380 5403
rect 7410 5437 7470 5463
rect 7410 5403 7428 5437
rect 7462 5403 7470 5437
rect 7410 5377 7470 5403
rect 5516 5297 5570 5323
rect 5516 5263 5524 5297
rect 5558 5263 5570 5297
rect 5516 5237 5570 5263
rect 5600 5297 5670 5323
rect 5600 5263 5618 5297
rect 5652 5263 5670 5297
rect 5600 5237 5670 5263
rect 5700 5237 5770 5323
rect 5800 5297 5870 5323
rect 5800 5263 5818 5297
rect 5852 5263 5870 5297
rect 5800 5237 5870 5263
rect 5900 5297 5970 5323
rect 5900 5263 5918 5297
rect 5952 5263 5970 5297
rect 5900 5237 5970 5263
rect 6000 5237 6070 5323
rect 6100 5237 6170 5323
rect 6200 5297 6270 5323
rect 6200 5263 6218 5297
rect 6252 5263 6270 5297
rect 6200 5237 6270 5263
rect 6300 5297 6370 5323
rect 6300 5263 6318 5297
rect 6352 5263 6370 5297
rect 6300 5237 6370 5263
rect 6400 5297 6454 5323
rect 6400 5263 6412 5297
rect 6446 5263 6454 5297
rect 6400 5237 6454 5263
rect 6512 5312 6570 5323
rect 6512 5278 6524 5312
rect 6558 5278 6570 5312
rect 6512 5237 6570 5278
rect 6600 5297 6670 5323
rect 6600 5263 6618 5297
rect 6652 5263 6670 5297
rect 6600 5237 6670 5263
rect 6700 5282 6758 5323
rect 6700 5248 6712 5282
rect 6746 5248 6758 5282
rect 6700 5237 6758 5248
rect 6820 5297 6880 5323
rect 6820 5263 6828 5297
rect 6862 5263 6880 5297
rect 6820 5237 6880 5263
rect 6910 5297 6980 5323
rect 6910 5263 6928 5297
rect 6962 5263 6980 5297
rect 6910 5237 6980 5263
rect 7010 5297 7080 5323
rect 7010 5263 7028 5297
rect 7062 5263 7080 5297
rect 7010 5237 7080 5263
rect 7110 5297 7180 5323
rect 7110 5263 7128 5297
rect 7162 5263 7180 5297
rect 7110 5237 7180 5263
rect 7210 5297 7280 5323
rect 7210 5263 7228 5297
rect 7262 5263 7280 5297
rect 7210 5237 7280 5263
rect 7310 5297 7380 5323
rect 7310 5263 7328 5297
rect 7362 5263 7380 5297
rect 7310 5237 7380 5263
rect 7410 5297 7470 5323
rect 7410 5263 7428 5297
rect 7462 5263 7470 5297
rect 7410 5237 7470 5263
rect 4816 5157 4870 5183
rect 4816 5123 4824 5157
rect 4858 5123 4870 5157
rect 4816 5097 4870 5123
rect 4900 5157 4970 5183
rect 4900 5123 4918 5157
rect 4952 5123 4970 5157
rect 4900 5097 4970 5123
rect 5000 5157 5070 5183
rect 5000 5123 5018 5157
rect 5052 5123 5070 5157
rect 5000 5097 5070 5123
rect 5100 5157 5170 5183
rect 5100 5123 5118 5157
rect 5152 5123 5170 5157
rect 5100 5097 5170 5123
rect 5200 5157 5270 5183
rect 5200 5123 5218 5157
rect 5252 5123 5270 5157
rect 5200 5097 5270 5123
rect 5300 5097 5370 5183
rect 5400 5097 5470 5183
rect 5500 5157 5570 5183
rect 5500 5123 5518 5157
rect 5552 5123 5570 5157
rect 5500 5097 5570 5123
rect 5600 5157 5670 5183
rect 5600 5123 5618 5157
rect 5652 5123 5670 5157
rect 5600 5097 5670 5123
rect 5700 5157 5754 5183
rect 5700 5123 5712 5157
rect 5746 5123 5754 5157
rect 5700 5097 5754 5123
rect 2916 4787 2970 4813
rect 2916 4753 2924 4787
rect 2958 4753 2970 4787
rect 2916 4727 2970 4753
rect 3000 4787 3070 4813
rect 3000 4753 3018 4787
rect 3052 4753 3070 4787
rect 3000 4727 3070 4753
rect 3100 4727 3170 4813
rect 3200 4727 3270 4813
rect 3300 4727 3370 4813
rect 3400 4787 3470 4813
rect 3400 4753 3418 4787
rect 3452 4753 3470 4787
rect 3400 4727 3470 4753
rect 3500 4787 3570 4813
rect 3500 4753 3518 4787
rect 3552 4753 3570 4787
rect 3500 4727 3570 4753
rect 3600 4787 3670 4813
rect 3600 4753 3618 4787
rect 3652 4753 3670 4787
rect 3600 4727 3670 4753
rect 3700 4727 3770 4813
rect 3800 4727 3870 4813
rect 3900 4727 3970 4813
rect 4000 4727 4070 4813
rect 4100 4727 4170 4813
rect 4200 4787 4270 4813
rect 4200 4753 4218 4787
rect 4252 4753 4270 4787
rect 4200 4727 4270 4753
rect 4300 4787 4370 4813
rect 4300 4753 4318 4787
rect 4352 4753 4370 4787
rect 4300 4727 4370 4753
rect 4400 4727 4470 4813
rect 4500 4787 4570 4813
rect 4500 4753 4518 4787
rect 4552 4753 4570 4787
rect 4500 4727 4570 4753
rect 4600 4787 4654 4813
rect 4600 4753 4612 4787
rect 4646 4753 4654 4787
rect 4600 4727 4654 4753
rect 2116 4647 2170 4673
rect 2116 4613 2124 4647
rect 2158 4613 2170 4647
rect 2116 4587 2170 4613
rect 2200 4647 2270 4673
rect 2200 4613 2218 4647
rect 2252 4613 2270 4647
rect 2200 4587 2270 4613
rect 2300 4587 2370 4673
rect 2400 4587 2470 4673
rect 2500 4647 2570 4673
rect 2500 4613 2518 4647
rect 2552 4613 2570 4647
rect 2500 4587 2570 4613
rect 2600 4647 2670 4673
rect 2600 4613 2618 4647
rect 2652 4613 2670 4647
rect 2600 4587 2670 4613
rect 2700 4587 2770 4673
rect 2800 4647 2870 4673
rect 2800 4613 2818 4647
rect 2852 4613 2870 4647
rect 2800 4587 2870 4613
rect 2900 4647 2970 4673
rect 2900 4613 2918 4647
rect 2952 4613 2970 4647
rect 2900 4587 2970 4613
rect 3000 4647 3070 4673
rect 3000 4613 3018 4647
rect 3052 4613 3070 4647
rect 3000 4587 3070 4613
rect 3100 4647 3170 4673
rect 3100 4613 3118 4647
rect 3152 4613 3170 4647
rect 3100 4587 3170 4613
rect 3200 4647 3254 4673
rect 3200 4613 3212 4647
rect 3246 4613 3254 4647
rect 3200 4587 3254 4613
rect 1716 4507 1770 4533
rect 1716 4473 1724 4507
rect 1758 4473 1770 4507
rect 1716 4447 1770 4473
rect 1800 4507 1870 4533
rect 1800 4473 1818 4507
rect 1852 4473 1870 4507
rect 1800 4447 1870 4473
rect 1900 4447 1970 4533
rect 2000 4507 2070 4533
rect 2000 4473 2018 4507
rect 2052 4473 2070 4507
rect 2000 4447 2070 4473
rect 2100 4507 2170 4533
rect 2100 4473 2118 4507
rect 2152 4473 2170 4507
rect 2100 4447 2170 4473
rect 2200 4447 2270 4533
rect 2300 4507 2370 4533
rect 2300 4473 2318 4507
rect 2352 4473 2370 4507
rect 2300 4447 2370 4473
rect 2400 4507 2454 4533
rect 2400 4473 2412 4507
rect 2446 4473 2454 4507
rect 2400 4447 2454 4473
rect 816 4367 870 4393
rect 816 4333 824 4367
rect 858 4333 870 4367
rect 816 4307 870 4333
rect 900 4367 970 4393
rect 900 4333 918 4367
rect 952 4333 970 4367
rect 900 4307 970 4333
rect 1000 4367 1070 4393
rect 1000 4333 1018 4367
rect 1052 4333 1070 4367
rect 1000 4307 1070 4333
rect 1100 4307 1170 4393
rect 1200 4307 1270 4393
rect 1300 4307 1370 4393
rect 1400 4307 1470 4393
rect 1500 4307 1570 4393
rect 1600 4367 1670 4393
rect 1600 4333 1618 4367
rect 1652 4333 1670 4367
rect 1600 4307 1670 4333
rect 1700 4367 1770 4393
rect 1700 4333 1718 4367
rect 1752 4333 1770 4367
rect 1700 4307 1770 4333
rect 1800 4307 1870 4393
rect 1900 4307 1970 4393
rect 2000 4367 2070 4393
rect 2000 4333 2018 4367
rect 2052 4333 2070 4367
rect 2000 4307 2070 4333
rect 2100 4367 2170 4393
rect 2100 4333 2118 4367
rect 2152 4333 2170 4367
rect 2100 4307 2170 4333
rect 2200 4307 2270 4393
rect 2300 4367 2370 4393
rect 2300 4333 2318 4367
rect 2352 4333 2370 4367
rect 2300 4307 2370 4333
rect 2400 4367 2454 4393
rect 2400 4333 2412 4367
rect 2446 4333 2454 4367
rect 2400 4307 2454 4333
rect 416 4227 470 4253
rect 416 4193 424 4227
rect 458 4193 470 4227
rect 416 4167 470 4193
rect 500 4227 570 4253
rect 500 4193 518 4227
rect 552 4193 570 4227
rect 500 4167 570 4193
rect 600 4167 670 4253
rect 700 4167 770 4253
rect 800 4167 870 4253
rect 900 4227 970 4253
rect 900 4193 918 4227
rect 952 4193 970 4227
rect 900 4167 970 4193
rect 1000 4227 1070 4253
rect 1000 4193 1018 4227
rect 1052 4193 1070 4227
rect 1000 4167 1070 4193
rect 1100 4227 1170 4253
rect 1100 4193 1118 4227
rect 1152 4193 1170 4227
rect 1100 4167 1170 4193
rect 1200 4227 1270 4253
rect 1200 4193 1218 4227
rect 1252 4193 1270 4227
rect 1200 4167 1270 4193
rect 1300 4227 1370 4253
rect 1300 4193 1318 4227
rect 1352 4193 1370 4227
rect 1300 4167 1370 4193
rect 1400 4227 1454 4253
rect 1400 4193 1412 4227
rect 1446 4193 1454 4227
rect 1400 4167 1454 4193
rect 16 4087 70 4113
rect 16 4053 24 4087
rect 58 4053 70 4087
rect 16 4027 70 4053
rect 100 4087 170 4113
rect 100 4053 118 4087
rect 152 4053 170 4087
rect 100 4027 170 4053
rect 200 4027 270 4113
rect 300 4087 370 4113
rect 300 4053 318 4087
rect 352 4053 370 4087
rect 300 4027 370 4053
rect 400 4087 454 4113
rect 400 4053 412 4087
rect 446 4053 454 4087
rect 400 4027 454 4053
rect 516 4087 570 4113
rect 516 4053 524 4087
rect 558 4053 570 4087
rect 516 4027 570 4053
rect 600 4087 654 4113
rect 600 4053 612 4087
rect 646 4053 654 4087
rect 600 4027 654 4053
rect 16 3887 70 3973
rect 100 3887 170 3973
rect 200 3947 270 3973
rect 200 3913 218 3947
rect 252 3913 270 3947
rect 200 3887 270 3913
rect 300 3947 370 3973
rect 300 3913 318 3947
rect 352 3913 370 3947
rect 300 3887 370 3913
rect 400 3947 470 3973
rect 400 3913 418 3947
rect 452 3913 470 3947
rect 400 3887 470 3913
rect 500 3947 554 3973
rect 500 3913 512 3947
rect 546 3913 554 3947
rect 500 3887 554 3913
rect 3316 4647 3370 4673
rect 3316 4613 3324 4647
rect 3358 4613 3370 4647
rect 3316 4587 3370 4613
rect 3400 4647 3470 4673
rect 3400 4613 3418 4647
rect 3452 4613 3470 4647
rect 3400 4587 3470 4613
rect 3500 4647 3570 4673
rect 3500 4613 3518 4647
rect 3552 4613 3570 4647
rect 3500 4587 3570 4613
rect 3600 4587 3670 4673
rect 3700 4647 3770 4673
rect 3700 4613 3718 4647
rect 3752 4613 3770 4647
rect 3700 4587 3770 4613
rect 3800 4647 3870 4673
rect 3800 4613 3818 4647
rect 3852 4613 3870 4647
rect 3800 4587 3870 4613
rect 3900 4647 3970 4673
rect 3900 4613 3918 4647
rect 3952 4613 3970 4647
rect 3900 4587 3970 4613
rect 4000 4587 4070 4673
rect 4100 4647 4170 4673
rect 4100 4613 4118 4647
rect 4152 4613 4170 4647
rect 4100 4587 4170 4613
rect 4200 4647 4270 4673
rect 4200 4613 4218 4647
rect 4252 4613 4270 4647
rect 4200 4587 4270 4613
rect 4300 4647 4370 4673
rect 4300 4613 4318 4647
rect 4352 4613 4370 4647
rect 4300 4587 4370 4613
rect 4400 4647 4470 4673
rect 4400 4613 4418 4647
rect 4452 4613 4470 4647
rect 4400 4587 4470 4613
rect 4500 4647 4554 4673
rect 4500 4613 4512 4647
rect 4546 4613 4554 4647
rect 4500 4587 4554 4613
rect 2516 4507 2570 4533
rect 2516 4473 2524 4507
rect 2558 4473 2570 4507
rect 2516 4447 2570 4473
rect 2600 4507 2670 4533
rect 2600 4473 2618 4507
rect 2652 4473 2670 4507
rect 2600 4447 2670 4473
rect 2700 4447 2770 4533
rect 2800 4507 2870 4533
rect 2800 4473 2818 4507
rect 2852 4473 2870 4507
rect 2800 4447 2870 4473
rect 2900 4507 2970 4533
rect 2900 4473 2918 4507
rect 2952 4473 2970 4507
rect 2900 4447 2970 4473
rect 3000 4507 3070 4533
rect 3000 4473 3018 4507
rect 3052 4473 3070 4507
rect 3000 4447 3070 4473
rect 3100 4447 3170 4533
rect 3200 4507 3270 4533
rect 3200 4473 3218 4507
rect 3252 4473 3270 4507
rect 3200 4447 3270 4473
rect 3300 4507 3354 4533
rect 3300 4473 3312 4507
rect 3346 4473 3354 4507
rect 3300 4447 3354 4473
rect 2516 4367 2570 4393
rect 2516 4333 2524 4367
rect 2558 4333 2570 4367
rect 2516 4307 2570 4333
rect 2600 4367 2670 4393
rect 2600 4333 2618 4367
rect 2652 4333 2670 4367
rect 2600 4307 2670 4333
rect 2700 4367 2770 4393
rect 2700 4333 2718 4367
rect 2752 4333 2770 4367
rect 2700 4307 2770 4333
rect 2800 4367 2854 4393
rect 2800 4333 2812 4367
rect 2846 4333 2854 4367
rect 2800 4307 2854 4333
rect 2916 4367 2970 4393
rect 2916 4333 2924 4367
rect 2958 4333 2970 4367
rect 2916 4307 2970 4333
rect 3000 4367 3070 4393
rect 3000 4333 3018 4367
rect 3052 4333 3070 4367
rect 3000 4307 3070 4333
rect 3100 4367 3170 4393
rect 3100 4333 3118 4367
rect 3152 4333 3170 4367
rect 3100 4307 3170 4333
rect 3200 4367 3254 4393
rect 3200 4333 3212 4367
rect 3246 4333 3254 4367
rect 3200 4307 3254 4333
rect 3416 4507 3470 4533
rect 3416 4473 3424 4507
rect 3458 4473 3470 4507
rect 3416 4447 3470 4473
rect 3500 4507 3570 4533
rect 3500 4473 3518 4507
rect 3552 4473 3570 4507
rect 3500 4447 3570 4473
rect 3600 4447 3670 4533
rect 3700 4507 3770 4533
rect 3700 4473 3718 4507
rect 3752 4473 3770 4507
rect 3700 4447 3770 4473
rect 3800 4507 3870 4533
rect 3800 4473 3818 4507
rect 3852 4473 3870 4507
rect 3800 4447 3870 4473
rect 3900 4447 3970 4533
rect 4000 4447 4070 4533
rect 4100 4507 4170 4533
rect 4100 4473 4118 4507
rect 4152 4473 4170 4507
rect 4100 4447 4170 4473
rect 4200 4507 4270 4533
rect 4200 4473 4218 4507
rect 4252 4473 4270 4507
rect 4200 4447 4270 4473
rect 4300 4507 4354 4533
rect 4300 4473 4312 4507
rect 4346 4473 4354 4507
rect 4300 4447 4354 4473
rect 4716 4787 4770 4813
rect 4716 4753 4724 4787
rect 4758 4753 4770 4787
rect 4716 4727 4770 4753
rect 4800 4787 4870 4813
rect 4800 4753 4818 4787
rect 4852 4753 4870 4787
rect 4800 4727 4870 4753
rect 4900 4727 4970 4813
rect 5000 4727 5070 4813
rect 5100 4787 5170 4813
rect 5100 4753 5118 4787
rect 5152 4753 5170 4787
rect 5100 4727 5170 4753
rect 5200 4787 5270 4813
rect 5200 4753 5218 4787
rect 5252 4753 5270 4787
rect 5200 4727 5270 4753
rect 5300 4787 5370 4813
rect 5300 4753 5318 4787
rect 5352 4753 5370 4787
rect 5300 4727 5370 4753
rect 5400 4787 5454 4813
rect 5400 4753 5412 4787
rect 5446 4753 5454 4787
rect 5400 4727 5454 4753
rect 5816 5157 5870 5183
rect 5816 5123 5824 5157
rect 5858 5123 5870 5157
rect 5816 5097 5870 5123
rect 5900 5157 5970 5183
rect 5900 5123 5918 5157
rect 5952 5123 5970 5157
rect 5900 5097 5970 5123
rect 6000 5097 6070 5183
rect 6100 5097 6170 5183
rect 6200 5097 6270 5183
rect 6300 5097 6370 5183
rect 6400 5097 6454 5183
rect 6512 5172 6570 5183
rect 6512 5138 6524 5172
rect 6558 5138 6570 5172
rect 6512 5097 6570 5138
rect 6600 5157 6670 5183
rect 6600 5123 6618 5157
rect 6652 5123 6670 5157
rect 6600 5097 6670 5123
rect 6700 5142 6758 5183
rect 6700 5108 6712 5142
rect 6746 5108 6758 5142
rect 6700 5097 6758 5108
rect 6820 5157 6880 5183
rect 6820 5123 6828 5157
rect 6862 5123 6880 5157
rect 6820 5097 6880 5123
rect 6910 5157 6980 5183
rect 6910 5123 6928 5157
rect 6962 5123 6980 5157
rect 6910 5097 6980 5123
rect 7010 5157 7080 5183
rect 7010 5123 7028 5157
rect 7062 5123 7080 5157
rect 7010 5097 7080 5123
rect 7110 5157 7180 5183
rect 7110 5123 7128 5157
rect 7162 5123 7180 5157
rect 7110 5097 7180 5123
rect 7210 5157 7280 5183
rect 7210 5123 7228 5157
rect 7262 5123 7280 5157
rect 7210 5097 7280 5123
rect 7310 5157 7380 5183
rect 7310 5123 7328 5157
rect 7362 5123 7380 5157
rect 7310 5097 7380 5123
rect 7410 5157 7470 5183
rect 7410 5123 7428 5157
rect 7462 5123 7470 5157
rect 7410 5097 7470 5123
rect 5516 4787 5570 4813
rect 5516 4753 5524 4787
rect 5558 4753 5570 4787
rect 5516 4727 5570 4753
rect 5600 4787 5670 4813
rect 5600 4753 5618 4787
rect 5652 4753 5670 4787
rect 5600 4727 5670 4753
rect 5700 4727 5770 4813
rect 5800 4787 5870 4813
rect 5800 4753 5818 4787
rect 5852 4753 5870 4787
rect 5800 4727 5870 4753
rect 5900 4787 5954 4813
rect 5900 4753 5912 4787
rect 5946 4753 5954 4787
rect 5900 4727 5954 4753
rect 6016 4787 6070 4813
rect 6016 4753 6024 4787
rect 6058 4753 6070 4787
rect 6016 4727 6070 4753
rect 6100 4787 6154 4813
rect 6100 4753 6112 4787
rect 6146 4753 6154 4787
rect 6100 4727 6154 4753
rect 4616 4647 4670 4673
rect 4616 4613 4624 4647
rect 4658 4613 4670 4647
rect 4616 4587 4670 4613
rect 4700 4647 4770 4673
rect 4700 4613 4718 4647
rect 4752 4613 4770 4647
rect 4700 4587 4770 4613
rect 4800 4587 4870 4673
rect 4900 4587 4970 4673
rect 5000 4647 5070 4673
rect 5000 4613 5018 4647
rect 5052 4613 5070 4647
rect 5000 4587 5070 4613
rect 5100 4647 5170 4673
rect 5100 4613 5118 4647
rect 5152 4613 5170 4647
rect 5100 4587 5170 4613
rect 5200 4647 5270 4673
rect 5200 4613 5218 4647
rect 5252 4613 5270 4647
rect 5200 4587 5270 4613
rect 5300 4647 5370 4673
rect 5300 4613 5318 4647
rect 5352 4613 5370 4647
rect 5300 4587 5370 4613
rect 5400 4647 5470 4673
rect 5400 4613 5418 4647
rect 5452 4613 5470 4647
rect 5400 4587 5470 4613
rect 5500 4587 5570 4673
rect 5600 4587 5670 4673
rect 5700 4647 5770 4673
rect 5700 4613 5718 4647
rect 5752 4613 5770 4647
rect 5700 4587 5770 4613
rect 5800 4647 5870 4673
rect 5800 4613 5818 4647
rect 5852 4613 5870 4647
rect 5800 4587 5870 4613
rect 5900 4647 5970 4673
rect 5900 4613 5918 4647
rect 5952 4613 5970 4647
rect 5900 4587 5970 4613
rect 6000 4647 6054 4673
rect 6000 4613 6012 4647
rect 6046 4613 6054 4647
rect 6000 4587 6054 4613
rect 4416 4507 4470 4533
rect 4416 4473 4424 4507
rect 4458 4473 4470 4507
rect 4416 4447 4470 4473
rect 4500 4507 4570 4533
rect 4500 4473 4518 4507
rect 4552 4473 4570 4507
rect 4500 4447 4570 4473
rect 4600 4507 4670 4533
rect 4600 4473 4618 4507
rect 4652 4473 4670 4507
rect 4600 4447 4670 4473
rect 4700 4447 4770 4533
rect 4800 4447 4870 4533
rect 4900 4447 4970 4533
rect 5000 4507 5070 4533
rect 5000 4473 5018 4507
rect 5052 4473 5070 4507
rect 5000 4447 5070 4473
rect 5100 4507 5170 4533
rect 5100 4473 5118 4507
rect 5152 4473 5170 4507
rect 5100 4447 5170 4473
rect 5200 4507 5254 4533
rect 5200 4473 5212 4507
rect 5246 4473 5254 4507
rect 5200 4447 5254 4473
rect 3316 4367 3370 4393
rect 3316 4333 3324 4367
rect 3358 4333 3370 4367
rect 3316 4307 3370 4333
rect 3400 4367 3470 4393
rect 3400 4333 3418 4367
rect 3452 4333 3470 4367
rect 3400 4307 3470 4333
rect 3500 4367 3570 4393
rect 3500 4333 3518 4367
rect 3552 4333 3570 4367
rect 3500 4307 3570 4333
rect 3600 4367 3670 4393
rect 3600 4333 3618 4367
rect 3652 4333 3670 4367
rect 3600 4307 3670 4333
rect 3700 4307 3770 4393
rect 3800 4307 3870 4393
rect 3900 4307 3970 4393
rect 4000 4367 4070 4393
rect 4000 4333 4018 4367
rect 4052 4333 4070 4367
rect 4000 4307 4070 4333
rect 4100 4367 4170 4393
rect 4100 4333 4118 4367
rect 4152 4333 4170 4367
rect 4100 4307 4170 4333
rect 4200 4367 4270 4393
rect 4200 4333 4218 4367
rect 4252 4333 4270 4367
rect 4200 4307 4270 4333
rect 4300 4307 4370 4393
rect 4400 4307 4470 4393
rect 4500 4307 4570 4393
rect 4600 4307 4670 4393
rect 4700 4307 4770 4393
rect 4800 4367 4870 4393
rect 4800 4333 4818 4367
rect 4852 4333 4870 4367
rect 4800 4307 4870 4333
rect 4900 4367 4970 4393
rect 4900 4333 4918 4367
rect 4952 4333 4970 4367
rect 4900 4307 4970 4333
rect 5000 4367 5054 4393
rect 5000 4333 5012 4367
rect 5046 4333 5054 4367
rect 5000 4307 5054 4333
rect 1516 4227 1570 4253
rect 1516 4193 1524 4227
rect 1558 4193 1570 4227
rect 1516 4167 1570 4193
rect 1600 4227 1670 4253
rect 1600 4193 1618 4227
rect 1652 4193 1670 4227
rect 1600 4167 1670 4193
rect 1700 4167 1770 4253
rect 1800 4167 1870 4253
rect 1900 4227 1970 4253
rect 1900 4193 1918 4227
rect 1952 4193 1970 4227
rect 1900 4167 1970 4193
rect 2000 4227 2070 4253
rect 2000 4193 2018 4227
rect 2052 4193 2070 4227
rect 2000 4167 2070 4193
rect 2100 4227 2170 4253
rect 2100 4193 2118 4227
rect 2152 4193 2170 4227
rect 2100 4167 2170 4193
rect 2200 4227 2270 4253
rect 2200 4193 2218 4227
rect 2252 4193 2270 4227
rect 2200 4167 2270 4193
rect 2300 4167 2370 4253
rect 2400 4167 2470 4253
rect 2500 4227 2570 4253
rect 2500 4193 2518 4227
rect 2552 4193 2570 4227
rect 2500 4167 2570 4193
rect 2600 4227 2670 4253
rect 2600 4193 2618 4227
rect 2652 4193 2670 4227
rect 2600 4167 2670 4193
rect 2700 4167 2770 4253
rect 2800 4227 2870 4253
rect 2800 4193 2818 4227
rect 2852 4193 2870 4227
rect 2800 4167 2870 4193
rect 2900 4227 2970 4253
rect 2900 4193 2918 4227
rect 2952 4193 2970 4227
rect 2900 4167 2970 4193
rect 3000 4227 3070 4253
rect 3000 4193 3018 4227
rect 3052 4193 3070 4227
rect 3000 4167 3070 4193
rect 3100 4167 3170 4253
rect 3200 4227 3270 4253
rect 3200 4193 3218 4227
rect 3252 4193 3270 4227
rect 3200 4167 3270 4193
rect 3300 4227 3370 4253
rect 3300 4193 3318 4227
rect 3352 4193 3370 4227
rect 3300 4167 3370 4193
rect 3400 4227 3454 4253
rect 3400 4193 3412 4227
rect 3446 4193 3454 4227
rect 3400 4167 3454 4193
rect 716 4087 770 4113
rect 716 4053 724 4087
rect 758 4053 770 4087
rect 716 4027 770 4053
rect 800 4087 870 4113
rect 800 4053 818 4087
rect 852 4053 870 4087
rect 800 4027 870 4053
rect 900 4087 970 4113
rect 900 4053 918 4087
rect 952 4053 970 4087
rect 900 4027 970 4053
rect 1000 4027 1070 4113
rect 1100 4027 1170 4113
rect 1200 4027 1270 4113
rect 1300 4087 1370 4113
rect 1300 4053 1318 4087
rect 1352 4053 1370 4087
rect 1300 4027 1370 4053
rect 1400 4087 1470 4113
rect 1400 4053 1418 4087
rect 1452 4053 1470 4087
rect 1400 4027 1470 4053
rect 1500 4087 1554 4113
rect 1500 4053 1512 4087
rect 1546 4053 1554 4087
rect 1500 4027 1554 4053
rect 1616 4087 1670 4113
rect 1616 4053 1624 4087
rect 1658 4053 1670 4087
rect 1616 4027 1670 4053
rect 1700 4087 1754 4113
rect 1700 4053 1712 4087
rect 1746 4053 1754 4087
rect 1700 4027 1754 4053
rect 1816 4087 1870 4113
rect 1816 4053 1824 4087
rect 1858 4053 1870 4087
rect 1816 4027 1870 4053
rect 1900 4087 1954 4113
rect 1900 4053 1912 4087
rect 1946 4053 1954 4087
rect 1900 4027 1954 4053
rect 2016 4087 2070 4113
rect 2016 4053 2024 4087
rect 2058 4053 2070 4087
rect 2016 4027 2070 4053
rect 2100 4087 2170 4113
rect 2100 4053 2118 4087
rect 2152 4053 2170 4087
rect 2100 4027 2170 4053
rect 2200 4087 2254 4113
rect 2200 4053 2212 4087
rect 2246 4053 2254 4087
rect 2200 4027 2254 4053
rect 616 3947 670 3973
rect 616 3913 624 3947
rect 658 3913 670 3947
rect 616 3887 670 3913
rect 700 3947 770 3973
rect 700 3913 718 3947
rect 752 3913 770 3947
rect 700 3887 770 3913
rect 800 3887 870 3973
rect 900 3887 970 3973
rect 1000 3887 1070 3973
rect 1100 3947 1170 3973
rect 1100 3913 1118 3947
rect 1152 3913 1170 3947
rect 1100 3887 1170 3913
rect 1200 3947 1270 3973
rect 1200 3913 1218 3947
rect 1252 3913 1270 3947
rect 1200 3887 1270 3913
rect 1300 3887 1370 3973
rect 1400 3887 1470 3973
rect 1500 3947 1570 3973
rect 1500 3913 1518 3947
rect 1552 3913 1570 3947
rect 1500 3887 1570 3913
rect 1600 3947 1670 3973
rect 1600 3913 1618 3947
rect 1652 3913 1670 3947
rect 1600 3887 1670 3913
rect 1700 3887 1770 3973
rect 1800 3887 1870 3973
rect 1900 3947 1970 3973
rect 1900 3913 1918 3947
rect 1952 3913 1970 3947
rect 1900 3887 1970 3913
rect 2000 3947 2070 3973
rect 2000 3913 2018 3947
rect 2052 3913 2070 3947
rect 2000 3887 2070 3913
rect 2100 3947 2154 3973
rect 2100 3913 2112 3947
rect 2146 3913 2154 3947
rect 2100 3887 2154 3913
rect 16 3747 70 3833
rect 100 3807 170 3833
rect 100 3773 118 3807
rect 152 3773 170 3807
rect 100 3747 170 3773
rect 200 3807 270 3833
rect 200 3773 218 3807
rect 252 3773 270 3807
rect 200 3747 270 3773
rect 300 3807 370 3833
rect 300 3773 318 3807
rect 352 3773 370 3807
rect 300 3747 370 3773
rect 400 3807 470 3833
rect 400 3773 418 3807
rect 452 3773 470 3807
rect 400 3747 470 3773
rect 500 3807 570 3833
rect 500 3773 518 3807
rect 552 3773 570 3807
rect 500 3747 570 3773
rect 600 3747 670 3833
rect 700 3747 770 3833
rect 800 3807 870 3833
rect 800 3773 818 3807
rect 852 3773 870 3807
rect 800 3747 870 3773
rect 900 3807 970 3833
rect 900 3773 918 3807
rect 952 3773 970 3807
rect 900 3747 970 3773
rect 1000 3807 1070 3833
rect 1000 3773 1018 3807
rect 1052 3773 1070 3807
rect 1000 3747 1070 3773
rect 1100 3807 1170 3833
rect 1100 3773 1118 3807
rect 1152 3773 1170 3807
rect 1100 3747 1170 3773
rect 1200 3807 1254 3833
rect 1200 3773 1212 3807
rect 1246 3773 1254 3807
rect 1200 3747 1254 3773
rect 16 3517 70 3603
rect 100 3577 170 3603
rect 100 3543 118 3577
rect 152 3543 170 3577
rect 100 3517 170 3543
rect 200 3577 254 3603
rect 200 3543 212 3577
rect 246 3543 254 3577
rect 200 3517 254 3543
rect 1316 3807 1370 3833
rect 1316 3773 1324 3807
rect 1358 3773 1370 3807
rect 1316 3747 1370 3773
rect 1400 3807 1454 3833
rect 1400 3773 1412 3807
rect 1446 3773 1454 3807
rect 1400 3747 1454 3773
rect 316 3577 370 3603
rect 316 3543 324 3577
rect 358 3543 370 3577
rect 316 3517 370 3543
rect 400 3577 470 3603
rect 400 3543 418 3577
rect 452 3543 470 3577
rect 400 3517 470 3543
rect 500 3577 570 3603
rect 500 3543 518 3577
rect 552 3543 570 3577
rect 500 3517 570 3543
rect 600 3577 670 3603
rect 600 3543 618 3577
rect 652 3543 670 3577
rect 600 3517 670 3543
rect 700 3577 770 3603
rect 700 3543 718 3577
rect 752 3543 770 3577
rect 700 3517 770 3543
rect 800 3577 870 3603
rect 800 3543 818 3577
rect 852 3543 870 3577
rect 800 3517 870 3543
rect 900 3517 970 3603
rect 1000 3577 1070 3603
rect 1000 3543 1018 3577
rect 1052 3543 1070 3577
rect 1000 3517 1070 3543
rect 1100 3577 1170 3603
rect 1100 3543 1118 3577
rect 1152 3543 1170 3577
rect 1100 3517 1170 3543
rect 1200 3577 1270 3603
rect 1200 3543 1218 3577
rect 1252 3543 1270 3577
rect 1200 3517 1270 3543
rect 1300 3577 1354 3603
rect 1300 3543 1312 3577
rect 1346 3543 1354 3577
rect 1300 3517 1354 3543
rect 16 3377 70 3463
rect 100 3377 170 3463
rect 200 3377 270 3463
rect 300 3437 370 3463
rect 300 3403 318 3437
rect 352 3403 370 3437
rect 300 3377 370 3403
rect 400 3437 470 3463
rect 400 3403 418 3437
rect 452 3403 470 3437
rect 400 3377 470 3403
rect 500 3437 554 3463
rect 500 3403 512 3437
rect 546 3403 554 3437
rect 500 3377 554 3403
rect 616 3437 670 3463
rect 616 3403 624 3437
rect 658 3403 670 3437
rect 616 3377 670 3403
rect 700 3437 754 3463
rect 700 3403 712 3437
rect 746 3403 754 3437
rect 700 3377 754 3403
rect 1516 3807 1570 3833
rect 1516 3773 1524 3807
rect 1558 3773 1570 3807
rect 1516 3747 1570 3773
rect 1600 3807 1670 3833
rect 1600 3773 1618 3807
rect 1652 3773 1670 3807
rect 1600 3747 1670 3773
rect 1700 3807 1754 3833
rect 1700 3773 1712 3807
rect 1746 3773 1754 3807
rect 1700 3747 1754 3773
rect 1416 3577 1470 3603
rect 1416 3543 1424 3577
rect 1458 3543 1470 3577
rect 1416 3517 1470 3543
rect 1500 3577 1554 3603
rect 1500 3543 1512 3577
rect 1546 3543 1554 3577
rect 1500 3517 1554 3543
rect 2316 4087 2370 4113
rect 2316 4053 2324 4087
rect 2358 4053 2370 4087
rect 2316 4027 2370 4053
rect 2400 4087 2454 4113
rect 2400 4053 2412 4087
rect 2446 4053 2454 4087
rect 2400 4027 2454 4053
rect 2516 4087 2570 4113
rect 2516 4053 2524 4087
rect 2558 4053 2570 4087
rect 2516 4027 2570 4053
rect 2600 4087 2670 4113
rect 2600 4053 2618 4087
rect 2652 4053 2670 4087
rect 2600 4027 2670 4053
rect 2700 4027 2770 4113
rect 2800 4027 2870 4113
rect 2900 4027 2970 4113
rect 3000 4027 3070 4113
rect 3100 4087 3170 4113
rect 3100 4053 3118 4087
rect 3152 4053 3170 4087
rect 3100 4027 3170 4053
rect 3200 4087 3254 4113
rect 3200 4053 3212 4087
rect 3246 4053 3254 4087
rect 3200 4027 3254 4053
rect 2216 3947 2270 3973
rect 2216 3913 2224 3947
rect 2258 3913 2270 3947
rect 2216 3887 2270 3913
rect 2300 3947 2370 3973
rect 2300 3913 2318 3947
rect 2352 3913 2370 3947
rect 2300 3887 2370 3913
rect 2400 3947 2470 3973
rect 2400 3913 2418 3947
rect 2452 3913 2470 3947
rect 2400 3887 2470 3913
rect 2500 3947 2570 3973
rect 2500 3913 2518 3947
rect 2552 3913 2570 3947
rect 2500 3887 2570 3913
rect 2600 3887 2670 3973
rect 2700 3887 2770 3973
rect 2800 3947 2870 3973
rect 2800 3913 2818 3947
rect 2852 3913 2870 3947
rect 2800 3887 2870 3913
rect 2900 3947 2970 3973
rect 2900 3913 2918 3947
rect 2952 3913 2970 3947
rect 2900 3887 2970 3913
rect 3000 3887 3070 3973
rect 3100 3947 3170 3973
rect 3100 3913 3118 3947
rect 3152 3913 3170 3947
rect 3100 3887 3170 3913
rect 3200 3947 3254 3973
rect 3200 3913 3212 3947
rect 3246 3913 3254 3947
rect 3200 3887 3254 3913
rect 3316 4087 3370 4113
rect 3316 4053 3324 4087
rect 3358 4053 3370 4087
rect 3316 4027 3370 4053
rect 3400 4087 3454 4113
rect 3400 4053 3412 4087
rect 3446 4053 3454 4087
rect 3400 4027 3454 4053
rect 3516 4227 3570 4253
rect 3516 4193 3524 4227
rect 3558 4193 3570 4227
rect 3516 4167 3570 4193
rect 3600 4227 3654 4253
rect 3600 4193 3612 4227
rect 3646 4193 3654 4227
rect 3600 4167 3654 4193
rect 3716 4227 3770 4253
rect 3716 4193 3724 4227
rect 3758 4193 3770 4227
rect 3716 4167 3770 4193
rect 3800 4227 3870 4253
rect 3800 4193 3818 4227
rect 3852 4193 3870 4227
rect 3800 4167 3870 4193
rect 3900 4227 3970 4253
rect 3900 4193 3918 4227
rect 3952 4193 3970 4227
rect 3900 4167 3970 4193
rect 4000 4167 4070 4253
rect 4100 4167 4170 4253
rect 4200 4167 4270 4253
rect 4300 4227 4370 4253
rect 4300 4193 4318 4227
rect 4352 4193 4370 4227
rect 4300 4167 4370 4193
rect 4400 4227 4454 4253
rect 4400 4193 4412 4227
rect 4446 4193 4454 4227
rect 4400 4167 4454 4193
rect 4516 4227 4570 4253
rect 4516 4193 4524 4227
rect 4558 4193 4570 4227
rect 4516 4167 4570 4193
rect 4600 4227 4670 4253
rect 4600 4193 4618 4227
rect 4652 4193 4670 4227
rect 4600 4167 4670 4193
rect 4700 4167 4770 4253
rect 4800 4167 4870 4253
rect 4900 4227 4970 4253
rect 4900 4193 4918 4227
rect 4952 4193 4970 4227
rect 4900 4167 4970 4193
rect 5000 4227 5054 4253
rect 5000 4193 5012 4227
rect 5046 4193 5054 4227
rect 5000 4167 5054 4193
rect 3516 4087 3570 4113
rect 3516 4053 3524 4087
rect 3558 4053 3570 4087
rect 3516 4027 3570 4053
rect 3600 4087 3670 4113
rect 3600 4053 3618 4087
rect 3652 4053 3670 4087
rect 3600 4027 3670 4053
rect 3700 4027 3770 4113
rect 3800 4027 3870 4113
rect 3900 4087 3970 4113
rect 3900 4053 3918 4087
rect 3952 4053 3970 4087
rect 3900 4027 3970 4053
rect 4000 4087 4070 4113
rect 4000 4053 4018 4087
rect 4052 4053 4070 4087
rect 4000 4027 4070 4053
rect 4100 4027 4170 4113
rect 4200 4087 4270 4113
rect 4200 4053 4218 4087
rect 4252 4053 4270 4087
rect 4200 4027 4270 4053
rect 4300 4087 4370 4113
rect 4300 4053 4318 4087
rect 4352 4053 4370 4087
rect 4300 4027 4370 4053
rect 4400 4027 4470 4113
rect 4500 4087 4570 4113
rect 4500 4053 4518 4087
rect 4552 4053 4570 4087
rect 4500 4027 4570 4053
rect 4600 4087 4670 4113
rect 4600 4053 4618 4087
rect 4652 4053 4670 4087
rect 4600 4027 4670 4053
rect 4700 4087 4754 4113
rect 4700 4053 4712 4087
rect 4746 4053 4754 4087
rect 4700 4027 4754 4053
rect 3316 3947 3370 3973
rect 3316 3913 3324 3947
rect 3358 3913 3370 3947
rect 3316 3887 3370 3913
rect 3400 3947 3470 3973
rect 3400 3913 3418 3947
rect 3452 3913 3470 3947
rect 3400 3887 3470 3913
rect 3500 3947 3570 3973
rect 3500 3913 3518 3947
rect 3552 3913 3570 3947
rect 3500 3887 3570 3913
rect 3600 3887 3670 3973
rect 3700 3887 3770 3973
rect 3800 3887 3870 3973
rect 3900 3887 3970 3973
rect 4000 3947 4070 3973
rect 4000 3913 4018 3947
rect 4052 3913 4070 3947
rect 4000 3887 4070 3913
rect 4100 3947 4154 3973
rect 4100 3913 4112 3947
rect 4146 3913 4154 3947
rect 4100 3887 4154 3913
rect 1816 3807 1870 3833
rect 1816 3773 1824 3807
rect 1858 3773 1870 3807
rect 1816 3747 1870 3773
rect 1900 3807 1970 3833
rect 1900 3773 1918 3807
rect 1952 3773 1970 3807
rect 1900 3747 1970 3773
rect 2000 3747 2070 3833
rect 2100 3807 2170 3833
rect 2100 3773 2118 3807
rect 2152 3773 2170 3807
rect 2100 3747 2170 3773
rect 2200 3807 2270 3833
rect 2200 3773 2218 3807
rect 2252 3773 2270 3807
rect 2200 3747 2270 3773
rect 2300 3807 2370 3833
rect 2300 3773 2318 3807
rect 2352 3773 2370 3807
rect 2300 3747 2370 3773
rect 2400 3747 2470 3833
rect 2500 3747 2570 3833
rect 2600 3807 2670 3833
rect 2600 3773 2618 3807
rect 2652 3773 2670 3807
rect 2600 3747 2670 3773
rect 2700 3807 2770 3833
rect 2700 3773 2718 3807
rect 2752 3773 2770 3807
rect 2700 3747 2770 3773
rect 2800 3807 2870 3833
rect 2800 3773 2818 3807
rect 2852 3773 2870 3807
rect 2800 3747 2870 3773
rect 2900 3807 2970 3833
rect 2900 3773 2918 3807
rect 2952 3773 2970 3807
rect 2900 3747 2970 3773
rect 3000 3747 3070 3833
rect 3100 3747 3170 3833
rect 3200 3807 3270 3833
rect 3200 3773 3218 3807
rect 3252 3773 3270 3807
rect 3200 3747 3270 3773
rect 3300 3807 3370 3833
rect 3300 3773 3318 3807
rect 3352 3773 3370 3807
rect 3300 3747 3370 3773
rect 3400 3807 3454 3833
rect 3400 3773 3412 3807
rect 3446 3773 3454 3807
rect 3400 3747 3454 3773
rect 1616 3577 1670 3603
rect 1616 3543 1624 3577
rect 1658 3543 1670 3577
rect 1616 3517 1670 3543
rect 1700 3577 1770 3603
rect 1700 3543 1718 3577
rect 1752 3543 1770 3577
rect 1700 3517 1770 3543
rect 1800 3577 1870 3603
rect 1800 3543 1818 3577
rect 1852 3543 1870 3577
rect 1800 3517 1870 3543
rect 1900 3577 1970 3603
rect 1900 3543 1918 3577
rect 1952 3543 1970 3577
rect 1900 3517 1970 3543
rect 2000 3517 2070 3603
rect 2100 3577 2170 3603
rect 2100 3543 2118 3577
rect 2152 3543 2170 3577
rect 2100 3517 2170 3543
rect 2200 3577 2254 3603
rect 2200 3543 2212 3577
rect 2246 3543 2254 3577
rect 2200 3517 2254 3543
rect 816 3437 870 3463
rect 816 3403 824 3437
rect 858 3403 870 3437
rect 816 3377 870 3403
rect 900 3437 970 3463
rect 900 3403 918 3437
rect 952 3403 970 3437
rect 900 3377 970 3403
rect 1000 3437 1070 3463
rect 1000 3403 1018 3437
rect 1052 3403 1070 3437
rect 1000 3377 1070 3403
rect 1100 3377 1170 3463
rect 1200 3437 1270 3463
rect 1200 3403 1218 3437
rect 1252 3403 1270 3437
rect 1200 3377 1270 3403
rect 1300 3437 1370 3463
rect 1300 3403 1318 3437
rect 1352 3403 1370 3437
rect 1300 3377 1370 3403
rect 1400 3377 1470 3463
rect 1500 3437 1570 3463
rect 1500 3403 1518 3437
rect 1552 3403 1570 3437
rect 1500 3377 1570 3403
rect 1600 3437 1670 3463
rect 1600 3403 1618 3437
rect 1652 3403 1670 3437
rect 1600 3377 1670 3403
rect 1700 3437 1770 3463
rect 1700 3403 1718 3437
rect 1752 3403 1770 3437
rect 1700 3377 1770 3403
rect 1800 3437 1870 3463
rect 1800 3403 1818 3437
rect 1852 3403 1870 3437
rect 1800 3377 1870 3403
rect 1900 3437 1954 3463
rect 1900 3403 1912 3437
rect 1946 3403 1954 3437
rect 1900 3377 1954 3403
rect 16 3297 70 3323
rect 16 3263 24 3297
rect 58 3263 70 3297
rect 16 3237 70 3263
rect 100 3297 170 3323
rect 100 3263 118 3297
rect 152 3263 170 3297
rect 100 3237 170 3263
rect 200 3297 270 3323
rect 200 3263 218 3297
rect 252 3263 270 3297
rect 200 3237 270 3263
rect 300 3297 370 3323
rect 300 3263 318 3297
rect 352 3263 370 3297
rect 300 3237 370 3263
rect 400 3237 470 3323
rect 500 3237 570 3323
rect 600 3237 670 3323
rect 700 3297 770 3323
rect 700 3263 718 3297
rect 752 3263 770 3297
rect 700 3237 770 3263
rect 800 3297 870 3323
rect 800 3263 818 3297
rect 852 3263 870 3297
rect 800 3237 870 3263
rect 900 3297 970 3323
rect 900 3263 918 3297
rect 952 3263 970 3297
rect 900 3237 970 3263
rect 1000 3237 1070 3323
rect 1100 3297 1170 3323
rect 1100 3263 1118 3297
rect 1152 3263 1170 3297
rect 1100 3237 1170 3263
rect 1200 3297 1254 3323
rect 1200 3263 1212 3297
rect 1246 3263 1254 3297
rect 1200 3237 1254 3263
rect 16 3097 70 3183
rect 100 3097 170 3183
rect 200 3157 270 3183
rect 200 3123 218 3157
rect 252 3123 270 3157
rect 200 3097 270 3123
rect 300 3157 370 3183
rect 300 3123 318 3157
rect 352 3123 370 3157
rect 300 3097 370 3123
rect 400 3157 454 3183
rect 400 3123 412 3157
rect 446 3123 454 3157
rect 400 3097 454 3123
rect 516 3157 570 3183
rect 516 3123 524 3157
rect 558 3123 570 3157
rect 516 3097 570 3123
rect 600 3157 670 3183
rect 600 3123 618 3157
rect 652 3123 670 3157
rect 600 3097 670 3123
rect 700 3157 770 3183
rect 700 3123 718 3157
rect 752 3123 770 3157
rect 700 3097 770 3123
rect 800 3097 870 3183
rect 900 3157 970 3183
rect 900 3123 918 3157
rect 952 3123 970 3157
rect 900 3097 970 3123
rect 1000 3157 1070 3183
rect 1000 3123 1018 3157
rect 1052 3123 1070 3157
rect 1000 3097 1070 3123
rect 1100 3157 1154 3183
rect 1100 3123 1112 3157
rect 1146 3123 1154 3157
rect 1100 3097 1154 3123
rect 4216 3947 4270 3973
rect 4216 3913 4224 3947
rect 4258 3913 4270 3947
rect 4216 3887 4270 3913
rect 4300 3947 4370 3973
rect 4300 3913 4318 3947
rect 4352 3913 4370 3947
rect 4300 3887 4370 3913
rect 4400 3947 4470 3973
rect 4400 3913 4418 3947
rect 4452 3913 4470 3947
rect 4400 3887 4470 3913
rect 4500 3947 4554 3973
rect 4500 3913 4512 3947
rect 4546 3913 4554 3947
rect 4500 3887 4554 3913
rect 5316 4507 5370 4533
rect 5316 4473 5324 4507
rect 5358 4473 5370 4507
rect 5316 4447 5370 4473
rect 5400 4507 5470 4533
rect 5400 4473 5418 4507
rect 5452 4473 5470 4507
rect 5400 4447 5470 4473
rect 5500 4507 5570 4533
rect 5500 4473 5518 4507
rect 5552 4473 5570 4507
rect 5500 4447 5570 4473
rect 5600 4507 5670 4533
rect 5600 4473 5618 4507
rect 5652 4473 5670 4507
rect 5600 4447 5670 4473
rect 5700 4507 5754 4533
rect 5700 4473 5712 4507
rect 5746 4473 5754 4507
rect 5700 4447 5754 4473
rect 5116 4367 5170 4393
rect 5116 4333 5124 4367
rect 5158 4333 5170 4367
rect 5116 4307 5170 4333
rect 5200 4367 5270 4393
rect 5200 4333 5218 4367
rect 5252 4333 5270 4367
rect 5200 4307 5270 4333
rect 5300 4367 5370 4393
rect 5300 4333 5318 4367
rect 5352 4333 5370 4367
rect 5300 4307 5370 4333
rect 5400 4367 5454 4393
rect 5400 4333 5412 4367
rect 5446 4333 5454 4367
rect 5400 4307 5454 4333
rect 5116 4227 5170 4253
rect 5116 4193 5124 4227
rect 5158 4193 5170 4227
rect 5116 4167 5170 4193
rect 5200 4227 5270 4253
rect 5200 4193 5218 4227
rect 5252 4193 5270 4227
rect 5200 4167 5270 4193
rect 5300 4227 5370 4253
rect 5300 4193 5318 4227
rect 5352 4193 5370 4227
rect 5300 4167 5370 4193
rect 5400 4227 5454 4253
rect 5400 4193 5412 4227
rect 5446 4193 5454 4227
rect 5400 4167 5454 4193
rect 6216 4787 6270 4813
rect 6216 4753 6224 4787
rect 6258 4753 6270 4787
rect 6216 4727 6270 4753
rect 6300 4787 6370 4813
rect 6300 4753 6318 4787
rect 6352 4753 6370 4787
rect 6300 4727 6370 4753
rect 6400 4727 6454 4813
rect 6512 4802 6570 4813
rect 6512 4768 6524 4802
rect 6558 4768 6570 4802
rect 6512 4727 6570 4768
rect 6600 4787 6670 4813
rect 6600 4753 6618 4787
rect 6652 4753 6670 4787
rect 6600 4727 6670 4753
rect 6700 4772 6758 4813
rect 6700 4738 6712 4772
rect 6746 4738 6758 4772
rect 6700 4727 6758 4738
rect 6820 4787 6880 4813
rect 6820 4753 6828 4787
rect 6862 4753 6880 4787
rect 6820 4727 6880 4753
rect 6910 4787 6980 4813
rect 6910 4753 6928 4787
rect 6962 4753 6980 4787
rect 6910 4727 6980 4753
rect 7010 4787 7080 4813
rect 7010 4753 7028 4787
rect 7062 4753 7080 4787
rect 7010 4727 7080 4753
rect 7110 4787 7180 4813
rect 7110 4753 7128 4787
rect 7162 4753 7180 4787
rect 7110 4727 7180 4753
rect 7210 4787 7280 4813
rect 7210 4753 7228 4787
rect 7262 4753 7280 4787
rect 7210 4727 7280 4753
rect 7310 4787 7380 4813
rect 7310 4753 7328 4787
rect 7362 4753 7380 4787
rect 7310 4727 7380 4753
rect 7410 4787 7470 4813
rect 7410 4753 7428 4787
rect 7462 4753 7470 4787
rect 7410 4727 7470 4753
rect 6116 4647 6170 4673
rect 6116 4613 6124 4647
rect 6158 4613 6170 4647
rect 6116 4587 6170 4613
rect 6200 4647 6254 4673
rect 6200 4613 6212 4647
rect 6246 4613 6254 4647
rect 6200 4587 6254 4613
rect 5816 4507 5870 4533
rect 5816 4473 5824 4507
rect 5858 4473 5870 4507
rect 5816 4447 5870 4473
rect 5900 4507 5970 4533
rect 5900 4473 5918 4507
rect 5952 4473 5970 4507
rect 5900 4447 5970 4473
rect 6000 4447 6070 4533
rect 6100 4507 6170 4533
rect 6100 4473 6118 4507
rect 6152 4473 6170 4507
rect 6100 4447 6170 4473
rect 6200 4507 6254 4533
rect 6200 4473 6212 4507
rect 6246 4473 6254 4507
rect 6200 4447 6254 4473
rect 5516 4367 5570 4393
rect 5516 4333 5524 4367
rect 5558 4333 5570 4367
rect 5516 4307 5570 4333
rect 5600 4367 5670 4393
rect 5600 4333 5618 4367
rect 5652 4333 5670 4367
rect 5600 4307 5670 4333
rect 5700 4307 5770 4393
rect 5800 4307 5870 4393
rect 5900 4367 5970 4393
rect 5900 4333 5918 4367
rect 5952 4333 5970 4367
rect 5900 4307 5970 4333
rect 6000 4367 6054 4393
rect 6000 4333 6012 4367
rect 6046 4333 6054 4367
rect 6000 4307 6054 4333
rect 5516 4227 5570 4253
rect 5516 4193 5524 4227
rect 5558 4193 5570 4227
rect 5516 4167 5570 4193
rect 5600 4227 5670 4253
rect 5600 4193 5618 4227
rect 5652 4193 5670 4227
rect 5600 4167 5670 4193
rect 5700 4227 5770 4253
rect 5700 4193 5718 4227
rect 5752 4193 5770 4227
rect 5700 4167 5770 4193
rect 5800 4227 5854 4253
rect 5800 4193 5812 4227
rect 5846 4193 5854 4227
rect 5800 4167 5854 4193
rect 4816 4087 4870 4113
rect 4816 4053 4824 4087
rect 4858 4053 4870 4087
rect 4816 4027 4870 4053
rect 4900 4087 4970 4113
rect 4900 4053 4918 4087
rect 4952 4053 4970 4087
rect 4900 4027 4970 4053
rect 5000 4087 5070 4113
rect 5000 4053 5018 4087
rect 5052 4053 5070 4087
rect 5000 4027 5070 4053
rect 5100 4027 5170 4113
rect 5200 4087 5270 4113
rect 5200 4053 5218 4087
rect 5252 4053 5270 4087
rect 5200 4027 5270 4053
rect 5300 4087 5370 4113
rect 5300 4053 5318 4087
rect 5352 4053 5370 4087
rect 5300 4027 5370 4053
rect 5400 4027 5470 4113
rect 5500 4087 5570 4113
rect 5500 4053 5518 4087
rect 5552 4053 5570 4087
rect 5500 4027 5570 4053
rect 5600 4087 5654 4113
rect 5600 4053 5612 4087
rect 5646 4053 5654 4087
rect 5600 4027 5654 4053
rect 6116 4367 6170 4393
rect 6116 4333 6124 4367
rect 6158 4333 6170 4367
rect 6116 4307 6170 4333
rect 6200 4367 6254 4393
rect 6200 4333 6212 4367
rect 6246 4333 6254 4367
rect 6200 4307 6254 4333
rect 6316 4647 6370 4673
rect 6316 4613 6324 4647
rect 6358 4613 6370 4647
rect 6316 4587 6370 4613
rect 6400 4647 6454 4673
rect 6400 4613 6412 4647
rect 6446 4613 6454 4647
rect 6400 4587 6454 4613
rect 6512 4662 6570 4673
rect 6512 4628 6524 4662
rect 6558 4628 6570 4662
rect 6512 4587 6570 4628
rect 6600 4647 6670 4673
rect 6600 4613 6618 4647
rect 6652 4613 6670 4647
rect 6600 4587 6670 4613
rect 6700 4632 6758 4673
rect 6700 4598 6712 4632
rect 6746 4598 6758 4632
rect 6700 4587 6758 4598
rect 6820 4647 6880 4673
rect 6820 4613 6828 4647
rect 6862 4613 6880 4647
rect 6820 4587 6880 4613
rect 6910 4647 6980 4673
rect 6910 4613 6928 4647
rect 6962 4613 6980 4647
rect 6910 4587 6980 4613
rect 7010 4647 7080 4673
rect 7010 4613 7028 4647
rect 7062 4613 7080 4647
rect 7010 4587 7080 4613
rect 7110 4647 7180 4673
rect 7110 4613 7128 4647
rect 7162 4613 7180 4647
rect 7110 4587 7180 4613
rect 7210 4647 7280 4673
rect 7210 4613 7228 4647
rect 7262 4613 7280 4647
rect 7210 4587 7280 4613
rect 7310 4647 7380 4673
rect 7310 4613 7328 4647
rect 7362 4613 7380 4647
rect 7310 4587 7380 4613
rect 7410 4647 7470 4673
rect 7410 4613 7428 4647
rect 7462 4613 7470 4647
rect 7410 4587 7470 4613
rect 6316 4507 6370 4533
rect 6316 4473 6324 4507
rect 6358 4473 6370 4507
rect 6316 4447 6370 4473
rect 6400 4507 6454 4533
rect 6400 4473 6412 4507
rect 6446 4473 6454 4507
rect 6400 4447 6454 4473
rect 6512 4522 6570 4533
rect 6512 4488 6524 4522
rect 6558 4488 6570 4522
rect 6512 4447 6570 4488
rect 6600 4507 6670 4533
rect 6600 4473 6618 4507
rect 6652 4473 6670 4507
rect 6600 4447 6670 4473
rect 6700 4492 6758 4533
rect 6700 4458 6712 4492
rect 6746 4458 6758 4492
rect 6700 4447 6758 4458
rect 6820 4507 6880 4533
rect 6820 4473 6828 4507
rect 6862 4473 6880 4507
rect 6820 4447 6880 4473
rect 6910 4507 6980 4533
rect 6910 4473 6928 4507
rect 6962 4473 6980 4507
rect 6910 4447 6980 4473
rect 7010 4507 7080 4533
rect 7010 4473 7028 4507
rect 7062 4473 7080 4507
rect 7010 4447 7080 4473
rect 7110 4507 7180 4533
rect 7110 4473 7128 4507
rect 7162 4473 7180 4507
rect 7110 4447 7180 4473
rect 7210 4507 7280 4533
rect 7210 4473 7228 4507
rect 7262 4473 7280 4507
rect 7210 4447 7280 4473
rect 7310 4507 7380 4533
rect 7310 4473 7328 4507
rect 7362 4473 7380 4507
rect 7310 4447 7380 4473
rect 7410 4507 7470 4533
rect 7410 4473 7428 4507
rect 7462 4473 7470 4507
rect 7410 4447 7470 4473
rect 6316 4367 6370 4393
rect 6316 4333 6324 4367
rect 6358 4333 6370 4367
rect 6316 4307 6370 4333
rect 6400 4367 6454 4393
rect 6400 4333 6412 4367
rect 6446 4333 6454 4367
rect 6400 4307 6454 4333
rect 6512 4382 6570 4393
rect 6512 4348 6524 4382
rect 6558 4348 6570 4382
rect 6512 4307 6570 4348
rect 6600 4367 6670 4393
rect 6600 4333 6618 4367
rect 6652 4333 6670 4367
rect 6600 4307 6670 4333
rect 6700 4352 6758 4393
rect 6700 4318 6712 4352
rect 6746 4318 6758 4352
rect 6700 4307 6758 4318
rect 6820 4367 6880 4393
rect 6820 4333 6828 4367
rect 6862 4333 6880 4367
rect 6820 4307 6880 4333
rect 6910 4367 6980 4393
rect 6910 4333 6928 4367
rect 6962 4333 6980 4367
rect 6910 4307 6980 4333
rect 7010 4367 7080 4393
rect 7010 4333 7028 4367
rect 7062 4333 7080 4367
rect 7010 4307 7080 4333
rect 7110 4367 7180 4393
rect 7110 4333 7128 4367
rect 7162 4333 7180 4367
rect 7110 4307 7180 4333
rect 7210 4367 7280 4393
rect 7210 4333 7228 4367
rect 7262 4333 7280 4367
rect 7210 4307 7280 4333
rect 7310 4367 7380 4393
rect 7310 4333 7328 4367
rect 7362 4333 7380 4367
rect 7310 4307 7380 4333
rect 7410 4367 7470 4393
rect 7410 4333 7428 4367
rect 7462 4333 7470 4367
rect 7410 4307 7470 4333
rect 5916 4227 5970 4253
rect 5916 4193 5924 4227
rect 5958 4193 5970 4227
rect 5916 4167 5970 4193
rect 6000 4227 6070 4253
rect 6000 4193 6018 4227
rect 6052 4193 6070 4227
rect 6000 4167 6070 4193
rect 6100 4227 6170 4253
rect 6100 4193 6118 4227
rect 6152 4193 6170 4227
rect 6100 4167 6170 4193
rect 6200 4167 6270 4253
rect 6300 4227 6370 4253
rect 6300 4193 6318 4227
rect 6352 4193 6370 4227
rect 6300 4167 6370 4193
rect 6400 4227 6454 4253
rect 6400 4193 6412 4227
rect 6446 4193 6454 4227
rect 6400 4167 6454 4193
rect 6512 4242 6570 4253
rect 6512 4208 6524 4242
rect 6558 4208 6570 4242
rect 6512 4167 6570 4208
rect 6600 4227 6670 4253
rect 6600 4193 6618 4227
rect 6652 4193 6670 4227
rect 6600 4167 6670 4193
rect 6700 4212 6758 4253
rect 6700 4178 6712 4212
rect 6746 4178 6758 4212
rect 6700 4167 6758 4178
rect 6820 4227 6880 4253
rect 6820 4193 6828 4227
rect 6862 4193 6880 4227
rect 6820 4167 6880 4193
rect 6910 4227 6980 4253
rect 6910 4193 6928 4227
rect 6962 4193 6980 4227
rect 6910 4167 6980 4193
rect 7010 4227 7080 4253
rect 7010 4193 7028 4227
rect 7062 4193 7080 4227
rect 7010 4167 7080 4193
rect 7110 4227 7180 4253
rect 7110 4193 7128 4227
rect 7162 4193 7180 4227
rect 7110 4167 7180 4193
rect 7210 4227 7280 4253
rect 7210 4193 7228 4227
rect 7262 4193 7280 4227
rect 7210 4167 7280 4193
rect 7310 4227 7380 4253
rect 7310 4193 7328 4227
rect 7362 4193 7380 4227
rect 7310 4167 7380 4193
rect 7410 4227 7470 4253
rect 7410 4193 7428 4227
rect 7462 4193 7470 4227
rect 7410 4167 7470 4193
rect 5716 4087 5770 4113
rect 5716 4053 5724 4087
rect 5758 4053 5770 4087
rect 5716 4027 5770 4053
rect 5800 4087 5870 4113
rect 5800 4053 5818 4087
rect 5852 4053 5870 4087
rect 5800 4027 5870 4053
rect 5900 4027 5970 4113
rect 6000 4027 6070 4113
rect 6100 4087 6170 4113
rect 6100 4053 6118 4087
rect 6152 4053 6170 4087
rect 6100 4027 6170 4053
rect 6200 4087 6270 4113
rect 6200 4053 6218 4087
rect 6252 4053 6270 4087
rect 6200 4027 6270 4053
rect 6300 4087 6370 4113
rect 6300 4053 6318 4087
rect 6352 4053 6370 4087
rect 6300 4027 6370 4053
rect 6400 4087 6454 4113
rect 6400 4053 6412 4087
rect 6446 4053 6454 4087
rect 6400 4027 6454 4053
rect 6512 4102 6570 4113
rect 6512 4068 6524 4102
rect 6558 4068 6570 4102
rect 6512 4027 6570 4068
rect 6600 4087 6670 4113
rect 6600 4053 6618 4087
rect 6652 4053 6670 4087
rect 6600 4027 6670 4053
rect 6700 4072 6758 4113
rect 6700 4038 6712 4072
rect 6746 4038 6758 4072
rect 6700 4027 6758 4038
rect 6820 4087 6880 4113
rect 6820 4053 6828 4087
rect 6862 4053 6880 4087
rect 6820 4027 6880 4053
rect 6910 4087 6980 4113
rect 6910 4053 6928 4087
rect 6962 4053 6980 4087
rect 6910 4027 6980 4053
rect 7010 4087 7080 4113
rect 7010 4053 7028 4087
rect 7062 4053 7080 4087
rect 7010 4027 7080 4053
rect 7110 4087 7180 4113
rect 7110 4053 7128 4087
rect 7162 4053 7180 4087
rect 7110 4027 7180 4053
rect 7210 4087 7280 4113
rect 7210 4053 7228 4087
rect 7262 4053 7280 4087
rect 7210 4027 7280 4053
rect 7310 4087 7380 4113
rect 7310 4053 7328 4087
rect 7362 4053 7380 4087
rect 7310 4027 7380 4053
rect 7410 4087 7470 4113
rect 7410 4053 7428 4087
rect 7462 4053 7470 4087
rect 7410 4027 7470 4053
rect 4616 3947 4670 3973
rect 4616 3913 4624 3947
rect 4658 3913 4670 3947
rect 4616 3887 4670 3913
rect 4700 3947 4770 3973
rect 4700 3913 4718 3947
rect 4752 3913 4770 3947
rect 4700 3887 4770 3913
rect 4800 3887 4870 3973
rect 4900 3887 4970 3973
rect 5000 3947 5070 3973
rect 5000 3913 5018 3947
rect 5052 3913 5070 3947
rect 5000 3887 5070 3913
rect 5100 3947 5170 3973
rect 5100 3913 5118 3947
rect 5152 3913 5170 3947
rect 5100 3887 5170 3913
rect 5200 3887 5270 3973
rect 5300 3887 5370 3973
rect 5400 3947 5470 3973
rect 5400 3913 5418 3947
rect 5452 3913 5470 3947
rect 5400 3887 5470 3913
rect 5500 3947 5570 3973
rect 5500 3913 5518 3947
rect 5552 3913 5570 3947
rect 5500 3887 5570 3913
rect 5600 3887 5670 3973
rect 5700 3947 5770 3973
rect 5700 3913 5718 3947
rect 5752 3913 5770 3947
rect 5700 3887 5770 3913
rect 5800 3947 5870 3973
rect 5800 3913 5818 3947
rect 5852 3913 5870 3947
rect 5800 3887 5870 3913
rect 5900 3947 5970 3973
rect 5900 3913 5918 3947
rect 5952 3913 5970 3947
rect 5900 3887 5970 3913
rect 6000 3947 6054 3973
rect 6000 3913 6012 3947
rect 6046 3913 6054 3947
rect 6000 3887 6054 3913
rect 3516 3807 3570 3833
rect 3516 3773 3524 3807
rect 3558 3773 3570 3807
rect 3516 3747 3570 3773
rect 3600 3807 3670 3833
rect 3600 3773 3618 3807
rect 3652 3773 3670 3807
rect 3600 3747 3670 3773
rect 3700 3807 3770 3833
rect 3700 3773 3718 3807
rect 3752 3773 3770 3807
rect 3700 3747 3770 3773
rect 3800 3747 3870 3833
rect 3900 3747 3970 3833
rect 4000 3747 4070 3833
rect 4100 3747 4170 3833
rect 4200 3747 4270 3833
rect 4300 3747 4370 3833
rect 4400 3747 4470 3833
rect 4500 3747 4570 3833
rect 4600 3807 4670 3833
rect 4600 3773 4618 3807
rect 4652 3773 4670 3807
rect 4600 3747 4670 3773
rect 4700 3807 4754 3833
rect 4700 3773 4712 3807
rect 4746 3773 4754 3807
rect 4700 3747 4754 3773
rect 2316 3577 2370 3603
rect 2316 3543 2324 3577
rect 2358 3543 2370 3577
rect 2316 3517 2370 3543
rect 2400 3577 2470 3603
rect 2400 3543 2418 3577
rect 2452 3543 2470 3577
rect 2400 3517 2470 3543
rect 2500 3577 2570 3603
rect 2500 3543 2518 3577
rect 2552 3543 2570 3577
rect 2500 3517 2570 3543
rect 2600 3577 2670 3603
rect 2600 3543 2618 3577
rect 2652 3543 2670 3577
rect 2600 3517 2670 3543
rect 2700 3577 2770 3603
rect 2700 3543 2718 3577
rect 2752 3543 2770 3577
rect 2700 3517 2770 3543
rect 2800 3517 2870 3603
rect 2900 3517 2970 3603
rect 3000 3577 3070 3603
rect 3000 3543 3018 3577
rect 3052 3543 3070 3577
rect 3000 3517 3070 3543
rect 3100 3577 3170 3603
rect 3100 3543 3118 3577
rect 3152 3543 3170 3577
rect 3100 3517 3170 3543
rect 3200 3517 3270 3603
rect 3300 3517 3370 3603
rect 3400 3577 3470 3603
rect 3400 3543 3418 3577
rect 3452 3543 3470 3577
rect 3400 3517 3470 3543
rect 3500 3577 3554 3603
rect 3500 3543 3512 3577
rect 3546 3543 3554 3577
rect 3500 3517 3554 3543
rect 2016 3437 2070 3463
rect 2016 3403 2024 3437
rect 2058 3403 2070 3437
rect 2016 3377 2070 3403
rect 2100 3437 2170 3463
rect 2100 3403 2118 3437
rect 2152 3403 2170 3437
rect 2100 3377 2170 3403
rect 2200 3437 2270 3463
rect 2200 3403 2218 3437
rect 2252 3403 2270 3437
rect 2200 3377 2270 3403
rect 2300 3437 2370 3463
rect 2300 3403 2318 3437
rect 2352 3403 2370 3437
rect 2300 3377 2370 3403
rect 2400 3437 2470 3463
rect 2400 3403 2418 3437
rect 2452 3403 2470 3437
rect 2400 3377 2470 3403
rect 2500 3437 2570 3463
rect 2500 3403 2518 3437
rect 2552 3403 2570 3437
rect 2500 3377 2570 3403
rect 2600 3437 2670 3463
rect 2600 3403 2618 3437
rect 2652 3403 2670 3437
rect 2600 3377 2670 3403
rect 2700 3437 2770 3463
rect 2700 3403 2718 3437
rect 2752 3403 2770 3437
rect 2700 3377 2770 3403
rect 2800 3437 2854 3463
rect 2800 3403 2812 3437
rect 2846 3403 2854 3437
rect 2800 3377 2854 3403
rect 1316 3297 1370 3323
rect 1316 3263 1324 3297
rect 1358 3263 1370 3297
rect 1316 3237 1370 3263
rect 1400 3297 1470 3323
rect 1400 3263 1418 3297
rect 1452 3263 1470 3297
rect 1400 3237 1470 3263
rect 1500 3297 1570 3323
rect 1500 3263 1518 3297
rect 1552 3263 1570 3297
rect 1500 3237 1570 3263
rect 1600 3237 1670 3323
rect 1700 3297 1770 3323
rect 1700 3263 1718 3297
rect 1752 3263 1770 3297
rect 1700 3237 1770 3263
rect 1800 3297 1870 3323
rect 1800 3263 1818 3297
rect 1852 3263 1870 3297
rect 1800 3237 1870 3263
rect 1900 3297 1970 3323
rect 1900 3263 1918 3297
rect 1952 3263 1970 3297
rect 1900 3237 1970 3263
rect 2000 3297 2070 3323
rect 2000 3263 2018 3297
rect 2052 3263 2070 3297
rect 2000 3237 2070 3263
rect 2100 3297 2170 3323
rect 2100 3263 2118 3297
rect 2152 3263 2170 3297
rect 2100 3237 2170 3263
rect 2200 3297 2270 3323
rect 2200 3263 2218 3297
rect 2252 3263 2270 3297
rect 2200 3237 2270 3263
rect 2300 3297 2370 3323
rect 2300 3263 2318 3297
rect 2352 3263 2370 3297
rect 2300 3237 2370 3263
rect 2400 3297 2470 3323
rect 2400 3263 2418 3297
rect 2452 3263 2470 3297
rect 2400 3237 2470 3263
rect 2500 3297 2570 3323
rect 2500 3263 2518 3297
rect 2552 3263 2570 3297
rect 2500 3237 2570 3263
rect 2600 3297 2670 3323
rect 2600 3263 2618 3297
rect 2652 3263 2670 3297
rect 2600 3237 2670 3263
rect 2700 3297 2754 3323
rect 2700 3263 2712 3297
rect 2746 3263 2754 3297
rect 2700 3237 2754 3263
rect 1216 3157 1270 3183
rect 1216 3123 1224 3157
rect 1258 3123 1270 3157
rect 1216 3097 1270 3123
rect 1300 3157 1370 3183
rect 1300 3123 1318 3157
rect 1352 3123 1370 3157
rect 1300 3097 1370 3123
rect 1400 3097 1470 3183
rect 1500 3097 1570 3183
rect 1600 3097 1670 3183
rect 1700 3157 1770 3183
rect 1700 3123 1718 3157
rect 1752 3123 1770 3157
rect 1700 3097 1770 3123
rect 1800 3157 1870 3183
rect 1800 3123 1818 3157
rect 1852 3123 1870 3157
rect 1800 3097 1870 3123
rect 1900 3157 1970 3183
rect 1900 3123 1918 3157
rect 1952 3123 1970 3157
rect 1900 3097 1970 3123
rect 2000 3157 2070 3183
rect 2000 3123 2018 3157
rect 2052 3123 2070 3157
rect 2000 3097 2070 3123
rect 2100 3157 2170 3183
rect 2100 3123 2118 3157
rect 2152 3123 2170 3157
rect 2100 3097 2170 3123
rect 2200 3097 2270 3183
rect 2300 3157 2370 3183
rect 2300 3123 2318 3157
rect 2352 3123 2370 3157
rect 2300 3097 2370 3123
rect 2400 3157 2454 3183
rect 2400 3123 2412 3157
rect 2446 3123 2454 3157
rect 2400 3097 2454 3123
rect 3616 3577 3670 3603
rect 3616 3543 3624 3577
rect 3658 3543 3670 3577
rect 3616 3517 3670 3543
rect 3700 3577 3754 3603
rect 3700 3543 3712 3577
rect 3746 3543 3754 3577
rect 3700 3517 3754 3543
rect 3816 3577 3870 3603
rect 3816 3543 3824 3577
rect 3858 3543 3870 3577
rect 3816 3517 3870 3543
rect 3900 3577 3970 3603
rect 3900 3543 3918 3577
rect 3952 3543 3970 3577
rect 3900 3517 3970 3543
rect 4000 3577 4070 3603
rect 4000 3543 4018 3577
rect 4052 3543 4070 3577
rect 4000 3517 4070 3543
rect 4100 3577 4170 3603
rect 4100 3543 4118 3577
rect 4152 3543 4170 3577
rect 4100 3517 4170 3543
rect 4200 3577 4254 3603
rect 4200 3543 4212 3577
rect 4246 3543 4254 3577
rect 4200 3517 4254 3543
rect 4816 3807 4870 3833
rect 4816 3773 4824 3807
rect 4858 3773 4870 3807
rect 4816 3747 4870 3773
rect 4900 3807 4970 3833
rect 4900 3773 4918 3807
rect 4952 3773 4970 3807
rect 4900 3747 4970 3773
rect 5000 3807 5070 3833
rect 5000 3773 5018 3807
rect 5052 3773 5070 3807
rect 5000 3747 5070 3773
rect 5100 3747 5170 3833
rect 5200 3747 5270 3833
rect 5300 3747 5370 3833
rect 5400 3807 5470 3833
rect 5400 3773 5418 3807
rect 5452 3773 5470 3807
rect 5400 3747 5470 3773
rect 5500 3807 5570 3833
rect 5500 3773 5518 3807
rect 5552 3773 5570 3807
rect 5500 3747 5570 3773
rect 5600 3807 5654 3833
rect 5600 3773 5612 3807
rect 5646 3773 5654 3807
rect 5600 3747 5654 3773
rect 4316 3577 4370 3603
rect 4316 3543 4324 3577
rect 4358 3543 4370 3577
rect 4316 3517 4370 3543
rect 4400 3577 4470 3603
rect 4400 3543 4418 3577
rect 4452 3543 4470 3577
rect 4400 3517 4470 3543
rect 4500 3517 4570 3603
rect 4600 3577 4670 3603
rect 4600 3543 4618 3577
rect 4652 3543 4670 3577
rect 4600 3517 4670 3543
rect 4700 3577 4754 3603
rect 4700 3543 4712 3577
rect 4746 3543 4754 3577
rect 4700 3517 4754 3543
rect 4816 3577 4870 3603
rect 4816 3543 4824 3577
rect 4858 3543 4870 3577
rect 4816 3517 4870 3543
rect 4900 3577 4970 3603
rect 4900 3543 4918 3577
rect 4952 3543 4970 3577
rect 4900 3517 4970 3543
rect 5000 3517 5070 3603
rect 5100 3577 5170 3603
rect 5100 3543 5118 3577
rect 5152 3543 5170 3577
rect 5100 3517 5170 3543
rect 5200 3577 5254 3603
rect 5200 3543 5212 3577
rect 5246 3543 5254 3577
rect 5200 3517 5254 3543
rect 6116 3947 6170 3973
rect 6116 3913 6124 3947
rect 6158 3913 6170 3947
rect 6116 3887 6170 3913
rect 6200 3947 6270 3973
rect 6200 3913 6218 3947
rect 6252 3913 6270 3947
rect 6200 3887 6270 3913
rect 6300 3947 6370 3973
rect 6300 3913 6318 3947
rect 6352 3913 6370 3947
rect 6300 3887 6370 3913
rect 6400 3887 6454 3973
rect 6512 3962 6570 3973
rect 6512 3928 6524 3962
rect 6558 3928 6570 3962
rect 6512 3887 6570 3928
rect 6600 3947 6670 3973
rect 6600 3913 6618 3947
rect 6652 3913 6670 3947
rect 6600 3887 6670 3913
rect 6700 3932 6758 3973
rect 6700 3898 6712 3932
rect 6746 3898 6758 3932
rect 6700 3887 6758 3898
rect 6820 3947 6880 3973
rect 6820 3913 6828 3947
rect 6862 3913 6880 3947
rect 6820 3887 6880 3913
rect 6910 3947 6980 3973
rect 6910 3913 6928 3947
rect 6962 3913 6980 3947
rect 6910 3887 6980 3913
rect 7010 3947 7080 3973
rect 7010 3913 7028 3947
rect 7062 3913 7080 3947
rect 7010 3887 7080 3913
rect 7110 3947 7180 3973
rect 7110 3913 7128 3947
rect 7162 3913 7180 3947
rect 7110 3887 7180 3913
rect 7210 3947 7280 3973
rect 7210 3913 7228 3947
rect 7262 3913 7280 3947
rect 7210 3887 7280 3913
rect 7310 3947 7380 3973
rect 7310 3913 7328 3947
rect 7362 3913 7380 3947
rect 7310 3887 7380 3913
rect 7410 3947 7470 3973
rect 7410 3913 7428 3947
rect 7462 3913 7470 3947
rect 7410 3887 7470 3913
rect 5716 3807 5770 3833
rect 5716 3773 5724 3807
rect 5758 3773 5770 3807
rect 5716 3747 5770 3773
rect 5800 3807 5870 3833
rect 5800 3773 5818 3807
rect 5852 3773 5870 3807
rect 5800 3747 5870 3773
rect 5900 3747 5970 3833
rect 6000 3807 6070 3833
rect 6000 3773 6018 3807
rect 6052 3773 6070 3807
rect 6000 3747 6070 3773
rect 6100 3807 6170 3833
rect 6100 3773 6118 3807
rect 6152 3773 6170 3807
rect 6100 3747 6170 3773
rect 6200 3807 6270 3833
rect 6200 3773 6218 3807
rect 6252 3773 6270 3807
rect 6200 3747 6270 3773
rect 6300 3807 6370 3833
rect 6300 3773 6318 3807
rect 6352 3773 6370 3807
rect 6300 3747 6370 3773
rect 6400 3747 6454 3833
rect 6512 3822 6570 3833
rect 6512 3788 6524 3822
rect 6558 3788 6570 3822
rect 6512 3747 6570 3788
rect 6600 3807 6670 3833
rect 6600 3773 6618 3807
rect 6652 3773 6670 3807
rect 6600 3747 6670 3773
rect 6700 3792 6758 3833
rect 6700 3758 6712 3792
rect 6746 3758 6758 3792
rect 6700 3747 6758 3758
rect 6820 3807 6880 3833
rect 6820 3773 6828 3807
rect 6862 3773 6880 3807
rect 6820 3747 6880 3773
rect 6910 3807 6980 3833
rect 6910 3773 6928 3807
rect 6962 3773 6980 3807
rect 6910 3747 6980 3773
rect 7010 3807 7080 3833
rect 7010 3773 7028 3807
rect 7062 3773 7080 3807
rect 7010 3747 7080 3773
rect 7110 3807 7180 3833
rect 7110 3773 7128 3807
rect 7162 3773 7180 3807
rect 7110 3747 7180 3773
rect 7210 3807 7280 3833
rect 7210 3773 7228 3807
rect 7262 3773 7280 3807
rect 7210 3747 7280 3773
rect 7310 3807 7380 3833
rect 7310 3773 7328 3807
rect 7362 3773 7380 3807
rect 7310 3747 7380 3773
rect 7410 3807 7470 3833
rect 7410 3773 7428 3807
rect 7462 3773 7470 3807
rect 7410 3747 7470 3773
rect 5316 3577 5370 3603
rect 5316 3543 5324 3577
rect 5358 3543 5370 3577
rect 5316 3517 5370 3543
rect 5400 3577 5470 3603
rect 5400 3543 5418 3577
rect 5452 3543 5470 3577
rect 5400 3517 5470 3543
rect 5500 3577 5570 3603
rect 5500 3543 5518 3577
rect 5552 3543 5570 3577
rect 5500 3517 5570 3543
rect 5600 3577 5670 3603
rect 5600 3543 5618 3577
rect 5652 3543 5670 3577
rect 5600 3517 5670 3543
rect 5700 3577 5770 3603
rect 5700 3543 5718 3577
rect 5752 3543 5770 3577
rect 5700 3517 5770 3543
rect 5800 3577 5870 3603
rect 5800 3543 5818 3577
rect 5852 3543 5870 3577
rect 5800 3517 5870 3543
rect 5900 3577 5970 3603
rect 5900 3543 5918 3577
rect 5952 3543 5970 3577
rect 5900 3517 5970 3543
rect 6000 3517 6070 3603
rect 6100 3517 6170 3603
rect 6200 3577 6270 3603
rect 6200 3543 6218 3577
rect 6252 3543 6270 3577
rect 6200 3517 6270 3543
rect 6300 3577 6370 3603
rect 6300 3543 6318 3577
rect 6352 3543 6370 3577
rect 6300 3517 6370 3543
rect 6400 3577 6454 3603
rect 6400 3543 6412 3577
rect 6446 3543 6454 3577
rect 6400 3517 6454 3543
rect 6512 3592 6570 3603
rect 6512 3558 6524 3592
rect 6558 3558 6570 3592
rect 6512 3517 6570 3558
rect 6600 3577 6670 3603
rect 6600 3543 6618 3577
rect 6652 3543 6670 3577
rect 6600 3517 6670 3543
rect 6700 3562 6758 3603
rect 6700 3528 6712 3562
rect 6746 3528 6758 3562
rect 6700 3517 6758 3528
rect 6820 3577 6880 3603
rect 6820 3543 6828 3577
rect 6862 3543 6880 3577
rect 6820 3517 6880 3543
rect 6910 3577 6980 3603
rect 6910 3543 6928 3577
rect 6962 3543 6980 3577
rect 6910 3517 6980 3543
rect 7010 3577 7080 3603
rect 7010 3543 7028 3577
rect 7062 3543 7080 3577
rect 7010 3517 7080 3543
rect 7110 3577 7180 3603
rect 7110 3543 7128 3577
rect 7162 3543 7180 3577
rect 7110 3517 7180 3543
rect 7210 3577 7280 3603
rect 7210 3543 7228 3577
rect 7262 3543 7280 3577
rect 7210 3517 7280 3543
rect 7310 3577 7380 3603
rect 7310 3543 7328 3577
rect 7362 3543 7380 3577
rect 7310 3517 7380 3543
rect 7410 3577 7470 3603
rect 7410 3543 7428 3577
rect 7462 3543 7470 3577
rect 7410 3517 7470 3543
rect 2916 3437 2970 3463
rect 2916 3403 2924 3437
rect 2958 3403 2970 3437
rect 2916 3377 2970 3403
rect 3000 3437 3070 3463
rect 3000 3403 3018 3437
rect 3052 3403 3070 3437
rect 3000 3377 3070 3403
rect 3100 3437 3170 3463
rect 3100 3403 3118 3437
rect 3152 3403 3170 3437
rect 3100 3377 3170 3403
rect 3200 3437 3270 3463
rect 3200 3403 3218 3437
rect 3252 3403 3270 3437
rect 3200 3377 3270 3403
rect 3300 3437 3370 3463
rect 3300 3403 3318 3437
rect 3352 3403 3370 3437
rect 3300 3377 3370 3403
rect 3400 3437 3470 3463
rect 3400 3403 3418 3437
rect 3452 3403 3470 3437
rect 3400 3377 3470 3403
rect 3500 3437 3570 3463
rect 3500 3403 3518 3437
rect 3552 3403 3570 3437
rect 3500 3377 3570 3403
rect 3600 3377 3670 3463
rect 3700 3377 3770 3463
rect 3800 3377 3870 3463
rect 3900 3437 3970 3463
rect 3900 3403 3918 3437
rect 3952 3403 3970 3437
rect 3900 3377 3970 3403
rect 4000 3437 4070 3463
rect 4000 3403 4018 3437
rect 4052 3403 4070 3437
rect 4000 3377 4070 3403
rect 4100 3437 4170 3463
rect 4100 3403 4118 3437
rect 4152 3403 4170 3437
rect 4100 3377 4170 3403
rect 4200 3437 4270 3463
rect 4200 3403 4218 3437
rect 4252 3403 4270 3437
rect 4200 3377 4270 3403
rect 4300 3377 4370 3463
rect 4400 3377 4470 3463
rect 4500 3377 4570 3463
rect 4600 3437 4670 3463
rect 4600 3403 4618 3437
rect 4652 3403 4670 3437
rect 4600 3377 4670 3403
rect 4700 3437 4770 3463
rect 4700 3403 4718 3437
rect 4752 3403 4770 3437
rect 4700 3377 4770 3403
rect 4800 3377 4870 3463
rect 4900 3377 4970 3463
rect 5000 3437 5070 3463
rect 5000 3403 5018 3437
rect 5052 3403 5070 3437
rect 5000 3377 5070 3403
rect 5100 3437 5170 3463
rect 5100 3403 5118 3437
rect 5152 3403 5170 3437
rect 5100 3377 5170 3403
rect 5200 3437 5270 3463
rect 5200 3403 5218 3437
rect 5252 3403 5270 3437
rect 5200 3377 5270 3403
rect 5300 3437 5370 3463
rect 5300 3403 5318 3437
rect 5352 3403 5370 3437
rect 5300 3377 5370 3403
rect 5400 3437 5470 3463
rect 5400 3403 5418 3437
rect 5452 3403 5470 3437
rect 5400 3377 5470 3403
rect 5500 3437 5570 3463
rect 5500 3403 5518 3437
rect 5552 3403 5570 3437
rect 5500 3377 5570 3403
rect 5600 3437 5670 3463
rect 5600 3403 5618 3437
rect 5652 3403 5670 3437
rect 5600 3377 5670 3403
rect 5700 3377 5770 3463
rect 5800 3437 5870 3463
rect 5800 3403 5818 3437
rect 5852 3403 5870 3437
rect 5800 3377 5870 3403
rect 5900 3437 5954 3463
rect 5900 3403 5912 3437
rect 5946 3403 5954 3437
rect 5900 3377 5954 3403
rect 2816 3297 2870 3323
rect 2816 3263 2824 3297
rect 2858 3263 2870 3297
rect 2816 3237 2870 3263
rect 2900 3297 2954 3323
rect 2900 3263 2912 3297
rect 2946 3263 2954 3297
rect 2900 3237 2954 3263
rect 3016 3297 3070 3323
rect 3016 3263 3024 3297
rect 3058 3263 3070 3297
rect 3016 3237 3070 3263
rect 3100 3297 3170 3323
rect 3100 3263 3118 3297
rect 3152 3263 3170 3297
rect 3100 3237 3170 3263
rect 3200 3237 3270 3323
rect 3300 3237 3370 3323
rect 3400 3237 3470 3323
rect 3500 3237 3570 3323
rect 3600 3297 3670 3323
rect 3600 3263 3618 3297
rect 3652 3263 3670 3297
rect 3600 3237 3670 3263
rect 3700 3297 3770 3323
rect 3700 3263 3718 3297
rect 3752 3263 3770 3297
rect 3700 3237 3770 3263
rect 3800 3297 3870 3323
rect 3800 3263 3818 3297
rect 3852 3263 3870 3297
rect 3800 3237 3870 3263
rect 3900 3297 3970 3323
rect 3900 3263 3918 3297
rect 3952 3263 3970 3297
rect 3900 3237 3970 3263
rect 4000 3237 4070 3323
rect 4100 3237 4170 3323
rect 4200 3297 4270 3323
rect 4200 3263 4218 3297
rect 4252 3263 4270 3297
rect 4200 3237 4270 3263
rect 4300 3297 4354 3323
rect 4300 3263 4312 3297
rect 4346 3263 4354 3297
rect 4300 3237 4354 3263
rect 2516 3157 2570 3183
rect 2516 3123 2524 3157
rect 2558 3123 2570 3157
rect 2516 3097 2570 3123
rect 2600 3157 2670 3183
rect 2600 3123 2618 3157
rect 2652 3123 2670 3157
rect 2600 3097 2670 3123
rect 2700 3097 2770 3183
rect 2800 3097 2870 3183
rect 2900 3097 2970 3183
rect 3000 3097 3070 3183
rect 3100 3157 3170 3183
rect 3100 3123 3118 3157
rect 3152 3123 3170 3157
rect 3100 3097 3170 3123
rect 3200 3157 3254 3183
rect 3200 3123 3212 3157
rect 3246 3123 3254 3157
rect 3200 3097 3254 3123
rect 3316 3157 3370 3183
rect 3316 3123 3324 3157
rect 3358 3123 3370 3157
rect 3316 3097 3370 3123
rect 3400 3157 3470 3183
rect 3400 3123 3418 3157
rect 3452 3123 3470 3157
rect 3400 3097 3470 3123
rect 3500 3157 3570 3183
rect 3500 3123 3518 3157
rect 3552 3123 3570 3157
rect 3500 3097 3570 3123
rect 3600 3157 3654 3183
rect 3600 3123 3612 3157
rect 3646 3123 3654 3157
rect 3600 3097 3654 3123
rect 16 2957 70 3043
rect 100 3017 170 3043
rect 100 2983 118 3017
rect 152 2983 170 3017
rect 100 2957 170 2983
rect 200 3017 270 3043
rect 200 2983 218 3017
rect 252 2983 270 3017
rect 200 2957 270 2983
rect 300 2957 370 3043
rect 400 3017 470 3043
rect 400 2983 418 3017
rect 452 2983 470 3017
rect 400 2957 470 2983
rect 500 3017 570 3043
rect 500 2983 518 3017
rect 552 2983 570 3017
rect 500 2957 570 2983
rect 600 3017 670 3043
rect 600 2983 618 3017
rect 652 2983 670 3017
rect 600 2957 670 2983
rect 700 3017 770 3043
rect 700 2983 718 3017
rect 752 2983 770 3017
rect 700 2957 770 2983
rect 800 3017 870 3043
rect 800 2983 818 3017
rect 852 2983 870 3017
rect 800 2957 870 2983
rect 900 2957 970 3043
rect 1000 3017 1070 3043
rect 1000 2983 1018 3017
rect 1052 2983 1070 3017
rect 1000 2957 1070 2983
rect 1100 3017 1170 3043
rect 1100 2983 1118 3017
rect 1152 2983 1170 3017
rect 1100 2957 1170 2983
rect 1200 2957 1270 3043
rect 1300 2957 1370 3043
rect 1400 2957 1470 3043
rect 1500 2957 1570 3043
rect 1600 3017 1670 3043
rect 1600 2983 1618 3017
rect 1652 2983 1670 3017
rect 1600 2957 1670 2983
rect 1700 3017 1770 3043
rect 1700 2983 1718 3017
rect 1752 2983 1770 3017
rect 1700 2957 1770 2983
rect 1800 2957 1870 3043
rect 1900 2957 1970 3043
rect 2000 3017 2070 3043
rect 2000 2983 2018 3017
rect 2052 2983 2070 3017
rect 2000 2957 2070 2983
rect 2100 3017 2170 3043
rect 2100 2983 2118 3017
rect 2152 2983 2170 3017
rect 2100 2957 2170 2983
rect 2200 2957 2270 3043
rect 2300 2957 2370 3043
rect 2400 2957 2470 3043
rect 2500 3017 2570 3043
rect 2500 2983 2518 3017
rect 2552 2983 2570 3017
rect 2500 2957 2570 2983
rect 2600 3017 2670 3043
rect 2600 2983 2618 3017
rect 2652 2983 2670 3017
rect 2600 2957 2670 2983
rect 2700 3017 2770 3043
rect 2700 2983 2718 3017
rect 2752 2983 2770 3017
rect 2700 2957 2770 2983
rect 2800 3017 2870 3043
rect 2800 2983 2818 3017
rect 2852 2983 2870 3017
rect 2800 2957 2870 2983
rect 2900 2957 2970 3043
rect 3000 2957 3070 3043
rect 3100 2957 3170 3043
rect 3200 3017 3270 3043
rect 3200 2983 3218 3017
rect 3252 2983 3270 3017
rect 3200 2957 3270 2983
rect 3300 3017 3354 3043
rect 3300 2983 3312 3017
rect 3346 2983 3354 3017
rect 3300 2957 3354 2983
rect 16 2817 70 2903
rect 100 2877 170 2903
rect 100 2843 118 2877
rect 152 2843 170 2877
rect 100 2817 170 2843
rect 200 2877 270 2903
rect 200 2843 218 2877
rect 252 2843 270 2877
rect 200 2817 270 2843
rect 300 2877 354 2903
rect 300 2843 312 2877
rect 346 2843 354 2877
rect 300 2817 354 2843
rect 416 2877 470 2903
rect 416 2843 424 2877
rect 458 2843 470 2877
rect 416 2817 470 2843
rect 500 2877 570 2903
rect 500 2843 518 2877
rect 552 2843 570 2877
rect 500 2817 570 2843
rect 600 2877 670 2903
rect 600 2843 618 2877
rect 652 2843 670 2877
rect 600 2817 670 2843
rect 700 2877 754 2903
rect 700 2843 712 2877
rect 746 2843 754 2877
rect 700 2817 754 2843
rect 816 2877 870 2903
rect 816 2843 824 2877
rect 858 2843 870 2877
rect 816 2817 870 2843
rect 900 2877 970 2903
rect 900 2843 918 2877
rect 952 2843 970 2877
rect 900 2817 970 2843
rect 1000 2877 1070 2903
rect 1000 2843 1018 2877
rect 1052 2843 1070 2877
rect 1000 2817 1070 2843
rect 1100 2877 1170 2903
rect 1100 2843 1118 2877
rect 1152 2843 1170 2877
rect 1100 2817 1170 2843
rect 1200 2877 1270 2903
rect 1200 2843 1218 2877
rect 1252 2843 1270 2877
rect 1200 2817 1270 2843
rect 1300 2877 1370 2903
rect 1300 2843 1318 2877
rect 1352 2843 1370 2877
rect 1300 2817 1370 2843
rect 1400 2877 1454 2903
rect 1400 2843 1412 2877
rect 1446 2843 1454 2877
rect 1400 2817 1454 2843
rect 16 2677 70 2763
rect 100 2737 170 2763
rect 100 2703 118 2737
rect 152 2703 170 2737
rect 100 2677 170 2703
rect 200 2737 270 2763
rect 200 2703 218 2737
rect 252 2703 270 2737
rect 200 2677 270 2703
rect 300 2737 370 2763
rect 300 2703 318 2737
rect 352 2703 370 2737
rect 300 2677 370 2703
rect 400 2677 470 2763
rect 500 2737 570 2763
rect 500 2703 518 2737
rect 552 2703 570 2737
rect 500 2677 570 2703
rect 600 2737 670 2763
rect 600 2703 618 2737
rect 652 2703 670 2737
rect 600 2677 670 2703
rect 700 2677 770 2763
rect 800 2737 870 2763
rect 800 2703 818 2737
rect 852 2703 870 2737
rect 800 2677 870 2703
rect 900 2737 970 2763
rect 900 2703 918 2737
rect 952 2703 970 2737
rect 900 2677 970 2703
rect 1000 2677 1070 2763
rect 1100 2737 1170 2763
rect 1100 2703 1118 2737
rect 1152 2703 1170 2737
rect 1100 2677 1170 2703
rect 1200 2737 1270 2763
rect 1200 2703 1218 2737
rect 1252 2703 1270 2737
rect 1200 2677 1270 2703
rect 1300 2737 1354 2763
rect 1300 2703 1312 2737
rect 1346 2703 1354 2737
rect 1300 2677 1354 2703
rect 1516 2877 1570 2903
rect 1516 2843 1524 2877
rect 1558 2843 1570 2877
rect 1516 2817 1570 2843
rect 1600 2877 1670 2903
rect 1600 2843 1618 2877
rect 1652 2843 1670 2877
rect 1600 2817 1670 2843
rect 1700 2817 1770 2903
rect 1800 2817 1870 2903
rect 1900 2877 1970 2903
rect 1900 2843 1918 2877
rect 1952 2843 1970 2877
rect 1900 2817 1970 2843
rect 2000 2877 2070 2903
rect 2000 2843 2018 2877
rect 2052 2843 2070 2877
rect 2000 2817 2070 2843
rect 2100 2877 2154 2903
rect 2100 2843 2112 2877
rect 2146 2843 2154 2877
rect 2100 2817 2154 2843
rect 1416 2737 1470 2763
rect 1416 2703 1424 2737
rect 1458 2703 1470 2737
rect 1416 2677 1470 2703
rect 1500 2737 1554 2763
rect 1500 2703 1512 2737
rect 1546 2703 1554 2737
rect 1500 2677 1554 2703
rect 16 2537 70 2623
rect 100 2537 170 2623
rect 200 2597 270 2623
rect 200 2563 218 2597
rect 252 2563 270 2597
rect 200 2537 270 2563
rect 300 2597 370 2623
rect 300 2563 318 2597
rect 352 2563 370 2597
rect 300 2537 370 2563
rect 400 2537 470 2623
rect 500 2597 570 2623
rect 500 2563 518 2597
rect 552 2563 570 2597
rect 500 2537 570 2563
rect 600 2597 670 2623
rect 600 2563 618 2597
rect 652 2563 670 2597
rect 600 2537 670 2563
rect 700 2597 770 2623
rect 700 2563 718 2597
rect 752 2563 770 2597
rect 700 2537 770 2563
rect 800 2537 870 2623
rect 900 2537 970 2623
rect 1000 2597 1070 2623
rect 1000 2563 1018 2597
rect 1052 2563 1070 2597
rect 1000 2537 1070 2563
rect 1100 2597 1170 2623
rect 1100 2563 1118 2597
rect 1152 2563 1170 2597
rect 1100 2537 1170 2563
rect 1200 2537 1270 2623
rect 1300 2537 1370 2623
rect 1400 2597 1470 2623
rect 1400 2563 1418 2597
rect 1452 2563 1470 2597
rect 1400 2537 1470 2563
rect 1500 2597 1554 2623
rect 1500 2563 1512 2597
rect 1546 2563 1554 2597
rect 1500 2537 1554 2563
rect 1616 2737 1670 2763
rect 1616 2703 1624 2737
rect 1658 2703 1670 2737
rect 1616 2677 1670 2703
rect 1700 2737 1770 2763
rect 1700 2703 1718 2737
rect 1752 2703 1770 2737
rect 1700 2677 1770 2703
rect 1800 2737 1870 2763
rect 1800 2703 1818 2737
rect 1852 2703 1870 2737
rect 1800 2677 1870 2703
rect 1900 2737 1970 2763
rect 1900 2703 1918 2737
rect 1952 2703 1970 2737
rect 1900 2677 1970 2703
rect 2000 2737 2054 2763
rect 2000 2703 2012 2737
rect 2046 2703 2054 2737
rect 2000 2677 2054 2703
rect 2216 2877 2270 2903
rect 2216 2843 2224 2877
rect 2258 2843 2270 2877
rect 2216 2817 2270 2843
rect 2300 2877 2354 2903
rect 2300 2843 2312 2877
rect 2346 2843 2354 2877
rect 2300 2817 2354 2843
rect 2416 2877 2470 2903
rect 2416 2843 2424 2877
rect 2458 2843 2470 2877
rect 2416 2817 2470 2843
rect 2500 2877 2554 2903
rect 2500 2843 2512 2877
rect 2546 2843 2554 2877
rect 2500 2817 2554 2843
rect 2616 2877 2670 2903
rect 2616 2843 2624 2877
rect 2658 2843 2670 2877
rect 2616 2817 2670 2843
rect 2700 2877 2770 2903
rect 2700 2843 2718 2877
rect 2752 2843 2770 2877
rect 2700 2817 2770 2843
rect 2800 2817 2870 2903
rect 2900 2877 2970 2903
rect 2900 2843 2918 2877
rect 2952 2843 2970 2877
rect 2900 2817 2970 2843
rect 3000 2877 3054 2903
rect 3000 2843 3012 2877
rect 3046 2843 3054 2877
rect 3000 2817 3054 2843
rect 2116 2737 2170 2763
rect 2116 2703 2124 2737
rect 2158 2703 2170 2737
rect 2116 2677 2170 2703
rect 2200 2737 2270 2763
rect 2200 2703 2218 2737
rect 2252 2703 2270 2737
rect 2200 2677 2270 2703
rect 2300 2677 2370 2763
rect 2400 2677 2470 2763
rect 2500 2737 2570 2763
rect 2500 2703 2518 2737
rect 2552 2703 2570 2737
rect 2500 2677 2570 2703
rect 2600 2737 2670 2763
rect 2600 2703 2618 2737
rect 2652 2703 2670 2737
rect 2600 2677 2670 2703
rect 2700 2737 2770 2763
rect 2700 2703 2718 2737
rect 2752 2703 2770 2737
rect 2700 2677 2770 2703
rect 2800 2737 2854 2763
rect 2800 2703 2812 2737
rect 2846 2703 2854 2737
rect 2800 2677 2854 2703
rect 1616 2597 1670 2623
rect 1616 2563 1624 2597
rect 1658 2563 1670 2597
rect 1616 2537 1670 2563
rect 1700 2597 1770 2623
rect 1700 2563 1718 2597
rect 1752 2563 1770 2597
rect 1700 2537 1770 2563
rect 1800 2597 1870 2623
rect 1800 2563 1818 2597
rect 1852 2563 1870 2597
rect 1800 2537 1870 2563
rect 1900 2537 1970 2623
rect 2000 2597 2070 2623
rect 2000 2563 2018 2597
rect 2052 2563 2070 2597
rect 2000 2537 2070 2563
rect 2100 2597 2154 2623
rect 2100 2563 2112 2597
rect 2146 2563 2154 2597
rect 2100 2537 2154 2563
rect 2216 2597 2270 2623
rect 2216 2563 2224 2597
rect 2258 2563 2270 2597
rect 2216 2537 2270 2563
rect 2300 2597 2370 2623
rect 2300 2563 2318 2597
rect 2352 2563 2370 2597
rect 2300 2537 2370 2563
rect 2400 2597 2454 2623
rect 2400 2563 2412 2597
rect 2446 2563 2454 2597
rect 2400 2537 2454 2563
rect 2516 2597 2570 2623
rect 2516 2563 2524 2597
rect 2558 2563 2570 2597
rect 2516 2537 2570 2563
rect 2600 2597 2654 2623
rect 2600 2563 2612 2597
rect 2646 2563 2654 2597
rect 2600 2537 2654 2563
rect 3716 3157 3770 3183
rect 3716 3123 3724 3157
rect 3758 3123 3770 3157
rect 3716 3097 3770 3123
rect 3800 3157 3870 3183
rect 3800 3123 3818 3157
rect 3852 3123 3870 3157
rect 3800 3097 3870 3123
rect 3900 3157 3970 3183
rect 3900 3123 3918 3157
rect 3952 3123 3970 3157
rect 3900 3097 3970 3123
rect 4000 3097 4070 3183
rect 4100 3157 4170 3183
rect 4100 3123 4118 3157
rect 4152 3123 4170 3157
rect 4100 3097 4170 3123
rect 4200 3157 4254 3183
rect 4200 3123 4212 3157
rect 4246 3123 4254 3157
rect 4200 3097 4254 3123
rect 3416 3017 3470 3043
rect 3416 2983 3424 3017
rect 3458 2983 3470 3017
rect 3416 2957 3470 2983
rect 3500 3017 3570 3043
rect 3500 2983 3518 3017
rect 3552 2983 3570 3017
rect 3500 2957 3570 2983
rect 3600 3017 3670 3043
rect 3600 2983 3618 3017
rect 3652 2983 3670 3017
rect 3600 2957 3670 2983
rect 3700 3017 3770 3043
rect 3700 2983 3718 3017
rect 3752 2983 3770 3017
rect 3700 2957 3770 2983
rect 3800 3017 3854 3043
rect 3800 2983 3812 3017
rect 3846 2983 3854 3017
rect 3800 2957 3854 2983
rect 3916 3017 3970 3043
rect 3916 2983 3924 3017
rect 3958 2983 3970 3017
rect 3916 2957 3970 2983
rect 4000 3017 4054 3043
rect 4000 2983 4012 3017
rect 4046 2983 4054 3017
rect 4000 2957 4054 2983
rect 4416 3297 4470 3323
rect 4416 3263 4424 3297
rect 4458 3263 4470 3297
rect 4416 3237 4470 3263
rect 4500 3297 4570 3323
rect 4500 3263 4518 3297
rect 4552 3263 4570 3297
rect 4500 3237 4570 3263
rect 4600 3297 4670 3323
rect 4600 3263 4618 3297
rect 4652 3263 4670 3297
rect 4600 3237 4670 3263
rect 4700 3297 4770 3323
rect 4700 3263 4718 3297
rect 4752 3263 4770 3297
rect 4700 3237 4770 3263
rect 4800 3297 4854 3323
rect 4800 3263 4812 3297
rect 4846 3263 4854 3297
rect 4800 3237 4854 3263
rect 4316 3157 4370 3183
rect 4316 3123 4324 3157
rect 4358 3123 4370 3157
rect 4316 3097 4370 3123
rect 4400 3157 4470 3183
rect 4400 3123 4418 3157
rect 4452 3123 4470 3157
rect 4400 3097 4470 3123
rect 4500 3157 4554 3183
rect 4500 3123 4512 3157
rect 4546 3123 4554 3157
rect 4500 3097 4554 3123
rect 4116 3017 4170 3043
rect 4116 2983 4124 3017
rect 4158 2983 4170 3017
rect 4116 2957 4170 2983
rect 4200 3017 4270 3043
rect 4200 2983 4218 3017
rect 4252 2983 4270 3017
rect 4200 2957 4270 2983
rect 4300 3017 4370 3043
rect 4300 2983 4318 3017
rect 4352 2983 4370 3017
rect 4300 2957 4370 2983
rect 4400 3017 4470 3043
rect 4400 2983 4418 3017
rect 4452 2983 4470 3017
rect 4400 2957 4470 2983
rect 4500 3017 4554 3043
rect 4500 2983 4512 3017
rect 4546 2983 4554 3017
rect 4500 2957 4554 2983
rect 4616 3157 4670 3183
rect 4616 3123 4624 3157
rect 4658 3123 4670 3157
rect 4616 3097 4670 3123
rect 4700 3157 4754 3183
rect 4700 3123 4712 3157
rect 4746 3123 4754 3157
rect 4700 3097 4754 3123
rect 4916 3297 4970 3323
rect 4916 3263 4924 3297
rect 4958 3263 4970 3297
rect 4916 3237 4970 3263
rect 5000 3297 5070 3323
rect 5000 3263 5018 3297
rect 5052 3263 5070 3297
rect 5000 3237 5070 3263
rect 5100 3237 5170 3323
rect 5200 3297 5270 3323
rect 5200 3263 5218 3297
rect 5252 3263 5270 3297
rect 5200 3237 5270 3263
rect 5300 3297 5370 3323
rect 5300 3263 5318 3297
rect 5352 3263 5370 3297
rect 5300 3237 5370 3263
rect 5400 3297 5470 3323
rect 5400 3263 5418 3297
rect 5452 3263 5470 3297
rect 5400 3237 5470 3263
rect 5500 3297 5554 3323
rect 5500 3263 5512 3297
rect 5546 3263 5554 3297
rect 5500 3237 5554 3263
rect 4816 3157 4870 3183
rect 4816 3123 4824 3157
rect 4858 3123 4870 3157
rect 4816 3097 4870 3123
rect 4900 3157 4970 3183
rect 4900 3123 4918 3157
rect 4952 3123 4970 3157
rect 4900 3097 4970 3123
rect 5000 3157 5054 3183
rect 5000 3123 5012 3157
rect 5046 3123 5054 3157
rect 5000 3097 5054 3123
rect 5116 3157 5170 3183
rect 5116 3123 5124 3157
rect 5158 3123 5170 3157
rect 5116 3097 5170 3123
rect 5200 3157 5270 3183
rect 5200 3123 5218 3157
rect 5252 3123 5270 3157
rect 5200 3097 5270 3123
rect 5300 3097 5370 3183
rect 5400 3157 5470 3183
rect 5400 3123 5418 3157
rect 5452 3123 5470 3157
rect 5400 3097 5470 3123
rect 5500 3157 5554 3183
rect 5500 3123 5512 3157
rect 5546 3123 5554 3157
rect 5500 3097 5554 3123
rect 6016 3437 6070 3463
rect 6016 3403 6024 3437
rect 6058 3403 6070 3437
rect 6016 3377 6070 3403
rect 6100 3437 6170 3463
rect 6100 3403 6118 3437
rect 6152 3403 6170 3437
rect 6100 3377 6170 3403
rect 6200 3437 6270 3463
rect 6200 3403 6218 3437
rect 6252 3403 6270 3437
rect 6200 3377 6270 3403
rect 6300 3437 6370 3463
rect 6300 3403 6318 3437
rect 6352 3403 6370 3437
rect 6300 3377 6370 3403
rect 6400 3377 6454 3463
rect 6512 3452 6570 3463
rect 6512 3418 6524 3452
rect 6558 3418 6570 3452
rect 6512 3377 6570 3418
rect 6600 3437 6670 3463
rect 6600 3403 6618 3437
rect 6652 3403 6670 3437
rect 6600 3377 6670 3403
rect 6700 3422 6758 3463
rect 6700 3388 6712 3422
rect 6746 3388 6758 3422
rect 6700 3377 6758 3388
rect 6820 3437 6880 3463
rect 6820 3403 6828 3437
rect 6862 3403 6880 3437
rect 6820 3377 6880 3403
rect 6910 3437 6980 3463
rect 6910 3403 6928 3437
rect 6962 3403 6980 3437
rect 6910 3377 6980 3403
rect 7010 3437 7080 3463
rect 7010 3403 7028 3437
rect 7062 3403 7080 3437
rect 7010 3377 7080 3403
rect 7110 3437 7180 3463
rect 7110 3403 7128 3437
rect 7162 3403 7180 3437
rect 7110 3377 7180 3403
rect 7210 3437 7280 3463
rect 7210 3403 7228 3437
rect 7262 3403 7280 3437
rect 7210 3377 7280 3403
rect 7310 3437 7380 3463
rect 7310 3403 7328 3437
rect 7362 3403 7380 3437
rect 7310 3377 7380 3403
rect 7410 3437 7470 3463
rect 7410 3403 7428 3437
rect 7462 3403 7470 3437
rect 7410 3377 7470 3403
rect 5616 3297 5670 3323
rect 5616 3263 5624 3297
rect 5658 3263 5670 3297
rect 5616 3237 5670 3263
rect 5700 3297 5770 3323
rect 5700 3263 5718 3297
rect 5752 3263 5770 3297
rect 5700 3237 5770 3263
rect 5800 3237 5870 3323
rect 5900 3297 5970 3323
rect 5900 3263 5918 3297
rect 5952 3263 5970 3297
rect 5900 3237 5970 3263
rect 6000 3297 6070 3323
rect 6000 3263 6018 3297
rect 6052 3263 6070 3297
rect 6000 3237 6070 3263
rect 6100 3297 6170 3323
rect 6100 3263 6118 3297
rect 6152 3263 6170 3297
rect 6100 3237 6170 3263
rect 6200 3297 6270 3323
rect 6200 3263 6218 3297
rect 6252 3263 6270 3297
rect 6200 3237 6270 3263
rect 6300 3297 6370 3323
rect 6300 3263 6318 3297
rect 6352 3263 6370 3297
rect 6300 3237 6370 3263
rect 6400 3237 6454 3323
rect 6512 3312 6570 3323
rect 6512 3278 6524 3312
rect 6558 3278 6570 3312
rect 6512 3237 6570 3278
rect 6600 3297 6670 3323
rect 6600 3263 6618 3297
rect 6652 3263 6670 3297
rect 6600 3237 6670 3263
rect 6700 3282 6758 3323
rect 6700 3248 6712 3282
rect 6746 3248 6758 3282
rect 6700 3237 6758 3248
rect 6820 3297 6880 3323
rect 6820 3263 6828 3297
rect 6862 3263 6880 3297
rect 6820 3237 6880 3263
rect 6910 3297 6980 3323
rect 6910 3263 6928 3297
rect 6962 3263 6980 3297
rect 6910 3237 6980 3263
rect 7010 3297 7080 3323
rect 7010 3263 7028 3297
rect 7062 3263 7080 3297
rect 7010 3237 7080 3263
rect 7110 3297 7180 3323
rect 7110 3263 7128 3297
rect 7162 3263 7180 3297
rect 7110 3237 7180 3263
rect 7210 3297 7280 3323
rect 7210 3263 7228 3297
rect 7262 3263 7280 3297
rect 7210 3237 7280 3263
rect 7310 3297 7380 3323
rect 7310 3263 7328 3297
rect 7362 3263 7380 3297
rect 7310 3237 7380 3263
rect 7410 3297 7470 3323
rect 7410 3263 7428 3297
rect 7462 3263 7470 3297
rect 7410 3237 7470 3263
rect 5616 3157 5670 3183
rect 5616 3123 5624 3157
rect 5658 3123 5670 3157
rect 5616 3097 5670 3123
rect 5700 3157 5754 3183
rect 5700 3123 5712 3157
rect 5746 3123 5754 3157
rect 5700 3097 5754 3123
rect 5816 3157 5870 3183
rect 5816 3123 5824 3157
rect 5858 3123 5870 3157
rect 5816 3097 5870 3123
rect 5900 3157 5970 3183
rect 5900 3123 5918 3157
rect 5952 3123 5970 3157
rect 5900 3097 5970 3123
rect 6000 3157 6070 3183
rect 6000 3123 6018 3157
rect 6052 3123 6070 3157
rect 6000 3097 6070 3123
rect 6100 3157 6170 3183
rect 6100 3123 6118 3157
rect 6152 3123 6170 3157
rect 6100 3097 6170 3123
rect 6200 3097 6270 3183
rect 6300 3097 6370 3183
rect 6400 3097 6454 3183
rect 6512 3172 6570 3183
rect 6512 3138 6524 3172
rect 6558 3138 6570 3172
rect 6512 3097 6570 3138
rect 6600 3157 6670 3183
rect 6600 3123 6618 3157
rect 6652 3123 6670 3157
rect 6600 3097 6670 3123
rect 6700 3142 6758 3183
rect 6700 3108 6712 3142
rect 6746 3108 6758 3142
rect 6700 3097 6758 3108
rect 6820 3157 6880 3183
rect 6820 3123 6828 3157
rect 6862 3123 6880 3157
rect 6820 3097 6880 3123
rect 6910 3157 6980 3183
rect 6910 3123 6928 3157
rect 6962 3123 6980 3157
rect 6910 3097 6980 3123
rect 7010 3157 7080 3183
rect 7010 3123 7028 3157
rect 7062 3123 7080 3157
rect 7010 3097 7080 3123
rect 7110 3157 7180 3183
rect 7110 3123 7128 3157
rect 7162 3123 7180 3157
rect 7110 3097 7180 3123
rect 7210 3157 7280 3183
rect 7210 3123 7228 3157
rect 7262 3123 7280 3157
rect 7210 3097 7280 3123
rect 7310 3157 7380 3183
rect 7310 3123 7328 3157
rect 7362 3123 7380 3157
rect 7310 3097 7380 3123
rect 7410 3157 7470 3183
rect 7410 3123 7428 3157
rect 7462 3123 7470 3157
rect 7410 3097 7470 3123
rect 4616 3017 4670 3043
rect 4616 2983 4624 3017
rect 4658 2983 4670 3017
rect 4616 2957 4670 2983
rect 4700 3017 4770 3043
rect 4700 2983 4718 3017
rect 4752 2983 4770 3017
rect 4700 2957 4770 2983
rect 4800 2957 4870 3043
rect 4900 3017 4970 3043
rect 4900 2983 4918 3017
rect 4952 2983 4970 3017
rect 4900 2957 4970 2983
rect 5000 3017 5070 3043
rect 5000 2983 5018 3017
rect 5052 2983 5070 3017
rect 5000 2957 5070 2983
rect 5100 3017 5170 3043
rect 5100 2983 5118 3017
rect 5152 2983 5170 3017
rect 5100 2957 5170 2983
rect 5200 2957 5270 3043
rect 5300 3017 5370 3043
rect 5300 2983 5318 3017
rect 5352 2983 5370 3017
rect 5300 2957 5370 2983
rect 5400 3017 5470 3043
rect 5400 2983 5418 3017
rect 5452 2983 5470 3017
rect 5400 2957 5470 2983
rect 5500 3017 5570 3043
rect 5500 2983 5518 3017
rect 5552 2983 5570 3017
rect 5500 2957 5570 2983
rect 5600 3017 5670 3043
rect 5600 2983 5618 3017
rect 5652 2983 5670 3017
rect 5600 2957 5670 2983
rect 5700 2957 5770 3043
rect 5800 3017 5870 3043
rect 5800 2983 5818 3017
rect 5852 2983 5870 3017
rect 5800 2957 5870 2983
rect 5900 3017 5954 3043
rect 5900 2983 5912 3017
rect 5946 2983 5954 3017
rect 5900 2957 5954 2983
rect 6016 3017 6070 3043
rect 6016 2983 6024 3017
rect 6058 2983 6070 3017
rect 6016 2957 6070 2983
rect 6100 3017 6170 3043
rect 6100 2983 6118 3017
rect 6152 2983 6170 3017
rect 6100 2957 6170 2983
rect 6200 3017 6270 3043
rect 6200 2983 6218 3017
rect 6252 2983 6270 3017
rect 6200 2957 6270 2983
rect 6300 2957 6370 3043
rect 6400 2957 6454 3043
rect 6512 3032 6570 3043
rect 6512 2998 6524 3032
rect 6558 2998 6570 3032
rect 6512 2957 6570 2998
rect 6600 3017 6670 3043
rect 6600 2983 6618 3017
rect 6652 2983 6670 3017
rect 6600 2957 6670 2983
rect 6700 3002 6758 3043
rect 6700 2968 6712 3002
rect 6746 2968 6758 3002
rect 6700 2957 6758 2968
rect 6820 3017 6880 3043
rect 6820 2983 6828 3017
rect 6862 2983 6880 3017
rect 6820 2957 6880 2983
rect 6910 3017 6980 3043
rect 6910 2983 6928 3017
rect 6962 2983 6980 3017
rect 6910 2957 6980 2983
rect 7010 3017 7080 3043
rect 7010 2983 7028 3017
rect 7062 2983 7080 3017
rect 7010 2957 7080 2983
rect 7110 3017 7180 3043
rect 7110 2983 7128 3017
rect 7162 2983 7180 3017
rect 7110 2957 7180 2983
rect 7210 3017 7280 3043
rect 7210 2983 7228 3017
rect 7262 2983 7280 3017
rect 7210 2957 7280 2983
rect 7310 3017 7380 3043
rect 7310 2983 7328 3017
rect 7362 2983 7380 3017
rect 7310 2957 7380 2983
rect 7410 3017 7470 3043
rect 7410 2983 7428 3017
rect 7462 2983 7470 3017
rect 7410 2957 7470 2983
rect 3116 2877 3170 2903
rect 3116 2843 3124 2877
rect 3158 2843 3170 2877
rect 3116 2817 3170 2843
rect 3200 2877 3270 2903
rect 3200 2843 3218 2877
rect 3252 2843 3270 2877
rect 3200 2817 3270 2843
rect 3300 2877 3370 2903
rect 3300 2843 3318 2877
rect 3352 2843 3370 2877
rect 3300 2817 3370 2843
rect 3400 2817 3470 2903
rect 3500 2817 3570 2903
rect 3600 2817 3670 2903
rect 3700 2817 3770 2903
rect 3800 2817 3870 2903
rect 3900 2877 3970 2903
rect 3900 2843 3918 2877
rect 3952 2843 3970 2877
rect 3900 2817 3970 2843
rect 4000 2877 4070 2903
rect 4000 2843 4018 2877
rect 4052 2843 4070 2877
rect 4000 2817 4070 2843
rect 4100 2817 4170 2903
rect 4200 2817 4270 2903
rect 4300 2817 4370 2903
rect 4400 2877 4470 2903
rect 4400 2843 4418 2877
rect 4452 2843 4470 2877
rect 4400 2817 4470 2843
rect 4500 2877 4570 2903
rect 4500 2843 4518 2877
rect 4552 2843 4570 2877
rect 4500 2817 4570 2843
rect 4600 2877 4670 2903
rect 4600 2843 4618 2877
rect 4652 2843 4670 2877
rect 4600 2817 4670 2843
rect 4700 2817 4770 2903
rect 4800 2877 4870 2903
rect 4800 2843 4818 2877
rect 4852 2843 4870 2877
rect 4800 2817 4870 2843
rect 4900 2877 4970 2903
rect 4900 2843 4918 2877
rect 4952 2843 4970 2877
rect 4900 2817 4970 2843
rect 5000 2877 5070 2903
rect 5000 2843 5018 2877
rect 5052 2843 5070 2877
rect 5000 2817 5070 2843
rect 5100 2877 5170 2903
rect 5100 2843 5118 2877
rect 5152 2843 5170 2877
rect 5100 2817 5170 2843
rect 5200 2877 5270 2903
rect 5200 2843 5218 2877
rect 5252 2843 5270 2877
rect 5200 2817 5270 2843
rect 5300 2817 5370 2903
rect 5400 2817 5470 2903
rect 5500 2877 5570 2903
rect 5500 2843 5518 2877
rect 5552 2843 5570 2877
rect 5500 2817 5570 2843
rect 5600 2877 5670 2903
rect 5600 2843 5618 2877
rect 5652 2843 5670 2877
rect 5600 2817 5670 2843
rect 5700 2817 5770 2903
rect 5800 2817 5870 2903
rect 5900 2877 5970 2903
rect 5900 2843 5918 2877
rect 5952 2843 5970 2877
rect 5900 2817 5970 2843
rect 6000 2877 6054 2903
rect 6000 2843 6012 2877
rect 6046 2843 6054 2877
rect 6000 2817 6054 2843
rect 2916 2737 2970 2763
rect 2916 2703 2924 2737
rect 2958 2703 2970 2737
rect 2916 2677 2970 2703
rect 3000 2737 3070 2763
rect 3000 2703 3018 2737
rect 3052 2703 3070 2737
rect 3000 2677 3070 2703
rect 3100 2737 3154 2763
rect 3100 2703 3112 2737
rect 3146 2703 3154 2737
rect 3100 2677 3154 2703
rect 3216 2737 3270 2763
rect 3216 2703 3224 2737
rect 3258 2703 3270 2737
rect 3216 2677 3270 2703
rect 3300 2737 3370 2763
rect 3300 2703 3318 2737
rect 3352 2703 3370 2737
rect 3300 2677 3370 2703
rect 3400 2737 3470 2763
rect 3400 2703 3418 2737
rect 3452 2703 3470 2737
rect 3400 2677 3470 2703
rect 3500 2677 3570 2763
rect 3600 2677 3670 2763
rect 3700 2677 3770 2763
rect 3800 2677 3870 2763
rect 3900 2737 3970 2763
rect 3900 2703 3918 2737
rect 3952 2703 3970 2737
rect 3900 2677 3970 2703
rect 4000 2737 4070 2763
rect 4000 2703 4018 2737
rect 4052 2703 4070 2737
rect 4000 2677 4070 2703
rect 4100 2737 4170 2763
rect 4100 2703 4118 2737
rect 4152 2703 4170 2737
rect 4100 2677 4170 2703
rect 4200 2677 4270 2763
rect 4300 2737 4370 2763
rect 4300 2703 4318 2737
rect 4352 2703 4370 2737
rect 4300 2677 4370 2703
rect 4400 2737 4454 2763
rect 4400 2703 4412 2737
rect 4446 2703 4454 2737
rect 4400 2677 4454 2703
rect 2716 2597 2770 2623
rect 2716 2563 2724 2597
rect 2758 2563 2770 2597
rect 2716 2537 2770 2563
rect 2800 2597 2870 2623
rect 2800 2563 2818 2597
rect 2852 2563 2870 2597
rect 2800 2537 2870 2563
rect 2900 2597 2970 2623
rect 2900 2563 2918 2597
rect 2952 2563 2970 2597
rect 2900 2537 2970 2563
rect 3000 2597 3070 2623
rect 3000 2563 3018 2597
rect 3052 2563 3070 2597
rect 3000 2537 3070 2563
rect 3100 2597 3170 2623
rect 3100 2563 3118 2597
rect 3152 2563 3170 2597
rect 3100 2537 3170 2563
rect 3200 2597 3254 2623
rect 3200 2563 3212 2597
rect 3246 2563 3254 2597
rect 3200 2537 3254 2563
rect 3316 2597 3370 2623
rect 3316 2563 3324 2597
rect 3358 2563 3370 2597
rect 3316 2537 3370 2563
rect 3400 2597 3454 2623
rect 3400 2563 3412 2597
rect 3446 2563 3454 2597
rect 3400 2537 3454 2563
rect 4516 2737 4570 2763
rect 4516 2703 4524 2737
rect 4558 2703 4570 2737
rect 4516 2677 4570 2703
rect 4600 2737 4654 2763
rect 4600 2703 4612 2737
rect 4646 2703 4654 2737
rect 4600 2677 4654 2703
rect 4716 2737 4770 2763
rect 4716 2703 4724 2737
rect 4758 2703 4770 2737
rect 4716 2677 4770 2703
rect 4800 2737 4870 2763
rect 4800 2703 4818 2737
rect 4852 2703 4870 2737
rect 4800 2677 4870 2703
rect 4900 2677 4970 2763
rect 5000 2737 5070 2763
rect 5000 2703 5018 2737
rect 5052 2703 5070 2737
rect 5000 2677 5070 2703
rect 5100 2737 5170 2763
rect 5100 2703 5118 2737
rect 5152 2703 5170 2737
rect 5100 2677 5170 2703
rect 5200 2677 5270 2763
rect 5300 2737 5370 2763
rect 5300 2703 5318 2737
rect 5352 2703 5370 2737
rect 5300 2677 5370 2703
rect 5400 2737 5454 2763
rect 5400 2703 5412 2737
rect 5446 2703 5454 2737
rect 5400 2677 5454 2703
rect 6116 2877 6170 2903
rect 6116 2843 6124 2877
rect 6158 2843 6170 2877
rect 6116 2817 6170 2843
rect 6200 2877 6270 2903
rect 6200 2843 6218 2877
rect 6252 2843 6270 2877
rect 6200 2817 6270 2843
rect 6300 2877 6370 2903
rect 6300 2843 6318 2877
rect 6352 2843 6370 2877
rect 6300 2817 6370 2843
rect 6400 2877 6454 2903
rect 6400 2843 6412 2877
rect 6446 2843 6454 2877
rect 6400 2817 6454 2843
rect 6512 2892 6570 2903
rect 6512 2858 6524 2892
rect 6558 2858 6570 2892
rect 6512 2817 6570 2858
rect 6600 2877 6670 2903
rect 6600 2843 6618 2877
rect 6652 2843 6670 2877
rect 6600 2817 6670 2843
rect 6700 2862 6758 2903
rect 6700 2828 6712 2862
rect 6746 2828 6758 2862
rect 6700 2817 6758 2828
rect 6820 2877 6880 2903
rect 6820 2843 6828 2877
rect 6862 2843 6880 2877
rect 6820 2817 6880 2843
rect 6910 2877 6980 2903
rect 6910 2843 6928 2877
rect 6962 2843 6980 2877
rect 6910 2817 6980 2843
rect 7010 2877 7080 2903
rect 7010 2843 7028 2877
rect 7062 2843 7080 2877
rect 7010 2817 7080 2843
rect 7110 2877 7180 2903
rect 7110 2843 7128 2877
rect 7162 2843 7180 2877
rect 7110 2817 7180 2843
rect 7210 2877 7280 2903
rect 7210 2843 7228 2877
rect 7262 2843 7280 2877
rect 7210 2817 7280 2843
rect 7310 2877 7380 2903
rect 7310 2843 7328 2877
rect 7362 2843 7380 2877
rect 7310 2817 7380 2843
rect 7410 2877 7470 2903
rect 7410 2843 7428 2877
rect 7462 2843 7470 2877
rect 7410 2817 7470 2843
rect 5516 2737 5570 2763
rect 5516 2703 5524 2737
rect 5558 2703 5570 2737
rect 5516 2677 5570 2703
rect 5600 2737 5670 2763
rect 5600 2703 5618 2737
rect 5652 2703 5670 2737
rect 5600 2677 5670 2703
rect 5700 2737 5770 2763
rect 5700 2703 5718 2737
rect 5752 2703 5770 2737
rect 5700 2677 5770 2703
rect 5800 2677 5870 2763
rect 5900 2677 5970 2763
rect 6000 2677 6070 2763
rect 6100 2737 6170 2763
rect 6100 2703 6118 2737
rect 6152 2703 6170 2737
rect 6100 2677 6170 2703
rect 6200 2737 6270 2763
rect 6200 2703 6218 2737
rect 6252 2703 6270 2737
rect 6200 2677 6270 2703
rect 6300 2737 6370 2763
rect 6300 2703 6318 2737
rect 6352 2703 6370 2737
rect 6300 2677 6370 2703
rect 6400 2677 6454 2763
rect 6512 2752 6570 2763
rect 6512 2718 6524 2752
rect 6558 2718 6570 2752
rect 6512 2677 6570 2718
rect 6600 2737 6670 2763
rect 6600 2703 6618 2737
rect 6652 2703 6670 2737
rect 6600 2677 6670 2703
rect 6700 2722 6758 2763
rect 6700 2688 6712 2722
rect 6746 2688 6758 2722
rect 6700 2677 6758 2688
rect 6820 2737 6880 2763
rect 6820 2703 6828 2737
rect 6862 2703 6880 2737
rect 6820 2677 6880 2703
rect 6910 2737 6980 2763
rect 6910 2703 6928 2737
rect 6962 2703 6980 2737
rect 6910 2677 6980 2703
rect 7010 2737 7080 2763
rect 7010 2703 7028 2737
rect 7062 2703 7080 2737
rect 7010 2677 7080 2703
rect 7110 2737 7180 2763
rect 7110 2703 7128 2737
rect 7162 2703 7180 2737
rect 7110 2677 7180 2703
rect 7210 2737 7280 2763
rect 7210 2703 7228 2737
rect 7262 2703 7280 2737
rect 7210 2677 7280 2703
rect 7310 2737 7380 2763
rect 7310 2703 7328 2737
rect 7362 2703 7380 2737
rect 7310 2677 7380 2703
rect 7410 2737 7470 2763
rect 7410 2703 7428 2737
rect 7462 2703 7470 2737
rect 7410 2677 7470 2703
rect 3516 2597 3570 2623
rect 3516 2563 3524 2597
rect 3558 2563 3570 2597
rect 3516 2537 3570 2563
rect 3600 2597 3670 2623
rect 3600 2563 3618 2597
rect 3652 2563 3670 2597
rect 3600 2537 3670 2563
rect 3700 2597 3770 2623
rect 3700 2563 3718 2597
rect 3752 2563 3770 2597
rect 3700 2537 3770 2563
rect 3800 2597 3870 2623
rect 3800 2563 3818 2597
rect 3852 2563 3870 2597
rect 3800 2537 3870 2563
rect 3900 2537 3970 2623
rect 4000 2597 4070 2623
rect 4000 2563 4018 2597
rect 4052 2563 4070 2597
rect 4000 2537 4070 2563
rect 4100 2597 4170 2623
rect 4100 2563 4118 2597
rect 4152 2563 4170 2597
rect 4100 2537 4170 2563
rect 4200 2597 4270 2623
rect 4200 2563 4218 2597
rect 4252 2563 4270 2597
rect 4200 2537 4270 2563
rect 4300 2537 4370 2623
rect 4400 2597 4470 2623
rect 4400 2563 4418 2597
rect 4452 2563 4470 2597
rect 4400 2537 4470 2563
rect 4500 2597 4570 2623
rect 4500 2563 4518 2597
rect 4552 2563 4570 2597
rect 4500 2537 4570 2563
rect 4600 2537 4670 2623
rect 4700 2597 4770 2623
rect 4700 2563 4718 2597
rect 4752 2563 4770 2597
rect 4700 2537 4770 2563
rect 4800 2597 4870 2623
rect 4800 2563 4818 2597
rect 4852 2563 4870 2597
rect 4800 2537 4870 2563
rect 4900 2537 4970 2623
rect 5000 2597 5070 2623
rect 5000 2563 5018 2597
rect 5052 2563 5070 2597
rect 5000 2537 5070 2563
rect 5100 2597 5170 2623
rect 5100 2563 5118 2597
rect 5152 2563 5170 2597
rect 5100 2537 5170 2563
rect 5200 2597 5270 2623
rect 5200 2563 5218 2597
rect 5252 2563 5270 2597
rect 5200 2537 5270 2563
rect 5300 2537 5370 2623
rect 5400 2597 5470 2623
rect 5400 2563 5418 2597
rect 5452 2563 5470 2597
rect 5400 2537 5470 2563
rect 5500 2597 5554 2623
rect 5500 2563 5512 2597
rect 5546 2563 5554 2597
rect 5500 2537 5554 2563
rect 5616 2597 5670 2623
rect 5616 2563 5624 2597
rect 5658 2563 5670 2597
rect 5616 2537 5670 2563
rect 5700 2597 5770 2623
rect 5700 2563 5718 2597
rect 5752 2563 5770 2597
rect 5700 2537 5770 2563
rect 5800 2537 5870 2623
rect 5900 2597 5970 2623
rect 5900 2563 5918 2597
rect 5952 2563 5970 2597
rect 5900 2537 5970 2563
rect 6000 2597 6070 2623
rect 6000 2563 6018 2597
rect 6052 2563 6070 2597
rect 6000 2537 6070 2563
rect 6100 2537 6170 2623
rect 6200 2597 6270 2623
rect 6200 2563 6218 2597
rect 6252 2563 6270 2597
rect 6200 2537 6270 2563
rect 6300 2597 6370 2623
rect 6300 2563 6318 2597
rect 6352 2563 6370 2597
rect 6300 2537 6370 2563
rect 6400 2537 6454 2623
rect 6512 2612 6570 2623
rect 6512 2578 6524 2612
rect 6558 2578 6570 2612
rect 6512 2537 6570 2578
rect 6600 2597 6670 2623
rect 6600 2563 6618 2597
rect 6652 2563 6670 2597
rect 6600 2537 6670 2563
rect 6700 2582 6758 2623
rect 6700 2548 6712 2582
rect 6746 2548 6758 2582
rect 6700 2537 6758 2548
rect 6820 2597 6880 2623
rect 6820 2563 6828 2597
rect 6862 2563 6880 2597
rect 6820 2537 6880 2563
rect 6910 2597 6980 2623
rect 6910 2563 6928 2597
rect 6962 2563 6980 2597
rect 6910 2537 6980 2563
rect 7010 2597 7080 2623
rect 7010 2563 7028 2597
rect 7062 2563 7080 2597
rect 7010 2537 7080 2563
rect 7110 2597 7180 2623
rect 7110 2563 7128 2597
rect 7162 2563 7180 2597
rect 7110 2537 7180 2563
rect 7210 2597 7280 2623
rect 7210 2563 7228 2597
rect 7262 2563 7280 2597
rect 7210 2537 7280 2563
rect 7310 2597 7380 2623
rect 7310 2563 7328 2597
rect 7362 2563 7380 2597
rect 7310 2537 7380 2563
rect 7410 2597 7470 2623
rect 7410 2563 7428 2597
rect 7462 2563 7470 2597
rect 7410 2537 7470 2563
rect 16 2307 70 2393
rect 100 2307 170 2393
rect 200 2307 270 2393
rect 300 2307 370 2393
rect 400 2367 470 2393
rect 400 2333 418 2367
rect 452 2333 470 2367
rect 400 2307 470 2333
rect 500 2367 570 2393
rect 500 2333 518 2367
rect 552 2333 570 2367
rect 500 2307 570 2333
rect 600 2307 670 2393
rect 700 2307 770 2393
rect 800 2367 870 2393
rect 800 2333 818 2367
rect 852 2333 870 2367
rect 800 2307 870 2333
rect 900 2367 970 2393
rect 900 2333 918 2367
rect 952 2333 970 2367
rect 900 2307 970 2333
rect 1000 2367 1070 2393
rect 1000 2333 1018 2367
rect 1052 2333 1070 2367
rect 1000 2307 1070 2333
rect 1100 2307 1170 2393
rect 1200 2307 1270 2393
rect 1300 2307 1370 2393
rect 1400 2307 1470 2393
rect 1500 2367 1570 2393
rect 1500 2333 1518 2367
rect 1552 2333 1570 2367
rect 1500 2307 1570 2333
rect 1600 2367 1670 2393
rect 1600 2333 1618 2367
rect 1652 2333 1670 2367
rect 1600 2307 1670 2333
rect 1700 2307 1770 2393
rect 1800 2367 1870 2393
rect 1800 2333 1818 2367
rect 1852 2333 1870 2367
rect 1800 2307 1870 2333
rect 1900 2367 1970 2393
rect 1900 2333 1918 2367
rect 1952 2333 1970 2367
rect 1900 2307 1970 2333
rect 2000 2367 2070 2393
rect 2000 2333 2018 2367
rect 2052 2333 2070 2367
rect 2000 2307 2070 2333
rect 2100 2367 2170 2393
rect 2100 2333 2118 2367
rect 2152 2333 2170 2367
rect 2100 2307 2170 2333
rect 2200 2307 2270 2393
rect 2300 2367 2370 2393
rect 2300 2333 2318 2367
rect 2352 2333 2370 2367
rect 2300 2307 2370 2333
rect 2400 2367 2470 2393
rect 2400 2333 2418 2367
rect 2452 2333 2470 2367
rect 2400 2307 2470 2333
rect 2500 2367 2570 2393
rect 2500 2333 2518 2367
rect 2552 2333 2570 2367
rect 2500 2307 2570 2333
rect 2600 2307 2670 2393
rect 2700 2367 2770 2393
rect 2700 2333 2718 2367
rect 2752 2333 2770 2367
rect 2700 2307 2770 2333
rect 2800 2367 2870 2393
rect 2800 2333 2818 2367
rect 2852 2333 2870 2367
rect 2800 2307 2870 2333
rect 2900 2307 2970 2393
rect 3000 2307 3070 2393
rect 3100 2307 3170 2393
rect 3200 2307 3270 2393
rect 3300 2367 3370 2393
rect 3300 2333 3318 2367
rect 3352 2333 3370 2367
rect 3300 2307 3370 2333
rect 3400 2367 3470 2393
rect 3400 2333 3418 2367
rect 3452 2333 3470 2367
rect 3400 2307 3470 2333
rect 3500 2307 3570 2393
rect 3600 2307 3670 2393
rect 3700 2307 3770 2393
rect 3800 2307 3870 2393
rect 3900 2307 3970 2393
rect 4000 2367 4070 2393
rect 4000 2333 4018 2367
rect 4052 2333 4070 2367
rect 4000 2307 4070 2333
rect 4100 2367 4170 2393
rect 4100 2333 4118 2367
rect 4152 2333 4170 2367
rect 4100 2307 4170 2333
rect 4200 2307 4270 2393
rect 4300 2367 4370 2393
rect 4300 2333 4318 2367
rect 4352 2333 4370 2367
rect 4300 2307 4370 2333
rect 4400 2367 4470 2393
rect 4400 2333 4418 2367
rect 4452 2333 4470 2367
rect 4400 2307 4470 2333
rect 4500 2307 4570 2393
rect 4600 2307 4670 2393
rect 4700 2367 4770 2393
rect 4700 2333 4718 2367
rect 4752 2333 4770 2367
rect 4700 2307 4770 2333
rect 4800 2367 4870 2393
rect 4800 2333 4818 2367
rect 4852 2333 4870 2367
rect 4800 2307 4870 2333
rect 4900 2367 4970 2393
rect 4900 2333 4918 2367
rect 4952 2333 4970 2367
rect 4900 2307 4970 2333
rect 5000 2367 5070 2393
rect 5000 2333 5018 2367
rect 5052 2333 5070 2367
rect 5000 2307 5070 2333
rect 5100 2307 5170 2393
rect 5200 2307 5270 2393
rect 5300 2367 5370 2393
rect 5300 2333 5318 2367
rect 5352 2333 5370 2367
rect 5300 2307 5370 2333
rect 5400 2367 5454 2393
rect 5400 2333 5412 2367
rect 5446 2333 5454 2367
rect 5400 2307 5454 2333
rect 16 2227 70 2253
rect 16 2193 24 2227
rect 58 2193 70 2227
rect 16 2167 70 2193
rect 100 2227 170 2253
rect 100 2193 118 2227
rect 152 2193 170 2227
rect 100 2167 170 2193
rect 200 2227 254 2253
rect 200 2193 212 2227
rect 246 2193 254 2227
rect 200 2167 254 2193
rect 316 2227 370 2253
rect 316 2193 324 2227
rect 358 2193 370 2227
rect 316 2167 370 2193
rect 400 2227 470 2253
rect 400 2193 418 2227
rect 452 2193 470 2227
rect 400 2167 470 2193
rect 500 2227 570 2253
rect 500 2193 518 2227
rect 552 2193 570 2227
rect 500 2167 570 2193
rect 600 2227 670 2253
rect 600 2193 618 2227
rect 652 2193 670 2227
rect 600 2167 670 2193
rect 700 2167 770 2253
rect 800 2167 870 2253
rect 900 2167 970 2253
rect 1000 2227 1070 2253
rect 1000 2193 1018 2227
rect 1052 2193 1070 2227
rect 1000 2167 1070 2193
rect 1100 2227 1170 2253
rect 1100 2193 1118 2227
rect 1152 2193 1170 2227
rect 1100 2167 1170 2193
rect 1200 2227 1270 2253
rect 1200 2193 1218 2227
rect 1252 2193 1270 2227
rect 1200 2167 1270 2193
rect 1300 2227 1354 2253
rect 1300 2193 1312 2227
rect 1346 2193 1354 2227
rect 1300 2167 1354 2193
rect 16 2087 70 2113
rect 16 2053 24 2087
rect 58 2053 70 2087
rect 16 2027 70 2053
rect 100 2087 170 2113
rect 100 2053 118 2087
rect 152 2053 170 2087
rect 100 2027 170 2053
rect 200 2087 270 2113
rect 200 2053 218 2087
rect 252 2053 270 2087
rect 200 2027 270 2053
rect 300 2087 354 2113
rect 300 2053 312 2087
rect 346 2053 354 2087
rect 300 2027 354 2053
rect 16 1887 70 1973
rect 100 1887 170 1973
rect 200 1947 270 1973
rect 200 1913 218 1947
rect 252 1913 270 1947
rect 200 1887 270 1913
rect 300 1947 354 1973
rect 300 1913 312 1947
rect 346 1913 354 1947
rect 300 1887 354 1913
rect 416 2087 470 2113
rect 416 2053 424 2087
rect 458 2053 470 2087
rect 416 2027 470 2053
rect 500 2087 570 2113
rect 500 2053 518 2087
rect 552 2053 570 2087
rect 500 2027 570 2053
rect 600 2087 670 2113
rect 600 2053 618 2087
rect 652 2053 670 2087
rect 600 2027 670 2053
rect 700 2027 770 2113
rect 800 2087 870 2113
rect 800 2053 818 2087
rect 852 2053 870 2087
rect 800 2027 870 2053
rect 900 2087 970 2113
rect 900 2053 918 2087
rect 952 2053 970 2087
rect 900 2027 970 2053
rect 1000 2027 1070 2113
rect 1100 2027 1170 2113
rect 1200 2087 1270 2113
rect 1200 2053 1218 2087
rect 1252 2053 1270 2087
rect 1200 2027 1270 2053
rect 1300 2087 1354 2113
rect 1300 2053 1312 2087
rect 1346 2053 1354 2087
rect 1300 2027 1354 2053
rect 1416 2227 1470 2253
rect 1416 2193 1424 2227
rect 1458 2193 1470 2227
rect 1416 2167 1470 2193
rect 1500 2227 1554 2253
rect 1500 2193 1512 2227
rect 1546 2193 1554 2227
rect 1500 2167 1554 2193
rect 1416 2087 1470 2113
rect 1416 2053 1424 2087
rect 1458 2053 1470 2087
rect 1416 2027 1470 2053
rect 1500 2087 1554 2113
rect 1500 2053 1512 2087
rect 1546 2053 1554 2087
rect 1500 2027 1554 2053
rect 416 1947 470 1973
rect 416 1913 424 1947
rect 458 1913 470 1947
rect 416 1887 470 1913
rect 500 1947 570 1973
rect 500 1913 518 1947
rect 552 1913 570 1947
rect 500 1887 570 1913
rect 600 1887 670 1973
rect 700 1947 770 1973
rect 700 1913 718 1947
rect 752 1913 770 1947
rect 700 1887 770 1913
rect 800 1947 870 1973
rect 800 1913 818 1947
rect 852 1913 870 1947
rect 800 1887 870 1913
rect 900 1947 970 1973
rect 900 1913 918 1947
rect 952 1913 970 1947
rect 900 1887 970 1913
rect 1000 1947 1070 1973
rect 1000 1913 1018 1947
rect 1052 1913 1070 1947
rect 1000 1887 1070 1913
rect 1100 1947 1170 1973
rect 1100 1913 1118 1947
rect 1152 1913 1170 1947
rect 1100 1887 1170 1913
rect 1200 1947 1270 1973
rect 1200 1913 1218 1947
rect 1252 1913 1270 1947
rect 1200 1887 1270 1913
rect 1300 1947 1370 1973
rect 1300 1913 1318 1947
rect 1352 1913 1370 1947
rect 1300 1887 1370 1913
rect 1400 1947 1454 1973
rect 1400 1913 1412 1947
rect 1446 1913 1454 1947
rect 1400 1887 1454 1913
rect 16 1747 70 1833
rect 100 1807 170 1833
rect 100 1773 118 1807
rect 152 1773 170 1807
rect 100 1747 170 1773
rect 200 1807 270 1833
rect 200 1773 218 1807
rect 252 1773 270 1807
rect 200 1747 270 1773
rect 300 1747 370 1833
rect 400 1747 470 1833
rect 500 1747 570 1833
rect 600 1747 670 1833
rect 700 1807 770 1833
rect 700 1773 718 1807
rect 752 1773 770 1807
rect 700 1747 770 1773
rect 800 1807 870 1833
rect 800 1773 818 1807
rect 852 1773 870 1807
rect 800 1747 870 1773
rect 900 1807 954 1833
rect 900 1773 912 1807
rect 946 1773 954 1807
rect 900 1747 954 1773
rect 16 1667 70 1693
rect 16 1633 24 1667
rect 58 1633 70 1667
rect 16 1607 70 1633
rect 100 1667 154 1693
rect 100 1633 112 1667
rect 146 1633 154 1667
rect 100 1607 154 1633
rect 16 1527 70 1553
rect 16 1493 24 1527
rect 58 1493 70 1527
rect 16 1467 70 1493
rect 100 1527 154 1553
rect 100 1493 112 1527
rect 146 1493 154 1527
rect 100 1467 154 1493
rect 216 1667 270 1693
rect 216 1633 224 1667
rect 258 1633 270 1667
rect 216 1607 270 1633
rect 300 1667 370 1693
rect 300 1633 318 1667
rect 352 1633 370 1667
rect 300 1607 370 1633
rect 400 1667 470 1693
rect 400 1633 418 1667
rect 452 1633 470 1667
rect 400 1607 470 1633
rect 500 1607 570 1693
rect 600 1667 670 1693
rect 600 1633 618 1667
rect 652 1633 670 1667
rect 600 1607 670 1633
rect 700 1667 754 1693
rect 700 1633 712 1667
rect 746 1633 754 1667
rect 700 1607 754 1633
rect 216 1527 270 1553
rect 216 1493 224 1527
rect 258 1493 270 1527
rect 216 1467 270 1493
rect 300 1527 370 1553
rect 300 1493 318 1527
rect 352 1493 370 1527
rect 300 1467 370 1493
rect 400 1527 454 1553
rect 400 1493 412 1527
rect 446 1493 454 1527
rect 400 1467 454 1493
rect 16 1327 70 1413
rect 100 1387 170 1413
rect 100 1353 118 1387
rect 152 1353 170 1387
rect 100 1327 170 1353
rect 200 1387 254 1413
rect 200 1353 212 1387
rect 246 1353 254 1387
rect 200 1327 254 1353
rect 816 1667 870 1693
rect 816 1633 824 1667
rect 858 1633 870 1667
rect 816 1607 870 1633
rect 900 1667 954 1693
rect 900 1633 912 1667
rect 946 1633 954 1667
rect 900 1607 954 1633
rect 1616 2227 1670 2253
rect 1616 2193 1624 2227
rect 1658 2193 1670 2227
rect 1616 2167 1670 2193
rect 1700 2227 1770 2253
rect 1700 2193 1718 2227
rect 1752 2193 1770 2227
rect 1700 2167 1770 2193
rect 1800 2227 1854 2253
rect 1800 2193 1812 2227
rect 1846 2193 1854 2227
rect 1800 2167 1854 2193
rect 1616 2087 1670 2113
rect 1616 2053 1624 2087
rect 1658 2053 1670 2087
rect 1616 2027 1670 2053
rect 1700 2087 1770 2113
rect 1700 2053 1718 2087
rect 1752 2053 1770 2087
rect 1700 2027 1770 2053
rect 1800 2087 1854 2113
rect 1800 2053 1812 2087
rect 1846 2053 1854 2087
rect 1800 2027 1854 2053
rect 1916 2227 1970 2253
rect 1916 2193 1924 2227
rect 1958 2193 1970 2227
rect 1916 2167 1970 2193
rect 2000 2227 2070 2253
rect 2000 2193 2018 2227
rect 2052 2193 2070 2227
rect 2000 2167 2070 2193
rect 2100 2227 2170 2253
rect 2100 2193 2118 2227
rect 2152 2193 2170 2227
rect 2100 2167 2170 2193
rect 2200 2227 2254 2253
rect 2200 2193 2212 2227
rect 2246 2193 2254 2227
rect 2200 2167 2254 2193
rect 1916 2087 1970 2113
rect 1916 2053 1924 2087
rect 1958 2053 1970 2087
rect 1916 2027 1970 2053
rect 2000 2087 2070 2113
rect 2000 2053 2018 2087
rect 2052 2053 2070 2087
rect 2000 2027 2070 2053
rect 2100 2087 2170 2113
rect 2100 2053 2118 2087
rect 2152 2053 2170 2087
rect 2100 2027 2170 2053
rect 2200 2087 2254 2113
rect 2200 2053 2212 2087
rect 2246 2053 2254 2087
rect 2200 2027 2254 2053
rect 2316 2227 2370 2253
rect 2316 2193 2324 2227
rect 2358 2193 2370 2227
rect 2316 2167 2370 2193
rect 2400 2227 2470 2253
rect 2400 2193 2418 2227
rect 2452 2193 2470 2227
rect 2400 2167 2470 2193
rect 2500 2167 2570 2253
rect 2600 2227 2670 2253
rect 2600 2193 2618 2227
rect 2652 2193 2670 2227
rect 2600 2167 2670 2193
rect 2700 2227 2770 2253
rect 2700 2193 2718 2227
rect 2752 2193 2770 2227
rect 2700 2167 2770 2193
rect 2800 2227 2854 2253
rect 2800 2193 2812 2227
rect 2846 2193 2854 2227
rect 2800 2167 2854 2193
rect 2316 2087 2370 2113
rect 2316 2053 2324 2087
rect 2358 2053 2370 2087
rect 2316 2027 2370 2053
rect 2400 2087 2454 2113
rect 2400 2053 2412 2087
rect 2446 2053 2454 2087
rect 2400 2027 2454 2053
rect 1516 1947 1570 1973
rect 1516 1913 1524 1947
rect 1558 1913 1570 1947
rect 1516 1887 1570 1913
rect 1600 1947 1670 1973
rect 1600 1913 1618 1947
rect 1652 1913 1670 1947
rect 1600 1887 1670 1913
rect 1700 1947 1770 1973
rect 1700 1913 1718 1947
rect 1752 1913 1770 1947
rect 1700 1887 1770 1913
rect 1800 1947 1870 1973
rect 1800 1913 1818 1947
rect 1852 1913 1870 1947
rect 1800 1887 1870 1913
rect 1900 1947 1970 1973
rect 1900 1913 1918 1947
rect 1952 1913 1970 1947
rect 1900 1887 1970 1913
rect 2000 1947 2070 1973
rect 2000 1913 2018 1947
rect 2052 1913 2070 1947
rect 2000 1887 2070 1913
rect 2100 1887 2170 1973
rect 2200 1887 2270 1973
rect 2300 1947 2370 1973
rect 2300 1913 2318 1947
rect 2352 1913 2370 1947
rect 2300 1887 2370 1913
rect 2400 1947 2454 1973
rect 2400 1913 2412 1947
rect 2446 1913 2454 1947
rect 2400 1887 2454 1913
rect 1016 1807 1070 1833
rect 1016 1773 1024 1807
rect 1058 1773 1070 1807
rect 1016 1747 1070 1773
rect 1100 1807 1170 1833
rect 1100 1773 1118 1807
rect 1152 1773 1170 1807
rect 1100 1747 1170 1773
rect 1200 1747 1270 1833
rect 1300 1747 1370 1833
rect 1400 1807 1470 1833
rect 1400 1773 1418 1807
rect 1452 1773 1470 1807
rect 1400 1747 1470 1773
rect 1500 1807 1570 1833
rect 1500 1773 1518 1807
rect 1552 1773 1570 1807
rect 1500 1747 1570 1773
rect 1600 1747 1670 1833
rect 1700 1807 1770 1833
rect 1700 1773 1718 1807
rect 1752 1773 1770 1807
rect 1700 1747 1770 1773
rect 1800 1807 1854 1833
rect 1800 1773 1812 1807
rect 1846 1773 1854 1807
rect 1800 1747 1854 1773
rect 1016 1667 1070 1693
rect 1016 1633 1024 1667
rect 1058 1633 1070 1667
rect 1016 1607 1070 1633
rect 1100 1667 1170 1693
rect 1100 1633 1118 1667
rect 1152 1633 1170 1667
rect 1100 1607 1170 1633
rect 1200 1667 1270 1693
rect 1200 1633 1218 1667
rect 1252 1633 1270 1667
rect 1200 1607 1270 1633
rect 1300 1667 1370 1693
rect 1300 1633 1318 1667
rect 1352 1633 1370 1667
rect 1300 1607 1370 1633
rect 1400 1667 1470 1693
rect 1400 1633 1418 1667
rect 1452 1633 1470 1667
rect 1400 1607 1470 1633
rect 1500 1667 1554 1693
rect 1500 1633 1512 1667
rect 1546 1633 1554 1667
rect 1500 1607 1554 1633
rect 1616 1667 1670 1693
rect 1616 1633 1624 1667
rect 1658 1633 1670 1667
rect 1616 1607 1670 1633
rect 1700 1667 1754 1693
rect 1700 1633 1712 1667
rect 1746 1633 1754 1667
rect 1700 1607 1754 1633
rect 516 1527 570 1553
rect 516 1493 524 1527
rect 558 1493 570 1527
rect 516 1467 570 1493
rect 600 1527 670 1553
rect 600 1493 618 1527
rect 652 1493 670 1527
rect 600 1467 670 1493
rect 700 1467 770 1553
rect 800 1527 870 1553
rect 800 1493 818 1527
rect 852 1493 870 1527
rect 800 1467 870 1493
rect 900 1527 970 1553
rect 900 1493 918 1527
rect 952 1493 970 1527
rect 900 1467 970 1493
rect 1000 1467 1070 1553
rect 1100 1527 1170 1553
rect 1100 1493 1118 1527
rect 1152 1493 1170 1527
rect 1100 1467 1170 1493
rect 1200 1527 1270 1553
rect 1200 1493 1218 1527
rect 1252 1493 1270 1527
rect 1200 1467 1270 1493
rect 1300 1527 1370 1553
rect 1300 1493 1318 1527
rect 1352 1493 1370 1527
rect 1300 1467 1370 1493
rect 1400 1467 1470 1553
rect 1500 1527 1570 1553
rect 1500 1493 1518 1527
rect 1552 1493 1570 1527
rect 1500 1467 1570 1493
rect 1600 1527 1654 1553
rect 1600 1493 1612 1527
rect 1646 1493 1654 1527
rect 1600 1467 1654 1493
rect 316 1387 370 1413
rect 316 1353 324 1387
rect 358 1353 370 1387
rect 316 1327 370 1353
rect 400 1387 470 1413
rect 400 1353 418 1387
rect 452 1353 470 1387
rect 400 1327 470 1353
rect 500 1387 554 1413
rect 500 1353 512 1387
rect 546 1353 554 1387
rect 500 1327 554 1353
rect 16 1097 70 1183
rect 100 1097 170 1183
rect 200 1157 270 1183
rect 200 1123 218 1157
rect 252 1123 270 1157
rect 200 1097 270 1123
rect 300 1157 354 1183
rect 300 1123 312 1157
rect 346 1123 354 1157
rect 300 1097 354 1123
rect 616 1387 670 1413
rect 616 1353 624 1387
rect 658 1353 670 1387
rect 616 1327 670 1353
rect 700 1387 770 1413
rect 700 1353 718 1387
rect 752 1353 770 1387
rect 700 1327 770 1353
rect 800 1327 870 1413
rect 900 1327 970 1413
rect 1000 1387 1070 1413
rect 1000 1353 1018 1387
rect 1052 1353 1070 1387
rect 1000 1327 1070 1353
rect 1100 1387 1170 1413
rect 1100 1353 1118 1387
rect 1152 1353 1170 1387
rect 1100 1327 1170 1353
rect 1200 1327 1270 1413
rect 1300 1387 1370 1413
rect 1300 1353 1318 1387
rect 1352 1353 1370 1387
rect 1300 1327 1370 1353
rect 1400 1387 1470 1413
rect 1400 1353 1418 1387
rect 1452 1353 1470 1387
rect 1400 1327 1470 1353
rect 1500 1387 1554 1413
rect 1500 1353 1512 1387
rect 1546 1353 1554 1387
rect 1500 1327 1554 1353
rect 416 1157 470 1183
rect 416 1123 424 1157
rect 458 1123 470 1157
rect 416 1097 470 1123
rect 500 1157 554 1183
rect 500 1123 512 1157
rect 546 1123 554 1157
rect 500 1097 554 1123
rect 616 1157 670 1183
rect 616 1123 624 1157
rect 658 1123 670 1157
rect 616 1097 670 1123
rect 700 1157 754 1183
rect 700 1123 712 1157
rect 746 1123 754 1157
rect 700 1097 754 1123
rect 816 1157 870 1183
rect 816 1123 824 1157
rect 858 1123 870 1157
rect 816 1097 870 1123
rect 900 1157 970 1183
rect 900 1123 918 1157
rect 952 1123 970 1157
rect 900 1097 970 1123
rect 1000 1157 1070 1183
rect 1000 1123 1018 1157
rect 1052 1123 1070 1157
rect 1000 1097 1070 1123
rect 1100 1157 1170 1183
rect 1100 1123 1118 1157
rect 1152 1123 1170 1157
rect 1100 1097 1170 1123
rect 1200 1157 1254 1183
rect 1200 1123 1212 1157
rect 1246 1123 1254 1157
rect 1200 1097 1254 1123
rect 16 957 70 1043
rect 100 1017 170 1043
rect 100 983 118 1017
rect 152 983 170 1017
rect 100 957 170 983
rect 200 1017 270 1043
rect 200 983 218 1017
rect 252 983 270 1017
rect 200 957 270 983
rect 300 957 370 1043
rect 400 957 470 1043
rect 500 1017 570 1043
rect 500 983 518 1017
rect 552 983 570 1017
rect 500 957 570 983
rect 600 1017 670 1043
rect 600 983 618 1017
rect 652 983 670 1017
rect 600 957 670 983
rect 700 957 770 1043
rect 800 1017 870 1043
rect 800 983 818 1017
rect 852 983 870 1017
rect 800 957 870 983
rect 900 1017 954 1043
rect 900 983 912 1017
rect 946 983 954 1017
rect 900 957 954 983
rect 1016 1017 1070 1043
rect 1016 983 1024 1017
rect 1058 983 1070 1017
rect 1016 957 1070 983
rect 1100 1017 1154 1043
rect 1100 983 1112 1017
rect 1146 983 1154 1017
rect 1100 957 1154 983
rect 16 817 70 903
rect 100 817 170 903
rect 200 817 270 903
rect 300 817 370 903
rect 400 817 470 903
rect 500 817 570 903
rect 600 817 670 903
rect 700 817 770 903
rect 800 817 870 903
rect 900 877 970 903
rect 900 843 918 877
rect 952 843 970 877
rect 900 817 970 843
rect 1000 877 1054 903
rect 1000 843 1012 877
rect 1046 843 1054 877
rect 1000 817 1054 843
rect 16 737 70 763
rect 16 703 24 737
rect 58 703 70 737
rect 16 677 70 703
rect 100 737 170 763
rect 100 703 118 737
rect 152 703 170 737
rect 100 677 170 703
rect 200 737 270 763
rect 200 703 218 737
rect 252 703 270 737
rect 200 677 270 703
rect 300 737 370 763
rect 300 703 318 737
rect 352 703 370 737
rect 300 677 370 703
rect 400 677 470 763
rect 500 677 570 763
rect 600 737 670 763
rect 600 703 618 737
rect 652 703 670 737
rect 600 677 670 703
rect 700 737 770 763
rect 700 703 718 737
rect 752 703 770 737
rect 700 677 770 703
rect 800 737 870 763
rect 800 703 818 737
rect 852 703 870 737
rect 800 677 870 703
rect 900 737 954 763
rect 900 703 912 737
rect 946 703 954 737
rect 900 677 954 703
rect 16 537 70 623
rect 100 537 170 623
rect 200 597 270 623
rect 200 563 218 597
rect 252 563 270 597
rect 200 537 270 563
rect 300 597 370 623
rect 300 563 318 597
rect 352 563 370 597
rect 300 537 370 563
rect 400 597 470 623
rect 400 563 418 597
rect 452 563 470 597
rect 400 537 470 563
rect 500 597 554 623
rect 500 563 512 597
rect 546 563 554 597
rect 500 537 554 563
rect 16 397 70 483
rect 100 457 170 483
rect 100 423 118 457
rect 152 423 170 457
rect 100 397 170 423
rect 200 457 254 483
rect 200 423 212 457
rect 246 423 254 457
rect 200 397 254 423
rect 316 457 370 483
rect 316 423 324 457
rect 358 423 370 457
rect 316 397 370 423
rect 400 457 454 483
rect 400 423 412 457
rect 446 423 454 457
rect 400 397 454 423
rect 2916 2227 2970 2253
rect 2916 2193 2924 2227
rect 2958 2193 2970 2227
rect 2916 2167 2970 2193
rect 3000 2227 3070 2253
rect 3000 2193 3018 2227
rect 3052 2193 3070 2227
rect 3000 2167 3070 2193
rect 3100 2227 3170 2253
rect 3100 2193 3118 2227
rect 3152 2193 3170 2227
rect 3100 2167 3170 2193
rect 3200 2227 3270 2253
rect 3200 2193 3218 2227
rect 3252 2193 3270 2227
rect 3200 2167 3270 2193
rect 3300 2227 3370 2253
rect 3300 2193 3318 2227
rect 3352 2193 3370 2227
rect 3300 2167 3370 2193
rect 3400 2227 3470 2253
rect 3400 2193 3418 2227
rect 3452 2193 3470 2227
rect 3400 2167 3470 2193
rect 3500 2227 3554 2253
rect 3500 2193 3512 2227
rect 3546 2193 3554 2227
rect 3500 2167 3554 2193
rect 2516 2087 2570 2113
rect 2516 2053 2524 2087
rect 2558 2053 2570 2087
rect 2516 2027 2570 2053
rect 2600 2087 2670 2113
rect 2600 2053 2618 2087
rect 2652 2053 2670 2087
rect 2600 2027 2670 2053
rect 2700 2087 2770 2113
rect 2700 2053 2718 2087
rect 2752 2053 2770 2087
rect 2700 2027 2770 2053
rect 2800 2087 2870 2113
rect 2800 2053 2818 2087
rect 2852 2053 2870 2087
rect 2800 2027 2870 2053
rect 2900 2087 2970 2113
rect 2900 2053 2918 2087
rect 2952 2053 2970 2087
rect 2900 2027 2970 2053
rect 3000 2027 3070 2113
rect 3100 2027 3170 2113
rect 3200 2087 3270 2113
rect 3200 2053 3218 2087
rect 3252 2053 3270 2087
rect 3200 2027 3270 2053
rect 3300 2087 3354 2113
rect 3300 2053 3312 2087
rect 3346 2053 3354 2087
rect 3300 2027 3354 2053
rect 2516 1947 2570 1973
rect 2516 1913 2524 1947
rect 2558 1913 2570 1947
rect 2516 1887 2570 1913
rect 2600 1947 2670 1973
rect 2600 1913 2618 1947
rect 2652 1913 2670 1947
rect 2600 1887 2670 1913
rect 2700 1887 2770 1973
rect 2800 1887 2870 1973
rect 2900 1947 2970 1973
rect 2900 1913 2918 1947
rect 2952 1913 2970 1947
rect 2900 1887 2970 1913
rect 3000 1947 3054 1973
rect 3000 1913 3012 1947
rect 3046 1913 3054 1947
rect 3000 1887 3054 1913
rect 3616 2227 3670 2253
rect 3616 2193 3624 2227
rect 3658 2193 3670 2227
rect 3616 2167 3670 2193
rect 3700 2227 3770 2253
rect 3700 2193 3718 2227
rect 3752 2193 3770 2227
rect 3700 2167 3770 2193
rect 3800 2227 3870 2253
rect 3800 2193 3818 2227
rect 3852 2193 3870 2227
rect 3800 2167 3870 2193
rect 3900 2167 3970 2253
rect 4000 2227 4070 2253
rect 4000 2193 4018 2227
rect 4052 2193 4070 2227
rect 4000 2167 4070 2193
rect 4100 2227 4170 2253
rect 4100 2193 4118 2227
rect 4152 2193 4170 2227
rect 4100 2167 4170 2193
rect 4200 2227 4254 2253
rect 4200 2193 4212 2227
rect 4246 2193 4254 2227
rect 4200 2167 4254 2193
rect 3416 2087 3470 2113
rect 3416 2053 3424 2087
rect 3458 2053 3470 2087
rect 3416 2027 3470 2053
rect 3500 2087 3570 2113
rect 3500 2053 3518 2087
rect 3552 2053 3570 2087
rect 3500 2027 3570 2053
rect 3600 2087 3654 2113
rect 3600 2053 3612 2087
rect 3646 2053 3654 2087
rect 3600 2027 3654 2053
rect 3716 2087 3770 2113
rect 3716 2053 3724 2087
rect 3758 2053 3770 2087
rect 3716 2027 3770 2053
rect 3800 2087 3870 2113
rect 3800 2053 3818 2087
rect 3852 2053 3870 2087
rect 3800 2027 3870 2053
rect 3900 2087 3954 2113
rect 3900 2053 3912 2087
rect 3946 2053 3954 2087
rect 3900 2027 3954 2053
rect 3116 1947 3170 1973
rect 3116 1913 3124 1947
rect 3158 1913 3170 1947
rect 3116 1887 3170 1913
rect 3200 1947 3270 1973
rect 3200 1913 3218 1947
rect 3252 1913 3270 1947
rect 3200 1887 3270 1913
rect 3300 1887 3370 1973
rect 3400 1887 3470 1973
rect 3500 1947 3570 1973
rect 3500 1913 3518 1947
rect 3552 1913 3570 1947
rect 3500 1887 3570 1913
rect 3600 1947 3670 1973
rect 3600 1913 3618 1947
rect 3652 1913 3670 1947
rect 3600 1887 3670 1913
rect 3700 1947 3770 1973
rect 3700 1913 3718 1947
rect 3752 1913 3770 1947
rect 3700 1887 3770 1913
rect 3800 1947 3854 1973
rect 3800 1913 3812 1947
rect 3846 1913 3854 1947
rect 3800 1887 3854 1913
rect 1916 1807 1970 1833
rect 1916 1773 1924 1807
rect 1958 1773 1970 1807
rect 1916 1747 1970 1773
rect 2000 1807 2070 1833
rect 2000 1773 2018 1807
rect 2052 1773 2070 1807
rect 2000 1747 2070 1773
rect 2100 1747 2170 1833
rect 2200 1807 2270 1833
rect 2200 1773 2218 1807
rect 2252 1773 2270 1807
rect 2200 1747 2270 1773
rect 2300 1807 2370 1833
rect 2300 1773 2318 1807
rect 2352 1773 2370 1807
rect 2300 1747 2370 1773
rect 2400 1747 2470 1833
rect 2500 1747 2570 1833
rect 2600 1807 2670 1833
rect 2600 1773 2618 1807
rect 2652 1773 2670 1807
rect 2600 1747 2670 1773
rect 2700 1807 2770 1833
rect 2700 1773 2718 1807
rect 2752 1773 2770 1807
rect 2700 1747 2770 1773
rect 2800 1807 2870 1833
rect 2800 1773 2818 1807
rect 2852 1773 2870 1807
rect 2800 1747 2870 1773
rect 2900 1807 2970 1833
rect 2900 1773 2918 1807
rect 2952 1773 2970 1807
rect 2900 1747 2970 1773
rect 3000 1807 3070 1833
rect 3000 1773 3018 1807
rect 3052 1773 3070 1807
rect 3000 1747 3070 1773
rect 3100 1747 3170 1833
rect 3200 1747 3270 1833
rect 3300 1807 3370 1833
rect 3300 1773 3318 1807
rect 3352 1773 3370 1807
rect 3300 1747 3370 1773
rect 3400 1807 3454 1833
rect 3400 1773 3412 1807
rect 3446 1773 3454 1807
rect 3400 1747 3454 1773
rect 1816 1667 1870 1693
rect 1816 1633 1824 1667
rect 1858 1633 1870 1667
rect 1816 1607 1870 1633
rect 1900 1667 1954 1693
rect 1900 1633 1912 1667
rect 1946 1633 1954 1667
rect 1900 1607 1954 1633
rect 2016 1667 2070 1693
rect 2016 1633 2024 1667
rect 2058 1633 2070 1667
rect 2016 1607 2070 1633
rect 2100 1667 2170 1693
rect 2100 1633 2118 1667
rect 2152 1633 2170 1667
rect 2100 1607 2170 1633
rect 2200 1667 2270 1693
rect 2200 1633 2218 1667
rect 2252 1633 2270 1667
rect 2200 1607 2270 1633
rect 2300 1607 2370 1693
rect 2400 1607 2470 1693
rect 2500 1667 2570 1693
rect 2500 1633 2518 1667
rect 2552 1633 2570 1667
rect 2500 1607 2570 1633
rect 2600 1667 2654 1693
rect 2600 1633 2612 1667
rect 2646 1633 2654 1667
rect 2600 1607 2654 1633
rect 2716 1667 2770 1693
rect 2716 1633 2724 1667
rect 2758 1633 2770 1667
rect 2716 1607 2770 1633
rect 2800 1667 2870 1693
rect 2800 1633 2818 1667
rect 2852 1633 2870 1667
rect 2800 1607 2870 1633
rect 2900 1667 2970 1693
rect 2900 1633 2918 1667
rect 2952 1633 2970 1667
rect 2900 1607 2970 1633
rect 3000 1667 3070 1693
rect 3000 1633 3018 1667
rect 3052 1633 3070 1667
rect 3000 1607 3070 1633
rect 3100 1667 3170 1693
rect 3100 1633 3118 1667
rect 3152 1633 3170 1667
rect 3100 1607 3170 1633
rect 3200 1607 3270 1693
rect 3300 1667 3370 1693
rect 3300 1633 3318 1667
rect 3352 1633 3370 1667
rect 3300 1607 3370 1633
rect 3400 1667 3454 1693
rect 3400 1633 3412 1667
rect 3446 1633 3454 1667
rect 3400 1607 3454 1633
rect 3516 1807 3570 1833
rect 3516 1773 3524 1807
rect 3558 1773 3570 1807
rect 3516 1747 3570 1773
rect 3600 1807 3654 1833
rect 3600 1773 3612 1807
rect 3646 1773 3654 1807
rect 3600 1747 3654 1773
rect 4316 2227 4370 2253
rect 4316 2193 4324 2227
rect 4358 2193 4370 2227
rect 4316 2167 4370 2193
rect 4400 2227 4454 2253
rect 4400 2193 4412 2227
rect 4446 2193 4454 2227
rect 4400 2167 4454 2193
rect 4016 2087 4070 2113
rect 4016 2053 4024 2087
rect 4058 2053 4070 2087
rect 4016 2027 4070 2053
rect 4100 2087 4170 2113
rect 4100 2053 4118 2087
rect 4152 2053 4170 2087
rect 4100 2027 4170 2053
rect 4200 2027 4270 2113
rect 4300 2087 4370 2113
rect 4300 2053 4318 2087
rect 4352 2053 4370 2087
rect 4300 2027 4370 2053
rect 4400 2087 4454 2113
rect 4400 2053 4412 2087
rect 4446 2053 4454 2087
rect 4400 2027 4454 2053
rect 3916 1947 3970 1973
rect 3916 1913 3924 1947
rect 3958 1913 3970 1947
rect 3916 1887 3970 1913
rect 4000 1947 4070 1973
rect 4000 1913 4018 1947
rect 4052 1913 4070 1947
rect 4000 1887 4070 1913
rect 4100 1947 4170 1973
rect 4100 1913 4118 1947
rect 4152 1913 4170 1947
rect 4100 1887 4170 1913
rect 4200 1947 4270 1973
rect 4200 1913 4218 1947
rect 4252 1913 4270 1947
rect 4200 1887 4270 1913
rect 4300 1947 4370 1973
rect 4300 1913 4318 1947
rect 4352 1913 4370 1947
rect 4300 1887 4370 1913
rect 4400 1947 4454 1973
rect 4400 1913 4412 1947
rect 4446 1913 4454 1947
rect 4400 1887 4454 1913
rect 3716 1807 3770 1833
rect 3716 1773 3724 1807
rect 3758 1773 3770 1807
rect 3716 1747 3770 1773
rect 3800 1807 3870 1833
rect 3800 1773 3818 1807
rect 3852 1773 3870 1807
rect 3800 1747 3870 1773
rect 3900 1807 3954 1833
rect 3900 1773 3912 1807
rect 3946 1773 3954 1807
rect 3900 1747 3954 1773
rect 3516 1667 3570 1693
rect 3516 1633 3524 1667
rect 3558 1633 3570 1667
rect 3516 1607 3570 1633
rect 3600 1667 3670 1693
rect 3600 1633 3618 1667
rect 3652 1633 3670 1667
rect 3600 1607 3670 1633
rect 3700 1667 3754 1693
rect 3700 1633 3712 1667
rect 3746 1633 3754 1667
rect 3700 1607 3754 1633
rect 5516 2367 5570 2393
rect 5516 2333 5524 2367
rect 5558 2333 5570 2367
rect 5516 2307 5570 2333
rect 5600 2367 5670 2393
rect 5600 2333 5618 2367
rect 5652 2333 5670 2367
rect 5600 2307 5670 2333
rect 5700 2367 5770 2393
rect 5700 2333 5718 2367
rect 5752 2333 5770 2367
rect 5700 2307 5770 2333
rect 5800 2307 5870 2393
rect 5900 2367 5970 2393
rect 5900 2333 5918 2367
rect 5952 2333 5970 2367
rect 5900 2307 5970 2333
rect 6000 2367 6070 2393
rect 6000 2333 6018 2367
rect 6052 2333 6070 2367
rect 6000 2307 6070 2333
rect 6100 2307 6170 2393
rect 6200 2307 6270 2393
rect 6300 2367 6370 2393
rect 6300 2333 6318 2367
rect 6352 2333 6370 2367
rect 6300 2307 6370 2333
rect 6400 2367 6454 2393
rect 6400 2333 6412 2367
rect 6446 2333 6454 2367
rect 6400 2307 6454 2333
rect 6512 2382 6570 2393
rect 6512 2348 6524 2382
rect 6558 2348 6570 2382
rect 6512 2307 6570 2348
rect 6600 2367 6670 2393
rect 6600 2333 6618 2367
rect 6652 2333 6670 2367
rect 6600 2307 6670 2333
rect 6700 2352 6758 2393
rect 6700 2318 6712 2352
rect 6746 2318 6758 2352
rect 6700 2307 6758 2318
rect 6820 2367 6880 2393
rect 6820 2333 6828 2367
rect 6862 2333 6880 2367
rect 6820 2307 6880 2333
rect 6910 2367 6980 2393
rect 6910 2333 6928 2367
rect 6962 2333 6980 2367
rect 6910 2307 6980 2333
rect 7010 2367 7080 2393
rect 7010 2333 7028 2367
rect 7062 2333 7080 2367
rect 7010 2307 7080 2333
rect 7110 2367 7180 2393
rect 7110 2333 7128 2367
rect 7162 2333 7180 2367
rect 7110 2307 7180 2333
rect 7210 2367 7280 2393
rect 7210 2333 7228 2367
rect 7262 2333 7280 2367
rect 7210 2307 7280 2333
rect 7310 2367 7380 2393
rect 7310 2333 7328 2367
rect 7362 2333 7380 2367
rect 7310 2307 7380 2333
rect 7410 2367 7470 2393
rect 7410 2333 7428 2367
rect 7462 2333 7470 2367
rect 7410 2307 7470 2333
rect 4516 2227 4570 2253
rect 4516 2193 4524 2227
rect 4558 2193 4570 2227
rect 4516 2167 4570 2193
rect 4600 2227 4670 2253
rect 4600 2193 4618 2227
rect 4652 2193 4670 2227
rect 4600 2167 4670 2193
rect 4700 2227 4770 2253
rect 4700 2193 4718 2227
rect 4752 2193 4770 2227
rect 4700 2167 4770 2193
rect 4800 2167 4870 2253
rect 4900 2227 4970 2253
rect 4900 2193 4918 2227
rect 4952 2193 4970 2227
rect 4900 2167 4970 2193
rect 5000 2227 5070 2253
rect 5000 2193 5018 2227
rect 5052 2193 5070 2227
rect 5000 2167 5070 2193
rect 5100 2227 5170 2253
rect 5100 2193 5118 2227
rect 5152 2193 5170 2227
rect 5100 2167 5170 2193
rect 5200 2167 5270 2253
rect 5300 2167 5370 2253
rect 5400 2227 5470 2253
rect 5400 2193 5418 2227
rect 5452 2193 5470 2227
rect 5400 2167 5470 2193
rect 5500 2227 5570 2253
rect 5500 2193 5518 2227
rect 5552 2193 5570 2227
rect 5500 2167 5570 2193
rect 5600 2227 5670 2253
rect 5600 2193 5618 2227
rect 5652 2193 5670 2227
rect 5600 2167 5670 2193
rect 5700 2227 5770 2253
rect 5700 2193 5718 2227
rect 5752 2193 5770 2227
rect 5700 2167 5770 2193
rect 5800 2227 5870 2253
rect 5800 2193 5818 2227
rect 5852 2193 5870 2227
rect 5800 2167 5870 2193
rect 5900 2227 5970 2253
rect 5900 2193 5918 2227
rect 5952 2193 5970 2227
rect 5900 2167 5970 2193
rect 6000 2167 6070 2253
rect 6100 2167 6170 2253
rect 6200 2227 6270 2253
rect 6200 2193 6218 2227
rect 6252 2193 6270 2227
rect 6200 2167 6270 2193
rect 6300 2227 6370 2253
rect 6300 2193 6318 2227
rect 6352 2193 6370 2227
rect 6300 2167 6370 2193
rect 6400 2227 6454 2253
rect 6400 2193 6412 2227
rect 6446 2193 6454 2227
rect 6400 2167 6454 2193
rect 6512 2242 6570 2253
rect 6512 2208 6524 2242
rect 6558 2208 6570 2242
rect 6512 2167 6570 2208
rect 6600 2227 6670 2253
rect 6600 2193 6618 2227
rect 6652 2193 6670 2227
rect 6600 2167 6670 2193
rect 6700 2212 6758 2253
rect 6700 2178 6712 2212
rect 6746 2178 6758 2212
rect 6700 2167 6758 2178
rect 6820 2227 6880 2253
rect 6820 2193 6828 2227
rect 6862 2193 6880 2227
rect 6820 2167 6880 2193
rect 6910 2227 6980 2253
rect 6910 2193 6928 2227
rect 6962 2193 6980 2227
rect 6910 2167 6980 2193
rect 7010 2227 7080 2253
rect 7010 2193 7028 2227
rect 7062 2193 7080 2227
rect 7010 2167 7080 2193
rect 7110 2227 7180 2253
rect 7110 2193 7128 2227
rect 7162 2193 7180 2227
rect 7110 2167 7180 2193
rect 7210 2227 7280 2253
rect 7210 2193 7228 2227
rect 7262 2193 7280 2227
rect 7210 2167 7280 2193
rect 7310 2227 7380 2253
rect 7310 2193 7328 2227
rect 7362 2193 7380 2227
rect 7310 2167 7380 2193
rect 7410 2227 7470 2253
rect 7410 2193 7428 2227
rect 7462 2193 7470 2227
rect 7410 2167 7470 2193
rect 4516 2087 4570 2113
rect 4516 2053 4524 2087
rect 4558 2053 4570 2087
rect 4516 2027 4570 2053
rect 4600 2087 4670 2113
rect 4600 2053 4618 2087
rect 4652 2053 4670 2087
rect 4600 2027 4670 2053
rect 4700 2087 4770 2113
rect 4700 2053 4718 2087
rect 4752 2053 4770 2087
rect 4700 2027 4770 2053
rect 4800 2027 4870 2113
rect 4900 2087 4970 2113
rect 4900 2053 4918 2087
rect 4952 2053 4970 2087
rect 4900 2027 4970 2053
rect 5000 2087 5070 2113
rect 5000 2053 5018 2087
rect 5052 2053 5070 2087
rect 5000 2027 5070 2053
rect 5100 2027 5170 2113
rect 5200 2027 5270 2113
rect 5300 2087 5370 2113
rect 5300 2053 5318 2087
rect 5352 2053 5370 2087
rect 5300 2027 5370 2053
rect 5400 2087 5470 2113
rect 5400 2053 5418 2087
rect 5452 2053 5470 2087
rect 5400 2027 5470 2053
rect 5500 2087 5570 2113
rect 5500 2053 5518 2087
rect 5552 2053 5570 2087
rect 5500 2027 5570 2053
rect 5600 2087 5670 2113
rect 5600 2053 5618 2087
rect 5652 2053 5670 2087
rect 5600 2027 5670 2053
rect 5700 2027 5770 2113
rect 5800 2087 5870 2113
rect 5800 2053 5818 2087
rect 5852 2053 5870 2087
rect 5800 2027 5870 2053
rect 5900 2087 5970 2113
rect 5900 2053 5918 2087
rect 5952 2053 5970 2087
rect 5900 2027 5970 2053
rect 6000 2027 6070 2113
rect 6100 2087 6170 2113
rect 6100 2053 6118 2087
rect 6152 2053 6170 2087
rect 6100 2027 6170 2053
rect 6200 2087 6270 2113
rect 6200 2053 6218 2087
rect 6252 2053 6270 2087
rect 6200 2027 6270 2053
rect 6300 2087 6370 2113
rect 6300 2053 6318 2087
rect 6352 2053 6370 2087
rect 6300 2027 6370 2053
rect 6400 2027 6454 2113
rect 6512 2102 6570 2113
rect 6512 2068 6524 2102
rect 6558 2068 6570 2102
rect 6512 2027 6570 2068
rect 6600 2087 6670 2113
rect 6600 2053 6618 2087
rect 6652 2053 6670 2087
rect 6600 2027 6670 2053
rect 6700 2072 6758 2113
rect 6700 2038 6712 2072
rect 6746 2038 6758 2072
rect 6700 2027 6758 2038
rect 6820 2087 6880 2113
rect 6820 2053 6828 2087
rect 6862 2053 6880 2087
rect 6820 2027 6880 2053
rect 6910 2087 6980 2113
rect 6910 2053 6928 2087
rect 6962 2053 6980 2087
rect 6910 2027 6980 2053
rect 7010 2087 7080 2113
rect 7010 2053 7028 2087
rect 7062 2053 7080 2087
rect 7010 2027 7080 2053
rect 7110 2087 7180 2113
rect 7110 2053 7128 2087
rect 7162 2053 7180 2087
rect 7110 2027 7180 2053
rect 7210 2087 7280 2113
rect 7210 2053 7228 2087
rect 7262 2053 7280 2087
rect 7210 2027 7280 2053
rect 7310 2087 7380 2113
rect 7310 2053 7328 2087
rect 7362 2053 7380 2087
rect 7310 2027 7380 2053
rect 7410 2087 7470 2113
rect 7410 2053 7428 2087
rect 7462 2053 7470 2087
rect 7410 2027 7470 2053
rect 4516 1947 4570 1973
rect 4516 1913 4524 1947
rect 4558 1913 4570 1947
rect 4516 1887 4570 1913
rect 4600 1947 4670 1973
rect 4600 1913 4618 1947
rect 4652 1913 4670 1947
rect 4600 1887 4670 1913
rect 4700 1947 4770 1973
rect 4700 1913 4718 1947
rect 4752 1913 4770 1947
rect 4700 1887 4770 1913
rect 4800 1947 4870 1973
rect 4800 1913 4818 1947
rect 4852 1913 4870 1947
rect 4800 1887 4870 1913
rect 4900 1947 4954 1973
rect 4900 1913 4912 1947
rect 4946 1913 4954 1947
rect 4900 1887 4954 1913
rect 4016 1807 4070 1833
rect 4016 1773 4024 1807
rect 4058 1773 4070 1807
rect 4016 1747 4070 1773
rect 4100 1807 4170 1833
rect 4100 1773 4118 1807
rect 4152 1773 4170 1807
rect 4100 1747 4170 1773
rect 4200 1747 4270 1833
rect 4300 1807 4370 1833
rect 4300 1773 4318 1807
rect 4352 1773 4370 1807
rect 4300 1747 4370 1773
rect 4400 1807 4470 1833
rect 4400 1773 4418 1807
rect 4452 1773 4470 1807
rect 4400 1747 4470 1773
rect 4500 1807 4570 1833
rect 4500 1773 4518 1807
rect 4552 1773 4570 1807
rect 4500 1747 4570 1773
rect 4600 1747 4670 1833
rect 4700 1807 4770 1833
rect 4700 1773 4718 1807
rect 4752 1773 4770 1807
rect 4700 1747 4770 1773
rect 4800 1807 4854 1833
rect 4800 1773 4812 1807
rect 4846 1773 4854 1807
rect 4800 1747 4854 1773
rect 3816 1667 3870 1693
rect 3816 1633 3824 1667
rect 3858 1633 3870 1667
rect 3816 1607 3870 1633
rect 3900 1667 3970 1693
rect 3900 1633 3918 1667
rect 3952 1633 3970 1667
rect 3900 1607 3970 1633
rect 4000 1667 4070 1693
rect 4000 1633 4018 1667
rect 4052 1633 4070 1667
rect 4000 1607 4070 1633
rect 4100 1607 4170 1693
rect 4200 1667 4270 1693
rect 4200 1633 4218 1667
rect 4252 1633 4270 1667
rect 4200 1607 4270 1633
rect 4300 1667 4370 1693
rect 4300 1633 4318 1667
rect 4352 1633 4370 1667
rect 4300 1607 4370 1633
rect 4400 1667 4454 1693
rect 4400 1633 4412 1667
rect 4446 1633 4454 1667
rect 4400 1607 4454 1633
rect 1716 1527 1770 1553
rect 1716 1493 1724 1527
rect 1758 1493 1770 1527
rect 1716 1467 1770 1493
rect 1800 1527 1870 1553
rect 1800 1493 1818 1527
rect 1852 1493 1870 1527
rect 1800 1467 1870 1493
rect 1900 1527 1970 1553
rect 1900 1493 1918 1527
rect 1952 1493 1970 1527
rect 1900 1467 1970 1493
rect 2000 1527 2070 1553
rect 2000 1493 2018 1527
rect 2052 1493 2070 1527
rect 2000 1467 2070 1493
rect 2100 1527 2170 1553
rect 2100 1493 2118 1527
rect 2152 1493 2170 1527
rect 2100 1467 2170 1493
rect 2200 1527 2270 1553
rect 2200 1493 2218 1527
rect 2252 1493 2270 1527
rect 2200 1467 2270 1493
rect 2300 1467 2370 1553
rect 2400 1527 2470 1553
rect 2400 1493 2418 1527
rect 2452 1493 2470 1527
rect 2400 1467 2470 1493
rect 2500 1527 2570 1553
rect 2500 1493 2518 1527
rect 2552 1493 2570 1527
rect 2500 1467 2570 1493
rect 2600 1527 2670 1553
rect 2600 1493 2618 1527
rect 2652 1493 2670 1527
rect 2600 1467 2670 1493
rect 2700 1527 2770 1553
rect 2700 1493 2718 1527
rect 2752 1493 2770 1527
rect 2700 1467 2770 1493
rect 2800 1467 2870 1553
rect 2900 1467 2970 1553
rect 3000 1527 3070 1553
rect 3000 1493 3018 1527
rect 3052 1493 3070 1527
rect 3000 1467 3070 1493
rect 3100 1527 3170 1553
rect 3100 1493 3118 1527
rect 3152 1493 3170 1527
rect 3100 1467 3170 1493
rect 3200 1527 3270 1553
rect 3200 1493 3218 1527
rect 3252 1493 3270 1527
rect 3200 1467 3270 1493
rect 3300 1527 3370 1553
rect 3300 1493 3318 1527
rect 3352 1493 3370 1527
rect 3300 1467 3370 1493
rect 3400 1527 3470 1553
rect 3400 1493 3418 1527
rect 3452 1493 3470 1527
rect 3400 1467 3470 1493
rect 3500 1467 3570 1553
rect 3600 1527 3670 1553
rect 3600 1493 3618 1527
rect 3652 1493 3670 1527
rect 3600 1467 3670 1493
rect 3700 1527 3770 1553
rect 3700 1493 3718 1527
rect 3752 1493 3770 1527
rect 3700 1467 3770 1493
rect 3800 1467 3870 1553
rect 3900 1527 3970 1553
rect 3900 1493 3918 1527
rect 3952 1493 3970 1527
rect 3900 1467 3970 1493
rect 4000 1527 4070 1553
rect 4000 1493 4018 1527
rect 4052 1493 4070 1527
rect 4000 1467 4070 1493
rect 4100 1527 4154 1553
rect 4100 1493 4112 1527
rect 4146 1493 4154 1527
rect 4100 1467 4154 1493
rect 1616 1387 1670 1413
rect 1616 1353 1624 1387
rect 1658 1353 1670 1387
rect 1616 1327 1670 1353
rect 1700 1387 1754 1413
rect 1700 1353 1712 1387
rect 1746 1353 1754 1387
rect 1700 1327 1754 1353
rect 1816 1387 1870 1413
rect 1816 1353 1824 1387
rect 1858 1353 1870 1387
rect 1816 1327 1870 1353
rect 1900 1387 1970 1413
rect 1900 1353 1918 1387
rect 1952 1353 1970 1387
rect 1900 1327 1970 1353
rect 2000 1327 2070 1413
rect 2100 1327 2170 1413
rect 2200 1387 2270 1413
rect 2200 1353 2218 1387
rect 2252 1353 2270 1387
rect 2200 1327 2270 1353
rect 2300 1387 2370 1413
rect 2300 1353 2318 1387
rect 2352 1353 2370 1387
rect 2300 1327 2370 1353
rect 2400 1387 2470 1413
rect 2400 1353 2418 1387
rect 2452 1353 2470 1387
rect 2400 1327 2470 1353
rect 2500 1327 2570 1413
rect 2600 1327 2670 1413
rect 2700 1387 2770 1413
rect 2700 1353 2718 1387
rect 2752 1353 2770 1387
rect 2700 1327 2770 1353
rect 2800 1387 2870 1413
rect 2800 1353 2818 1387
rect 2852 1353 2870 1387
rect 2800 1327 2870 1353
rect 2900 1387 2954 1413
rect 2900 1353 2912 1387
rect 2946 1353 2954 1387
rect 2900 1327 2954 1353
rect 1316 1157 1370 1183
rect 1316 1123 1324 1157
rect 1358 1123 1370 1157
rect 1316 1097 1370 1123
rect 1400 1157 1470 1183
rect 1400 1123 1418 1157
rect 1452 1123 1470 1157
rect 1400 1097 1470 1123
rect 1500 1097 1570 1183
rect 1600 1157 1670 1183
rect 1600 1123 1618 1157
rect 1652 1123 1670 1157
rect 1600 1097 1670 1123
rect 1700 1157 1770 1183
rect 1700 1123 1718 1157
rect 1752 1123 1770 1157
rect 1700 1097 1770 1123
rect 1800 1157 1870 1183
rect 1800 1123 1818 1157
rect 1852 1123 1870 1157
rect 1800 1097 1870 1123
rect 1900 1157 1970 1183
rect 1900 1123 1918 1157
rect 1952 1123 1970 1157
rect 1900 1097 1970 1123
rect 2000 1097 2070 1183
rect 2100 1157 2170 1183
rect 2100 1123 2118 1157
rect 2152 1123 2170 1157
rect 2100 1097 2170 1123
rect 2200 1157 2270 1183
rect 2200 1123 2218 1157
rect 2252 1123 2270 1157
rect 2200 1097 2270 1123
rect 2300 1157 2370 1183
rect 2300 1123 2318 1157
rect 2352 1123 2370 1157
rect 2300 1097 2370 1123
rect 2400 1157 2470 1183
rect 2400 1123 2418 1157
rect 2452 1123 2470 1157
rect 2400 1097 2470 1123
rect 2500 1157 2554 1183
rect 2500 1123 2512 1157
rect 2546 1123 2554 1157
rect 2500 1097 2554 1123
rect 1216 1017 1270 1043
rect 1216 983 1224 1017
rect 1258 983 1270 1017
rect 1216 957 1270 983
rect 1300 1017 1370 1043
rect 1300 983 1318 1017
rect 1352 983 1370 1017
rect 1300 957 1370 983
rect 1400 957 1470 1043
rect 1500 1017 1570 1043
rect 1500 983 1518 1017
rect 1552 983 1570 1017
rect 1500 957 1570 983
rect 1600 1017 1670 1043
rect 1600 983 1618 1017
rect 1652 983 1670 1017
rect 1600 957 1670 983
rect 1700 957 1770 1043
rect 1800 1017 1870 1043
rect 1800 983 1818 1017
rect 1852 983 1870 1017
rect 1800 957 1870 983
rect 1900 1017 1970 1043
rect 1900 983 1918 1017
rect 1952 983 1970 1017
rect 1900 957 1970 983
rect 2000 1017 2070 1043
rect 2000 983 2018 1017
rect 2052 983 2070 1017
rect 2000 957 2070 983
rect 2100 1017 2154 1043
rect 2100 983 2112 1017
rect 2146 983 2154 1017
rect 2100 957 2154 983
rect 1116 877 1170 903
rect 1116 843 1124 877
rect 1158 843 1170 877
rect 1116 817 1170 843
rect 1200 877 1270 903
rect 1200 843 1218 877
rect 1252 843 1270 877
rect 1200 817 1270 843
rect 1300 877 1370 903
rect 1300 843 1318 877
rect 1352 843 1370 877
rect 1300 817 1370 843
rect 1400 817 1470 903
rect 1500 877 1570 903
rect 1500 843 1518 877
rect 1552 843 1570 877
rect 1500 817 1570 843
rect 1600 877 1670 903
rect 1600 843 1618 877
rect 1652 843 1670 877
rect 1600 817 1670 843
rect 1700 877 1754 903
rect 1700 843 1712 877
rect 1746 843 1754 877
rect 1700 817 1754 843
rect 2216 1017 2270 1043
rect 2216 983 2224 1017
rect 2258 983 2270 1017
rect 2216 957 2270 983
rect 2300 1017 2370 1043
rect 2300 983 2318 1017
rect 2352 983 2370 1017
rect 2300 957 2370 983
rect 2400 1017 2454 1043
rect 2400 983 2412 1017
rect 2446 983 2454 1017
rect 2400 957 2454 983
rect 2616 1157 2670 1183
rect 2616 1123 2624 1157
rect 2658 1123 2670 1157
rect 2616 1097 2670 1123
rect 2700 1157 2754 1183
rect 2700 1123 2712 1157
rect 2746 1123 2754 1157
rect 2700 1097 2754 1123
rect 3016 1387 3070 1413
rect 3016 1353 3024 1387
rect 3058 1353 3070 1387
rect 3016 1327 3070 1353
rect 3100 1387 3170 1413
rect 3100 1353 3118 1387
rect 3152 1353 3170 1387
rect 3100 1327 3170 1353
rect 3200 1327 3270 1413
rect 3300 1387 3370 1413
rect 3300 1353 3318 1387
rect 3352 1353 3370 1387
rect 3300 1327 3370 1353
rect 3400 1387 3470 1413
rect 3400 1353 3418 1387
rect 3452 1353 3470 1387
rect 3400 1327 3470 1353
rect 3500 1387 3554 1413
rect 3500 1353 3512 1387
rect 3546 1353 3554 1387
rect 3500 1327 3554 1353
rect 3616 1387 3670 1413
rect 3616 1353 3624 1387
rect 3658 1353 3670 1387
rect 3616 1327 3670 1353
rect 3700 1387 3770 1413
rect 3700 1353 3718 1387
rect 3752 1353 3770 1387
rect 3700 1327 3770 1353
rect 3800 1387 3854 1413
rect 3800 1353 3812 1387
rect 3846 1353 3854 1387
rect 3800 1327 3854 1353
rect 4216 1527 4270 1553
rect 4216 1493 4224 1527
rect 4258 1493 4270 1527
rect 4216 1467 4270 1493
rect 4300 1527 4370 1553
rect 4300 1493 4318 1527
rect 4352 1493 4370 1527
rect 4300 1467 4370 1493
rect 4400 1527 4454 1553
rect 4400 1493 4412 1527
rect 4446 1493 4454 1527
rect 4400 1467 4454 1493
rect 5016 1947 5070 1973
rect 5016 1913 5024 1947
rect 5058 1913 5070 1947
rect 5016 1887 5070 1913
rect 5100 1947 5154 1973
rect 5100 1913 5112 1947
rect 5146 1913 5154 1947
rect 5100 1887 5154 1913
rect 5216 1947 5270 1973
rect 5216 1913 5224 1947
rect 5258 1913 5270 1947
rect 5216 1887 5270 1913
rect 5300 1947 5354 1973
rect 5300 1913 5312 1947
rect 5346 1913 5354 1947
rect 5300 1887 5354 1913
rect 5416 1947 5470 1973
rect 5416 1913 5424 1947
rect 5458 1913 5470 1947
rect 5416 1887 5470 1913
rect 5500 1947 5570 1973
rect 5500 1913 5518 1947
rect 5552 1913 5570 1947
rect 5500 1887 5570 1913
rect 5600 1947 5670 1973
rect 5600 1913 5618 1947
rect 5652 1913 5670 1947
rect 5600 1887 5670 1913
rect 5700 1947 5754 1973
rect 5700 1913 5712 1947
rect 5746 1913 5754 1947
rect 5700 1887 5754 1913
rect 5816 1947 5870 1973
rect 5816 1913 5824 1947
rect 5858 1913 5870 1947
rect 5816 1887 5870 1913
rect 5900 1947 5970 1973
rect 5900 1913 5918 1947
rect 5952 1913 5970 1947
rect 5900 1887 5970 1913
rect 6000 1947 6054 1973
rect 6000 1913 6012 1947
rect 6046 1913 6054 1947
rect 6000 1887 6054 1913
rect 6116 1947 6170 1973
rect 6116 1913 6124 1947
rect 6158 1913 6170 1947
rect 6116 1887 6170 1913
rect 6200 1947 6270 1973
rect 6200 1913 6218 1947
rect 6252 1913 6270 1947
rect 6200 1887 6270 1913
rect 6300 1887 6370 1973
rect 6400 1887 6454 1973
rect 6512 1962 6570 1973
rect 6512 1928 6524 1962
rect 6558 1928 6570 1962
rect 6512 1887 6570 1928
rect 6600 1947 6670 1973
rect 6600 1913 6618 1947
rect 6652 1913 6670 1947
rect 6600 1887 6670 1913
rect 6700 1932 6758 1973
rect 6700 1898 6712 1932
rect 6746 1898 6758 1932
rect 6700 1887 6758 1898
rect 6820 1947 6880 1973
rect 6820 1913 6828 1947
rect 6862 1913 6880 1947
rect 6820 1887 6880 1913
rect 6910 1947 6980 1973
rect 6910 1913 6928 1947
rect 6962 1913 6980 1947
rect 6910 1887 6980 1913
rect 7010 1947 7080 1973
rect 7010 1913 7028 1947
rect 7062 1913 7080 1947
rect 7010 1887 7080 1913
rect 7110 1947 7180 1973
rect 7110 1913 7128 1947
rect 7162 1913 7180 1947
rect 7110 1887 7180 1913
rect 7210 1947 7280 1973
rect 7210 1913 7228 1947
rect 7262 1913 7280 1947
rect 7210 1887 7280 1913
rect 7310 1947 7380 1973
rect 7310 1913 7328 1947
rect 7362 1913 7380 1947
rect 7310 1887 7380 1913
rect 7410 1947 7470 1973
rect 7410 1913 7428 1947
rect 7462 1913 7470 1947
rect 7410 1887 7470 1913
rect 4916 1807 4970 1833
rect 4916 1773 4924 1807
rect 4958 1773 4970 1807
rect 4916 1747 4970 1773
rect 5000 1807 5070 1833
rect 5000 1773 5018 1807
rect 5052 1773 5070 1807
rect 5000 1747 5070 1773
rect 5100 1747 5170 1833
rect 5200 1747 5270 1833
rect 5300 1807 5370 1833
rect 5300 1773 5318 1807
rect 5352 1773 5370 1807
rect 5300 1747 5370 1773
rect 5400 1807 5470 1833
rect 5400 1773 5418 1807
rect 5452 1773 5470 1807
rect 5400 1747 5470 1773
rect 5500 1807 5570 1833
rect 5500 1773 5518 1807
rect 5552 1773 5570 1807
rect 5500 1747 5570 1773
rect 5600 1747 5670 1833
rect 5700 1807 5770 1833
rect 5700 1773 5718 1807
rect 5752 1773 5770 1807
rect 5700 1747 5770 1773
rect 5800 1807 5870 1833
rect 5800 1773 5818 1807
rect 5852 1773 5870 1807
rect 5800 1747 5870 1773
rect 5900 1747 5970 1833
rect 6000 1747 6070 1833
rect 6100 1807 6170 1833
rect 6100 1773 6118 1807
rect 6152 1773 6170 1807
rect 6100 1747 6170 1773
rect 6200 1807 6270 1833
rect 6200 1773 6218 1807
rect 6252 1773 6270 1807
rect 6200 1747 6270 1773
rect 6300 1807 6370 1833
rect 6300 1773 6318 1807
rect 6352 1773 6370 1807
rect 6300 1747 6370 1773
rect 6400 1747 6454 1833
rect 6512 1822 6570 1833
rect 6512 1788 6524 1822
rect 6558 1788 6570 1822
rect 6512 1747 6570 1788
rect 6600 1807 6670 1833
rect 6600 1773 6618 1807
rect 6652 1773 6670 1807
rect 6600 1747 6670 1773
rect 6700 1792 6758 1833
rect 6700 1758 6712 1792
rect 6746 1758 6758 1792
rect 6700 1747 6758 1758
rect 6820 1807 6880 1833
rect 6820 1773 6828 1807
rect 6862 1773 6880 1807
rect 6820 1747 6880 1773
rect 6910 1807 6980 1833
rect 6910 1773 6928 1807
rect 6962 1773 6980 1807
rect 6910 1747 6980 1773
rect 7010 1807 7080 1833
rect 7010 1773 7028 1807
rect 7062 1773 7080 1807
rect 7010 1747 7080 1773
rect 7110 1807 7180 1833
rect 7110 1773 7128 1807
rect 7162 1773 7180 1807
rect 7110 1747 7180 1773
rect 7210 1807 7280 1833
rect 7210 1773 7228 1807
rect 7262 1773 7280 1807
rect 7210 1747 7280 1773
rect 7310 1807 7380 1833
rect 7310 1773 7328 1807
rect 7362 1773 7380 1807
rect 7310 1747 7380 1773
rect 7410 1807 7470 1833
rect 7410 1773 7428 1807
rect 7462 1773 7470 1807
rect 7410 1747 7470 1773
rect 4516 1667 4570 1693
rect 4516 1633 4524 1667
rect 4558 1633 4570 1667
rect 4516 1607 4570 1633
rect 4600 1667 4670 1693
rect 4600 1633 4618 1667
rect 4652 1633 4670 1667
rect 4600 1607 4670 1633
rect 4700 1607 4770 1693
rect 4800 1667 4870 1693
rect 4800 1633 4818 1667
rect 4852 1633 4870 1667
rect 4800 1607 4870 1633
rect 4900 1667 4970 1693
rect 4900 1633 4918 1667
rect 4952 1633 4970 1667
rect 4900 1607 4970 1633
rect 5000 1667 5070 1693
rect 5000 1633 5018 1667
rect 5052 1633 5070 1667
rect 5000 1607 5070 1633
rect 5100 1667 5170 1693
rect 5100 1633 5118 1667
rect 5152 1633 5170 1667
rect 5100 1607 5170 1633
rect 5200 1667 5270 1693
rect 5200 1633 5218 1667
rect 5252 1633 5270 1667
rect 5200 1607 5270 1633
rect 5300 1667 5354 1693
rect 5300 1633 5312 1667
rect 5346 1633 5354 1667
rect 5300 1607 5354 1633
rect 4516 1527 4570 1553
rect 4516 1493 4524 1527
rect 4558 1493 4570 1527
rect 4516 1467 4570 1493
rect 4600 1527 4670 1553
rect 4600 1493 4618 1527
rect 4652 1493 4670 1527
rect 4600 1467 4670 1493
rect 4700 1467 4770 1553
rect 4800 1467 4870 1553
rect 4900 1527 4970 1553
rect 4900 1493 4918 1527
rect 4952 1493 4970 1527
rect 4900 1467 4970 1493
rect 5000 1527 5054 1553
rect 5000 1493 5012 1527
rect 5046 1493 5054 1527
rect 5000 1467 5054 1493
rect 3916 1387 3970 1413
rect 3916 1353 3924 1387
rect 3958 1353 3970 1387
rect 3916 1327 3970 1353
rect 4000 1387 4070 1413
rect 4000 1353 4018 1387
rect 4052 1353 4070 1387
rect 4000 1327 4070 1353
rect 4100 1387 4170 1413
rect 4100 1353 4118 1387
rect 4152 1353 4170 1387
rect 4100 1327 4170 1353
rect 4200 1387 4270 1413
rect 4200 1353 4218 1387
rect 4252 1353 4270 1387
rect 4200 1327 4270 1353
rect 4300 1327 4370 1413
rect 4400 1327 4470 1413
rect 4500 1327 4570 1413
rect 4600 1327 4670 1413
rect 4700 1387 4770 1413
rect 4700 1353 4718 1387
rect 4752 1353 4770 1387
rect 4700 1327 4770 1353
rect 4800 1387 4854 1413
rect 4800 1353 4812 1387
rect 4846 1353 4854 1387
rect 4800 1327 4854 1353
rect 2816 1157 2870 1183
rect 2816 1123 2824 1157
rect 2858 1123 2870 1157
rect 2816 1097 2870 1123
rect 2900 1157 2970 1183
rect 2900 1123 2918 1157
rect 2952 1123 2970 1157
rect 2900 1097 2970 1123
rect 3000 1097 3070 1183
rect 3100 1157 3170 1183
rect 3100 1123 3118 1157
rect 3152 1123 3170 1157
rect 3100 1097 3170 1123
rect 3200 1157 3270 1183
rect 3200 1123 3218 1157
rect 3252 1123 3270 1157
rect 3200 1097 3270 1123
rect 3300 1157 3370 1183
rect 3300 1123 3318 1157
rect 3352 1123 3370 1157
rect 3300 1097 3370 1123
rect 3400 1097 3470 1183
rect 3500 1097 3570 1183
rect 3600 1157 3670 1183
rect 3600 1123 3618 1157
rect 3652 1123 3670 1157
rect 3600 1097 3670 1123
rect 3700 1157 3770 1183
rect 3700 1123 3718 1157
rect 3752 1123 3770 1157
rect 3700 1097 3770 1123
rect 3800 1097 3870 1183
rect 3900 1097 3970 1183
rect 4000 1097 4070 1183
rect 4100 1157 4170 1183
rect 4100 1123 4118 1157
rect 4152 1123 4170 1157
rect 4100 1097 4170 1123
rect 4200 1157 4254 1183
rect 4200 1123 4212 1157
rect 4246 1123 4254 1157
rect 4200 1097 4254 1123
rect 2516 1017 2570 1043
rect 2516 983 2524 1017
rect 2558 983 2570 1017
rect 2516 957 2570 983
rect 2600 1017 2670 1043
rect 2600 983 2618 1017
rect 2652 983 2670 1017
rect 2600 957 2670 983
rect 2700 1017 2770 1043
rect 2700 983 2718 1017
rect 2752 983 2770 1017
rect 2700 957 2770 983
rect 2800 1017 2870 1043
rect 2800 983 2818 1017
rect 2852 983 2870 1017
rect 2800 957 2870 983
rect 2900 957 2970 1043
rect 3000 1017 3070 1043
rect 3000 983 3018 1017
rect 3052 983 3070 1017
rect 3000 957 3070 983
rect 3100 1017 3170 1043
rect 3100 983 3118 1017
rect 3152 983 3170 1017
rect 3100 957 3170 983
rect 3200 1017 3270 1043
rect 3200 983 3218 1017
rect 3252 983 3270 1017
rect 3200 957 3270 983
rect 3300 957 3370 1043
rect 3400 1017 3470 1043
rect 3400 983 3418 1017
rect 3452 983 3470 1017
rect 3400 957 3470 983
rect 3500 1017 3570 1043
rect 3500 983 3518 1017
rect 3552 983 3570 1017
rect 3500 957 3570 983
rect 3600 957 3670 1043
rect 3700 1017 3770 1043
rect 3700 983 3718 1017
rect 3752 983 3770 1017
rect 3700 957 3770 983
rect 3800 1017 3870 1043
rect 3800 983 3818 1017
rect 3852 983 3870 1017
rect 3800 957 3870 983
rect 3900 957 3970 1043
rect 4000 957 4070 1043
rect 4100 1017 4170 1043
rect 4100 983 4118 1017
rect 4152 983 4170 1017
rect 4100 957 4170 983
rect 4200 1017 4254 1043
rect 4200 983 4212 1017
rect 4246 983 4254 1017
rect 4200 957 4254 983
rect 4916 1387 4970 1413
rect 4916 1353 4924 1387
rect 4958 1353 4970 1387
rect 4916 1327 4970 1353
rect 5000 1387 5054 1413
rect 5000 1353 5012 1387
rect 5046 1353 5054 1387
rect 5000 1327 5054 1353
rect 5116 1527 5170 1553
rect 5116 1493 5124 1527
rect 5158 1493 5170 1527
rect 5116 1467 5170 1493
rect 5200 1527 5254 1553
rect 5200 1493 5212 1527
rect 5246 1493 5254 1527
rect 5200 1467 5254 1493
rect 5416 1667 5470 1693
rect 5416 1633 5424 1667
rect 5458 1633 5470 1667
rect 5416 1607 5470 1633
rect 5500 1667 5570 1693
rect 5500 1633 5518 1667
rect 5552 1633 5570 1667
rect 5500 1607 5570 1633
rect 5600 1667 5670 1693
rect 5600 1633 5618 1667
rect 5652 1633 5670 1667
rect 5600 1607 5670 1633
rect 5700 1667 5754 1693
rect 5700 1633 5712 1667
rect 5746 1633 5754 1667
rect 5700 1607 5754 1633
rect 5316 1527 5370 1553
rect 5316 1493 5324 1527
rect 5358 1493 5370 1527
rect 5316 1467 5370 1493
rect 5400 1527 5454 1553
rect 5400 1493 5412 1527
rect 5446 1493 5454 1527
rect 5400 1467 5454 1493
rect 5516 1527 5570 1553
rect 5516 1493 5524 1527
rect 5558 1493 5570 1527
rect 5516 1467 5570 1493
rect 5600 1527 5670 1553
rect 5600 1493 5618 1527
rect 5652 1493 5670 1527
rect 5600 1467 5670 1493
rect 5700 1527 5754 1553
rect 5700 1493 5712 1527
rect 5746 1493 5754 1527
rect 5700 1467 5754 1493
rect 5816 1667 5870 1693
rect 5816 1633 5824 1667
rect 5858 1633 5870 1667
rect 5816 1607 5870 1633
rect 5900 1667 5954 1693
rect 5900 1633 5912 1667
rect 5946 1633 5954 1667
rect 5900 1607 5954 1633
rect 5816 1527 5870 1553
rect 5816 1493 5824 1527
rect 5858 1493 5870 1527
rect 5816 1467 5870 1493
rect 5900 1527 5954 1553
rect 5900 1493 5912 1527
rect 5946 1493 5954 1527
rect 5900 1467 5954 1493
rect 6016 1667 6070 1693
rect 6016 1633 6024 1667
rect 6058 1633 6070 1667
rect 6016 1607 6070 1633
rect 6100 1667 6170 1693
rect 6100 1633 6118 1667
rect 6152 1633 6170 1667
rect 6100 1607 6170 1633
rect 6200 1667 6270 1693
rect 6200 1633 6218 1667
rect 6252 1633 6270 1667
rect 6200 1607 6270 1633
rect 6300 1607 6370 1693
rect 6400 1607 6454 1693
rect 6512 1682 6570 1693
rect 6512 1648 6524 1682
rect 6558 1648 6570 1682
rect 6512 1607 6570 1648
rect 6600 1667 6670 1693
rect 6600 1633 6618 1667
rect 6652 1633 6670 1667
rect 6600 1607 6670 1633
rect 6700 1652 6758 1693
rect 6700 1618 6712 1652
rect 6746 1618 6758 1652
rect 6700 1607 6758 1618
rect 6820 1667 6880 1693
rect 6820 1633 6828 1667
rect 6862 1633 6880 1667
rect 6820 1607 6880 1633
rect 6910 1667 6980 1693
rect 6910 1633 6928 1667
rect 6962 1633 6980 1667
rect 6910 1607 6980 1633
rect 7010 1667 7080 1693
rect 7010 1633 7028 1667
rect 7062 1633 7080 1667
rect 7010 1607 7080 1633
rect 7110 1667 7180 1693
rect 7110 1633 7128 1667
rect 7162 1633 7180 1667
rect 7110 1607 7180 1633
rect 7210 1667 7280 1693
rect 7210 1633 7228 1667
rect 7262 1633 7280 1667
rect 7210 1607 7280 1633
rect 7310 1667 7380 1693
rect 7310 1633 7328 1667
rect 7362 1633 7380 1667
rect 7310 1607 7380 1633
rect 7410 1667 7470 1693
rect 7410 1633 7428 1667
rect 7462 1633 7470 1667
rect 7410 1607 7470 1633
rect 6016 1527 6070 1553
rect 6016 1493 6024 1527
rect 6058 1493 6070 1527
rect 6016 1467 6070 1493
rect 6100 1527 6170 1553
rect 6100 1493 6118 1527
rect 6152 1493 6170 1527
rect 6100 1467 6170 1493
rect 6200 1527 6254 1553
rect 6200 1493 6212 1527
rect 6246 1493 6254 1527
rect 6200 1467 6254 1493
rect 5116 1387 5170 1413
rect 5116 1353 5124 1387
rect 5158 1353 5170 1387
rect 5116 1327 5170 1353
rect 5200 1387 5270 1413
rect 5200 1353 5218 1387
rect 5252 1353 5270 1387
rect 5200 1327 5270 1353
rect 5300 1327 5370 1413
rect 5400 1327 5470 1413
rect 5500 1387 5570 1413
rect 5500 1353 5518 1387
rect 5552 1353 5570 1387
rect 5500 1327 5570 1353
rect 5600 1387 5670 1413
rect 5600 1353 5618 1387
rect 5652 1353 5670 1387
rect 5600 1327 5670 1353
rect 5700 1387 5770 1413
rect 5700 1353 5718 1387
rect 5752 1353 5770 1387
rect 5700 1327 5770 1353
rect 5800 1327 5870 1413
rect 5900 1387 5970 1413
rect 5900 1353 5918 1387
rect 5952 1353 5970 1387
rect 5900 1327 5970 1353
rect 6000 1387 6070 1413
rect 6000 1353 6018 1387
rect 6052 1353 6070 1387
rect 6000 1327 6070 1353
rect 6100 1387 6154 1413
rect 6100 1353 6112 1387
rect 6146 1353 6154 1387
rect 6100 1327 6154 1353
rect 4316 1157 4370 1183
rect 4316 1123 4324 1157
rect 4358 1123 4370 1157
rect 4316 1097 4370 1123
rect 4400 1157 4470 1183
rect 4400 1123 4418 1157
rect 4452 1123 4470 1157
rect 4400 1097 4470 1123
rect 4500 1097 4570 1183
rect 4600 1097 4670 1183
rect 4700 1157 4770 1183
rect 4700 1123 4718 1157
rect 4752 1123 4770 1157
rect 4700 1097 4770 1123
rect 4800 1157 4870 1183
rect 4800 1123 4818 1157
rect 4852 1123 4870 1157
rect 4800 1097 4870 1123
rect 4900 1157 4970 1183
rect 4900 1123 4918 1157
rect 4952 1123 4970 1157
rect 4900 1097 4970 1123
rect 5000 1097 5070 1183
rect 5100 1157 5170 1183
rect 5100 1123 5118 1157
rect 5152 1123 5170 1157
rect 5100 1097 5170 1123
rect 5200 1157 5270 1183
rect 5200 1123 5218 1157
rect 5252 1123 5270 1157
rect 5200 1097 5270 1123
rect 5300 1157 5370 1183
rect 5300 1123 5318 1157
rect 5352 1123 5370 1157
rect 5300 1097 5370 1123
rect 5400 1157 5454 1183
rect 5400 1123 5412 1157
rect 5446 1123 5454 1157
rect 5400 1097 5454 1123
rect 4316 1017 4370 1043
rect 4316 983 4324 1017
rect 4358 983 4370 1017
rect 4316 957 4370 983
rect 4400 1017 4470 1043
rect 4400 983 4418 1017
rect 4452 983 4470 1017
rect 4400 957 4470 983
rect 4500 1017 4570 1043
rect 4500 983 4518 1017
rect 4552 983 4570 1017
rect 4500 957 4570 983
rect 4600 1017 4670 1043
rect 4600 983 4618 1017
rect 4652 983 4670 1017
rect 4600 957 4670 983
rect 4700 1017 4770 1043
rect 4700 983 4718 1017
rect 4752 983 4770 1017
rect 4700 957 4770 983
rect 4800 1017 4854 1043
rect 4800 983 4812 1017
rect 4846 983 4854 1017
rect 4800 957 4854 983
rect 1816 877 1870 903
rect 1816 843 1824 877
rect 1858 843 1870 877
rect 1816 817 1870 843
rect 1900 877 1970 903
rect 1900 843 1918 877
rect 1952 843 1970 877
rect 1900 817 1970 843
rect 2000 877 2070 903
rect 2000 843 2018 877
rect 2052 843 2070 877
rect 2000 817 2070 843
rect 2100 877 2170 903
rect 2100 843 2118 877
rect 2152 843 2170 877
rect 2100 817 2170 843
rect 2200 877 2270 903
rect 2200 843 2218 877
rect 2252 843 2270 877
rect 2200 817 2270 843
rect 2300 877 2370 903
rect 2300 843 2318 877
rect 2352 843 2370 877
rect 2300 817 2370 843
rect 2400 877 2470 903
rect 2400 843 2418 877
rect 2452 843 2470 877
rect 2400 817 2470 843
rect 2500 877 2570 903
rect 2500 843 2518 877
rect 2552 843 2570 877
rect 2500 817 2570 843
rect 2600 817 2670 903
rect 2700 817 2770 903
rect 2800 877 2870 903
rect 2800 843 2818 877
rect 2852 843 2870 877
rect 2800 817 2870 843
rect 2900 877 2970 903
rect 2900 843 2918 877
rect 2952 843 2970 877
rect 2900 817 2970 843
rect 3000 817 3070 903
rect 3100 877 3170 903
rect 3100 843 3118 877
rect 3152 843 3170 877
rect 3100 817 3170 843
rect 3200 877 3270 903
rect 3200 843 3218 877
rect 3252 843 3270 877
rect 3200 817 3270 843
rect 3300 877 3370 903
rect 3300 843 3318 877
rect 3352 843 3370 877
rect 3300 817 3370 843
rect 3400 817 3470 903
rect 3500 817 3570 903
rect 3600 817 3670 903
rect 3700 817 3770 903
rect 3800 817 3870 903
rect 3900 877 3970 903
rect 3900 843 3918 877
rect 3952 843 3970 877
rect 3900 817 3970 843
rect 4000 877 4070 903
rect 4000 843 4018 877
rect 4052 843 4070 877
rect 4000 817 4070 843
rect 4100 877 4170 903
rect 4100 843 4118 877
rect 4152 843 4170 877
rect 4100 817 4170 843
rect 4200 877 4270 903
rect 4200 843 4218 877
rect 4252 843 4270 877
rect 4200 817 4270 843
rect 4300 877 4354 903
rect 4300 843 4312 877
rect 4346 843 4354 877
rect 4300 817 4354 843
rect 1016 737 1070 763
rect 1016 703 1024 737
rect 1058 703 1070 737
rect 1016 677 1070 703
rect 1100 737 1170 763
rect 1100 703 1118 737
rect 1152 703 1170 737
rect 1100 677 1170 703
rect 1200 677 1270 763
rect 1300 677 1370 763
rect 1400 677 1470 763
rect 1500 677 1570 763
rect 1600 677 1670 763
rect 1700 677 1770 763
rect 1800 737 1870 763
rect 1800 703 1818 737
rect 1852 703 1870 737
rect 1800 677 1870 703
rect 1900 737 1970 763
rect 1900 703 1918 737
rect 1952 703 1970 737
rect 1900 677 1970 703
rect 2000 737 2054 763
rect 2000 703 2012 737
rect 2046 703 2054 737
rect 2000 677 2054 703
rect 616 597 670 623
rect 616 563 624 597
rect 658 563 670 597
rect 616 537 670 563
rect 700 597 770 623
rect 700 563 718 597
rect 752 563 770 597
rect 700 537 770 563
rect 800 537 870 623
rect 900 597 970 623
rect 900 563 918 597
rect 952 563 970 597
rect 900 537 970 563
rect 1000 597 1054 623
rect 1000 563 1012 597
rect 1046 563 1054 597
rect 1000 537 1054 563
rect 2116 737 2170 763
rect 2116 703 2124 737
rect 2158 703 2170 737
rect 2116 677 2170 703
rect 2200 737 2254 763
rect 2200 703 2212 737
rect 2246 703 2254 737
rect 2200 677 2254 703
rect 4416 877 4470 903
rect 4416 843 4424 877
rect 4458 843 4470 877
rect 4416 817 4470 843
rect 4500 877 4554 903
rect 4500 843 4512 877
rect 4546 843 4554 877
rect 4500 817 4554 843
rect 2316 737 2370 763
rect 2316 703 2324 737
rect 2358 703 2370 737
rect 2316 677 2370 703
rect 2400 737 2470 763
rect 2400 703 2418 737
rect 2452 703 2470 737
rect 2400 677 2470 703
rect 2500 677 2570 763
rect 2600 677 2670 763
rect 2700 737 2770 763
rect 2700 703 2718 737
rect 2752 703 2770 737
rect 2700 677 2770 703
rect 2800 737 2870 763
rect 2800 703 2818 737
rect 2852 703 2870 737
rect 2800 677 2870 703
rect 2900 737 2970 763
rect 2900 703 2918 737
rect 2952 703 2970 737
rect 2900 677 2970 703
rect 3000 737 3070 763
rect 3000 703 3018 737
rect 3052 703 3070 737
rect 3000 677 3070 703
rect 3100 737 3170 763
rect 3100 703 3118 737
rect 3152 703 3170 737
rect 3100 677 3170 703
rect 3200 737 3270 763
rect 3200 703 3218 737
rect 3252 703 3270 737
rect 3200 677 3270 703
rect 3300 677 3370 763
rect 3400 677 3470 763
rect 3500 737 3570 763
rect 3500 703 3518 737
rect 3552 703 3570 737
rect 3500 677 3570 703
rect 3600 737 3670 763
rect 3600 703 3618 737
rect 3652 703 3670 737
rect 3600 677 3670 703
rect 3700 677 3770 763
rect 3800 677 3870 763
rect 3900 737 3970 763
rect 3900 703 3918 737
rect 3952 703 3970 737
rect 3900 677 3970 703
rect 4000 737 4070 763
rect 4000 703 4018 737
rect 4052 703 4070 737
rect 4000 677 4070 703
rect 4100 737 4170 763
rect 4100 703 4118 737
rect 4152 703 4170 737
rect 4100 677 4170 703
rect 4200 677 4270 763
rect 4300 737 4370 763
rect 4300 703 4318 737
rect 4352 703 4370 737
rect 4300 677 4370 703
rect 4400 737 4454 763
rect 4400 703 4412 737
rect 4446 703 4454 737
rect 4400 677 4454 703
rect 1116 597 1170 623
rect 1116 563 1124 597
rect 1158 563 1170 597
rect 1116 537 1170 563
rect 1200 597 1270 623
rect 1200 563 1218 597
rect 1252 563 1270 597
rect 1200 537 1270 563
rect 1300 537 1370 623
rect 1400 537 1470 623
rect 1500 597 1570 623
rect 1500 563 1518 597
rect 1552 563 1570 597
rect 1500 537 1570 563
rect 1600 597 1670 623
rect 1600 563 1618 597
rect 1652 563 1670 597
rect 1600 537 1670 563
rect 1700 537 1770 623
rect 1800 597 1870 623
rect 1800 563 1818 597
rect 1852 563 1870 597
rect 1800 537 1870 563
rect 1900 597 1970 623
rect 1900 563 1918 597
rect 1952 563 1970 597
rect 1900 537 1970 563
rect 2000 597 2070 623
rect 2000 563 2018 597
rect 2052 563 2070 597
rect 2000 537 2070 563
rect 2100 597 2170 623
rect 2100 563 2118 597
rect 2152 563 2170 597
rect 2100 537 2170 563
rect 2200 537 2270 623
rect 2300 537 2370 623
rect 2400 537 2470 623
rect 2500 597 2570 623
rect 2500 563 2518 597
rect 2552 563 2570 597
rect 2500 537 2570 563
rect 2600 597 2670 623
rect 2600 563 2618 597
rect 2652 563 2670 597
rect 2600 537 2670 563
rect 2700 597 2770 623
rect 2700 563 2718 597
rect 2752 563 2770 597
rect 2700 537 2770 563
rect 2800 537 2870 623
rect 2900 537 2970 623
rect 3000 537 3070 623
rect 3100 597 3170 623
rect 3100 563 3118 597
rect 3152 563 3170 597
rect 3100 537 3170 563
rect 3200 597 3270 623
rect 3200 563 3218 597
rect 3252 563 3270 597
rect 3200 537 3270 563
rect 3300 537 3370 623
rect 3400 537 3470 623
rect 3500 597 3570 623
rect 3500 563 3518 597
rect 3552 563 3570 597
rect 3500 537 3570 563
rect 3600 597 3670 623
rect 3600 563 3618 597
rect 3652 563 3670 597
rect 3600 537 3670 563
rect 3700 597 3754 623
rect 3700 563 3712 597
rect 3746 563 3754 597
rect 3700 537 3754 563
rect 516 457 570 483
rect 516 423 524 457
rect 558 423 570 457
rect 516 397 570 423
rect 600 457 670 483
rect 600 423 618 457
rect 652 423 670 457
rect 600 397 670 423
rect 700 457 770 483
rect 700 423 718 457
rect 752 423 770 457
rect 700 397 770 423
rect 800 457 870 483
rect 800 423 818 457
rect 852 423 870 457
rect 800 397 870 423
rect 900 457 970 483
rect 900 423 918 457
rect 952 423 970 457
rect 900 397 970 423
rect 1000 457 1070 483
rect 1000 423 1018 457
rect 1052 423 1070 457
rect 1000 397 1070 423
rect 1100 397 1170 483
rect 1200 457 1270 483
rect 1200 423 1218 457
rect 1252 423 1270 457
rect 1200 397 1270 423
rect 1300 457 1370 483
rect 1300 423 1318 457
rect 1352 423 1370 457
rect 1300 397 1370 423
rect 1400 457 1454 483
rect 1400 423 1412 457
rect 1446 423 1454 457
rect 1400 397 1454 423
rect 16 257 70 343
rect 100 317 170 343
rect 100 283 118 317
rect 152 283 170 317
rect 100 257 170 283
rect 200 317 270 343
rect 200 283 218 317
rect 252 283 270 317
rect 200 257 270 283
rect 300 257 370 343
rect 400 317 470 343
rect 400 283 418 317
rect 452 283 470 317
rect 400 257 470 283
rect 500 317 570 343
rect 500 283 518 317
rect 552 283 570 317
rect 500 257 570 283
rect 600 317 654 343
rect 600 283 612 317
rect 646 283 654 317
rect 600 257 654 283
rect 1516 457 1570 483
rect 1516 423 1524 457
rect 1558 423 1570 457
rect 1516 397 1570 423
rect 1600 457 1670 483
rect 1600 423 1618 457
rect 1652 423 1670 457
rect 1600 397 1670 423
rect 1700 397 1770 483
rect 1800 457 1870 483
rect 1800 423 1818 457
rect 1852 423 1870 457
rect 1800 397 1870 423
rect 1900 457 1970 483
rect 1900 423 1918 457
rect 1952 423 1970 457
rect 1900 397 1970 423
rect 2000 457 2070 483
rect 2000 423 2018 457
rect 2052 423 2070 457
rect 2000 397 2070 423
rect 2100 397 2170 483
rect 2200 457 2270 483
rect 2200 423 2218 457
rect 2252 423 2270 457
rect 2200 397 2270 423
rect 2300 457 2370 483
rect 2300 423 2318 457
rect 2352 423 2370 457
rect 2300 397 2370 423
rect 2400 397 2470 483
rect 2500 397 2570 483
rect 2600 397 2670 483
rect 2700 457 2770 483
rect 2700 423 2718 457
rect 2752 423 2770 457
rect 2700 397 2770 423
rect 2800 457 2870 483
rect 2800 423 2818 457
rect 2852 423 2870 457
rect 2800 397 2870 423
rect 2900 457 2970 483
rect 2900 423 2918 457
rect 2952 423 2970 457
rect 2900 397 2970 423
rect 3000 457 3054 483
rect 3000 423 3012 457
rect 3046 423 3054 457
rect 3000 397 3054 423
rect 716 317 770 343
rect 716 283 724 317
rect 758 283 770 317
rect 716 257 770 283
rect 800 317 870 343
rect 800 283 818 317
rect 852 283 870 317
rect 800 257 870 283
rect 900 317 970 343
rect 900 283 918 317
rect 952 283 970 317
rect 900 257 970 283
rect 1000 257 1070 343
rect 1100 257 1170 343
rect 1200 257 1270 343
rect 1300 257 1370 343
rect 1400 317 1470 343
rect 1400 283 1418 317
rect 1452 283 1470 317
rect 1400 257 1470 283
rect 1500 317 1554 343
rect 1500 283 1512 317
rect 1546 283 1554 317
rect 1500 257 1554 283
rect 16 177 70 203
rect 16 143 24 177
rect 58 143 70 177
rect 16 117 70 143
rect 100 177 170 203
rect 100 143 118 177
rect 152 143 170 177
rect 100 117 170 143
rect 200 177 270 203
rect 200 143 218 177
rect 252 143 270 177
rect 200 117 270 143
rect 300 177 370 203
rect 300 143 318 177
rect 352 143 370 177
rect 300 117 370 143
rect 400 177 470 203
rect 400 143 418 177
rect 452 143 470 177
rect 400 117 470 143
rect 500 117 570 203
rect 600 177 670 203
rect 600 143 618 177
rect 652 143 670 177
rect 600 117 670 143
rect 700 177 770 203
rect 700 143 718 177
rect 752 143 770 177
rect 700 117 770 143
rect 800 177 854 203
rect 800 143 812 177
rect 846 143 854 177
rect 800 117 854 143
rect 1616 317 1670 343
rect 1616 283 1624 317
rect 1658 283 1670 317
rect 1616 257 1670 283
rect 1700 317 1770 343
rect 1700 283 1718 317
rect 1752 283 1770 317
rect 1700 257 1770 283
rect 1800 257 1870 343
rect 1900 257 1970 343
rect 2000 317 2070 343
rect 2000 283 2018 317
rect 2052 283 2070 317
rect 2000 257 2070 283
rect 2100 317 2170 343
rect 2100 283 2118 317
rect 2152 283 2170 317
rect 2100 257 2170 283
rect 2200 317 2254 343
rect 2200 283 2212 317
rect 2246 283 2254 317
rect 2200 257 2254 283
rect 916 177 970 203
rect 916 143 924 177
rect 958 143 970 177
rect 916 117 970 143
rect 1000 177 1070 203
rect 1000 143 1018 177
rect 1052 143 1070 177
rect 1000 117 1070 143
rect 1100 117 1170 203
rect 1200 117 1270 203
rect 1300 177 1370 203
rect 1300 143 1318 177
rect 1352 143 1370 177
rect 1300 117 1370 143
rect 1400 177 1470 203
rect 1400 143 1418 177
rect 1452 143 1470 177
rect 1400 117 1470 143
rect 1500 177 1570 203
rect 1500 143 1518 177
rect 1552 143 1570 177
rect 1500 117 1570 143
rect 1600 117 1670 203
rect 1700 177 1770 203
rect 1700 143 1718 177
rect 1752 143 1770 177
rect 1700 117 1770 143
rect 1800 177 1870 203
rect 1800 143 1818 177
rect 1852 143 1870 177
rect 1800 117 1870 143
rect 1900 177 1954 203
rect 1900 143 1912 177
rect 1946 143 1954 177
rect 1900 117 1954 143
rect 2316 317 2370 343
rect 2316 283 2324 317
rect 2358 283 2370 317
rect 2316 257 2370 283
rect 2400 317 2454 343
rect 2400 283 2412 317
rect 2446 283 2454 317
rect 2400 257 2454 283
rect 2516 317 2570 343
rect 2516 283 2524 317
rect 2558 283 2570 317
rect 2516 257 2570 283
rect 2600 317 2654 343
rect 2600 283 2612 317
rect 2646 283 2654 317
rect 2600 257 2654 283
rect 2716 317 2770 343
rect 2716 283 2724 317
rect 2758 283 2770 317
rect 2716 257 2770 283
rect 2800 317 2854 343
rect 2800 283 2812 317
rect 2846 283 2854 317
rect 2800 257 2854 283
rect 3116 457 3170 483
rect 3116 423 3124 457
rect 3158 423 3170 457
rect 3116 397 3170 423
rect 3200 457 3254 483
rect 3200 423 3212 457
rect 3246 423 3254 457
rect 3200 397 3254 423
rect 3316 457 3370 483
rect 3316 423 3324 457
rect 3358 423 3370 457
rect 3316 397 3370 423
rect 3400 457 3470 483
rect 3400 423 3418 457
rect 3452 423 3470 457
rect 3400 397 3470 423
rect 3500 457 3554 483
rect 3500 423 3512 457
rect 3546 423 3554 457
rect 3500 397 3554 423
rect 2916 317 2970 343
rect 2916 283 2924 317
rect 2958 283 2970 317
rect 2916 257 2970 283
rect 3000 317 3070 343
rect 3000 283 3018 317
rect 3052 283 3070 317
rect 3000 257 3070 283
rect 3100 317 3170 343
rect 3100 283 3118 317
rect 3152 283 3170 317
rect 3100 257 3170 283
rect 3200 257 3270 343
rect 3300 317 3370 343
rect 3300 283 3318 317
rect 3352 283 3370 317
rect 3300 257 3370 283
rect 3400 317 3470 343
rect 3400 283 3418 317
rect 3452 283 3470 317
rect 3400 257 3470 283
rect 3500 317 3554 343
rect 3500 283 3512 317
rect 3546 283 3554 317
rect 3500 257 3554 283
rect 2016 177 2070 203
rect 2016 143 2024 177
rect 2058 143 2070 177
rect 2016 117 2070 143
rect 2100 177 2170 203
rect 2100 143 2118 177
rect 2152 143 2170 177
rect 2100 117 2170 143
rect 2200 177 2270 203
rect 2200 143 2218 177
rect 2252 143 2270 177
rect 2200 117 2270 143
rect 2300 117 2370 203
rect 2400 177 2470 203
rect 2400 143 2418 177
rect 2452 143 2470 177
rect 2400 117 2470 143
rect 2500 177 2570 203
rect 2500 143 2518 177
rect 2552 143 2570 177
rect 2500 117 2570 143
rect 2600 177 2670 203
rect 2600 143 2618 177
rect 2652 143 2670 177
rect 2600 117 2670 143
rect 2700 117 2770 203
rect 2800 117 2870 203
rect 2900 117 2970 203
rect 3000 177 3070 203
rect 3000 143 3018 177
rect 3052 143 3070 177
rect 3000 117 3070 143
rect 3100 177 3170 203
rect 3100 143 3118 177
rect 3152 143 3170 177
rect 3100 117 3170 143
rect 3200 177 3270 203
rect 3200 143 3218 177
rect 3252 143 3270 177
rect 3200 117 3270 143
rect 3300 117 3370 203
rect 3400 177 3470 203
rect 3400 143 3418 177
rect 3452 143 3470 177
rect 3400 117 3470 143
rect 3500 177 3554 203
rect 3500 143 3512 177
rect 3546 143 3554 177
rect 3500 117 3554 143
rect 3616 457 3670 483
rect 3616 423 3624 457
rect 3658 423 3670 457
rect 3616 397 3670 423
rect 3700 457 3754 483
rect 3700 423 3712 457
rect 3746 423 3754 457
rect 3700 397 3754 423
rect 3816 597 3870 623
rect 3816 563 3824 597
rect 3858 563 3870 597
rect 3816 537 3870 563
rect 3900 597 3970 623
rect 3900 563 3918 597
rect 3952 563 3970 597
rect 3900 537 3970 563
rect 4000 597 4054 623
rect 4000 563 4012 597
rect 4046 563 4054 597
rect 4000 537 4054 563
rect 4116 597 4170 623
rect 4116 563 4124 597
rect 4158 563 4170 597
rect 4116 537 4170 563
rect 4200 597 4254 623
rect 4200 563 4212 597
rect 4246 563 4254 597
rect 4200 537 4254 563
rect 4916 1017 4970 1043
rect 4916 983 4924 1017
rect 4958 983 4970 1017
rect 4916 957 4970 983
rect 5000 1017 5054 1043
rect 5000 983 5012 1017
rect 5046 983 5054 1017
rect 5000 957 5054 983
rect 5516 1157 5570 1183
rect 5516 1123 5524 1157
rect 5558 1123 5570 1157
rect 5516 1097 5570 1123
rect 5600 1157 5670 1183
rect 5600 1123 5618 1157
rect 5652 1123 5670 1157
rect 5600 1097 5670 1123
rect 5700 1157 5770 1183
rect 5700 1123 5718 1157
rect 5752 1123 5770 1157
rect 5700 1097 5770 1123
rect 5800 1157 5870 1183
rect 5800 1123 5818 1157
rect 5852 1123 5870 1157
rect 5800 1097 5870 1123
rect 5900 1157 5954 1183
rect 5900 1123 5912 1157
rect 5946 1123 5954 1157
rect 5900 1097 5954 1123
rect 6316 1527 6370 1553
rect 6316 1493 6324 1527
rect 6358 1493 6370 1527
rect 6316 1467 6370 1493
rect 6400 1527 6454 1553
rect 6400 1493 6412 1527
rect 6446 1493 6454 1527
rect 6400 1467 6454 1493
rect 6512 1542 6570 1553
rect 6512 1508 6524 1542
rect 6558 1508 6570 1542
rect 6512 1467 6570 1508
rect 6600 1527 6670 1553
rect 6600 1493 6618 1527
rect 6652 1493 6670 1527
rect 6600 1467 6670 1493
rect 6700 1512 6758 1553
rect 6700 1478 6712 1512
rect 6746 1478 6758 1512
rect 6700 1467 6758 1478
rect 6820 1527 6880 1553
rect 6820 1493 6828 1527
rect 6862 1493 6880 1527
rect 6820 1467 6880 1493
rect 6910 1527 6980 1553
rect 6910 1493 6928 1527
rect 6962 1493 6980 1527
rect 6910 1467 6980 1493
rect 7010 1527 7080 1553
rect 7010 1493 7028 1527
rect 7062 1493 7080 1527
rect 7010 1467 7080 1493
rect 7110 1527 7180 1553
rect 7110 1493 7128 1527
rect 7162 1493 7180 1527
rect 7110 1467 7180 1493
rect 7210 1527 7280 1553
rect 7210 1493 7228 1527
rect 7262 1493 7280 1527
rect 7210 1467 7280 1493
rect 7310 1527 7380 1553
rect 7310 1493 7328 1527
rect 7362 1493 7380 1527
rect 7310 1467 7380 1493
rect 7410 1527 7470 1553
rect 7410 1493 7428 1527
rect 7462 1493 7470 1527
rect 7410 1467 7470 1493
rect 6216 1387 6270 1413
rect 6216 1353 6224 1387
rect 6258 1353 6270 1387
rect 6216 1327 6270 1353
rect 6300 1387 6370 1413
rect 6300 1353 6318 1387
rect 6352 1353 6370 1387
rect 6300 1327 6370 1353
rect 6400 1327 6454 1413
rect 6512 1402 6570 1413
rect 6512 1368 6524 1402
rect 6558 1368 6570 1402
rect 6512 1327 6570 1368
rect 6600 1387 6670 1413
rect 6600 1353 6618 1387
rect 6652 1353 6670 1387
rect 6600 1327 6670 1353
rect 6700 1372 6758 1413
rect 6700 1338 6712 1372
rect 6746 1338 6758 1372
rect 6700 1327 6758 1338
rect 6820 1387 6880 1413
rect 6820 1353 6828 1387
rect 6862 1353 6880 1387
rect 6820 1327 6880 1353
rect 6910 1387 6980 1413
rect 6910 1353 6928 1387
rect 6962 1353 6980 1387
rect 6910 1327 6980 1353
rect 7010 1387 7080 1413
rect 7010 1353 7028 1387
rect 7062 1353 7080 1387
rect 7010 1327 7080 1353
rect 7110 1387 7180 1413
rect 7110 1353 7128 1387
rect 7162 1353 7180 1387
rect 7110 1327 7180 1353
rect 7210 1387 7280 1413
rect 7210 1353 7228 1387
rect 7262 1353 7280 1387
rect 7210 1327 7280 1353
rect 7310 1387 7380 1413
rect 7310 1353 7328 1387
rect 7362 1353 7380 1387
rect 7310 1327 7380 1353
rect 7410 1387 7470 1413
rect 7410 1353 7428 1387
rect 7462 1353 7470 1387
rect 7410 1327 7470 1353
rect 6016 1157 6070 1183
rect 6016 1123 6024 1157
rect 6058 1123 6070 1157
rect 6016 1097 6070 1123
rect 6100 1157 6170 1183
rect 6100 1123 6118 1157
rect 6152 1123 6170 1157
rect 6100 1097 6170 1123
rect 6200 1157 6270 1183
rect 6200 1123 6218 1157
rect 6252 1123 6270 1157
rect 6200 1097 6270 1123
rect 6300 1157 6370 1183
rect 6300 1123 6318 1157
rect 6352 1123 6370 1157
rect 6300 1097 6370 1123
rect 6400 1157 6454 1183
rect 6400 1123 6412 1157
rect 6446 1123 6454 1157
rect 6400 1097 6454 1123
rect 6512 1172 6570 1183
rect 6512 1138 6524 1172
rect 6558 1138 6570 1172
rect 6512 1097 6570 1138
rect 6600 1157 6670 1183
rect 6600 1123 6618 1157
rect 6652 1123 6670 1157
rect 6600 1097 6670 1123
rect 6700 1142 6758 1183
rect 6700 1108 6712 1142
rect 6746 1108 6758 1142
rect 6700 1097 6758 1108
rect 6820 1157 6880 1183
rect 6820 1123 6828 1157
rect 6862 1123 6880 1157
rect 6820 1097 6880 1123
rect 6910 1157 6980 1183
rect 6910 1123 6928 1157
rect 6962 1123 6980 1157
rect 6910 1097 6980 1123
rect 7010 1157 7080 1183
rect 7010 1123 7028 1157
rect 7062 1123 7080 1157
rect 7010 1097 7080 1123
rect 7110 1157 7180 1183
rect 7110 1123 7128 1157
rect 7162 1123 7180 1157
rect 7110 1097 7180 1123
rect 7210 1157 7280 1183
rect 7210 1123 7228 1157
rect 7262 1123 7280 1157
rect 7210 1097 7280 1123
rect 7310 1157 7380 1183
rect 7310 1123 7328 1157
rect 7362 1123 7380 1157
rect 7310 1097 7380 1123
rect 7410 1157 7470 1183
rect 7410 1123 7428 1157
rect 7462 1123 7470 1157
rect 7410 1097 7470 1123
rect 5116 1017 5170 1043
rect 5116 983 5124 1017
rect 5158 983 5170 1017
rect 5116 957 5170 983
rect 5200 1017 5270 1043
rect 5200 983 5218 1017
rect 5252 983 5270 1017
rect 5200 957 5270 983
rect 5300 1017 5370 1043
rect 5300 983 5318 1017
rect 5352 983 5370 1017
rect 5300 957 5370 983
rect 5400 1017 5470 1043
rect 5400 983 5418 1017
rect 5452 983 5470 1017
rect 5400 957 5470 983
rect 5500 1017 5570 1043
rect 5500 983 5518 1017
rect 5552 983 5570 1017
rect 5500 957 5570 983
rect 5600 957 5670 1043
rect 5700 1017 5770 1043
rect 5700 983 5718 1017
rect 5752 983 5770 1017
rect 5700 957 5770 983
rect 5800 1017 5870 1043
rect 5800 983 5818 1017
rect 5852 983 5870 1017
rect 5800 957 5870 983
rect 5900 957 5970 1043
rect 6000 957 6070 1043
rect 6100 1017 6170 1043
rect 6100 983 6118 1017
rect 6152 983 6170 1017
rect 6100 957 6170 983
rect 6200 1017 6254 1043
rect 6200 983 6212 1017
rect 6246 983 6254 1017
rect 6200 957 6254 983
rect 6316 1017 6370 1043
rect 6316 983 6324 1017
rect 6358 983 6370 1017
rect 6316 957 6370 983
rect 6400 1017 6454 1043
rect 6400 983 6412 1017
rect 6446 983 6454 1017
rect 6400 957 6454 983
rect 6512 1032 6570 1043
rect 6512 998 6524 1032
rect 6558 998 6570 1032
rect 6512 957 6570 998
rect 6600 1017 6670 1043
rect 6600 983 6618 1017
rect 6652 983 6670 1017
rect 6600 957 6670 983
rect 6700 1002 6758 1043
rect 6700 968 6712 1002
rect 6746 968 6758 1002
rect 6700 957 6758 968
rect 6820 1017 6880 1043
rect 6820 983 6828 1017
rect 6862 983 6880 1017
rect 6820 957 6880 983
rect 6910 1017 6980 1043
rect 6910 983 6928 1017
rect 6962 983 6980 1017
rect 6910 957 6980 983
rect 7010 1017 7080 1043
rect 7010 983 7028 1017
rect 7062 983 7080 1017
rect 7010 957 7080 983
rect 7110 1017 7180 1043
rect 7110 983 7128 1017
rect 7162 983 7180 1017
rect 7110 957 7180 983
rect 7210 1017 7280 1043
rect 7210 983 7228 1017
rect 7262 983 7280 1017
rect 7210 957 7280 983
rect 7310 1017 7380 1043
rect 7310 983 7328 1017
rect 7362 983 7380 1017
rect 7310 957 7380 983
rect 7410 1017 7470 1043
rect 7410 983 7428 1017
rect 7462 983 7470 1017
rect 7410 957 7470 983
rect 4616 877 4670 903
rect 4616 843 4624 877
rect 4658 843 4670 877
rect 4616 817 4670 843
rect 4700 877 4770 903
rect 4700 843 4718 877
rect 4752 843 4770 877
rect 4700 817 4770 843
rect 4800 877 4870 903
rect 4800 843 4818 877
rect 4852 843 4870 877
rect 4800 817 4870 843
rect 4900 817 4970 903
rect 5000 877 5070 903
rect 5000 843 5018 877
rect 5052 843 5070 877
rect 5000 817 5070 843
rect 5100 877 5170 903
rect 5100 843 5118 877
rect 5152 843 5170 877
rect 5100 817 5170 843
rect 5200 877 5270 903
rect 5200 843 5218 877
rect 5252 843 5270 877
rect 5200 817 5270 843
rect 5300 877 5370 903
rect 5300 843 5318 877
rect 5352 843 5370 877
rect 5300 817 5370 843
rect 5400 817 5470 903
rect 5500 817 5570 903
rect 5600 877 5670 903
rect 5600 843 5618 877
rect 5652 843 5670 877
rect 5600 817 5670 843
rect 5700 877 5770 903
rect 5700 843 5718 877
rect 5752 843 5770 877
rect 5700 817 5770 843
rect 5800 817 5870 903
rect 5900 817 5970 903
rect 6000 877 6070 903
rect 6000 843 6018 877
rect 6052 843 6070 877
rect 6000 817 6070 843
rect 6100 877 6170 903
rect 6100 843 6118 877
rect 6152 843 6170 877
rect 6100 817 6170 843
rect 6200 817 6270 903
rect 6300 817 6370 903
rect 6400 817 6454 903
rect 6512 892 6570 903
rect 6512 858 6524 892
rect 6558 858 6570 892
rect 6512 817 6570 858
rect 6600 877 6670 903
rect 6600 843 6618 877
rect 6652 843 6670 877
rect 6600 817 6670 843
rect 6700 862 6758 903
rect 6700 828 6712 862
rect 6746 828 6758 862
rect 6700 817 6758 828
rect 6820 877 6880 903
rect 6820 843 6828 877
rect 6862 843 6880 877
rect 6820 817 6880 843
rect 6910 877 6980 903
rect 6910 843 6928 877
rect 6962 843 6980 877
rect 6910 817 6980 843
rect 7010 877 7080 903
rect 7010 843 7028 877
rect 7062 843 7080 877
rect 7010 817 7080 843
rect 7110 877 7180 903
rect 7110 843 7128 877
rect 7162 843 7180 877
rect 7110 817 7180 843
rect 7210 877 7280 903
rect 7210 843 7228 877
rect 7262 843 7280 877
rect 7210 817 7280 843
rect 7310 877 7380 903
rect 7310 843 7328 877
rect 7362 843 7380 877
rect 7310 817 7380 843
rect 7410 877 7470 903
rect 7410 843 7428 877
rect 7462 843 7470 877
rect 7410 817 7470 843
rect 4516 737 4570 763
rect 4516 703 4524 737
rect 4558 703 4570 737
rect 4516 677 4570 703
rect 4600 737 4670 763
rect 4600 703 4618 737
rect 4652 703 4670 737
rect 4600 677 4670 703
rect 4700 677 4770 763
rect 4800 737 4870 763
rect 4800 703 4818 737
rect 4852 703 4870 737
rect 4800 677 4870 703
rect 4900 737 4970 763
rect 4900 703 4918 737
rect 4952 703 4970 737
rect 4900 677 4970 703
rect 5000 737 5070 763
rect 5000 703 5018 737
rect 5052 703 5070 737
rect 5000 677 5070 703
rect 5100 677 5170 763
rect 5200 677 5270 763
rect 5300 737 5370 763
rect 5300 703 5318 737
rect 5352 703 5370 737
rect 5300 677 5370 703
rect 5400 737 5470 763
rect 5400 703 5418 737
rect 5452 703 5470 737
rect 5400 677 5470 703
rect 5500 737 5554 763
rect 5500 703 5512 737
rect 5546 703 5554 737
rect 5500 677 5554 703
rect 4316 597 4370 623
rect 4316 563 4324 597
rect 4358 563 4370 597
rect 4316 537 4370 563
rect 4400 597 4470 623
rect 4400 563 4418 597
rect 4452 563 4470 597
rect 4400 537 4470 563
rect 4500 597 4570 623
rect 4500 563 4518 597
rect 4552 563 4570 597
rect 4500 537 4570 563
rect 4600 597 4654 623
rect 4600 563 4612 597
rect 4646 563 4654 597
rect 4600 537 4654 563
rect 4716 597 4770 623
rect 4716 563 4724 597
rect 4758 563 4770 597
rect 4716 537 4770 563
rect 4800 597 4870 623
rect 4800 563 4818 597
rect 4852 563 4870 597
rect 4800 537 4870 563
rect 4900 537 4970 623
rect 5000 597 5070 623
rect 5000 563 5018 597
rect 5052 563 5070 597
rect 5000 537 5070 563
rect 5100 597 5170 623
rect 5100 563 5118 597
rect 5152 563 5170 597
rect 5100 537 5170 563
rect 5200 597 5254 623
rect 5200 563 5212 597
rect 5246 563 5254 597
rect 5200 537 5254 563
rect 5616 737 5670 763
rect 5616 703 5624 737
rect 5658 703 5670 737
rect 5616 677 5670 703
rect 5700 737 5754 763
rect 5700 703 5712 737
rect 5746 703 5754 737
rect 5700 677 5754 703
rect 5816 737 5870 763
rect 5816 703 5824 737
rect 5858 703 5870 737
rect 5816 677 5870 703
rect 5900 737 5970 763
rect 5900 703 5918 737
rect 5952 703 5970 737
rect 5900 677 5970 703
rect 6000 737 6070 763
rect 6000 703 6018 737
rect 6052 703 6070 737
rect 6000 677 6070 703
rect 6100 677 6170 763
rect 6200 737 6270 763
rect 6200 703 6218 737
rect 6252 703 6270 737
rect 6200 677 6270 703
rect 6300 737 6370 763
rect 6300 703 6318 737
rect 6352 703 6370 737
rect 6300 677 6370 703
rect 6400 677 6454 763
rect 6512 752 6570 763
rect 6512 718 6524 752
rect 6558 718 6570 752
rect 6512 677 6570 718
rect 6600 737 6670 763
rect 6600 703 6618 737
rect 6652 703 6670 737
rect 6600 677 6670 703
rect 6700 722 6758 763
rect 6700 688 6712 722
rect 6746 688 6758 722
rect 6700 677 6758 688
rect 6820 737 6880 763
rect 6820 703 6828 737
rect 6862 703 6880 737
rect 6820 677 6880 703
rect 6910 737 6980 763
rect 6910 703 6928 737
rect 6962 703 6980 737
rect 6910 677 6980 703
rect 7010 737 7080 763
rect 7010 703 7028 737
rect 7062 703 7080 737
rect 7010 677 7080 703
rect 7110 737 7180 763
rect 7110 703 7128 737
rect 7162 703 7180 737
rect 7110 677 7180 703
rect 7210 737 7280 763
rect 7210 703 7228 737
rect 7262 703 7280 737
rect 7210 677 7280 703
rect 7310 737 7380 763
rect 7310 703 7328 737
rect 7362 703 7380 737
rect 7310 677 7380 703
rect 7410 737 7470 763
rect 7410 703 7428 737
rect 7462 703 7470 737
rect 7410 677 7470 703
rect 5316 597 5370 623
rect 5316 563 5324 597
rect 5358 563 5370 597
rect 5316 537 5370 563
rect 5400 597 5470 623
rect 5400 563 5418 597
rect 5452 563 5470 597
rect 5400 537 5470 563
rect 5500 537 5570 623
rect 5600 537 5670 623
rect 5700 597 5770 623
rect 5700 563 5718 597
rect 5752 563 5770 597
rect 5700 537 5770 563
rect 5800 597 5870 623
rect 5800 563 5818 597
rect 5852 563 5870 597
rect 5800 537 5870 563
rect 5900 597 5970 623
rect 5900 563 5918 597
rect 5952 563 5970 597
rect 5900 537 5970 563
rect 6000 597 6054 623
rect 6000 563 6012 597
rect 6046 563 6054 597
rect 6000 537 6054 563
rect 3816 457 3870 483
rect 3816 423 3824 457
rect 3858 423 3870 457
rect 3816 397 3870 423
rect 3900 457 3970 483
rect 3900 423 3918 457
rect 3952 423 3970 457
rect 3900 397 3970 423
rect 4000 457 4070 483
rect 4000 423 4018 457
rect 4052 423 4070 457
rect 4000 397 4070 423
rect 4100 397 4170 483
rect 4200 397 4270 483
rect 4300 457 4370 483
rect 4300 423 4318 457
rect 4352 423 4370 457
rect 4300 397 4370 423
rect 4400 457 4470 483
rect 4400 423 4418 457
rect 4452 423 4470 457
rect 4400 397 4470 423
rect 4500 457 4570 483
rect 4500 423 4518 457
rect 4552 423 4570 457
rect 4500 397 4570 423
rect 4600 457 4670 483
rect 4600 423 4618 457
rect 4652 423 4670 457
rect 4600 397 4670 423
rect 4700 397 4770 483
rect 4800 457 4870 483
rect 4800 423 4818 457
rect 4852 423 4870 457
rect 4800 397 4870 423
rect 4900 457 4970 483
rect 4900 423 4918 457
rect 4952 423 4970 457
rect 4900 397 4970 423
rect 5000 457 5070 483
rect 5000 423 5018 457
rect 5052 423 5070 457
rect 5000 397 5070 423
rect 5100 457 5170 483
rect 5100 423 5118 457
rect 5152 423 5170 457
rect 5100 397 5170 423
rect 5200 457 5270 483
rect 5200 423 5218 457
rect 5252 423 5270 457
rect 5200 397 5270 423
rect 5300 457 5370 483
rect 5300 423 5318 457
rect 5352 423 5370 457
rect 5300 397 5370 423
rect 5400 457 5470 483
rect 5400 423 5418 457
rect 5452 423 5470 457
rect 5400 397 5470 423
rect 5500 457 5554 483
rect 5500 423 5512 457
rect 5546 423 5554 457
rect 5500 397 5554 423
rect 6116 597 6170 623
rect 6116 563 6124 597
rect 6158 563 6170 597
rect 6116 537 6170 563
rect 6200 597 6270 623
rect 6200 563 6218 597
rect 6252 563 6270 597
rect 6200 537 6270 563
rect 6300 597 6370 623
rect 6300 563 6318 597
rect 6352 563 6370 597
rect 6300 537 6370 563
rect 6400 597 6454 623
rect 6400 563 6412 597
rect 6446 563 6454 597
rect 6400 537 6454 563
rect 6512 612 6570 623
rect 6512 578 6524 612
rect 6558 578 6570 612
rect 6512 537 6570 578
rect 6600 597 6670 623
rect 6600 563 6618 597
rect 6652 563 6670 597
rect 6600 537 6670 563
rect 6700 582 6758 623
rect 6700 548 6712 582
rect 6746 548 6758 582
rect 6700 537 6758 548
rect 6820 597 6880 623
rect 6820 563 6828 597
rect 6862 563 6880 597
rect 6820 537 6880 563
rect 6910 597 6980 623
rect 6910 563 6928 597
rect 6962 563 6980 597
rect 6910 537 6980 563
rect 7010 597 7080 623
rect 7010 563 7028 597
rect 7062 563 7080 597
rect 7010 537 7080 563
rect 7110 597 7180 623
rect 7110 563 7128 597
rect 7162 563 7180 597
rect 7110 537 7180 563
rect 7210 597 7280 623
rect 7210 563 7228 597
rect 7262 563 7280 597
rect 7210 537 7280 563
rect 7310 597 7380 623
rect 7310 563 7328 597
rect 7362 563 7380 597
rect 7310 537 7380 563
rect 7410 597 7470 623
rect 7410 563 7428 597
rect 7462 563 7470 597
rect 7410 537 7470 563
rect 5616 457 5670 483
rect 5616 423 5624 457
rect 5658 423 5670 457
rect 5616 397 5670 423
rect 5700 457 5770 483
rect 5700 423 5718 457
rect 5752 423 5770 457
rect 5700 397 5770 423
rect 5800 397 5870 483
rect 5900 397 5970 483
rect 6000 457 6070 483
rect 6000 423 6018 457
rect 6052 423 6070 457
rect 6000 397 6070 423
rect 6100 457 6170 483
rect 6100 423 6118 457
rect 6152 423 6170 457
rect 6100 397 6170 423
rect 6200 457 6254 483
rect 6200 423 6212 457
rect 6246 423 6254 457
rect 6200 397 6254 423
rect 3616 317 3670 343
rect 3616 283 3624 317
rect 3658 283 3670 317
rect 3616 257 3670 283
rect 3700 317 3770 343
rect 3700 283 3718 317
rect 3752 283 3770 317
rect 3700 257 3770 283
rect 3800 317 3870 343
rect 3800 283 3818 317
rect 3852 283 3870 317
rect 3800 257 3870 283
rect 3900 317 3970 343
rect 3900 283 3918 317
rect 3952 283 3970 317
rect 3900 257 3970 283
rect 4000 257 4070 343
rect 4100 317 4170 343
rect 4100 283 4118 317
rect 4152 283 4170 317
rect 4100 257 4170 283
rect 4200 317 4270 343
rect 4200 283 4218 317
rect 4252 283 4270 317
rect 4200 257 4270 283
rect 4300 317 4370 343
rect 4300 283 4318 317
rect 4352 283 4370 317
rect 4300 257 4370 283
rect 4400 317 4470 343
rect 4400 283 4418 317
rect 4452 283 4470 317
rect 4400 257 4470 283
rect 4500 317 4570 343
rect 4500 283 4518 317
rect 4552 283 4570 317
rect 4500 257 4570 283
rect 4600 317 4670 343
rect 4600 283 4618 317
rect 4652 283 4670 317
rect 4600 257 4670 283
rect 4700 317 4770 343
rect 4700 283 4718 317
rect 4752 283 4770 317
rect 4700 257 4770 283
rect 4800 257 4870 343
rect 4900 257 4970 343
rect 5000 257 5070 343
rect 5100 317 5170 343
rect 5100 283 5118 317
rect 5152 283 5170 317
rect 5100 257 5170 283
rect 5200 317 5270 343
rect 5200 283 5218 317
rect 5252 283 5270 317
rect 5200 257 5270 283
rect 5300 257 5370 343
rect 5400 257 5470 343
rect 5500 317 5570 343
rect 5500 283 5518 317
rect 5552 283 5570 317
rect 5500 257 5570 283
rect 5600 317 5654 343
rect 5600 283 5612 317
rect 5646 283 5654 317
rect 5600 257 5654 283
rect 3616 177 3670 203
rect 3616 143 3624 177
rect 3658 143 3670 177
rect 3616 117 3670 143
rect 3700 177 3770 203
rect 3700 143 3718 177
rect 3752 143 3770 177
rect 3700 117 3770 143
rect 3800 117 3870 203
rect 3900 177 3970 203
rect 3900 143 3918 177
rect 3952 143 3970 177
rect 3900 117 3970 143
rect 4000 177 4070 203
rect 4000 143 4018 177
rect 4052 143 4070 177
rect 4000 117 4070 143
rect 4100 117 4170 203
rect 4200 117 4270 203
rect 4300 117 4370 203
rect 4400 177 4470 203
rect 4400 143 4418 177
rect 4452 143 4470 177
rect 4400 117 4470 143
rect 4500 177 4570 203
rect 4500 143 4518 177
rect 4552 143 4570 177
rect 4500 117 4570 143
rect 4600 177 4670 203
rect 4600 143 4618 177
rect 4652 143 4670 177
rect 4600 117 4670 143
rect 4700 177 4754 203
rect 4700 143 4712 177
rect 4746 143 4754 177
rect 4700 117 4754 143
rect 6316 457 6370 483
rect 6316 423 6324 457
rect 6358 423 6370 457
rect 6316 397 6370 423
rect 6400 457 6454 483
rect 6400 423 6412 457
rect 6446 423 6454 457
rect 6400 397 6454 423
rect 6512 472 6570 483
rect 6512 438 6524 472
rect 6558 438 6570 472
rect 6512 397 6570 438
rect 6600 457 6670 483
rect 6600 423 6618 457
rect 6652 423 6670 457
rect 6600 397 6670 423
rect 6700 442 6758 483
rect 6700 408 6712 442
rect 6746 408 6758 442
rect 6700 397 6758 408
rect 6820 457 6880 483
rect 6820 423 6828 457
rect 6862 423 6880 457
rect 6820 397 6880 423
rect 6910 457 6980 483
rect 6910 423 6928 457
rect 6962 423 6980 457
rect 6910 397 6980 423
rect 7010 457 7080 483
rect 7010 423 7028 457
rect 7062 423 7080 457
rect 7010 397 7080 423
rect 7110 457 7180 483
rect 7110 423 7128 457
rect 7162 423 7180 457
rect 7110 397 7180 423
rect 7210 457 7280 483
rect 7210 423 7228 457
rect 7262 423 7280 457
rect 7210 397 7280 423
rect 7310 457 7380 483
rect 7310 423 7328 457
rect 7362 423 7380 457
rect 7310 397 7380 423
rect 7410 457 7470 483
rect 7410 423 7428 457
rect 7462 423 7470 457
rect 7410 397 7470 423
rect 5716 317 5770 343
rect 5716 283 5724 317
rect 5758 283 5770 317
rect 5716 257 5770 283
rect 5800 317 5870 343
rect 5800 283 5818 317
rect 5852 283 5870 317
rect 5800 257 5870 283
rect 5900 317 5970 343
rect 5900 283 5918 317
rect 5952 283 5970 317
rect 5900 257 5970 283
rect 6000 317 6070 343
rect 6000 283 6018 317
rect 6052 283 6070 317
rect 6000 257 6070 283
rect 6100 317 6170 343
rect 6100 283 6118 317
rect 6152 283 6170 317
rect 6100 257 6170 283
rect 6200 317 6270 343
rect 6200 283 6218 317
rect 6252 283 6270 317
rect 6200 257 6270 283
rect 6300 317 6370 343
rect 6300 283 6318 317
rect 6352 283 6370 317
rect 6300 257 6370 283
rect 6400 317 6454 343
rect 6400 283 6412 317
rect 6446 283 6454 317
rect 6400 257 6454 283
rect 6512 332 6570 343
rect 6512 298 6524 332
rect 6558 298 6570 332
rect 6512 257 6570 298
rect 6600 317 6670 343
rect 6600 283 6618 317
rect 6652 283 6670 317
rect 6600 257 6670 283
rect 6700 302 6758 343
rect 6700 268 6712 302
rect 6746 268 6758 302
rect 6700 257 6758 268
rect 6820 317 6880 343
rect 6820 283 6828 317
rect 6862 283 6880 317
rect 6820 257 6880 283
rect 6910 317 6980 343
rect 6910 283 6928 317
rect 6962 283 6980 317
rect 6910 257 6980 283
rect 7010 317 7080 343
rect 7010 283 7028 317
rect 7062 283 7080 317
rect 7010 257 7080 283
rect 7110 317 7180 343
rect 7110 283 7128 317
rect 7162 283 7180 317
rect 7110 257 7180 283
rect 7210 317 7280 343
rect 7210 283 7228 317
rect 7262 283 7280 317
rect 7210 257 7280 283
rect 7310 317 7380 343
rect 7310 283 7328 317
rect 7362 283 7380 317
rect 7310 257 7380 283
rect 7410 317 7470 343
rect 7410 283 7428 317
rect 7462 283 7470 317
rect 7410 257 7470 283
rect 4816 177 4870 203
rect 4816 143 4824 177
rect 4858 143 4870 177
rect 4816 117 4870 143
rect 4900 177 4970 203
rect 4900 143 4918 177
rect 4952 143 4970 177
rect 4900 117 4970 143
rect 5000 177 5070 203
rect 5000 143 5018 177
rect 5052 143 5070 177
rect 5000 117 5070 143
rect 5100 177 5170 203
rect 5100 143 5118 177
rect 5152 143 5170 177
rect 5100 117 5170 143
rect 5200 177 5270 203
rect 5200 143 5218 177
rect 5252 143 5270 177
rect 5200 117 5270 143
rect 5300 117 5370 203
rect 5400 177 5470 203
rect 5400 143 5418 177
rect 5452 143 5470 177
rect 5400 117 5470 143
rect 5500 177 5570 203
rect 5500 143 5518 177
rect 5552 143 5570 177
rect 5500 117 5570 143
rect 5600 117 5670 203
rect 5700 177 5770 203
rect 5700 143 5718 177
rect 5752 143 5770 177
rect 5700 117 5770 143
rect 5800 177 5870 203
rect 5800 143 5818 177
rect 5852 143 5870 177
rect 5800 117 5870 143
rect 5900 117 5970 203
rect 6000 177 6070 203
rect 6000 143 6018 177
rect 6052 143 6070 177
rect 6000 117 6070 143
rect 6100 177 6154 203
rect 6100 143 6112 177
rect 6146 143 6154 177
rect 6100 117 6154 143
rect 6216 177 6270 203
rect 6216 143 6224 177
rect 6258 143 6270 177
rect 6216 117 6270 143
rect 6300 177 6370 203
rect 6300 143 6318 177
rect 6352 143 6370 177
rect 6300 117 6370 143
rect 6400 177 6454 203
rect 6400 143 6412 177
rect 6446 143 6454 177
rect 6400 117 6454 143
rect 6512 192 6570 203
rect 6512 158 6524 192
rect 6558 158 6570 192
rect 6512 117 6570 158
rect 6600 177 6670 203
rect 6600 143 6618 177
rect 6652 143 6670 177
rect 6600 117 6670 143
rect 6700 162 6758 203
rect 6700 128 6712 162
rect 6746 128 6758 162
rect 6700 117 6758 128
rect 6820 177 6880 203
rect 6820 143 6828 177
rect 6862 143 6880 177
rect 6820 117 6880 143
rect 6910 177 6980 203
rect 6910 143 6928 177
rect 6962 143 6980 177
rect 6910 117 6980 143
rect 7010 177 7080 203
rect 7010 143 7028 177
rect 7062 143 7080 177
rect 7010 117 7080 143
rect 7110 177 7180 203
rect 7110 143 7128 177
rect 7162 143 7180 177
rect 7110 117 7180 143
rect 7210 177 7280 203
rect 7210 143 7228 177
rect 7262 143 7280 177
rect 7210 117 7280 143
rect 7310 177 7380 203
rect 7310 143 7328 177
rect 7362 143 7380 177
rect 7310 117 7380 143
rect 7410 177 7470 203
rect 7410 143 7428 177
rect 7462 143 7470 177
rect 7410 117 7470 143
rect 8140 -8 8290 29
rect 8140 -42 8162 -8
rect 8196 -42 8230 -8
rect 8264 -42 8290 -8
rect 8140 -60 8290 -42
rect 9252 -8 9402 29
rect 9252 -42 9278 -8
rect 9312 -42 9346 -8
rect 9380 -42 9402 -8
rect 9252 -60 9402 -42
rect 8140 -108 8290 -90
rect -94 -149 -30 -126
rect -94 -183 -82 -149
rect -48 -183 -30 -149
rect -94 -210 -30 -183
rect 0 -149 70 -126
rect 0 -183 18 -149
rect 52 -183 70 -149
rect 0 -210 70 -183
rect 100 -149 170 -126
rect 100 -183 118 -149
rect 152 -183 170 -149
rect 100 -210 170 -183
rect 200 -149 270 -126
rect 200 -183 218 -149
rect 252 -183 270 -149
rect 200 -210 270 -183
rect 300 -149 370 -126
rect 300 -183 318 -149
rect 352 -183 370 -149
rect 300 -210 370 -183
rect 400 -149 470 -126
rect 400 -183 418 -149
rect 452 -183 470 -149
rect 400 -210 470 -183
rect 500 -149 570 -126
rect 500 -183 518 -149
rect 552 -183 570 -149
rect 500 -210 570 -183
rect 600 -149 670 -126
rect 600 -183 618 -149
rect 652 -183 670 -149
rect 600 -210 670 -183
rect 700 -149 770 -126
rect 700 -183 718 -149
rect 752 -183 770 -149
rect 700 -210 770 -183
rect 800 -149 870 -126
rect 800 -183 818 -149
rect 852 -183 870 -149
rect 800 -210 870 -183
rect 900 -149 970 -126
rect 900 -183 918 -149
rect 952 -183 970 -149
rect 900 -210 970 -183
rect 1000 -149 1070 -126
rect 1000 -183 1018 -149
rect 1052 -183 1070 -149
rect 1000 -210 1070 -183
rect 1100 -149 1170 -126
rect 1100 -183 1118 -149
rect 1152 -183 1170 -149
rect 1100 -210 1170 -183
rect 1200 -149 1270 -126
rect 1200 -183 1218 -149
rect 1252 -183 1270 -149
rect 1200 -210 1270 -183
rect 1300 -149 1370 -126
rect 1300 -183 1318 -149
rect 1352 -183 1370 -149
rect 1300 -210 1370 -183
rect 1400 -149 1470 -126
rect 1400 -183 1418 -149
rect 1452 -183 1470 -149
rect 1400 -210 1470 -183
rect 1500 -149 1570 -126
rect 1500 -183 1518 -149
rect 1552 -183 1570 -149
rect 1500 -210 1570 -183
rect 1600 -149 1670 -126
rect 1600 -183 1618 -149
rect 1652 -183 1670 -149
rect 1600 -210 1670 -183
rect 1700 -149 1770 -126
rect 1700 -183 1718 -149
rect 1752 -183 1770 -149
rect 1700 -210 1770 -183
rect 1800 -149 1870 -126
rect 1800 -183 1818 -149
rect 1852 -183 1870 -149
rect 1800 -210 1870 -183
rect 1900 -149 1970 -126
rect 1900 -183 1918 -149
rect 1952 -183 1970 -149
rect 1900 -210 1970 -183
rect 2000 -149 2070 -126
rect 2000 -183 2018 -149
rect 2052 -183 2070 -149
rect 2000 -210 2070 -183
rect 2100 -149 2170 -126
rect 2100 -183 2118 -149
rect 2152 -183 2170 -149
rect 2100 -210 2170 -183
rect 2200 -149 2270 -126
rect 2200 -183 2218 -149
rect 2252 -183 2270 -149
rect 2200 -210 2270 -183
rect 2300 -149 2370 -126
rect 2300 -183 2318 -149
rect 2352 -183 2370 -149
rect 2300 -210 2370 -183
rect 2400 -149 2470 -126
rect 2400 -183 2418 -149
rect 2452 -183 2470 -149
rect 2400 -210 2470 -183
rect 2500 -149 2570 -126
rect 2500 -183 2518 -149
rect 2552 -183 2570 -149
rect 2500 -210 2570 -183
rect 2600 -149 2670 -126
rect 2600 -183 2618 -149
rect 2652 -183 2670 -149
rect 2600 -210 2670 -183
rect 2700 -149 2770 -126
rect 2700 -183 2718 -149
rect 2752 -183 2770 -149
rect 2700 -210 2770 -183
rect 2800 -149 2870 -126
rect 2800 -183 2818 -149
rect 2852 -183 2870 -149
rect 2800 -210 2870 -183
rect 2900 -149 2970 -126
rect 2900 -183 2918 -149
rect 2952 -183 2970 -149
rect 2900 -210 2970 -183
rect 3000 -149 3070 -126
rect 3000 -183 3018 -149
rect 3052 -183 3070 -149
rect 3000 -210 3070 -183
rect 3100 -149 3170 -126
rect 3100 -183 3118 -149
rect 3152 -183 3170 -149
rect 3100 -210 3170 -183
rect 3200 -149 3270 -126
rect 3200 -183 3218 -149
rect 3252 -183 3270 -149
rect 3200 -210 3270 -183
rect 3300 -149 3370 -126
rect 3300 -183 3318 -149
rect 3352 -183 3370 -149
rect 3300 -210 3370 -183
rect 3400 -149 3470 -126
rect 3400 -183 3418 -149
rect 3452 -183 3470 -149
rect 3400 -210 3470 -183
rect 3500 -149 3570 -126
rect 3500 -183 3518 -149
rect 3552 -183 3570 -149
rect 3500 -210 3570 -183
rect 3600 -149 3670 -126
rect 3600 -183 3618 -149
rect 3652 -183 3670 -149
rect 3600 -210 3670 -183
rect 3700 -149 3770 -126
rect 3700 -183 3718 -149
rect 3752 -183 3770 -149
rect 3700 -210 3770 -183
rect 3800 -149 3870 -126
rect 3800 -183 3818 -149
rect 3852 -183 3870 -149
rect 3800 -210 3870 -183
rect 3900 -149 3970 -126
rect 3900 -183 3918 -149
rect 3952 -183 3970 -149
rect 3900 -210 3970 -183
rect 4000 -149 4070 -126
rect 4000 -183 4018 -149
rect 4052 -183 4070 -149
rect 4000 -210 4070 -183
rect 4100 -149 4170 -126
rect 4100 -183 4118 -149
rect 4152 -183 4170 -149
rect 4100 -210 4170 -183
rect 4200 -149 4270 -126
rect 4200 -183 4218 -149
rect 4252 -183 4270 -149
rect 4200 -210 4270 -183
rect 4300 -149 4370 -126
rect 4300 -183 4318 -149
rect 4352 -183 4370 -149
rect 4300 -210 4370 -183
rect 4400 -149 4470 -126
rect 4400 -183 4418 -149
rect 4452 -183 4470 -149
rect 4400 -210 4470 -183
rect 4500 -149 4570 -126
rect 4500 -183 4518 -149
rect 4552 -183 4570 -149
rect 4500 -210 4570 -183
rect 4600 -149 4670 -126
rect 4600 -183 4618 -149
rect 4652 -183 4670 -149
rect 4600 -210 4670 -183
rect 4700 -149 4770 -126
rect 4700 -183 4718 -149
rect 4752 -183 4770 -149
rect 4700 -210 4770 -183
rect 4800 -149 4870 -126
rect 4800 -183 4818 -149
rect 4852 -183 4870 -149
rect 4800 -210 4870 -183
rect 4900 -149 4970 -126
rect 4900 -183 4918 -149
rect 4952 -183 4970 -149
rect 4900 -210 4970 -183
rect 5000 -149 5070 -126
rect 5000 -183 5018 -149
rect 5052 -183 5070 -149
rect 5000 -210 5070 -183
rect 5100 -149 5170 -126
rect 5100 -183 5118 -149
rect 5152 -183 5170 -149
rect 5100 -210 5170 -183
rect 5200 -149 5270 -126
rect 5200 -183 5218 -149
rect 5252 -183 5270 -149
rect 5200 -210 5270 -183
rect 5300 -149 5370 -126
rect 5300 -183 5318 -149
rect 5352 -183 5370 -149
rect 5300 -210 5370 -183
rect 5400 -149 5470 -126
rect 5400 -183 5418 -149
rect 5452 -183 5470 -149
rect 5400 -210 5470 -183
rect 5500 -149 5570 -126
rect 5500 -183 5518 -149
rect 5552 -183 5570 -149
rect 5500 -210 5570 -183
rect 5600 -149 5670 -126
rect 5600 -183 5618 -149
rect 5652 -183 5670 -149
rect 5600 -210 5670 -183
rect 5700 -149 5770 -126
rect 5700 -183 5718 -149
rect 5752 -183 5770 -149
rect 5700 -210 5770 -183
rect 5800 -149 5870 -126
rect 5800 -183 5818 -149
rect 5852 -183 5870 -149
rect 5800 -210 5870 -183
rect 5900 -149 5970 -126
rect 5900 -183 5918 -149
rect 5952 -183 5970 -149
rect 5900 -210 5970 -183
rect 6000 -149 6070 -126
rect 6000 -183 6018 -149
rect 6052 -183 6070 -149
rect 6000 -210 6070 -183
rect 6100 -149 6170 -126
rect 6100 -183 6118 -149
rect 6152 -183 6170 -149
rect 6100 -210 6170 -183
rect 6200 -149 6270 -126
rect 6200 -183 6218 -149
rect 6252 -183 6270 -149
rect 6200 -210 6270 -183
rect 6300 -149 6364 -126
rect 6300 -183 6318 -149
rect 6352 -183 6364 -149
rect 8140 -142 8162 -108
rect 8196 -142 8230 -108
rect 8264 -142 8290 -108
rect 8140 -160 8290 -142
rect 9252 -108 9402 -90
rect 9252 -142 9278 -108
rect 9312 -142 9346 -108
rect 9380 -142 9402 -108
rect 9252 -160 9402 -142
rect 6300 -210 6364 -183
rect 8140 -208 8290 -190
rect 8140 -242 8162 -208
rect 8196 -242 8230 -208
rect 8264 -242 8290 -208
rect 8140 -260 8290 -242
rect 9252 -208 9402 -190
rect 9252 -242 9278 -208
rect 9312 -242 9346 -208
rect 9380 -242 9402 -208
rect 9252 -260 9402 -242
rect 8140 -308 8290 -290
rect 8140 -342 8162 -308
rect 8196 -342 8230 -308
rect 8264 -342 8290 -308
rect 8140 -360 8290 -342
rect 9252 -308 9402 -290
rect 9252 -342 9278 -308
rect 9312 -342 9346 -308
rect 9380 -342 9402 -308
rect 9252 -360 9402 -342
rect 8140 -408 8290 -390
rect 8140 -442 8162 -408
rect 8196 -442 8230 -408
rect 8264 -442 8290 -408
rect 8140 -460 8290 -442
rect 9252 -408 9402 -390
rect 9252 -442 9278 -408
rect 9312 -442 9346 -408
rect 9380 -442 9402 -408
rect 9252 -460 9402 -442
rect 8140 -508 8290 -490
rect 8140 -542 8162 -508
rect 8196 -542 8230 -508
rect 8264 -542 8290 -508
rect 8140 -560 8290 -542
rect 9252 -508 9402 -490
rect 9252 -542 9278 -508
rect 9312 -542 9346 -508
rect 9380 -542 9402 -508
rect 9252 -560 9402 -542
rect 8140 -608 8290 -590
rect 8140 -642 8162 -608
rect 8196 -642 8230 -608
rect 8264 -642 8290 -608
rect 8140 -660 8290 -642
rect 9252 -608 9402 -590
rect 9252 -642 9278 -608
rect 9312 -642 9346 -608
rect 9380 -642 9402 -608
rect 9252 -660 9402 -642
rect 8140 -708 8290 -690
rect 8140 -742 8162 -708
rect 8196 -742 8230 -708
rect 8264 -742 8290 -708
rect 8140 -760 8290 -742
rect 9252 -708 9402 -690
rect 9252 -742 9278 -708
rect 9312 -742 9346 -708
rect 9380 -742 9402 -708
rect 9252 -760 9402 -742
rect 8140 -808 8290 -790
rect 8140 -842 8162 -808
rect 8196 -842 8230 -808
rect 8264 -842 8290 -808
rect -10 -858 108 -846
rect -10 -892 -2 -858
rect 32 -892 66 -858
rect 100 -892 108 -858
rect -10 -910 108 -892
rect 162 -858 280 -846
rect 162 -892 170 -858
rect 204 -892 238 -858
rect 272 -892 280 -858
rect 162 -910 280 -892
rect 390 -858 508 -846
rect 390 -892 398 -858
rect 432 -892 466 -858
rect 500 -892 508 -858
rect 390 -910 508 -892
rect 562 -858 680 -846
rect 562 -892 570 -858
rect 604 -892 638 -858
rect 672 -892 680 -858
rect 562 -910 680 -892
rect 790 -858 908 -846
rect 790 -892 798 -858
rect 832 -892 866 -858
rect 900 -892 908 -858
rect -10 -958 108 -940
rect -10 -992 -2 -958
rect 32 -992 66 -958
rect 100 -992 108 -958
rect -10 -1010 108 -992
rect 162 -958 280 -940
rect 162 -992 170 -958
rect 204 -992 238 -958
rect 272 -992 280 -958
rect 162 -1010 280 -992
rect 390 -958 508 -940
rect 390 -992 398 -958
rect 432 -992 466 -958
rect 500 -992 508 -958
rect 390 -1010 508 -992
rect 562 -958 680 -940
rect 790 -910 908 -892
rect 962 -858 1080 -846
rect 962 -892 970 -858
rect 1004 -892 1038 -858
rect 1072 -892 1080 -858
rect 962 -910 1080 -892
rect 1190 -858 1308 -846
rect 1190 -892 1198 -858
rect 1232 -892 1266 -858
rect 1300 -892 1308 -858
rect 1190 -910 1308 -892
rect 1362 -858 1480 -846
rect 1362 -892 1370 -858
rect 1404 -892 1438 -858
rect 1472 -892 1480 -858
rect 1362 -910 1480 -892
rect 1590 -858 1708 -846
rect 1590 -892 1598 -858
rect 1632 -892 1666 -858
rect 1700 -892 1708 -858
rect 562 -992 570 -958
rect 604 -992 638 -958
rect 672 -992 680 -958
rect 562 -1010 680 -992
rect 790 -958 908 -940
rect 790 -992 798 -958
rect 832 -992 866 -958
rect 900 -992 908 -958
rect -10 -1058 108 -1040
rect -10 -1092 -2 -1058
rect 32 -1092 66 -1058
rect 100 -1092 108 -1058
rect -10 -1110 108 -1092
rect 162 -1058 280 -1040
rect 162 -1092 170 -1058
rect 204 -1092 238 -1058
rect 272 -1092 280 -1058
rect 162 -1110 280 -1092
rect 390 -1058 508 -1040
rect 390 -1092 398 -1058
rect 432 -1092 466 -1058
rect 500 -1092 508 -1058
rect 390 -1110 508 -1092
rect 562 -1058 680 -1040
rect 790 -1010 908 -992
rect 962 -958 1080 -940
rect 962 -992 970 -958
rect 1004 -992 1038 -958
rect 1072 -992 1080 -958
rect 962 -1010 1080 -992
rect 1190 -958 1308 -940
rect 1190 -992 1198 -958
rect 1232 -992 1266 -958
rect 1300 -992 1308 -958
rect 1190 -1010 1308 -992
rect 1362 -958 1480 -940
rect 1590 -910 1708 -892
rect 1762 -858 1880 -846
rect 1762 -892 1770 -858
rect 1804 -892 1838 -858
rect 1872 -892 1880 -858
rect 1762 -910 1880 -892
rect 1990 -858 2108 -846
rect 1990 -892 1998 -858
rect 2032 -892 2066 -858
rect 2100 -892 2108 -858
rect 1990 -910 2108 -892
rect 2162 -858 2280 -846
rect 2162 -892 2170 -858
rect 2204 -892 2238 -858
rect 2272 -892 2280 -858
rect 2162 -910 2280 -892
rect 2390 -858 2508 -846
rect 2390 -892 2398 -858
rect 2432 -892 2466 -858
rect 2500 -892 2508 -858
rect 1362 -992 1370 -958
rect 1404 -992 1438 -958
rect 1472 -992 1480 -958
rect 1362 -1010 1480 -992
rect 1590 -958 1708 -940
rect 1590 -992 1598 -958
rect 1632 -992 1666 -958
rect 1700 -992 1708 -958
rect 562 -1092 570 -1058
rect 604 -1092 638 -1058
rect 672 -1092 680 -1058
rect 562 -1110 680 -1092
rect 790 -1058 908 -1040
rect 790 -1092 798 -1058
rect 832 -1092 866 -1058
rect 900 -1092 908 -1058
rect -10 -1158 108 -1140
rect -10 -1192 -2 -1158
rect 32 -1192 66 -1158
rect 100 -1192 108 -1158
rect -10 -1210 108 -1192
rect 162 -1158 280 -1140
rect 162 -1192 170 -1158
rect 204 -1192 238 -1158
rect 272 -1192 280 -1158
rect 162 -1210 280 -1192
rect 390 -1158 508 -1140
rect 390 -1192 398 -1158
rect 432 -1192 466 -1158
rect 500 -1192 508 -1158
rect 390 -1210 508 -1192
rect 562 -1158 680 -1140
rect 790 -1110 908 -1092
rect 962 -1058 1080 -1040
rect 962 -1092 970 -1058
rect 1004 -1092 1038 -1058
rect 1072 -1092 1080 -1058
rect 962 -1110 1080 -1092
rect 1190 -1058 1308 -1040
rect 1190 -1092 1198 -1058
rect 1232 -1092 1266 -1058
rect 1300 -1092 1308 -1058
rect 1190 -1110 1308 -1092
rect 1362 -1058 1480 -1040
rect 1590 -1010 1708 -992
rect 1762 -958 1880 -940
rect 1762 -992 1770 -958
rect 1804 -992 1838 -958
rect 1872 -992 1880 -958
rect 1762 -1010 1880 -992
rect 1990 -958 2108 -940
rect 1990 -992 1998 -958
rect 2032 -992 2066 -958
rect 2100 -992 2108 -958
rect 1990 -1010 2108 -992
rect 2162 -958 2280 -940
rect 2390 -910 2508 -892
rect 2562 -858 2680 -846
rect 2562 -892 2570 -858
rect 2604 -892 2638 -858
rect 2672 -892 2680 -858
rect 2562 -910 2680 -892
rect 2790 -858 2908 -846
rect 2790 -892 2798 -858
rect 2832 -892 2866 -858
rect 2900 -892 2908 -858
rect 2790 -910 2908 -892
rect 2962 -858 3080 -846
rect 2962 -892 2970 -858
rect 3004 -892 3038 -858
rect 3072 -892 3080 -858
rect 2962 -910 3080 -892
rect 3190 -858 3308 -846
rect 3190 -892 3198 -858
rect 3232 -892 3266 -858
rect 3300 -892 3308 -858
rect 2162 -992 2170 -958
rect 2204 -992 2238 -958
rect 2272 -992 2280 -958
rect 2162 -1010 2280 -992
rect 2390 -958 2508 -940
rect 2390 -992 2398 -958
rect 2432 -992 2466 -958
rect 2500 -992 2508 -958
rect 1362 -1092 1370 -1058
rect 1404 -1092 1438 -1058
rect 1472 -1092 1480 -1058
rect 1362 -1110 1480 -1092
rect 1590 -1058 1708 -1040
rect 1590 -1092 1598 -1058
rect 1632 -1092 1666 -1058
rect 1700 -1092 1708 -1058
rect 562 -1192 570 -1158
rect 604 -1192 638 -1158
rect 672 -1192 680 -1158
rect 562 -1210 680 -1192
rect 790 -1158 908 -1140
rect 790 -1192 798 -1158
rect 832 -1192 866 -1158
rect 900 -1192 908 -1158
rect -10 -1258 108 -1240
rect -10 -1292 -2 -1258
rect 32 -1292 66 -1258
rect 100 -1292 108 -1258
rect -10 -1310 108 -1292
rect 162 -1258 280 -1240
rect 162 -1292 170 -1258
rect 204 -1292 238 -1258
rect 272 -1292 280 -1258
rect 162 -1310 280 -1292
rect 390 -1258 508 -1240
rect 390 -1292 398 -1258
rect 432 -1292 466 -1258
rect 500 -1292 508 -1258
rect 390 -1310 508 -1292
rect 562 -1258 680 -1240
rect 790 -1210 908 -1192
rect 962 -1158 1080 -1140
rect 962 -1192 970 -1158
rect 1004 -1192 1038 -1158
rect 1072 -1192 1080 -1158
rect 962 -1210 1080 -1192
rect 1190 -1158 1308 -1140
rect 1190 -1192 1198 -1158
rect 1232 -1192 1266 -1158
rect 1300 -1192 1308 -1158
rect 1190 -1210 1308 -1192
rect 1362 -1158 1480 -1140
rect 1590 -1110 1708 -1092
rect 1762 -1058 1880 -1040
rect 1762 -1092 1770 -1058
rect 1804 -1092 1838 -1058
rect 1872 -1092 1880 -1058
rect 1762 -1110 1880 -1092
rect 1990 -1058 2108 -1040
rect 1990 -1092 1998 -1058
rect 2032 -1092 2066 -1058
rect 2100 -1092 2108 -1058
rect 1990 -1110 2108 -1092
rect 2162 -1058 2280 -1040
rect 2390 -1010 2508 -992
rect 2562 -958 2680 -940
rect 2562 -992 2570 -958
rect 2604 -992 2638 -958
rect 2672 -992 2680 -958
rect 2562 -1010 2680 -992
rect 2790 -958 2908 -940
rect 2790 -992 2798 -958
rect 2832 -992 2866 -958
rect 2900 -992 2908 -958
rect 2790 -1010 2908 -992
rect 2962 -958 3080 -940
rect 3190 -910 3308 -892
rect 3362 -858 3480 -846
rect 3362 -892 3370 -858
rect 3404 -892 3438 -858
rect 3472 -892 3480 -858
rect 3362 -910 3480 -892
rect 3590 -858 3708 -846
rect 3590 -892 3598 -858
rect 3632 -892 3666 -858
rect 3700 -892 3708 -858
rect 3590 -910 3708 -892
rect 3762 -858 3880 -846
rect 3762 -892 3770 -858
rect 3804 -892 3838 -858
rect 3872 -892 3880 -858
rect 3762 -910 3880 -892
rect 3990 -858 4108 -846
rect 3990 -892 3998 -858
rect 4032 -892 4066 -858
rect 4100 -892 4108 -858
rect 2962 -992 2970 -958
rect 3004 -992 3038 -958
rect 3072 -992 3080 -958
rect 2962 -1010 3080 -992
rect 3190 -958 3308 -940
rect 3190 -992 3198 -958
rect 3232 -992 3266 -958
rect 3300 -992 3308 -958
rect 2162 -1092 2170 -1058
rect 2204 -1092 2238 -1058
rect 2272 -1092 2280 -1058
rect 2162 -1110 2280 -1092
rect 2390 -1058 2508 -1040
rect 2390 -1092 2398 -1058
rect 2432 -1092 2466 -1058
rect 2500 -1092 2508 -1058
rect 1362 -1192 1370 -1158
rect 1404 -1192 1438 -1158
rect 1472 -1192 1480 -1158
rect 1362 -1210 1480 -1192
rect 1590 -1158 1708 -1140
rect 1590 -1192 1598 -1158
rect 1632 -1192 1666 -1158
rect 1700 -1192 1708 -1158
rect 562 -1292 570 -1258
rect 604 -1292 638 -1258
rect 672 -1292 680 -1258
rect 562 -1310 680 -1292
rect 790 -1258 908 -1240
rect 790 -1292 798 -1258
rect 832 -1292 866 -1258
rect 900 -1292 908 -1258
rect -10 -1358 108 -1340
rect -10 -1392 -2 -1358
rect 32 -1392 66 -1358
rect 100 -1392 108 -1358
rect -10 -1410 108 -1392
rect 162 -1358 280 -1340
rect 162 -1392 170 -1358
rect 204 -1392 238 -1358
rect 272 -1392 280 -1358
rect 162 -1410 280 -1392
rect 390 -1358 508 -1340
rect 390 -1392 398 -1358
rect 432 -1392 466 -1358
rect 500 -1392 508 -1358
rect 390 -1410 508 -1392
rect 562 -1358 680 -1340
rect 790 -1310 908 -1292
rect 962 -1258 1080 -1240
rect 962 -1292 970 -1258
rect 1004 -1292 1038 -1258
rect 1072 -1292 1080 -1258
rect 962 -1310 1080 -1292
rect 1190 -1258 1308 -1240
rect 1190 -1292 1198 -1258
rect 1232 -1292 1266 -1258
rect 1300 -1292 1308 -1258
rect 1190 -1310 1308 -1292
rect 1362 -1258 1480 -1240
rect 1590 -1210 1708 -1192
rect 1762 -1158 1880 -1140
rect 1762 -1192 1770 -1158
rect 1804 -1192 1838 -1158
rect 1872 -1192 1880 -1158
rect 1762 -1210 1880 -1192
rect 1990 -1158 2108 -1140
rect 1990 -1192 1998 -1158
rect 2032 -1192 2066 -1158
rect 2100 -1192 2108 -1158
rect 1990 -1210 2108 -1192
rect 2162 -1158 2280 -1140
rect 2390 -1110 2508 -1092
rect 2562 -1058 2680 -1040
rect 2562 -1092 2570 -1058
rect 2604 -1092 2638 -1058
rect 2672 -1092 2680 -1058
rect 2562 -1110 2680 -1092
rect 2790 -1058 2908 -1040
rect 2790 -1092 2798 -1058
rect 2832 -1092 2866 -1058
rect 2900 -1092 2908 -1058
rect 2790 -1110 2908 -1092
rect 2962 -1058 3080 -1040
rect 3190 -1010 3308 -992
rect 3362 -958 3480 -940
rect 3362 -992 3370 -958
rect 3404 -992 3438 -958
rect 3472 -992 3480 -958
rect 3362 -1010 3480 -992
rect 3590 -958 3708 -940
rect 3590 -992 3598 -958
rect 3632 -992 3666 -958
rect 3700 -992 3708 -958
rect 3590 -1010 3708 -992
rect 3762 -958 3880 -940
rect 3990 -910 4108 -892
rect 4162 -858 4280 -846
rect 4162 -892 4170 -858
rect 4204 -892 4238 -858
rect 4272 -892 4280 -858
rect 4162 -910 4280 -892
rect 4390 -858 4508 -846
rect 4390 -892 4398 -858
rect 4432 -892 4466 -858
rect 4500 -892 4508 -858
rect 4390 -910 4508 -892
rect 4562 -858 4680 -846
rect 4562 -892 4570 -858
rect 4604 -892 4638 -858
rect 4672 -892 4680 -858
rect 4562 -910 4680 -892
rect 4790 -858 4908 -846
rect 4790 -892 4798 -858
rect 4832 -892 4866 -858
rect 4900 -892 4908 -858
rect 3762 -992 3770 -958
rect 3804 -992 3838 -958
rect 3872 -992 3880 -958
rect 3762 -1010 3880 -992
rect 3990 -958 4108 -940
rect 3990 -992 3998 -958
rect 4032 -992 4066 -958
rect 4100 -992 4108 -958
rect 2962 -1092 2970 -1058
rect 3004 -1092 3038 -1058
rect 3072 -1092 3080 -1058
rect 2962 -1110 3080 -1092
rect 3190 -1058 3308 -1040
rect 3190 -1092 3198 -1058
rect 3232 -1092 3266 -1058
rect 3300 -1092 3308 -1058
rect 2162 -1192 2170 -1158
rect 2204 -1192 2238 -1158
rect 2272 -1192 2280 -1158
rect 2162 -1210 2280 -1192
rect 2390 -1158 2508 -1140
rect 2390 -1192 2398 -1158
rect 2432 -1192 2466 -1158
rect 2500 -1192 2508 -1158
rect 1362 -1292 1370 -1258
rect 1404 -1292 1438 -1258
rect 1472 -1292 1480 -1258
rect 1362 -1310 1480 -1292
rect 1590 -1258 1708 -1240
rect 1590 -1292 1598 -1258
rect 1632 -1292 1666 -1258
rect 1700 -1292 1708 -1258
rect 562 -1392 570 -1358
rect 604 -1392 638 -1358
rect 672 -1392 680 -1358
rect 562 -1410 680 -1392
rect 790 -1358 908 -1340
rect 790 -1392 798 -1358
rect 832 -1392 866 -1358
rect 900 -1392 908 -1358
rect -10 -1458 108 -1440
rect -10 -1492 -2 -1458
rect 32 -1492 66 -1458
rect 100 -1492 108 -1458
rect -10 -1510 108 -1492
rect 162 -1458 280 -1440
rect 162 -1492 170 -1458
rect 204 -1492 238 -1458
rect 272 -1492 280 -1458
rect 162 -1510 280 -1492
rect 390 -1458 508 -1440
rect 390 -1492 398 -1458
rect 432 -1492 466 -1458
rect 500 -1492 508 -1458
rect 390 -1510 508 -1492
rect 562 -1458 680 -1440
rect 790 -1410 908 -1392
rect 962 -1358 1080 -1340
rect 962 -1392 970 -1358
rect 1004 -1392 1038 -1358
rect 1072 -1392 1080 -1358
rect 962 -1410 1080 -1392
rect 1190 -1358 1308 -1340
rect 1190 -1392 1198 -1358
rect 1232 -1392 1266 -1358
rect 1300 -1392 1308 -1358
rect 1190 -1410 1308 -1392
rect 1362 -1358 1480 -1340
rect 1590 -1310 1708 -1292
rect 1762 -1258 1880 -1240
rect 1762 -1292 1770 -1258
rect 1804 -1292 1838 -1258
rect 1872 -1292 1880 -1258
rect 1762 -1310 1880 -1292
rect 1990 -1258 2108 -1240
rect 1990 -1292 1998 -1258
rect 2032 -1292 2066 -1258
rect 2100 -1292 2108 -1258
rect 1990 -1310 2108 -1292
rect 2162 -1258 2280 -1240
rect 2390 -1210 2508 -1192
rect 2562 -1158 2680 -1140
rect 2562 -1192 2570 -1158
rect 2604 -1192 2638 -1158
rect 2672 -1192 2680 -1158
rect 2562 -1210 2680 -1192
rect 2790 -1158 2908 -1140
rect 2790 -1192 2798 -1158
rect 2832 -1192 2866 -1158
rect 2900 -1192 2908 -1158
rect 2790 -1210 2908 -1192
rect 2962 -1158 3080 -1140
rect 3190 -1110 3308 -1092
rect 3362 -1058 3480 -1040
rect 3362 -1092 3370 -1058
rect 3404 -1092 3438 -1058
rect 3472 -1092 3480 -1058
rect 3362 -1110 3480 -1092
rect 3590 -1058 3708 -1040
rect 3590 -1092 3598 -1058
rect 3632 -1092 3666 -1058
rect 3700 -1092 3708 -1058
rect 3590 -1110 3708 -1092
rect 3762 -1058 3880 -1040
rect 3990 -1010 4108 -992
rect 4162 -958 4280 -940
rect 4162 -992 4170 -958
rect 4204 -992 4238 -958
rect 4272 -992 4280 -958
rect 4162 -1010 4280 -992
rect 4390 -958 4508 -940
rect 4390 -992 4398 -958
rect 4432 -992 4466 -958
rect 4500 -992 4508 -958
rect 4390 -1010 4508 -992
rect 4562 -958 4680 -940
rect 4790 -910 4908 -892
rect 4962 -858 5080 -846
rect 4962 -892 4970 -858
rect 5004 -892 5038 -858
rect 5072 -892 5080 -858
rect 4962 -910 5080 -892
rect 5190 -858 5308 -846
rect 5190 -892 5198 -858
rect 5232 -892 5266 -858
rect 5300 -892 5308 -858
rect 5190 -910 5308 -892
rect 5362 -858 5480 -846
rect 5362 -892 5370 -858
rect 5404 -892 5438 -858
rect 5472 -892 5480 -858
rect 5362 -910 5480 -892
rect 5590 -858 5708 -846
rect 5590 -892 5598 -858
rect 5632 -892 5666 -858
rect 5700 -892 5708 -858
rect 4562 -992 4570 -958
rect 4604 -992 4638 -958
rect 4672 -992 4680 -958
rect 4562 -1010 4680 -992
rect 4790 -958 4908 -940
rect 4790 -992 4798 -958
rect 4832 -992 4866 -958
rect 4900 -992 4908 -958
rect 3762 -1092 3770 -1058
rect 3804 -1092 3838 -1058
rect 3872 -1092 3880 -1058
rect 3762 -1110 3880 -1092
rect 3990 -1058 4108 -1040
rect 3990 -1092 3998 -1058
rect 4032 -1092 4066 -1058
rect 4100 -1092 4108 -1058
rect 2962 -1192 2970 -1158
rect 3004 -1192 3038 -1158
rect 3072 -1192 3080 -1158
rect 2962 -1210 3080 -1192
rect 3190 -1158 3308 -1140
rect 3190 -1192 3198 -1158
rect 3232 -1192 3266 -1158
rect 3300 -1192 3308 -1158
rect 2162 -1292 2170 -1258
rect 2204 -1292 2238 -1258
rect 2272 -1292 2280 -1258
rect 2162 -1310 2280 -1292
rect 2390 -1258 2508 -1240
rect 2390 -1292 2398 -1258
rect 2432 -1292 2466 -1258
rect 2500 -1292 2508 -1258
rect 1362 -1392 1370 -1358
rect 1404 -1392 1438 -1358
rect 1472 -1392 1480 -1358
rect 1362 -1410 1480 -1392
rect 1590 -1358 1708 -1340
rect 1590 -1392 1598 -1358
rect 1632 -1392 1666 -1358
rect 1700 -1392 1708 -1358
rect 562 -1492 570 -1458
rect 604 -1492 638 -1458
rect 672 -1492 680 -1458
rect 562 -1510 680 -1492
rect 790 -1458 908 -1440
rect 790 -1492 798 -1458
rect 832 -1492 866 -1458
rect 900 -1492 908 -1458
rect -10 -1558 108 -1540
rect -10 -1592 -2 -1558
rect 32 -1592 66 -1558
rect 100 -1592 108 -1558
rect -10 -1610 108 -1592
rect 162 -1558 280 -1540
rect 162 -1592 170 -1558
rect 204 -1592 238 -1558
rect 272 -1592 280 -1558
rect 162 -1610 280 -1592
rect 390 -1558 508 -1540
rect 390 -1592 398 -1558
rect 432 -1592 466 -1558
rect 500 -1592 508 -1558
rect 390 -1610 508 -1592
rect 562 -1558 680 -1540
rect 790 -1510 908 -1492
rect 962 -1458 1080 -1440
rect 962 -1492 970 -1458
rect 1004 -1492 1038 -1458
rect 1072 -1492 1080 -1458
rect 962 -1510 1080 -1492
rect 1190 -1458 1308 -1440
rect 1190 -1492 1198 -1458
rect 1232 -1492 1266 -1458
rect 1300 -1492 1308 -1458
rect 1190 -1510 1308 -1492
rect 1362 -1458 1480 -1440
rect 1590 -1410 1708 -1392
rect 1762 -1358 1880 -1340
rect 1762 -1392 1770 -1358
rect 1804 -1392 1838 -1358
rect 1872 -1392 1880 -1358
rect 1762 -1410 1880 -1392
rect 1990 -1358 2108 -1340
rect 1990 -1392 1998 -1358
rect 2032 -1392 2066 -1358
rect 2100 -1392 2108 -1358
rect 1990 -1410 2108 -1392
rect 2162 -1358 2280 -1340
rect 2390 -1310 2508 -1292
rect 2562 -1258 2680 -1240
rect 2562 -1292 2570 -1258
rect 2604 -1292 2638 -1258
rect 2672 -1292 2680 -1258
rect 2562 -1310 2680 -1292
rect 2790 -1258 2908 -1240
rect 2790 -1292 2798 -1258
rect 2832 -1292 2866 -1258
rect 2900 -1292 2908 -1258
rect 2790 -1310 2908 -1292
rect 2962 -1258 3080 -1240
rect 3190 -1210 3308 -1192
rect 3362 -1158 3480 -1140
rect 3362 -1192 3370 -1158
rect 3404 -1192 3438 -1158
rect 3472 -1192 3480 -1158
rect 3362 -1210 3480 -1192
rect 3590 -1158 3708 -1140
rect 3590 -1192 3598 -1158
rect 3632 -1192 3666 -1158
rect 3700 -1192 3708 -1158
rect 3590 -1210 3708 -1192
rect 3762 -1158 3880 -1140
rect 3990 -1110 4108 -1092
rect 4162 -1058 4280 -1040
rect 4162 -1092 4170 -1058
rect 4204 -1092 4238 -1058
rect 4272 -1092 4280 -1058
rect 4162 -1110 4280 -1092
rect 4390 -1058 4508 -1040
rect 4390 -1092 4398 -1058
rect 4432 -1092 4466 -1058
rect 4500 -1092 4508 -1058
rect 4390 -1110 4508 -1092
rect 4562 -1058 4680 -1040
rect 4790 -1010 4908 -992
rect 4962 -958 5080 -940
rect 4962 -992 4970 -958
rect 5004 -992 5038 -958
rect 5072 -992 5080 -958
rect 4962 -1010 5080 -992
rect 5190 -958 5308 -940
rect 5190 -992 5198 -958
rect 5232 -992 5266 -958
rect 5300 -992 5308 -958
rect 5190 -1010 5308 -992
rect 5362 -958 5480 -940
rect 5590 -910 5708 -892
rect 5762 -858 5880 -846
rect 5762 -892 5770 -858
rect 5804 -892 5838 -858
rect 5872 -892 5880 -858
rect 5762 -910 5880 -892
rect 5990 -858 6108 -846
rect 5990 -892 5998 -858
rect 6032 -892 6066 -858
rect 6100 -892 6108 -858
rect 5990 -910 6108 -892
rect 6162 -858 6280 -846
rect 6162 -892 6170 -858
rect 6204 -892 6238 -858
rect 6272 -892 6280 -858
rect 8140 -860 8290 -842
rect 9252 -808 9402 -790
rect 9252 -842 9278 -808
rect 9312 -842 9346 -808
rect 9380 -842 9402 -808
rect 9252 -860 9402 -842
rect 6162 -910 6280 -892
rect 5362 -992 5370 -958
rect 5404 -992 5438 -958
rect 5472 -992 5480 -958
rect 5362 -1010 5480 -992
rect 5590 -958 5708 -940
rect 5590 -992 5598 -958
rect 5632 -992 5666 -958
rect 5700 -992 5708 -958
rect 4562 -1092 4570 -1058
rect 4604 -1092 4638 -1058
rect 4672 -1092 4680 -1058
rect 4562 -1110 4680 -1092
rect 4790 -1058 4908 -1040
rect 4790 -1092 4798 -1058
rect 4832 -1092 4866 -1058
rect 4900 -1092 4908 -1058
rect 3762 -1192 3770 -1158
rect 3804 -1192 3838 -1158
rect 3872 -1192 3880 -1158
rect 3762 -1210 3880 -1192
rect 3990 -1158 4108 -1140
rect 3990 -1192 3998 -1158
rect 4032 -1192 4066 -1158
rect 4100 -1192 4108 -1158
rect 2962 -1292 2970 -1258
rect 3004 -1292 3038 -1258
rect 3072 -1292 3080 -1258
rect 2962 -1310 3080 -1292
rect 3190 -1258 3308 -1240
rect 3190 -1292 3198 -1258
rect 3232 -1292 3266 -1258
rect 3300 -1292 3308 -1258
rect 2162 -1392 2170 -1358
rect 2204 -1392 2238 -1358
rect 2272 -1392 2280 -1358
rect 2162 -1410 2280 -1392
rect 2390 -1358 2508 -1340
rect 2390 -1392 2398 -1358
rect 2432 -1392 2466 -1358
rect 2500 -1392 2508 -1358
rect 1362 -1492 1370 -1458
rect 1404 -1492 1438 -1458
rect 1472 -1492 1480 -1458
rect 1362 -1510 1480 -1492
rect 1590 -1458 1708 -1440
rect 1590 -1492 1598 -1458
rect 1632 -1492 1666 -1458
rect 1700 -1492 1708 -1458
rect 562 -1592 570 -1558
rect 604 -1592 638 -1558
rect 672 -1592 680 -1558
rect 562 -1610 680 -1592
rect 790 -1558 908 -1540
rect 790 -1592 798 -1558
rect 832 -1592 866 -1558
rect 900 -1592 908 -1558
rect -10 -1658 108 -1640
rect -10 -1692 -2 -1658
rect 32 -1692 66 -1658
rect 100 -1692 108 -1658
rect -10 -1710 108 -1692
rect 162 -1658 280 -1640
rect 162 -1692 170 -1658
rect 204 -1692 238 -1658
rect 272 -1692 280 -1658
rect 162 -1710 280 -1692
rect 390 -1658 508 -1640
rect 390 -1692 398 -1658
rect 432 -1692 466 -1658
rect 500 -1692 508 -1658
rect 390 -1710 508 -1692
rect 562 -1658 680 -1640
rect 790 -1610 908 -1592
rect 962 -1558 1080 -1540
rect 962 -1592 970 -1558
rect 1004 -1592 1038 -1558
rect 1072 -1592 1080 -1558
rect 962 -1610 1080 -1592
rect 1190 -1558 1308 -1540
rect 1190 -1592 1198 -1558
rect 1232 -1592 1266 -1558
rect 1300 -1592 1308 -1558
rect 1190 -1610 1308 -1592
rect 1362 -1558 1480 -1540
rect 1590 -1510 1708 -1492
rect 1762 -1458 1880 -1440
rect 1762 -1492 1770 -1458
rect 1804 -1492 1838 -1458
rect 1872 -1492 1880 -1458
rect 1762 -1510 1880 -1492
rect 1990 -1458 2108 -1440
rect 1990 -1492 1998 -1458
rect 2032 -1492 2066 -1458
rect 2100 -1492 2108 -1458
rect 1990 -1510 2108 -1492
rect 2162 -1458 2280 -1440
rect 2390 -1410 2508 -1392
rect 2562 -1358 2680 -1340
rect 2562 -1392 2570 -1358
rect 2604 -1392 2638 -1358
rect 2672 -1392 2680 -1358
rect 2562 -1410 2680 -1392
rect 2790 -1358 2908 -1340
rect 2790 -1392 2798 -1358
rect 2832 -1392 2866 -1358
rect 2900 -1392 2908 -1358
rect 2790 -1410 2908 -1392
rect 2962 -1358 3080 -1340
rect 3190 -1310 3308 -1292
rect 3362 -1258 3480 -1240
rect 3362 -1292 3370 -1258
rect 3404 -1292 3438 -1258
rect 3472 -1292 3480 -1258
rect 3362 -1310 3480 -1292
rect 3590 -1258 3708 -1240
rect 3590 -1292 3598 -1258
rect 3632 -1292 3666 -1258
rect 3700 -1292 3708 -1258
rect 3590 -1310 3708 -1292
rect 3762 -1258 3880 -1240
rect 3990 -1210 4108 -1192
rect 4162 -1158 4280 -1140
rect 4162 -1192 4170 -1158
rect 4204 -1192 4238 -1158
rect 4272 -1192 4280 -1158
rect 4162 -1210 4280 -1192
rect 4390 -1158 4508 -1140
rect 4390 -1192 4398 -1158
rect 4432 -1192 4466 -1158
rect 4500 -1192 4508 -1158
rect 4390 -1210 4508 -1192
rect 4562 -1158 4680 -1140
rect 4790 -1110 4908 -1092
rect 4962 -1058 5080 -1040
rect 4962 -1092 4970 -1058
rect 5004 -1092 5038 -1058
rect 5072 -1092 5080 -1058
rect 4962 -1110 5080 -1092
rect 5190 -1058 5308 -1040
rect 5190 -1092 5198 -1058
rect 5232 -1092 5266 -1058
rect 5300 -1092 5308 -1058
rect 5190 -1110 5308 -1092
rect 5362 -1058 5480 -1040
rect 5590 -1010 5708 -992
rect 5762 -958 5880 -940
rect 5762 -992 5770 -958
rect 5804 -992 5838 -958
rect 5872 -992 5880 -958
rect 5762 -1010 5880 -992
rect 5990 -958 6108 -940
rect 5990 -992 5998 -958
rect 6032 -992 6066 -958
rect 6100 -992 6108 -958
rect 5990 -1010 6108 -992
rect 6162 -958 6280 -940
rect 8140 -908 8290 -890
rect 8140 -942 8162 -908
rect 8196 -942 8230 -908
rect 8264 -942 8290 -908
rect 6162 -992 6170 -958
rect 6204 -992 6238 -958
rect 6272 -992 6280 -958
rect 8140 -960 8290 -942
rect 9252 -908 9402 -890
rect 9252 -942 9278 -908
rect 9312 -942 9346 -908
rect 9380 -942 9402 -908
rect 9252 -960 9402 -942
rect 6162 -1010 6280 -992
rect 5362 -1092 5370 -1058
rect 5404 -1092 5438 -1058
rect 5472 -1092 5480 -1058
rect 5362 -1110 5480 -1092
rect 5590 -1058 5708 -1040
rect 5590 -1092 5598 -1058
rect 5632 -1092 5666 -1058
rect 5700 -1092 5708 -1058
rect 4562 -1192 4570 -1158
rect 4604 -1192 4638 -1158
rect 4672 -1192 4680 -1158
rect 4562 -1210 4680 -1192
rect 4790 -1158 4908 -1140
rect 4790 -1192 4798 -1158
rect 4832 -1192 4866 -1158
rect 4900 -1192 4908 -1158
rect 3762 -1292 3770 -1258
rect 3804 -1292 3838 -1258
rect 3872 -1292 3880 -1258
rect 3762 -1310 3880 -1292
rect 3990 -1258 4108 -1240
rect 3990 -1292 3998 -1258
rect 4032 -1292 4066 -1258
rect 4100 -1292 4108 -1258
rect 2962 -1392 2970 -1358
rect 3004 -1392 3038 -1358
rect 3072 -1392 3080 -1358
rect 2962 -1410 3080 -1392
rect 3190 -1358 3308 -1340
rect 3190 -1392 3198 -1358
rect 3232 -1392 3266 -1358
rect 3300 -1392 3308 -1358
rect 2162 -1492 2170 -1458
rect 2204 -1492 2238 -1458
rect 2272 -1492 2280 -1458
rect 2162 -1510 2280 -1492
rect 2390 -1458 2508 -1440
rect 2390 -1492 2398 -1458
rect 2432 -1492 2466 -1458
rect 2500 -1492 2508 -1458
rect 1362 -1592 1370 -1558
rect 1404 -1592 1438 -1558
rect 1472 -1592 1480 -1558
rect 1362 -1610 1480 -1592
rect 1590 -1558 1708 -1540
rect 1590 -1592 1598 -1558
rect 1632 -1592 1666 -1558
rect 1700 -1592 1708 -1558
rect 562 -1692 570 -1658
rect 604 -1692 638 -1658
rect 672 -1692 680 -1658
rect 562 -1710 680 -1692
rect 790 -1658 908 -1640
rect 790 -1692 798 -1658
rect 832 -1692 866 -1658
rect 900 -1692 908 -1658
rect -10 -1758 108 -1740
rect -10 -1792 -2 -1758
rect 32 -1792 66 -1758
rect 100 -1792 108 -1758
rect -10 -1810 108 -1792
rect 162 -1758 280 -1740
rect 162 -1792 170 -1758
rect 204 -1792 238 -1758
rect 272 -1792 280 -1758
rect 162 -1810 280 -1792
rect 390 -1758 508 -1740
rect 390 -1792 398 -1758
rect 432 -1792 466 -1758
rect 500 -1792 508 -1758
rect 390 -1810 508 -1792
rect 562 -1758 680 -1740
rect 790 -1710 908 -1692
rect 962 -1658 1080 -1640
rect 962 -1692 970 -1658
rect 1004 -1692 1038 -1658
rect 1072 -1692 1080 -1658
rect 962 -1710 1080 -1692
rect 1190 -1658 1308 -1640
rect 1190 -1692 1198 -1658
rect 1232 -1692 1266 -1658
rect 1300 -1692 1308 -1658
rect 1190 -1710 1308 -1692
rect 1362 -1658 1480 -1640
rect 1590 -1610 1708 -1592
rect 1762 -1558 1880 -1540
rect 1762 -1592 1770 -1558
rect 1804 -1592 1838 -1558
rect 1872 -1592 1880 -1558
rect 1762 -1610 1880 -1592
rect 1990 -1558 2108 -1540
rect 1990 -1592 1998 -1558
rect 2032 -1592 2066 -1558
rect 2100 -1592 2108 -1558
rect 1990 -1610 2108 -1592
rect 2162 -1558 2280 -1540
rect 2390 -1510 2508 -1492
rect 2562 -1458 2680 -1440
rect 2562 -1492 2570 -1458
rect 2604 -1492 2638 -1458
rect 2672 -1492 2680 -1458
rect 2562 -1510 2680 -1492
rect 2790 -1458 2908 -1440
rect 2790 -1492 2798 -1458
rect 2832 -1492 2866 -1458
rect 2900 -1492 2908 -1458
rect 2790 -1510 2908 -1492
rect 2962 -1458 3080 -1440
rect 3190 -1410 3308 -1392
rect 3362 -1358 3480 -1340
rect 3362 -1392 3370 -1358
rect 3404 -1392 3438 -1358
rect 3472 -1392 3480 -1358
rect 3362 -1410 3480 -1392
rect 3590 -1358 3708 -1340
rect 3590 -1392 3598 -1358
rect 3632 -1392 3666 -1358
rect 3700 -1392 3708 -1358
rect 3590 -1410 3708 -1392
rect 3762 -1358 3880 -1340
rect 3990 -1310 4108 -1292
rect 4162 -1258 4280 -1240
rect 4162 -1292 4170 -1258
rect 4204 -1292 4238 -1258
rect 4272 -1292 4280 -1258
rect 4162 -1310 4280 -1292
rect 4390 -1258 4508 -1240
rect 4390 -1292 4398 -1258
rect 4432 -1292 4466 -1258
rect 4500 -1292 4508 -1258
rect 4390 -1310 4508 -1292
rect 4562 -1258 4680 -1240
rect 4790 -1210 4908 -1192
rect 4962 -1158 5080 -1140
rect 4962 -1192 4970 -1158
rect 5004 -1192 5038 -1158
rect 5072 -1192 5080 -1158
rect 4962 -1210 5080 -1192
rect 5190 -1158 5308 -1140
rect 5190 -1192 5198 -1158
rect 5232 -1192 5266 -1158
rect 5300 -1192 5308 -1158
rect 5190 -1210 5308 -1192
rect 5362 -1158 5480 -1140
rect 5590 -1110 5708 -1092
rect 5762 -1058 5880 -1040
rect 5762 -1092 5770 -1058
rect 5804 -1092 5838 -1058
rect 5872 -1092 5880 -1058
rect 5762 -1110 5880 -1092
rect 5990 -1058 6108 -1040
rect 5990 -1092 5998 -1058
rect 6032 -1092 6066 -1058
rect 6100 -1092 6108 -1058
rect 5990 -1110 6108 -1092
rect 6162 -1058 6280 -1040
rect 8140 -1008 8290 -990
rect 8140 -1042 8162 -1008
rect 8196 -1042 8230 -1008
rect 8264 -1042 8290 -1008
rect 6162 -1092 6170 -1058
rect 6204 -1092 6238 -1058
rect 6272 -1092 6280 -1058
rect 8140 -1060 8290 -1042
rect 9252 -1008 9402 -990
rect 9252 -1042 9278 -1008
rect 9312 -1042 9346 -1008
rect 9380 -1042 9402 -1008
rect 9252 -1060 9402 -1042
rect 6162 -1110 6280 -1092
rect 5362 -1192 5370 -1158
rect 5404 -1192 5438 -1158
rect 5472 -1192 5480 -1158
rect 5362 -1210 5480 -1192
rect 5590 -1158 5708 -1140
rect 5590 -1192 5598 -1158
rect 5632 -1192 5666 -1158
rect 5700 -1192 5708 -1158
rect 4562 -1292 4570 -1258
rect 4604 -1292 4638 -1258
rect 4672 -1292 4680 -1258
rect 4562 -1310 4680 -1292
rect 4790 -1258 4908 -1240
rect 4790 -1292 4798 -1258
rect 4832 -1292 4866 -1258
rect 4900 -1292 4908 -1258
rect 3762 -1392 3770 -1358
rect 3804 -1392 3838 -1358
rect 3872 -1392 3880 -1358
rect 3762 -1410 3880 -1392
rect 3990 -1358 4108 -1340
rect 3990 -1392 3998 -1358
rect 4032 -1392 4066 -1358
rect 4100 -1392 4108 -1358
rect 2962 -1492 2970 -1458
rect 3004 -1492 3038 -1458
rect 3072 -1492 3080 -1458
rect 2962 -1510 3080 -1492
rect 3190 -1458 3308 -1440
rect 3190 -1492 3198 -1458
rect 3232 -1492 3266 -1458
rect 3300 -1492 3308 -1458
rect 2162 -1592 2170 -1558
rect 2204 -1592 2238 -1558
rect 2272 -1592 2280 -1558
rect 2162 -1610 2280 -1592
rect 2390 -1558 2508 -1540
rect 2390 -1592 2398 -1558
rect 2432 -1592 2466 -1558
rect 2500 -1592 2508 -1558
rect 1362 -1692 1370 -1658
rect 1404 -1692 1438 -1658
rect 1472 -1692 1480 -1658
rect 1362 -1710 1480 -1692
rect 1590 -1658 1708 -1640
rect 1590 -1692 1598 -1658
rect 1632 -1692 1666 -1658
rect 1700 -1692 1708 -1658
rect 562 -1792 570 -1758
rect 604 -1792 638 -1758
rect 672 -1792 680 -1758
rect 562 -1810 680 -1792
rect 790 -1758 908 -1740
rect 790 -1792 798 -1758
rect 832 -1792 866 -1758
rect 900 -1792 908 -1758
rect -10 -1858 108 -1840
rect -10 -1892 -2 -1858
rect 32 -1892 66 -1858
rect 100 -1892 108 -1858
rect -10 -1929 108 -1892
rect 162 -1858 280 -1840
rect 162 -1892 170 -1858
rect 204 -1892 238 -1858
rect 272 -1892 280 -1858
rect 162 -1929 280 -1892
rect 390 -1858 508 -1840
rect 390 -1892 398 -1858
rect 432 -1892 466 -1858
rect 500 -1892 508 -1858
rect 390 -1929 508 -1892
rect 562 -1858 680 -1840
rect 790 -1810 908 -1792
rect 962 -1758 1080 -1740
rect 962 -1792 970 -1758
rect 1004 -1792 1038 -1758
rect 1072 -1792 1080 -1758
rect 962 -1810 1080 -1792
rect 1190 -1758 1308 -1740
rect 1190 -1792 1198 -1758
rect 1232 -1792 1266 -1758
rect 1300 -1792 1308 -1758
rect 1190 -1810 1308 -1792
rect 1362 -1758 1480 -1740
rect 1590 -1710 1708 -1692
rect 1762 -1658 1880 -1640
rect 1762 -1692 1770 -1658
rect 1804 -1692 1838 -1658
rect 1872 -1692 1880 -1658
rect 1762 -1710 1880 -1692
rect 1990 -1658 2108 -1640
rect 1990 -1692 1998 -1658
rect 2032 -1692 2066 -1658
rect 2100 -1692 2108 -1658
rect 1990 -1710 2108 -1692
rect 2162 -1658 2280 -1640
rect 2390 -1610 2508 -1592
rect 2562 -1558 2680 -1540
rect 2562 -1592 2570 -1558
rect 2604 -1592 2638 -1558
rect 2672 -1592 2680 -1558
rect 2562 -1610 2680 -1592
rect 2790 -1558 2908 -1540
rect 2790 -1592 2798 -1558
rect 2832 -1592 2866 -1558
rect 2900 -1592 2908 -1558
rect 2790 -1610 2908 -1592
rect 2962 -1558 3080 -1540
rect 3190 -1510 3308 -1492
rect 3362 -1458 3480 -1440
rect 3362 -1492 3370 -1458
rect 3404 -1492 3438 -1458
rect 3472 -1492 3480 -1458
rect 3362 -1510 3480 -1492
rect 3590 -1458 3708 -1440
rect 3590 -1492 3598 -1458
rect 3632 -1492 3666 -1458
rect 3700 -1492 3708 -1458
rect 3590 -1510 3708 -1492
rect 3762 -1458 3880 -1440
rect 3990 -1410 4108 -1392
rect 4162 -1358 4280 -1340
rect 4162 -1392 4170 -1358
rect 4204 -1392 4238 -1358
rect 4272 -1392 4280 -1358
rect 4162 -1410 4280 -1392
rect 4390 -1358 4508 -1340
rect 4390 -1392 4398 -1358
rect 4432 -1392 4466 -1358
rect 4500 -1392 4508 -1358
rect 4390 -1410 4508 -1392
rect 4562 -1358 4680 -1340
rect 4790 -1310 4908 -1292
rect 4962 -1258 5080 -1240
rect 4962 -1292 4970 -1258
rect 5004 -1292 5038 -1258
rect 5072 -1292 5080 -1258
rect 4962 -1310 5080 -1292
rect 5190 -1258 5308 -1240
rect 5190 -1292 5198 -1258
rect 5232 -1292 5266 -1258
rect 5300 -1292 5308 -1258
rect 5190 -1310 5308 -1292
rect 5362 -1258 5480 -1240
rect 5590 -1210 5708 -1192
rect 5762 -1158 5880 -1140
rect 5762 -1192 5770 -1158
rect 5804 -1192 5838 -1158
rect 5872 -1192 5880 -1158
rect 5762 -1210 5880 -1192
rect 5990 -1158 6108 -1140
rect 5990 -1192 5998 -1158
rect 6032 -1192 6066 -1158
rect 6100 -1192 6108 -1158
rect 5990 -1210 6108 -1192
rect 6162 -1158 6280 -1140
rect 8140 -1108 8290 -1090
rect 8140 -1142 8162 -1108
rect 8196 -1142 8230 -1108
rect 8264 -1142 8290 -1108
rect 6162 -1192 6170 -1158
rect 6204 -1192 6238 -1158
rect 6272 -1192 6280 -1158
rect 8140 -1160 8290 -1142
rect 9252 -1108 9402 -1090
rect 9252 -1142 9278 -1108
rect 9312 -1142 9346 -1108
rect 9380 -1142 9402 -1108
rect 9252 -1160 9402 -1142
rect 6162 -1210 6280 -1192
rect 5362 -1292 5370 -1258
rect 5404 -1292 5438 -1258
rect 5472 -1292 5480 -1258
rect 5362 -1310 5480 -1292
rect 5590 -1258 5708 -1240
rect 5590 -1292 5598 -1258
rect 5632 -1292 5666 -1258
rect 5700 -1292 5708 -1258
rect 4562 -1392 4570 -1358
rect 4604 -1392 4638 -1358
rect 4672 -1392 4680 -1358
rect 4562 -1410 4680 -1392
rect 4790 -1358 4908 -1340
rect 4790 -1392 4798 -1358
rect 4832 -1392 4866 -1358
rect 4900 -1392 4908 -1358
rect 3762 -1492 3770 -1458
rect 3804 -1492 3838 -1458
rect 3872 -1492 3880 -1458
rect 3762 -1510 3880 -1492
rect 3990 -1458 4108 -1440
rect 3990 -1492 3998 -1458
rect 4032 -1492 4066 -1458
rect 4100 -1492 4108 -1458
rect 2962 -1592 2970 -1558
rect 3004 -1592 3038 -1558
rect 3072 -1592 3080 -1558
rect 2962 -1610 3080 -1592
rect 3190 -1558 3308 -1540
rect 3190 -1592 3198 -1558
rect 3232 -1592 3266 -1558
rect 3300 -1592 3308 -1558
rect 2162 -1692 2170 -1658
rect 2204 -1692 2238 -1658
rect 2272 -1692 2280 -1658
rect 2162 -1710 2280 -1692
rect 2390 -1658 2508 -1640
rect 2390 -1692 2398 -1658
rect 2432 -1692 2466 -1658
rect 2500 -1692 2508 -1658
rect 1362 -1792 1370 -1758
rect 1404 -1792 1438 -1758
rect 1472 -1792 1480 -1758
rect 1362 -1810 1480 -1792
rect 1590 -1758 1708 -1740
rect 1590 -1792 1598 -1758
rect 1632 -1792 1666 -1758
rect 1700 -1792 1708 -1758
rect 562 -1892 570 -1858
rect 604 -1892 638 -1858
rect 672 -1892 680 -1858
rect 562 -1929 680 -1892
rect 790 -1858 908 -1840
rect 790 -1892 798 -1858
rect 832 -1892 866 -1858
rect 900 -1892 908 -1858
rect 790 -1929 908 -1892
rect 962 -1858 1080 -1840
rect 962 -1892 970 -1858
rect 1004 -1892 1038 -1858
rect 1072 -1892 1080 -1858
rect 962 -1929 1080 -1892
rect 1190 -1858 1308 -1840
rect 1190 -1892 1198 -1858
rect 1232 -1892 1266 -1858
rect 1300 -1892 1308 -1858
rect 1190 -1929 1308 -1892
rect 1362 -1858 1480 -1840
rect 1590 -1810 1708 -1792
rect 1762 -1758 1880 -1740
rect 1762 -1792 1770 -1758
rect 1804 -1792 1838 -1758
rect 1872 -1792 1880 -1758
rect 1762 -1810 1880 -1792
rect 1990 -1758 2108 -1740
rect 1990 -1792 1998 -1758
rect 2032 -1792 2066 -1758
rect 2100 -1792 2108 -1758
rect 1990 -1810 2108 -1792
rect 2162 -1758 2280 -1740
rect 2390 -1710 2508 -1692
rect 2562 -1658 2680 -1640
rect 2562 -1692 2570 -1658
rect 2604 -1692 2638 -1658
rect 2672 -1692 2680 -1658
rect 2562 -1710 2680 -1692
rect 2790 -1658 2908 -1640
rect 2790 -1692 2798 -1658
rect 2832 -1692 2866 -1658
rect 2900 -1692 2908 -1658
rect 2790 -1710 2908 -1692
rect 2962 -1658 3080 -1640
rect 3190 -1610 3308 -1592
rect 3362 -1558 3480 -1540
rect 3362 -1592 3370 -1558
rect 3404 -1592 3438 -1558
rect 3472 -1592 3480 -1558
rect 3362 -1610 3480 -1592
rect 3590 -1558 3708 -1540
rect 3590 -1592 3598 -1558
rect 3632 -1592 3666 -1558
rect 3700 -1592 3708 -1558
rect 3590 -1610 3708 -1592
rect 3762 -1558 3880 -1540
rect 3990 -1510 4108 -1492
rect 4162 -1458 4280 -1440
rect 4162 -1492 4170 -1458
rect 4204 -1492 4238 -1458
rect 4272 -1492 4280 -1458
rect 4162 -1510 4280 -1492
rect 4390 -1458 4508 -1440
rect 4390 -1492 4398 -1458
rect 4432 -1492 4466 -1458
rect 4500 -1492 4508 -1458
rect 4390 -1510 4508 -1492
rect 4562 -1458 4680 -1440
rect 4790 -1410 4908 -1392
rect 4962 -1358 5080 -1340
rect 4962 -1392 4970 -1358
rect 5004 -1392 5038 -1358
rect 5072 -1392 5080 -1358
rect 4962 -1410 5080 -1392
rect 5190 -1358 5308 -1340
rect 5190 -1392 5198 -1358
rect 5232 -1392 5266 -1358
rect 5300 -1392 5308 -1358
rect 5190 -1410 5308 -1392
rect 5362 -1358 5480 -1340
rect 5590 -1310 5708 -1292
rect 5762 -1258 5880 -1240
rect 5762 -1292 5770 -1258
rect 5804 -1292 5838 -1258
rect 5872 -1292 5880 -1258
rect 5762 -1310 5880 -1292
rect 5990 -1258 6108 -1240
rect 5990 -1292 5998 -1258
rect 6032 -1292 6066 -1258
rect 6100 -1292 6108 -1258
rect 5990 -1310 6108 -1292
rect 6162 -1258 6280 -1240
rect 8140 -1208 8290 -1190
rect 8140 -1242 8162 -1208
rect 8196 -1242 8230 -1208
rect 8264 -1242 8290 -1208
rect 6162 -1292 6170 -1258
rect 6204 -1292 6238 -1258
rect 6272 -1292 6280 -1258
rect 8140 -1260 8290 -1242
rect 9252 -1208 9402 -1190
rect 9252 -1242 9278 -1208
rect 9312 -1242 9346 -1208
rect 9380 -1242 9402 -1208
rect 9252 -1260 9402 -1242
rect 6162 -1310 6280 -1292
rect 5362 -1392 5370 -1358
rect 5404 -1392 5438 -1358
rect 5472 -1392 5480 -1358
rect 5362 -1410 5480 -1392
rect 5590 -1358 5708 -1340
rect 5590 -1392 5598 -1358
rect 5632 -1392 5666 -1358
rect 5700 -1392 5708 -1358
rect 4562 -1492 4570 -1458
rect 4604 -1492 4638 -1458
rect 4672 -1492 4680 -1458
rect 4562 -1510 4680 -1492
rect 4790 -1458 4908 -1440
rect 4790 -1492 4798 -1458
rect 4832 -1492 4866 -1458
rect 4900 -1492 4908 -1458
rect 3762 -1592 3770 -1558
rect 3804 -1592 3838 -1558
rect 3872 -1592 3880 -1558
rect 3762 -1610 3880 -1592
rect 3990 -1558 4108 -1540
rect 3990 -1592 3998 -1558
rect 4032 -1592 4066 -1558
rect 4100 -1592 4108 -1558
rect 2962 -1692 2970 -1658
rect 3004 -1692 3038 -1658
rect 3072 -1692 3080 -1658
rect 2962 -1710 3080 -1692
rect 3190 -1658 3308 -1640
rect 3190 -1692 3198 -1658
rect 3232 -1692 3266 -1658
rect 3300 -1692 3308 -1658
rect 2162 -1792 2170 -1758
rect 2204 -1792 2238 -1758
rect 2272 -1792 2280 -1758
rect 2162 -1810 2280 -1792
rect 2390 -1758 2508 -1740
rect 2390 -1792 2398 -1758
rect 2432 -1792 2466 -1758
rect 2500 -1792 2508 -1758
rect 1362 -1892 1370 -1858
rect 1404 -1892 1438 -1858
rect 1472 -1892 1480 -1858
rect 1362 -1929 1480 -1892
rect 1590 -1858 1708 -1840
rect 1590 -1892 1598 -1858
rect 1632 -1892 1666 -1858
rect 1700 -1892 1708 -1858
rect 1590 -1929 1708 -1892
rect 1762 -1858 1880 -1840
rect 1762 -1892 1770 -1858
rect 1804 -1892 1838 -1858
rect 1872 -1892 1880 -1858
rect 1762 -1929 1880 -1892
rect 1990 -1858 2108 -1840
rect 1990 -1892 1998 -1858
rect 2032 -1892 2066 -1858
rect 2100 -1892 2108 -1858
rect 1990 -1929 2108 -1892
rect 2162 -1858 2280 -1840
rect 2390 -1810 2508 -1792
rect 2562 -1758 2680 -1740
rect 2562 -1792 2570 -1758
rect 2604 -1792 2638 -1758
rect 2672 -1792 2680 -1758
rect 2562 -1810 2680 -1792
rect 2790 -1758 2908 -1740
rect 2790 -1792 2798 -1758
rect 2832 -1792 2866 -1758
rect 2900 -1792 2908 -1758
rect 2790 -1810 2908 -1792
rect 2962 -1758 3080 -1740
rect 3190 -1710 3308 -1692
rect 3362 -1658 3480 -1640
rect 3362 -1692 3370 -1658
rect 3404 -1692 3438 -1658
rect 3472 -1692 3480 -1658
rect 3362 -1710 3480 -1692
rect 3590 -1658 3708 -1640
rect 3590 -1692 3598 -1658
rect 3632 -1692 3666 -1658
rect 3700 -1692 3708 -1658
rect 3590 -1710 3708 -1692
rect 3762 -1658 3880 -1640
rect 3990 -1610 4108 -1592
rect 4162 -1558 4280 -1540
rect 4162 -1592 4170 -1558
rect 4204 -1592 4238 -1558
rect 4272 -1592 4280 -1558
rect 4162 -1610 4280 -1592
rect 4390 -1558 4508 -1540
rect 4390 -1592 4398 -1558
rect 4432 -1592 4466 -1558
rect 4500 -1592 4508 -1558
rect 4390 -1610 4508 -1592
rect 4562 -1558 4680 -1540
rect 4790 -1510 4908 -1492
rect 4962 -1458 5080 -1440
rect 4962 -1492 4970 -1458
rect 5004 -1492 5038 -1458
rect 5072 -1492 5080 -1458
rect 4962 -1510 5080 -1492
rect 5190 -1458 5308 -1440
rect 5190 -1492 5198 -1458
rect 5232 -1492 5266 -1458
rect 5300 -1492 5308 -1458
rect 5190 -1510 5308 -1492
rect 5362 -1458 5480 -1440
rect 5590 -1410 5708 -1392
rect 5762 -1358 5880 -1340
rect 5762 -1392 5770 -1358
rect 5804 -1392 5838 -1358
rect 5872 -1392 5880 -1358
rect 5762 -1410 5880 -1392
rect 5990 -1358 6108 -1340
rect 5990 -1392 5998 -1358
rect 6032 -1392 6066 -1358
rect 6100 -1392 6108 -1358
rect 5990 -1410 6108 -1392
rect 6162 -1358 6280 -1340
rect 8140 -1308 8290 -1290
rect 8140 -1342 8162 -1308
rect 8196 -1342 8230 -1308
rect 8264 -1342 8290 -1308
rect 6162 -1392 6170 -1358
rect 6204 -1392 6238 -1358
rect 6272 -1392 6280 -1358
rect 8140 -1360 8290 -1342
rect 9252 -1308 9402 -1290
rect 9252 -1342 9278 -1308
rect 9312 -1342 9346 -1308
rect 9380 -1342 9402 -1308
rect 9252 -1360 9402 -1342
rect 6162 -1410 6280 -1392
rect 5362 -1492 5370 -1458
rect 5404 -1492 5438 -1458
rect 5472 -1492 5480 -1458
rect 5362 -1510 5480 -1492
rect 5590 -1458 5708 -1440
rect 5590 -1492 5598 -1458
rect 5632 -1492 5666 -1458
rect 5700 -1492 5708 -1458
rect 4562 -1592 4570 -1558
rect 4604 -1592 4638 -1558
rect 4672 -1592 4680 -1558
rect 4562 -1610 4680 -1592
rect 4790 -1558 4908 -1540
rect 4790 -1592 4798 -1558
rect 4832 -1592 4866 -1558
rect 4900 -1592 4908 -1558
rect 3762 -1692 3770 -1658
rect 3804 -1692 3838 -1658
rect 3872 -1692 3880 -1658
rect 3762 -1710 3880 -1692
rect 3990 -1658 4108 -1640
rect 3990 -1692 3998 -1658
rect 4032 -1692 4066 -1658
rect 4100 -1692 4108 -1658
rect 2962 -1792 2970 -1758
rect 3004 -1792 3038 -1758
rect 3072 -1792 3080 -1758
rect 2962 -1810 3080 -1792
rect 3190 -1758 3308 -1740
rect 3190 -1792 3198 -1758
rect 3232 -1792 3266 -1758
rect 3300 -1792 3308 -1758
rect 2162 -1892 2170 -1858
rect 2204 -1892 2238 -1858
rect 2272 -1892 2280 -1858
rect 2162 -1929 2280 -1892
rect 2390 -1858 2508 -1840
rect 2390 -1892 2398 -1858
rect 2432 -1892 2466 -1858
rect 2500 -1892 2508 -1858
rect 2390 -1929 2508 -1892
rect 2562 -1858 2680 -1840
rect 2562 -1892 2570 -1858
rect 2604 -1892 2638 -1858
rect 2672 -1892 2680 -1858
rect 2562 -1929 2680 -1892
rect 2790 -1858 2908 -1840
rect 2790 -1892 2798 -1858
rect 2832 -1892 2866 -1858
rect 2900 -1892 2908 -1858
rect 2790 -1929 2908 -1892
rect 2962 -1858 3080 -1840
rect 3190 -1810 3308 -1792
rect 3362 -1758 3480 -1740
rect 3362 -1792 3370 -1758
rect 3404 -1792 3438 -1758
rect 3472 -1792 3480 -1758
rect 3362 -1810 3480 -1792
rect 3590 -1758 3708 -1740
rect 3590 -1792 3598 -1758
rect 3632 -1792 3666 -1758
rect 3700 -1792 3708 -1758
rect 3590 -1810 3708 -1792
rect 3762 -1758 3880 -1740
rect 3990 -1710 4108 -1692
rect 4162 -1658 4280 -1640
rect 4162 -1692 4170 -1658
rect 4204 -1692 4238 -1658
rect 4272 -1692 4280 -1658
rect 4162 -1710 4280 -1692
rect 4390 -1658 4508 -1640
rect 4390 -1692 4398 -1658
rect 4432 -1692 4466 -1658
rect 4500 -1692 4508 -1658
rect 4390 -1710 4508 -1692
rect 4562 -1658 4680 -1640
rect 4790 -1610 4908 -1592
rect 4962 -1558 5080 -1540
rect 4962 -1592 4970 -1558
rect 5004 -1592 5038 -1558
rect 5072 -1592 5080 -1558
rect 4962 -1610 5080 -1592
rect 5190 -1558 5308 -1540
rect 5190 -1592 5198 -1558
rect 5232 -1592 5266 -1558
rect 5300 -1592 5308 -1558
rect 5190 -1610 5308 -1592
rect 5362 -1558 5480 -1540
rect 5590 -1510 5708 -1492
rect 5762 -1458 5880 -1440
rect 5762 -1492 5770 -1458
rect 5804 -1492 5838 -1458
rect 5872 -1492 5880 -1458
rect 5762 -1510 5880 -1492
rect 5990 -1458 6108 -1440
rect 5990 -1492 5998 -1458
rect 6032 -1492 6066 -1458
rect 6100 -1492 6108 -1458
rect 5990 -1510 6108 -1492
rect 6162 -1458 6280 -1440
rect 8140 -1408 8290 -1390
rect 8140 -1442 8162 -1408
rect 8196 -1442 8230 -1408
rect 8264 -1442 8290 -1408
rect 6162 -1492 6170 -1458
rect 6204 -1492 6238 -1458
rect 6272 -1492 6280 -1458
rect 8140 -1460 8290 -1442
rect 9252 -1408 9402 -1390
rect 9252 -1442 9278 -1408
rect 9312 -1442 9346 -1408
rect 9380 -1442 9402 -1408
rect 9252 -1460 9402 -1442
rect 6162 -1510 6280 -1492
rect 5362 -1592 5370 -1558
rect 5404 -1592 5438 -1558
rect 5472 -1592 5480 -1558
rect 5362 -1610 5480 -1592
rect 5590 -1558 5708 -1540
rect 5590 -1592 5598 -1558
rect 5632 -1592 5666 -1558
rect 5700 -1592 5708 -1558
rect 4562 -1692 4570 -1658
rect 4604 -1692 4638 -1658
rect 4672 -1692 4680 -1658
rect 4562 -1710 4680 -1692
rect 4790 -1658 4908 -1640
rect 4790 -1692 4798 -1658
rect 4832 -1692 4866 -1658
rect 4900 -1692 4908 -1658
rect 3762 -1792 3770 -1758
rect 3804 -1792 3838 -1758
rect 3872 -1792 3880 -1758
rect 3762 -1810 3880 -1792
rect 3990 -1758 4108 -1740
rect 3990 -1792 3998 -1758
rect 4032 -1792 4066 -1758
rect 4100 -1792 4108 -1758
rect 2962 -1892 2970 -1858
rect 3004 -1892 3038 -1858
rect 3072 -1892 3080 -1858
rect 2962 -1929 3080 -1892
rect 3190 -1858 3308 -1840
rect 3190 -1892 3198 -1858
rect 3232 -1892 3266 -1858
rect 3300 -1892 3308 -1858
rect 3190 -1929 3308 -1892
rect 3362 -1858 3480 -1840
rect 3362 -1892 3370 -1858
rect 3404 -1892 3438 -1858
rect 3472 -1892 3480 -1858
rect 3362 -1929 3480 -1892
rect 3590 -1858 3708 -1840
rect 3590 -1892 3598 -1858
rect 3632 -1892 3666 -1858
rect 3700 -1892 3708 -1858
rect 3590 -1929 3708 -1892
rect 3762 -1858 3880 -1840
rect 3990 -1810 4108 -1792
rect 4162 -1758 4280 -1740
rect 4162 -1792 4170 -1758
rect 4204 -1792 4238 -1758
rect 4272 -1792 4280 -1758
rect 4162 -1810 4280 -1792
rect 4390 -1758 4508 -1740
rect 4390 -1792 4398 -1758
rect 4432 -1792 4466 -1758
rect 4500 -1792 4508 -1758
rect 4390 -1810 4508 -1792
rect 4562 -1758 4680 -1740
rect 4790 -1710 4908 -1692
rect 4962 -1658 5080 -1640
rect 4962 -1692 4970 -1658
rect 5004 -1692 5038 -1658
rect 5072 -1692 5080 -1658
rect 4962 -1710 5080 -1692
rect 5190 -1658 5308 -1640
rect 5190 -1692 5198 -1658
rect 5232 -1692 5266 -1658
rect 5300 -1692 5308 -1658
rect 5190 -1710 5308 -1692
rect 5362 -1658 5480 -1640
rect 5590 -1610 5708 -1592
rect 5762 -1558 5880 -1540
rect 5762 -1592 5770 -1558
rect 5804 -1592 5838 -1558
rect 5872 -1592 5880 -1558
rect 5762 -1610 5880 -1592
rect 5990 -1558 6108 -1540
rect 5990 -1592 5998 -1558
rect 6032 -1592 6066 -1558
rect 6100 -1592 6108 -1558
rect 5990 -1610 6108 -1592
rect 6162 -1558 6280 -1540
rect 8140 -1508 8290 -1490
rect 8140 -1542 8162 -1508
rect 8196 -1542 8230 -1508
rect 8264 -1542 8290 -1508
rect 6162 -1592 6170 -1558
rect 6204 -1592 6238 -1558
rect 6272 -1592 6280 -1558
rect 8140 -1560 8290 -1542
rect 9252 -1508 9402 -1490
rect 9252 -1542 9278 -1508
rect 9312 -1542 9346 -1508
rect 9380 -1542 9402 -1508
rect 9252 -1560 9402 -1542
rect 6162 -1610 6280 -1592
rect 5362 -1692 5370 -1658
rect 5404 -1692 5438 -1658
rect 5472 -1692 5480 -1658
rect 5362 -1710 5480 -1692
rect 5590 -1658 5708 -1640
rect 5590 -1692 5598 -1658
rect 5632 -1692 5666 -1658
rect 5700 -1692 5708 -1658
rect 4562 -1792 4570 -1758
rect 4604 -1792 4638 -1758
rect 4672 -1792 4680 -1758
rect 4562 -1810 4680 -1792
rect 4790 -1758 4908 -1740
rect 4790 -1792 4798 -1758
rect 4832 -1792 4866 -1758
rect 4900 -1792 4908 -1758
rect 3762 -1892 3770 -1858
rect 3804 -1892 3838 -1858
rect 3872 -1892 3880 -1858
rect 3762 -1929 3880 -1892
rect 3990 -1858 4108 -1840
rect 3990 -1892 3998 -1858
rect 4032 -1892 4066 -1858
rect 4100 -1892 4108 -1858
rect 3990 -1929 4108 -1892
rect 4162 -1858 4280 -1840
rect 4162 -1892 4170 -1858
rect 4204 -1892 4238 -1858
rect 4272 -1892 4280 -1858
rect 4162 -1929 4280 -1892
rect 4390 -1858 4508 -1840
rect 4390 -1892 4398 -1858
rect 4432 -1892 4466 -1858
rect 4500 -1892 4508 -1858
rect 4390 -1929 4508 -1892
rect 4562 -1858 4680 -1840
rect 4790 -1810 4908 -1792
rect 4962 -1758 5080 -1740
rect 4962 -1792 4970 -1758
rect 5004 -1792 5038 -1758
rect 5072 -1792 5080 -1758
rect 4962 -1810 5080 -1792
rect 5190 -1758 5308 -1740
rect 5190 -1792 5198 -1758
rect 5232 -1792 5266 -1758
rect 5300 -1792 5308 -1758
rect 5190 -1810 5308 -1792
rect 5362 -1758 5480 -1740
rect 5590 -1710 5708 -1692
rect 5762 -1658 5880 -1640
rect 5762 -1692 5770 -1658
rect 5804 -1692 5838 -1658
rect 5872 -1692 5880 -1658
rect 5762 -1710 5880 -1692
rect 5990 -1658 6108 -1640
rect 5990 -1692 5998 -1658
rect 6032 -1692 6066 -1658
rect 6100 -1692 6108 -1658
rect 5990 -1710 6108 -1692
rect 6162 -1658 6280 -1640
rect 8140 -1608 8290 -1590
rect 8140 -1642 8162 -1608
rect 8196 -1642 8230 -1608
rect 8264 -1642 8290 -1608
rect 6162 -1692 6170 -1658
rect 6204 -1692 6238 -1658
rect 6272 -1692 6280 -1658
rect 8140 -1660 8290 -1642
rect 9252 -1608 9402 -1590
rect 9252 -1642 9278 -1608
rect 9312 -1642 9346 -1608
rect 9380 -1642 9402 -1608
rect 9252 -1660 9402 -1642
rect 6162 -1710 6280 -1692
rect 5362 -1792 5370 -1758
rect 5404 -1792 5438 -1758
rect 5472 -1792 5480 -1758
rect 5362 -1810 5480 -1792
rect 5590 -1758 5708 -1740
rect 5590 -1792 5598 -1758
rect 5632 -1792 5666 -1758
rect 5700 -1792 5708 -1758
rect 4562 -1892 4570 -1858
rect 4604 -1892 4638 -1858
rect 4672 -1892 4680 -1858
rect 4562 -1929 4680 -1892
rect 4790 -1858 4908 -1840
rect 4790 -1892 4798 -1858
rect 4832 -1892 4866 -1858
rect 4900 -1892 4908 -1858
rect 4790 -1929 4908 -1892
rect 4962 -1858 5080 -1840
rect 4962 -1892 4970 -1858
rect 5004 -1892 5038 -1858
rect 5072 -1892 5080 -1858
rect 4962 -1929 5080 -1892
rect 5190 -1858 5308 -1840
rect 5190 -1892 5198 -1858
rect 5232 -1892 5266 -1858
rect 5300 -1892 5308 -1858
rect 5190 -1929 5308 -1892
rect 5362 -1858 5480 -1840
rect 5590 -1810 5708 -1792
rect 5762 -1758 5880 -1740
rect 5762 -1792 5770 -1758
rect 5804 -1792 5838 -1758
rect 5872 -1792 5880 -1758
rect 5762 -1810 5880 -1792
rect 5990 -1758 6108 -1740
rect 5990 -1792 5998 -1758
rect 6032 -1792 6066 -1758
rect 6100 -1792 6108 -1758
rect 5990 -1810 6108 -1792
rect 6162 -1758 6280 -1740
rect 8140 -1708 8290 -1690
rect 8140 -1742 8162 -1708
rect 8196 -1742 8230 -1708
rect 8264 -1742 8290 -1708
rect 6162 -1792 6170 -1758
rect 6204 -1792 6238 -1758
rect 6272 -1792 6280 -1758
rect 8140 -1760 8290 -1742
rect 9252 -1708 9402 -1690
rect 9252 -1742 9278 -1708
rect 9312 -1742 9346 -1708
rect 9380 -1742 9402 -1708
rect 9252 -1760 9402 -1742
rect 6162 -1810 6280 -1792
rect 5362 -1892 5370 -1858
rect 5404 -1892 5438 -1858
rect 5472 -1892 5480 -1858
rect 5362 -1929 5480 -1892
rect 5590 -1858 5708 -1840
rect 5590 -1892 5598 -1858
rect 5632 -1892 5666 -1858
rect 5700 -1892 5708 -1858
rect 5590 -1929 5708 -1892
rect 5762 -1858 5880 -1840
rect 5762 -1892 5770 -1858
rect 5804 -1892 5838 -1858
rect 5872 -1892 5880 -1858
rect 5762 -1929 5880 -1892
rect 5990 -1858 6108 -1840
rect 5990 -1892 5998 -1858
rect 6032 -1892 6066 -1858
rect 6100 -1892 6108 -1858
rect 5990 -1929 6108 -1892
rect 6162 -1858 6280 -1840
rect 8140 -1808 8290 -1790
rect 8140 -1842 8162 -1808
rect 8196 -1842 8230 -1808
rect 8264 -1842 8290 -1808
rect 6162 -1892 6170 -1858
rect 6204 -1892 6238 -1858
rect 6272 -1892 6280 -1858
rect 6162 -1929 6280 -1892
rect 8140 -1879 8290 -1842
rect 9252 -1808 9402 -1790
rect 9252 -1842 9278 -1808
rect 9312 -1842 9346 -1808
rect 9380 -1842 9402 -1808
rect 9252 -1879 9402 -1842
<< pdiff >>
rect 8416 -8 8716 29
rect 8416 -42 8447 -8
rect 8481 -42 8515 -8
rect 8549 -42 8583 -8
rect 8617 -42 8651 -8
rect 8685 -42 8716 -8
rect 8416 -60 8716 -42
rect 8826 -8 9126 29
rect 8826 -42 8857 -8
rect 8891 -42 8925 -8
rect 8959 -42 8993 -8
rect 9027 -42 9061 -8
rect 9095 -42 9126 -8
rect 8826 -60 9126 -42
rect 8416 -108 8716 -90
rect 8416 -142 8447 -108
rect 8481 -142 8515 -108
rect 8549 -142 8583 -108
rect 8617 -142 8651 -108
rect 8685 -142 8716 -108
rect 8416 -160 8716 -142
rect 8826 -108 9126 -90
rect 8826 -142 8857 -108
rect 8891 -142 8925 -108
rect 8959 -142 8993 -108
rect 9027 -142 9061 -108
rect 9095 -142 9126 -108
rect 8826 -160 9126 -142
rect 8416 -208 8716 -190
rect 8416 -242 8447 -208
rect 8481 -242 8515 -208
rect 8549 -242 8583 -208
rect 8617 -242 8651 -208
rect 8685 -242 8716 -208
rect 8416 -260 8716 -242
rect 8826 -208 9126 -190
rect 8826 -242 8857 -208
rect 8891 -242 8925 -208
rect 8959 -242 8993 -208
rect 9027 -242 9061 -208
rect 9095 -242 9126 -208
rect 8826 -260 9126 -242
rect -94 -363 -30 -330
rect -94 -397 -82 -363
rect -48 -397 -30 -363
rect -94 -431 -30 -397
rect -94 -465 -82 -431
rect -48 -465 -30 -431
rect -94 -498 -30 -465
rect 0 -363 70 -330
rect 0 -397 18 -363
rect 52 -397 70 -363
rect 0 -431 70 -397
rect 0 -465 18 -431
rect 52 -465 70 -431
rect 0 -498 70 -465
rect 100 -363 170 -330
rect 100 -397 118 -363
rect 152 -397 170 -363
rect 100 -431 170 -397
rect 100 -465 118 -431
rect 152 -465 170 -431
rect 100 -498 170 -465
rect 200 -363 270 -330
rect 200 -397 218 -363
rect 252 -397 270 -363
rect 200 -431 270 -397
rect 200 -465 218 -431
rect 252 -465 270 -431
rect 200 -498 270 -465
rect 300 -363 370 -330
rect 300 -397 318 -363
rect 352 -397 370 -363
rect 300 -431 370 -397
rect 300 -465 318 -431
rect 352 -465 370 -431
rect 300 -498 370 -465
rect 400 -363 470 -330
rect 400 -397 418 -363
rect 452 -397 470 -363
rect 400 -431 470 -397
rect 400 -465 418 -431
rect 452 -465 470 -431
rect 400 -498 470 -465
rect 500 -363 570 -330
rect 500 -397 518 -363
rect 552 -397 570 -363
rect 500 -431 570 -397
rect 500 -465 518 -431
rect 552 -465 570 -431
rect 500 -498 570 -465
rect 600 -363 670 -330
rect 600 -397 618 -363
rect 652 -397 670 -363
rect 600 -431 670 -397
rect 600 -465 618 -431
rect 652 -465 670 -431
rect 600 -498 670 -465
rect 700 -363 770 -330
rect 700 -397 718 -363
rect 752 -397 770 -363
rect 700 -431 770 -397
rect 700 -465 718 -431
rect 752 -465 770 -431
rect 700 -498 770 -465
rect 800 -363 870 -330
rect 800 -397 818 -363
rect 852 -397 870 -363
rect 800 -431 870 -397
rect 800 -465 818 -431
rect 852 -465 870 -431
rect 800 -498 870 -465
rect 900 -363 970 -330
rect 900 -397 918 -363
rect 952 -397 970 -363
rect 900 -431 970 -397
rect 900 -465 918 -431
rect 952 -465 970 -431
rect 900 -498 970 -465
rect 1000 -363 1070 -330
rect 1000 -397 1018 -363
rect 1052 -397 1070 -363
rect 1000 -431 1070 -397
rect 1000 -465 1018 -431
rect 1052 -465 1070 -431
rect 1000 -498 1070 -465
rect 1100 -363 1170 -330
rect 1100 -397 1118 -363
rect 1152 -397 1170 -363
rect 1100 -431 1170 -397
rect 1100 -465 1118 -431
rect 1152 -465 1170 -431
rect 1100 -498 1170 -465
rect 1200 -363 1270 -330
rect 1200 -397 1218 -363
rect 1252 -397 1270 -363
rect 1200 -431 1270 -397
rect 1200 -465 1218 -431
rect 1252 -465 1270 -431
rect 1200 -498 1270 -465
rect 1300 -363 1370 -330
rect 1300 -397 1318 -363
rect 1352 -397 1370 -363
rect 1300 -431 1370 -397
rect 1300 -465 1318 -431
rect 1352 -465 1370 -431
rect 1300 -498 1370 -465
rect 1400 -363 1470 -330
rect 1400 -397 1418 -363
rect 1452 -397 1470 -363
rect 1400 -431 1470 -397
rect 1400 -465 1418 -431
rect 1452 -465 1470 -431
rect 1400 -498 1470 -465
rect 1500 -363 1570 -330
rect 1500 -397 1518 -363
rect 1552 -397 1570 -363
rect 1500 -431 1570 -397
rect 1500 -465 1518 -431
rect 1552 -465 1570 -431
rect 1500 -498 1570 -465
rect 1600 -363 1670 -330
rect 1600 -397 1618 -363
rect 1652 -397 1670 -363
rect 1600 -431 1670 -397
rect 1600 -465 1618 -431
rect 1652 -465 1670 -431
rect 1600 -498 1670 -465
rect 1700 -363 1770 -330
rect 1700 -397 1718 -363
rect 1752 -397 1770 -363
rect 1700 -431 1770 -397
rect 1700 -465 1718 -431
rect 1752 -465 1770 -431
rect 1700 -498 1770 -465
rect 1800 -363 1870 -330
rect 1800 -397 1818 -363
rect 1852 -397 1870 -363
rect 1800 -431 1870 -397
rect 1800 -465 1818 -431
rect 1852 -465 1870 -431
rect 1800 -498 1870 -465
rect 1900 -363 1970 -330
rect 1900 -397 1918 -363
rect 1952 -397 1970 -363
rect 1900 -431 1970 -397
rect 1900 -465 1918 -431
rect 1952 -465 1970 -431
rect 1900 -498 1970 -465
rect 2000 -363 2070 -330
rect 2000 -397 2018 -363
rect 2052 -397 2070 -363
rect 2000 -431 2070 -397
rect 2000 -465 2018 -431
rect 2052 -465 2070 -431
rect 2000 -498 2070 -465
rect 2100 -363 2170 -330
rect 2100 -397 2118 -363
rect 2152 -397 2170 -363
rect 2100 -431 2170 -397
rect 2100 -465 2118 -431
rect 2152 -465 2170 -431
rect 2100 -498 2170 -465
rect 2200 -363 2270 -330
rect 2200 -397 2218 -363
rect 2252 -397 2270 -363
rect 2200 -431 2270 -397
rect 2200 -465 2218 -431
rect 2252 -465 2270 -431
rect 2200 -498 2270 -465
rect 2300 -363 2370 -330
rect 2300 -397 2318 -363
rect 2352 -397 2370 -363
rect 2300 -431 2370 -397
rect 2300 -465 2318 -431
rect 2352 -465 2370 -431
rect 2300 -498 2370 -465
rect 2400 -363 2470 -330
rect 2400 -397 2418 -363
rect 2452 -397 2470 -363
rect 2400 -431 2470 -397
rect 2400 -465 2418 -431
rect 2452 -465 2470 -431
rect 2400 -498 2470 -465
rect 2500 -363 2570 -330
rect 2500 -397 2518 -363
rect 2552 -397 2570 -363
rect 2500 -431 2570 -397
rect 2500 -465 2518 -431
rect 2552 -465 2570 -431
rect 2500 -498 2570 -465
rect 2600 -363 2670 -330
rect 2600 -397 2618 -363
rect 2652 -397 2670 -363
rect 2600 -431 2670 -397
rect 2600 -465 2618 -431
rect 2652 -465 2670 -431
rect 2600 -498 2670 -465
rect 2700 -363 2770 -330
rect 2700 -397 2718 -363
rect 2752 -397 2770 -363
rect 2700 -431 2770 -397
rect 2700 -465 2718 -431
rect 2752 -465 2770 -431
rect 2700 -498 2770 -465
rect 2800 -363 2870 -330
rect 2800 -397 2818 -363
rect 2852 -397 2870 -363
rect 2800 -431 2870 -397
rect 2800 -465 2818 -431
rect 2852 -465 2870 -431
rect 2800 -498 2870 -465
rect 2900 -363 2970 -330
rect 2900 -397 2918 -363
rect 2952 -397 2970 -363
rect 2900 -431 2970 -397
rect 2900 -465 2918 -431
rect 2952 -465 2970 -431
rect 2900 -498 2970 -465
rect 3000 -363 3070 -330
rect 3000 -397 3018 -363
rect 3052 -397 3070 -363
rect 3000 -431 3070 -397
rect 3000 -465 3018 -431
rect 3052 -465 3070 -431
rect 3000 -498 3070 -465
rect 3100 -363 3170 -330
rect 3100 -397 3118 -363
rect 3152 -397 3170 -363
rect 3100 -431 3170 -397
rect 3100 -465 3118 -431
rect 3152 -465 3170 -431
rect 3100 -498 3170 -465
rect 3200 -363 3270 -330
rect 3200 -397 3218 -363
rect 3252 -397 3270 -363
rect 3200 -431 3270 -397
rect 3200 -465 3218 -431
rect 3252 -465 3270 -431
rect 3200 -498 3270 -465
rect 3300 -363 3370 -330
rect 3300 -397 3318 -363
rect 3352 -397 3370 -363
rect 3300 -431 3370 -397
rect 3300 -465 3318 -431
rect 3352 -465 3370 -431
rect 3300 -498 3370 -465
rect 3400 -363 3470 -330
rect 3400 -397 3418 -363
rect 3452 -397 3470 -363
rect 3400 -431 3470 -397
rect 3400 -465 3418 -431
rect 3452 -465 3470 -431
rect 3400 -498 3470 -465
rect 3500 -363 3570 -330
rect 3500 -397 3518 -363
rect 3552 -397 3570 -363
rect 3500 -431 3570 -397
rect 3500 -465 3518 -431
rect 3552 -465 3570 -431
rect 3500 -498 3570 -465
rect 3600 -363 3670 -330
rect 3600 -397 3618 -363
rect 3652 -397 3670 -363
rect 3600 -431 3670 -397
rect 3600 -465 3618 -431
rect 3652 -465 3670 -431
rect 3600 -498 3670 -465
rect 3700 -363 3770 -330
rect 3700 -397 3718 -363
rect 3752 -397 3770 -363
rect 3700 -431 3770 -397
rect 3700 -465 3718 -431
rect 3752 -465 3770 -431
rect 3700 -498 3770 -465
rect 3800 -363 3870 -330
rect 3800 -397 3818 -363
rect 3852 -397 3870 -363
rect 3800 -431 3870 -397
rect 3800 -465 3818 -431
rect 3852 -465 3870 -431
rect 3800 -498 3870 -465
rect 3900 -363 3970 -330
rect 3900 -397 3918 -363
rect 3952 -397 3970 -363
rect 3900 -431 3970 -397
rect 3900 -465 3918 -431
rect 3952 -465 3970 -431
rect 3900 -498 3970 -465
rect 4000 -363 4070 -330
rect 4000 -397 4018 -363
rect 4052 -397 4070 -363
rect 4000 -431 4070 -397
rect 4000 -465 4018 -431
rect 4052 -465 4070 -431
rect 4000 -498 4070 -465
rect 4100 -363 4170 -330
rect 4100 -397 4118 -363
rect 4152 -397 4170 -363
rect 4100 -431 4170 -397
rect 4100 -465 4118 -431
rect 4152 -465 4170 -431
rect 4100 -498 4170 -465
rect 4200 -363 4270 -330
rect 4200 -397 4218 -363
rect 4252 -397 4270 -363
rect 4200 -431 4270 -397
rect 4200 -465 4218 -431
rect 4252 -465 4270 -431
rect 4200 -498 4270 -465
rect 4300 -363 4370 -330
rect 4300 -397 4318 -363
rect 4352 -397 4370 -363
rect 4300 -431 4370 -397
rect 4300 -465 4318 -431
rect 4352 -465 4370 -431
rect 4300 -498 4370 -465
rect 4400 -363 4470 -330
rect 4400 -397 4418 -363
rect 4452 -397 4470 -363
rect 4400 -431 4470 -397
rect 4400 -465 4418 -431
rect 4452 -465 4470 -431
rect 4400 -498 4470 -465
rect 4500 -363 4570 -330
rect 4500 -397 4518 -363
rect 4552 -397 4570 -363
rect 4500 -431 4570 -397
rect 4500 -465 4518 -431
rect 4552 -465 4570 -431
rect 4500 -498 4570 -465
rect 4600 -363 4670 -330
rect 4600 -397 4618 -363
rect 4652 -397 4670 -363
rect 4600 -431 4670 -397
rect 4600 -465 4618 -431
rect 4652 -465 4670 -431
rect 4600 -498 4670 -465
rect 4700 -363 4770 -330
rect 4700 -397 4718 -363
rect 4752 -397 4770 -363
rect 4700 -431 4770 -397
rect 4700 -465 4718 -431
rect 4752 -465 4770 -431
rect 4700 -498 4770 -465
rect 4800 -363 4870 -330
rect 4800 -397 4818 -363
rect 4852 -397 4870 -363
rect 4800 -431 4870 -397
rect 4800 -465 4818 -431
rect 4852 -465 4870 -431
rect 4800 -498 4870 -465
rect 4900 -363 4970 -330
rect 4900 -397 4918 -363
rect 4952 -397 4970 -363
rect 4900 -431 4970 -397
rect 4900 -465 4918 -431
rect 4952 -465 4970 -431
rect 4900 -498 4970 -465
rect 5000 -363 5070 -330
rect 5000 -397 5018 -363
rect 5052 -397 5070 -363
rect 5000 -431 5070 -397
rect 5000 -465 5018 -431
rect 5052 -465 5070 -431
rect 5000 -498 5070 -465
rect 5100 -363 5170 -330
rect 5100 -397 5118 -363
rect 5152 -397 5170 -363
rect 5100 -431 5170 -397
rect 5100 -465 5118 -431
rect 5152 -465 5170 -431
rect 5100 -498 5170 -465
rect 5200 -363 5270 -330
rect 5200 -397 5218 -363
rect 5252 -397 5270 -363
rect 5200 -431 5270 -397
rect 5200 -465 5218 -431
rect 5252 -465 5270 -431
rect 5200 -498 5270 -465
rect 5300 -363 5370 -330
rect 5300 -397 5318 -363
rect 5352 -397 5370 -363
rect 5300 -431 5370 -397
rect 5300 -465 5318 -431
rect 5352 -465 5370 -431
rect 5300 -498 5370 -465
rect 5400 -363 5470 -330
rect 5400 -397 5418 -363
rect 5452 -397 5470 -363
rect 5400 -431 5470 -397
rect 5400 -465 5418 -431
rect 5452 -465 5470 -431
rect 5400 -498 5470 -465
rect 5500 -363 5570 -330
rect 5500 -397 5518 -363
rect 5552 -397 5570 -363
rect 5500 -431 5570 -397
rect 5500 -465 5518 -431
rect 5552 -465 5570 -431
rect 5500 -498 5570 -465
rect 5600 -363 5670 -330
rect 5600 -397 5618 -363
rect 5652 -397 5670 -363
rect 5600 -431 5670 -397
rect 5600 -465 5618 -431
rect 5652 -465 5670 -431
rect 5600 -498 5670 -465
rect 5700 -363 5770 -330
rect 5700 -397 5718 -363
rect 5752 -397 5770 -363
rect 5700 -431 5770 -397
rect 5700 -465 5718 -431
rect 5752 -465 5770 -431
rect 5700 -498 5770 -465
rect 5800 -363 5870 -330
rect 5800 -397 5818 -363
rect 5852 -397 5870 -363
rect 5800 -431 5870 -397
rect 5800 -465 5818 -431
rect 5852 -465 5870 -431
rect 5800 -498 5870 -465
rect 5900 -363 5970 -330
rect 5900 -397 5918 -363
rect 5952 -397 5970 -363
rect 5900 -431 5970 -397
rect 5900 -465 5918 -431
rect 5952 -465 5970 -431
rect 5900 -498 5970 -465
rect 6000 -363 6070 -330
rect 6000 -397 6018 -363
rect 6052 -397 6070 -363
rect 6000 -431 6070 -397
rect 6000 -465 6018 -431
rect 6052 -465 6070 -431
rect 6000 -498 6070 -465
rect 6100 -363 6170 -330
rect 6100 -397 6118 -363
rect 6152 -397 6170 -363
rect 6100 -431 6170 -397
rect 6100 -465 6118 -431
rect 6152 -465 6170 -431
rect 6100 -498 6170 -465
rect 6200 -363 6270 -330
rect 6200 -397 6218 -363
rect 6252 -397 6270 -363
rect 6200 -431 6270 -397
rect 6200 -465 6218 -431
rect 6252 -465 6270 -431
rect 6200 -498 6270 -465
rect 6300 -363 6364 -330
rect 8416 -308 8716 -290
rect 8416 -342 8447 -308
rect 8481 -342 8515 -308
rect 8549 -342 8583 -308
rect 8617 -342 8651 -308
rect 8685 -342 8716 -308
rect 8416 -360 8716 -342
rect 8826 -308 9126 -290
rect 8826 -342 8857 -308
rect 8891 -342 8925 -308
rect 8959 -342 8993 -308
rect 9027 -342 9061 -308
rect 9095 -342 9126 -308
rect 8826 -360 9126 -342
rect 6300 -397 6318 -363
rect 6352 -397 6364 -363
rect 6300 -431 6364 -397
rect 6300 -465 6318 -431
rect 6352 -465 6364 -431
rect 8416 -408 8716 -390
rect 8416 -442 8447 -408
rect 8481 -442 8515 -408
rect 8549 -442 8583 -408
rect 8617 -442 8651 -408
rect 8685 -442 8716 -408
rect 8416 -460 8716 -442
rect 8826 -408 9126 -390
rect 8826 -442 8857 -408
rect 8891 -442 8925 -408
rect 8959 -442 8993 -408
rect 9027 -442 9061 -408
rect 9095 -442 9126 -408
rect 8826 -460 9126 -442
rect 6300 -498 6364 -465
rect 8416 -508 8716 -490
rect 8416 -542 8447 -508
rect 8481 -542 8515 -508
rect 8549 -542 8583 -508
rect 8617 -542 8651 -508
rect 8685 -542 8716 -508
rect 8416 -560 8716 -542
rect 8826 -508 9126 -490
rect 8826 -542 8857 -508
rect 8891 -542 8925 -508
rect 8959 -542 8993 -508
rect 9027 -542 9061 -508
rect 9095 -542 9126 -508
rect 8826 -560 9126 -542
rect -38 -683 15 -658
rect -38 -717 -30 -683
rect 4 -717 15 -683
rect -38 -742 15 -717
rect 107 -683 163 -658
rect 107 -717 118 -683
rect 152 -717 163 -683
rect 107 -742 163 -717
rect 255 -683 308 -658
rect 255 -717 266 -683
rect 300 -717 308 -683
rect 255 -742 308 -717
rect 362 -683 415 -658
rect 362 -717 370 -683
rect 404 -717 415 -683
rect 362 -742 415 -717
rect 507 -683 563 -658
rect 507 -717 518 -683
rect 552 -717 563 -683
rect 507 -742 563 -717
rect 655 -683 708 -658
rect 655 -717 666 -683
rect 700 -717 708 -683
rect 655 -742 708 -717
rect 762 -683 815 -658
rect 762 -717 770 -683
rect 804 -717 815 -683
rect 762 -742 815 -717
rect 907 -683 963 -658
rect 907 -717 918 -683
rect 952 -717 963 -683
rect 907 -742 963 -717
rect 1055 -683 1108 -658
rect 1055 -717 1066 -683
rect 1100 -717 1108 -683
rect 1055 -742 1108 -717
rect 1162 -683 1215 -658
rect 1162 -717 1170 -683
rect 1204 -717 1215 -683
rect 1162 -742 1215 -717
rect 1307 -683 1363 -658
rect 1307 -717 1318 -683
rect 1352 -717 1363 -683
rect 1307 -742 1363 -717
rect 1455 -683 1508 -658
rect 1455 -717 1466 -683
rect 1500 -717 1508 -683
rect 1455 -742 1508 -717
rect 1562 -683 1615 -658
rect 1562 -717 1570 -683
rect 1604 -717 1615 -683
rect 1562 -742 1615 -717
rect 1707 -683 1763 -658
rect 1707 -717 1718 -683
rect 1752 -717 1763 -683
rect 1707 -742 1763 -717
rect 1855 -683 1908 -658
rect 1855 -717 1866 -683
rect 1900 -717 1908 -683
rect 1855 -742 1908 -717
rect 1962 -683 2015 -658
rect 1962 -717 1970 -683
rect 2004 -717 2015 -683
rect 1962 -742 2015 -717
rect 2107 -683 2163 -658
rect 2107 -717 2118 -683
rect 2152 -717 2163 -683
rect 2107 -742 2163 -717
rect 2255 -683 2308 -658
rect 2255 -717 2266 -683
rect 2300 -717 2308 -683
rect 2255 -742 2308 -717
rect 2362 -683 2415 -658
rect 2362 -717 2370 -683
rect 2404 -717 2415 -683
rect 2362 -742 2415 -717
rect 2507 -683 2563 -658
rect 2507 -717 2518 -683
rect 2552 -717 2563 -683
rect 2507 -742 2563 -717
rect 2655 -683 2708 -658
rect 2655 -717 2666 -683
rect 2700 -717 2708 -683
rect 2655 -742 2708 -717
rect 2762 -683 2815 -658
rect 2762 -717 2770 -683
rect 2804 -717 2815 -683
rect 2762 -742 2815 -717
rect 2907 -683 2963 -658
rect 2907 -717 2918 -683
rect 2952 -717 2963 -683
rect 2907 -742 2963 -717
rect 3055 -683 3108 -658
rect 3055 -717 3066 -683
rect 3100 -717 3108 -683
rect 3055 -742 3108 -717
rect 3162 -683 3215 -658
rect 3162 -717 3170 -683
rect 3204 -717 3215 -683
rect 3162 -742 3215 -717
rect 3307 -683 3363 -658
rect 3307 -717 3318 -683
rect 3352 -717 3363 -683
rect 3307 -742 3363 -717
rect 3455 -683 3508 -658
rect 3455 -717 3466 -683
rect 3500 -717 3508 -683
rect 3455 -742 3508 -717
rect 3562 -683 3615 -658
rect 3562 -717 3570 -683
rect 3604 -717 3615 -683
rect 3562 -742 3615 -717
rect 3707 -683 3763 -658
rect 3707 -717 3718 -683
rect 3752 -717 3763 -683
rect 3707 -742 3763 -717
rect 3855 -683 3908 -658
rect 3855 -717 3866 -683
rect 3900 -717 3908 -683
rect 3855 -742 3908 -717
rect 3962 -683 4015 -658
rect 3962 -717 3970 -683
rect 4004 -717 4015 -683
rect 3962 -742 4015 -717
rect 4107 -683 4163 -658
rect 4107 -717 4118 -683
rect 4152 -717 4163 -683
rect 4107 -742 4163 -717
rect 4255 -683 4308 -658
rect 4255 -717 4266 -683
rect 4300 -717 4308 -683
rect 4255 -742 4308 -717
rect 4362 -683 4415 -658
rect 4362 -717 4370 -683
rect 4404 -717 4415 -683
rect 4362 -742 4415 -717
rect 4507 -683 4563 -658
rect 4507 -717 4518 -683
rect 4552 -717 4563 -683
rect 4507 -742 4563 -717
rect 4655 -683 4708 -658
rect 4655 -717 4666 -683
rect 4700 -717 4708 -683
rect 4655 -742 4708 -717
rect 4762 -683 4815 -658
rect 4762 -717 4770 -683
rect 4804 -717 4815 -683
rect 4762 -742 4815 -717
rect 4907 -683 4963 -658
rect 4907 -717 4918 -683
rect 4952 -717 4963 -683
rect 4907 -742 4963 -717
rect 5055 -683 5108 -658
rect 5055 -717 5066 -683
rect 5100 -717 5108 -683
rect 5055 -742 5108 -717
rect 5162 -683 5215 -658
rect 5162 -717 5170 -683
rect 5204 -717 5215 -683
rect 5162 -742 5215 -717
rect 5307 -683 5363 -658
rect 5307 -717 5318 -683
rect 5352 -717 5363 -683
rect 5307 -742 5363 -717
rect 5455 -683 5508 -658
rect 5455 -717 5466 -683
rect 5500 -717 5508 -683
rect 5455 -742 5508 -717
rect 5562 -683 5615 -658
rect 5562 -717 5570 -683
rect 5604 -717 5615 -683
rect 5562 -742 5615 -717
rect 5707 -683 5763 -658
rect 5707 -717 5718 -683
rect 5752 -717 5763 -683
rect 5707 -742 5763 -717
rect 5855 -683 5908 -658
rect 5855 -717 5866 -683
rect 5900 -717 5908 -683
rect 5855 -742 5908 -717
rect 5962 -683 6015 -658
rect 5962 -717 5970 -683
rect 6004 -717 6015 -683
rect 5962 -742 6015 -717
rect 6107 -683 6163 -658
rect 6107 -717 6118 -683
rect 6152 -717 6163 -683
rect 6107 -742 6163 -717
rect 6255 -683 6308 -658
rect 8416 -608 8716 -590
rect 8416 -642 8447 -608
rect 8481 -642 8515 -608
rect 8549 -642 8583 -608
rect 8617 -642 8651 -608
rect 8685 -642 8716 -608
rect 8416 -660 8716 -642
rect 8826 -608 9126 -590
rect 8826 -642 8857 -608
rect 8891 -642 8925 -608
rect 8959 -642 8993 -608
rect 9027 -642 9061 -608
rect 9095 -642 9126 -608
rect 8826 -660 9126 -642
rect 6255 -717 6266 -683
rect 6300 -717 6308 -683
rect 6255 -742 6308 -717
rect 8416 -708 8716 -690
rect 8416 -742 8447 -708
rect 8481 -742 8515 -708
rect 8549 -742 8583 -708
rect 8617 -742 8651 -708
rect 8685 -742 8716 -708
rect 8416 -760 8716 -742
rect 8826 -708 9126 -690
rect 8826 -742 8857 -708
rect 8891 -742 8925 -708
rect 8959 -742 8993 -708
rect 9027 -742 9061 -708
rect 9095 -742 9126 -708
rect 8826 -760 9126 -742
rect 8416 -808 8716 -790
rect 8416 -842 8447 -808
rect 8481 -842 8515 -808
rect 8549 -842 8583 -808
rect 8617 -842 8651 -808
rect 8685 -842 8716 -808
rect 8416 -860 8716 -842
rect 8826 -808 9126 -790
rect 8826 -842 8857 -808
rect 8891 -842 8925 -808
rect 8959 -842 8993 -808
rect 9027 -842 9061 -808
rect 9095 -842 9126 -808
rect 8826 -860 9126 -842
rect 8416 -908 8716 -890
rect 8416 -942 8447 -908
rect 8481 -942 8515 -908
rect 8549 -942 8583 -908
rect 8617 -942 8651 -908
rect 8685 -942 8716 -908
rect 8416 -960 8716 -942
rect 8826 -908 9126 -890
rect 8826 -942 8857 -908
rect 8891 -942 8925 -908
rect 8959 -942 8993 -908
rect 9027 -942 9061 -908
rect 9095 -942 9126 -908
rect 8826 -960 9126 -942
rect 8416 -1008 8716 -990
rect 8416 -1042 8447 -1008
rect 8481 -1042 8515 -1008
rect 8549 -1042 8583 -1008
rect 8617 -1042 8651 -1008
rect 8685 -1042 8716 -1008
rect 8416 -1060 8716 -1042
rect 8826 -1008 9126 -990
rect 8826 -1042 8857 -1008
rect 8891 -1042 8925 -1008
rect 8959 -1042 8993 -1008
rect 9027 -1042 9061 -1008
rect 9095 -1042 9126 -1008
rect 8826 -1060 9126 -1042
rect 8416 -1108 8716 -1090
rect 8416 -1142 8447 -1108
rect 8481 -1142 8515 -1108
rect 8549 -1142 8583 -1108
rect 8617 -1142 8651 -1108
rect 8685 -1142 8716 -1108
rect 8416 -1160 8716 -1142
rect 8826 -1108 9126 -1090
rect 8826 -1142 8857 -1108
rect 8891 -1142 8925 -1108
rect 8959 -1142 8993 -1108
rect 9027 -1142 9061 -1108
rect 9095 -1142 9126 -1108
rect 8826 -1160 9126 -1142
rect 8416 -1208 8716 -1190
rect 8416 -1242 8447 -1208
rect 8481 -1242 8515 -1208
rect 8549 -1242 8583 -1208
rect 8617 -1242 8651 -1208
rect 8685 -1242 8716 -1208
rect 8416 -1260 8716 -1242
rect 8826 -1208 9126 -1190
rect 8826 -1242 8857 -1208
rect 8891 -1242 8925 -1208
rect 8959 -1242 8993 -1208
rect 9027 -1242 9061 -1208
rect 9095 -1242 9126 -1208
rect 8826 -1260 9126 -1242
rect 8416 -1308 8716 -1290
rect 8416 -1342 8447 -1308
rect 8481 -1342 8515 -1308
rect 8549 -1342 8583 -1308
rect 8617 -1342 8651 -1308
rect 8685 -1342 8716 -1308
rect 8416 -1360 8716 -1342
rect 8826 -1308 9126 -1290
rect 8826 -1342 8857 -1308
rect 8891 -1342 8925 -1308
rect 8959 -1342 8993 -1308
rect 9027 -1342 9061 -1308
rect 9095 -1342 9126 -1308
rect 8826 -1360 9126 -1342
rect 8416 -1408 8716 -1390
rect 8416 -1442 8447 -1408
rect 8481 -1442 8515 -1408
rect 8549 -1442 8583 -1408
rect 8617 -1442 8651 -1408
rect 8685 -1442 8716 -1408
rect 8416 -1460 8716 -1442
rect 8826 -1408 9126 -1390
rect 8826 -1442 8857 -1408
rect 8891 -1442 8925 -1408
rect 8959 -1442 8993 -1408
rect 9027 -1442 9061 -1408
rect 9095 -1442 9126 -1408
rect 8826 -1460 9126 -1442
rect 8416 -1508 8716 -1490
rect 8416 -1542 8447 -1508
rect 8481 -1542 8515 -1508
rect 8549 -1542 8583 -1508
rect 8617 -1542 8651 -1508
rect 8685 -1542 8716 -1508
rect 8416 -1560 8716 -1542
rect 8826 -1508 9126 -1490
rect 8826 -1542 8857 -1508
rect 8891 -1542 8925 -1508
rect 8959 -1542 8993 -1508
rect 9027 -1542 9061 -1508
rect 9095 -1542 9126 -1508
rect 8826 -1560 9126 -1542
rect 8416 -1608 8716 -1590
rect 8416 -1642 8447 -1608
rect 8481 -1642 8515 -1608
rect 8549 -1642 8583 -1608
rect 8617 -1642 8651 -1608
rect 8685 -1642 8716 -1608
rect 8416 -1660 8716 -1642
rect 8826 -1608 9126 -1590
rect 8826 -1642 8857 -1608
rect 8891 -1642 8925 -1608
rect 8959 -1642 8993 -1608
rect 9027 -1642 9061 -1608
rect 9095 -1642 9126 -1608
rect 8826 -1660 9126 -1642
rect 8416 -1708 8716 -1690
rect 8416 -1742 8447 -1708
rect 8481 -1742 8515 -1708
rect 8549 -1742 8583 -1708
rect 8617 -1742 8651 -1708
rect 8685 -1742 8716 -1708
rect 8416 -1760 8716 -1742
rect 8826 -1708 9126 -1690
rect 8826 -1742 8857 -1708
rect 8891 -1742 8925 -1708
rect 8959 -1742 8993 -1708
rect 9027 -1742 9061 -1708
rect 9095 -1742 9126 -1708
rect 8826 -1760 9126 -1742
rect 8416 -1808 8716 -1790
rect 8416 -1842 8447 -1808
rect 8481 -1842 8515 -1808
rect 8549 -1842 8583 -1808
rect 8617 -1842 8651 -1808
rect 8685 -1842 8716 -1808
rect 8416 -1879 8716 -1842
rect 8826 -1808 9126 -1790
rect 8826 -1842 8857 -1808
rect 8891 -1842 8925 -1808
rect 8959 -1842 8993 -1808
rect 9027 -1842 9061 -1808
rect 9095 -1842 9126 -1808
rect 8826 -1879 9126 -1842
<< ndiffc >>
rect 118 9733 152 9767
rect 218 9733 252 9767
rect 518 9733 552 9767
rect 618 9733 652 9767
rect 918 9733 952 9767
rect 1018 9733 1052 9767
rect 1118 9733 1152 9767
rect 1418 9733 1452 9767
rect 1512 9733 1546 9767
rect 218 9593 252 9627
rect 318 9593 352 9627
rect 518 9593 552 9627
rect 612 9593 646 9627
rect 118 9453 152 9487
rect 218 9453 252 9487
rect 318 9453 352 9487
rect 412 9453 446 9487
rect 1624 9733 1658 9767
rect 1718 9733 1752 9767
rect 1918 9733 1952 9767
rect 2018 9733 2052 9767
rect 2112 9733 2146 9767
rect 724 9593 758 9627
rect 818 9593 852 9627
rect 1218 9593 1252 9627
rect 1318 9593 1352 9627
rect 1418 9593 1452 9627
rect 1518 9593 1552 9627
rect 1618 9593 1652 9627
rect 1718 9593 1752 9627
rect 2018 9593 2052 9627
rect 2112 9593 2146 9627
rect 524 9453 558 9487
rect 618 9453 652 9487
rect 718 9453 752 9487
rect 818 9453 852 9487
rect 912 9453 946 9487
rect 1024 9453 1058 9487
rect 1112 9453 1146 9487
rect 1224 9453 1258 9487
rect 1318 9453 1352 9487
rect 1618 9453 1652 9487
rect 1712 9453 1746 9487
rect 418 9313 452 9347
rect 518 9313 552 9347
rect 618 9313 652 9347
rect 718 9313 752 9347
rect 918 9313 952 9347
rect 1018 9313 1052 9347
rect 1118 9313 1152 9347
rect 1218 9313 1252 9347
rect 1518 9313 1552 9347
rect 1618 9313 1652 9347
rect 1712 9313 1746 9347
rect 24 9173 58 9207
rect 118 9173 152 9207
rect 218 9173 252 9207
rect 318 9173 352 9207
rect 418 9173 452 9207
rect 618 9173 652 9207
rect 718 9173 752 9207
rect 818 9173 852 9207
rect 918 9173 952 9207
rect 1018 9173 1052 9207
rect 1218 9173 1252 9207
rect 1318 9173 1352 9207
rect 1418 9173 1452 9207
rect 1512 9173 1546 9207
rect 118 9033 152 9067
rect 218 9033 252 9067
rect 518 9033 552 9067
rect 612 9033 646 9067
rect 1824 9453 1858 9487
rect 1918 9453 1952 9487
rect 2012 9453 2046 9487
rect 2224 9733 2258 9767
rect 2318 9733 2352 9767
rect 2618 9733 2652 9767
rect 2712 9733 2746 9767
rect 2224 9593 2258 9627
rect 2312 9593 2346 9627
rect 2124 9453 2158 9487
rect 2218 9453 2252 9487
rect 2312 9453 2346 9487
rect 2824 9733 2858 9767
rect 2918 9733 2952 9767
rect 3118 9733 3152 9767
rect 3212 9733 3246 9767
rect 2424 9593 2458 9627
rect 2518 9593 2552 9627
rect 2818 9593 2852 9627
rect 2912 9593 2946 9627
rect 2424 9453 2458 9487
rect 2512 9453 2546 9487
rect 2624 9453 2658 9487
rect 2712 9453 2746 9487
rect 3324 9733 3358 9767
rect 3418 9733 3452 9767
rect 3512 9733 3546 9767
rect 3624 9733 3658 9767
rect 3718 9733 3752 9767
rect 3818 9733 3852 9767
rect 4018 9733 4052 9767
rect 4118 9733 4152 9767
rect 4218 9733 4252 9767
rect 4818 9733 4852 9767
rect 4918 9733 4952 9767
rect 5318 9733 5352 9767
rect 5412 9733 5446 9767
rect 3024 9593 3058 9627
rect 3118 9593 3152 9627
rect 3218 9593 3252 9627
rect 3318 9593 3352 9627
rect 3418 9593 3452 9627
rect 3518 9593 3552 9627
rect 3618 9593 3652 9627
rect 3918 9593 3952 9627
rect 4012 9593 4046 9627
rect 2824 9453 2858 9487
rect 2918 9453 2952 9487
rect 3418 9453 3452 9487
rect 3518 9453 3552 9487
rect 3618 9453 3652 9487
rect 3818 9453 3852 9487
rect 3918 9453 3952 9487
rect 4012 9453 4046 9487
rect 5524 9733 5558 9767
rect 5618 9733 5652 9767
rect 5712 9733 5746 9767
rect 5824 9733 5858 9767
rect 5912 9733 5946 9767
rect 4124 9593 4158 9627
rect 4218 9593 4252 9627
rect 4318 9593 4352 9627
rect 4618 9593 4652 9627
rect 4718 9593 4752 9627
rect 4818 9593 4852 9627
rect 4918 9593 4952 9627
rect 5518 9593 5552 9627
rect 5618 9593 5652 9627
rect 5718 9593 5752 9627
rect 5818 9593 5852 9627
rect 5912 9593 5946 9627
rect 4124 9453 4158 9487
rect 4218 9453 4252 9487
rect 4318 9453 4352 9487
rect 4418 9453 4452 9487
rect 4512 9453 4546 9487
rect 1824 9313 1858 9347
rect 1918 9313 1952 9347
rect 2018 9313 2052 9347
rect 2718 9313 2752 9347
rect 2818 9313 2852 9347
rect 2918 9313 2952 9347
rect 3218 9313 3252 9347
rect 3318 9313 3352 9347
rect 3518 9313 3552 9347
rect 3618 9313 3652 9347
rect 3718 9313 3752 9347
rect 3818 9313 3852 9347
rect 4018 9313 4052 9347
rect 4112 9313 4146 9347
rect 1624 9173 1658 9207
rect 1718 9173 1752 9207
rect 1818 9173 1852 9207
rect 2018 9173 2052 9207
rect 2118 9173 2152 9207
rect 2218 9173 2252 9207
rect 2318 9173 2352 9207
rect 2412 9173 2446 9207
rect 724 9033 758 9067
rect 818 9033 852 9067
rect 918 9033 952 9067
rect 1118 9033 1152 9067
rect 1218 9033 1252 9067
rect 1518 9033 1552 9067
rect 1618 9033 1652 9067
rect 1712 9033 1746 9067
rect 1824 9033 1858 9067
rect 1912 9033 1946 9067
rect 2524 9173 2558 9207
rect 2618 9173 2652 9207
rect 2718 9173 2752 9207
rect 3318 9173 3352 9207
rect 3418 9173 3452 9207
rect 3718 9173 3752 9207
rect 3818 9173 3852 9207
rect 3918 9173 3952 9207
rect 4012 9173 4046 9207
rect 2024 9033 2058 9067
rect 2118 9033 2152 9067
rect 2418 9033 2452 9067
rect 2518 9033 2552 9067
rect 2612 9033 2646 9067
rect 218 8893 252 8927
rect 318 8893 352 8927
rect 418 8893 452 8927
rect 918 8893 952 8927
rect 1018 8893 1052 8927
rect 1118 8893 1152 8927
rect 1218 8893 1252 8927
rect 1318 8893 1352 8927
rect 1418 8893 1452 8927
rect 1518 8893 1552 8927
rect 1918 8893 1952 8927
rect 2018 8893 2052 8927
rect 2118 8893 2152 8927
rect 2218 8893 2252 8927
rect 2518 8893 2552 8927
rect 2612 8893 2646 8927
rect 24 8753 58 8787
rect 118 8753 152 8787
rect 212 8753 246 8787
rect 324 8753 358 8787
rect 418 8753 452 8787
rect 618 8753 652 8787
rect 718 8753 752 8787
rect 918 8753 952 8787
rect 1018 8753 1052 8787
rect 1118 8753 1152 8787
rect 1218 8753 1252 8787
rect 1318 8753 1352 8787
rect 1518 8753 1552 8787
rect 1618 8753 1652 8787
rect 1718 8753 1752 8787
rect 1918 8753 1952 8787
rect 2018 8753 2052 8787
rect 2118 8753 2152 8787
rect 2218 8753 2252 8787
rect 2318 8753 2352 8787
rect 2418 8753 2452 8787
rect 2518 8753 2552 8787
rect 2612 8753 2646 8787
rect 218 8523 252 8557
rect 318 8523 352 8557
rect 518 8523 552 8557
rect 618 8523 652 8557
rect 718 8523 752 8557
rect 812 8523 846 8557
rect 924 8523 958 8557
rect 1012 8523 1046 8557
rect 2724 9033 2758 9067
rect 2812 9033 2846 9067
rect 2924 9033 2958 9067
rect 3018 9033 3052 9067
rect 3118 9033 3152 9067
rect 3212 9033 3246 9067
rect 4624 9453 4658 9487
rect 4718 9453 4752 9487
rect 4812 9453 4846 9487
rect 4924 9453 4958 9487
rect 5012 9453 5046 9487
rect 5124 9453 5158 9487
rect 5212 9453 5246 9487
rect 5324 9453 5358 9487
rect 5418 9453 5452 9487
rect 5518 9453 5552 9487
rect 5612 9453 5646 9487
rect 5724 9453 5758 9487
rect 5812 9453 5846 9487
rect 6024 9733 6058 9767
rect 6118 9733 6152 9767
rect 6218 9733 6252 9767
rect 6318 9733 6352 9767
rect 6412 9733 6446 9767
rect 6524 9748 6558 9782
rect 6618 9733 6652 9767
rect 6712 9718 6746 9752
rect 6828 9733 6862 9767
rect 6928 9733 6962 9767
rect 7028 9733 7062 9767
rect 7128 9733 7162 9767
rect 7228 9733 7262 9767
rect 7328 9733 7362 9767
rect 7428 9733 7462 9767
rect 6024 9593 6058 9627
rect 6118 9593 6152 9627
rect 6318 9593 6352 9627
rect 6412 9593 6446 9627
rect 6524 9608 6558 9642
rect 6618 9593 6652 9627
rect 6712 9578 6746 9612
rect 6828 9593 6862 9627
rect 6928 9593 6962 9627
rect 7028 9593 7062 9627
rect 7128 9593 7162 9627
rect 7228 9593 7262 9627
rect 7328 9593 7362 9627
rect 7428 9593 7462 9627
rect 5924 9453 5958 9487
rect 6018 9453 6052 9487
rect 6112 9453 6146 9487
rect 6224 9453 6258 9487
rect 6318 9453 6352 9487
rect 6412 9453 6446 9487
rect 6524 9468 6558 9502
rect 6618 9453 6652 9487
rect 6712 9438 6746 9472
rect 6828 9453 6862 9487
rect 6928 9453 6962 9487
rect 7028 9453 7062 9487
rect 7128 9453 7162 9487
rect 7228 9453 7262 9487
rect 7328 9453 7362 9487
rect 7428 9453 7462 9487
rect 4224 9313 4258 9347
rect 4318 9313 4352 9347
rect 4518 9313 4552 9347
rect 4618 9313 4652 9347
rect 4818 9313 4852 9347
rect 4918 9313 4952 9347
rect 5118 9313 5152 9347
rect 5218 9313 5252 9347
rect 5318 9313 5352 9347
rect 5418 9313 5452 9347
rect 5518 9313 5552 9347
rect 5818 9313 5852 9347
rect 5918 9313 5952 9347
rect 6118 9313 6152 9347
rect 6218 9313 6252 9347
rect 6318 9313 6352 9347
rect 6412 9313 6446 9347
rect 6524 9328 6558 9362
rect 6618 9313 6652 9347
rect 6712 9298 6746 9332
rect 6828 9313 6862 9347
rect 6928 9313 6962 9347
rect 7028 9313 7062 9347
rect 7128 9313 7162 9347
rect 7228 9313 7262 9347
rect 7328 9313 7362 9347
rect 7428 9313 7462 9347
rect 4124 9173 4158 9207
rect 4218 9173 4252 9207
rect 4418 9173 4452 9207
rect 4518 9173 4552 9207
rect 4918 9173 4952 9207
rect 5012 9173 5046 9207
rect 3324 9033 3358 9067
rect 3418 9033 3452 9067
rect 3518 9033 3552 9067
rect 3618 9033 3652 9067
rect 4018 9033 4052 9067
rect 4118 9033 4152 9067
rect 4218 9033 4252 9067
rect 4418 9033 4452 9067
rect 4512 9033 4546 9067
rect 2724 8893 2758 8927
rect 2818 8893 2852 8927
rect 3018 8893 3052 8927
rect 3118 8893 3152 8927
rect 3818 8893 3852 8927
rect 3918 8893 3952 8927
rect 4118 8893 4152 8927
rect 4218 8893 4252 8927
rect 4318 8893 4352 8927
rect 4412 8893 4446 8927
rect 2724 8753 2758 8787
rect 2818 8753 2852 8787
rect 3018 8753 3052 8787
rect 3112 8753 3146 8787
rect 1124 8523 1158 8557
rect 1218 8523 1252 8557
rect 1818 8523 1852 8557
rect 1918 8523 1952 8557
rect 2018 8523 2052 8557
rect 2118 8523 2152 8557
rect 2318 8523 2352 8557
rect 2418 8523 2452 8557
rect 2618 8523 2652 8557
rect 2712 8523 2746 8557
rect 24 8383 58 8417
rect 118 8383 152 8417
rect 418 8383 452 8417
rect 518 8383 552 8417
rect 618 8383 652 8417
rect 718 8383 752 8417
rect 818 8383 852 8417
rect 1118 8383 1152 8417
rect 1218 8383 1252 8417
rect 1312 8383 1346 8417
rect 118 8243 152 8277
rect 218 8243 252 8277
rect 318 8243 352 8277
rect 518 8243 552 8277
rect 612 8243 646 8277
rect 724 8243 758 8277
rect 812 8243 846 8277
rect 1424 8383 1458 8417
rect 1518 8383 1552 8417
rect 1618 8383 1652 8417
rect 1718 8383 1752 8417
rect 1812 8383 1846 8417
rect 1924 8383 1958 8417
rect 2012 8383 2046 8417
rect 924 8243 958 8277
rect 1018 8243 1052 8277
rect 1418 8243 1452 8277
rect 1518 8243 1552 8277
rect 1618 8243 1652 8277
rect 1818 8243 1852 8277
rect 1912 8243 1946 8277
rect 218 8103 252 8137
rect 318 8103 352 8137
rect 518 8103 552 8137
rect 618 8103 652 8137
rect 1018 8103 1052 8137
rect 1118 8103 1152 8137
rect 1212 8103 1246 8137
rect 118 7963 152 7997
rect 212 7963 246 7997
rect 324 7963 358 7997
rect 418 7963 452 7997
rect 618 7963 652 7997
rect 718 7963 752 7997
rect 818 7963 852 7997
rect 918 7963 952 7997
rect 1012 7963 1046 7997
rect 24 7823 58 7857
rect 118 7823 152 7857
rect 218 7823 252 7857
rect 318 7823 352 7857
rect 518 7823 552 7857
rect 612 7823 646 7857
rect 724 7823 758 7857
rect 812 7823 846 7857
rect 2124 8383 2158 8417
rect 2218 8383 2252 8417
rect 2312 8383 2346 8417
rect 2024 8243 2058 8277
rect 2118 8243 2152 8277
rect 2218 8243 2252 8277
rect 2312 8243 2346 8277
rect 4624 9033 4658 9067
rect 4712 9033 4746 9067
rect 4524 8893 4558 8927
rect 4612 8893 4646 8927
rect 5124 9173 5158 9207
rect 5218 9173 5252 9207
rect 5318 9173 5352 9207
rect 5412 9173 5446 9207
rect 4824 9033 4858 9067
rect 4918 9033 4952 9067
rect 5118 9033 5152 9067
rect 5212 9033 5246 9067
rect 4724 8893 4758 8927
rect 4812 8893 4846 8927
rect 5524 9173 5558 9207
rect 5618 9173 5652 9207
rect 5712 9173 5746 9207
rect 5824 9173 5858 9207
rect 5918 9173 5952 9207
rect 6118 9173 6152 9207
rect 6218 9173 6252 9207
rect 6318 9173 6352 9207
rect 6524 9188 6558 9222
rect 6618 9173 6652 9207
rect 6712 9158 6746 9192
rect 6828 9173 6862 9207
rect 6928 9173 6962 9207
rect 7028 9173 7062 9207
rect 7128 9173 7162 9207
rect 7228 9173 7262 9207
rect 7328 9173 7362 9207
rect 7428 9173 7462 9207
rect 5324 9033 5358 9067
rect 5418 9033 5452 9067
rect 5818 9033 5852 9067
rect 5918 9033 5952 9067
rect 6018 9033 6052 9067
rect 6218 9033 6252 9067
rect 6318 9033 6352 9067
rect 6412 9033 6446 9067
rect 6524 9048 6558 9082
rect 6618 9033 6652 9067
rect 6712 9018 6746 9052
rect 6828 9033 6862 9067
rect 6928 9033 6962 9067
rect 7028 9033 7062 9067
rect 7128 9033 7162 9067
rect 7228 9033 7262 9067
rect 7328 9033 7362 9067
rect 7428 9033 7462 9067
rect 4924 8893 4958 8927
rect 5018 8893 5052 8927
rect 5118 8893 5152 8927
rect 5218 8893 5252 8927
rect 5318 8893 5352 8927
rect 5518 8893 5552 8927
rect 5612 8893 5646 8927
rect 3224 8753 3258 8787
rect 3318 8753 3352 8787
rect 3418 8753 3452 8787
rect 3618 8753 3652 8787
rect 3718 8753 3752 8787
rect 3918 8753 3952 8787
rect 4018 8753 4052 8787
rect 4118 8753 4152 8787
rect 4518 8753 4552 8787
rect 4618 8753 4652 8787
rect 4718 8753 4752 8787
rect 5118 8753 5152 8787
rect 5218 8753 5252 8787
rect 5418 8753 5452 8787
rect 5512 8753 5546 8787
rect 2824 8523 2858 8557
rect 2918 8523 2952 8557
rect 3118 8523 3152 8557
rect 3218 8523 3252 8557
rect 3312 8523 3346 8557
rect 3424 8523 3458 8557
rect 3512 8523 3546 8557
rect 3624 8523 3658 8557
rect 3718 8523 3752 8557
rect 3918 8523 3952 8557
rect 4012 8523 4046 8557
rect 2424 8383 2458 8417
rect 2518 8383 2552 8417
rect 2618 8383 2652 8417
rect 2718 8383 2752 8417
rect 2818 8383 2852 8417
rect 3018 8383 3052 8417
rect 3118 8383 3152 8417
rect 3218 8383 3252 8417
rect 3418 8383 3452 8417
rect 3518 8383 3552 8417
rect 3618 8383 3652 8417
rect 3718 8383 3752 8417
rect 3812 8383 3846 8417
rect 2424 8243 2458 8277
rect 2512 8243 2546 8277
rect 2624 8243 2658 8277
rect 2718 8243 2752 8277
rect 2918 8243 2952 8277
rect 3018 8243 3052 8277
rect 3112 8243 3146 8277
rect 1324 8103 1358 8137
rect 1418 8103 1452 8137
rect 1518 8103 1552 8137
rect 1918 8103 1952 8137
rect 2018 8103 2052 8137
rect 2118 8103 2152 8137
rect 2218 8103 2252 8137
rect 2318 8103 2352 8137
rect 2518 8103 2552 8137
rect 2612 8103 2646 8137
rect 1124 7963 1158 7997
rect 1218 7963 1252 7997
rect 1312 7963 1346 7997
rect 1424 7963 1458 7997
rect 1518 7963 1552 7997
rect 1618 7963 1652 7997
rect 1712 7963 1746 7997
rect 924 7823 958 7857
rect 1018 7823 1052 7857
rect 1118 7823 1152 7857
rect 1218 7823 1252 7857
rect 1318 7823 1352 7857
rect 1412 7823 1446 7857
rect 1524 7823 1558 7857
rect 1612 7823 1646 7857
rect 24 7683 58 7717
rect 118 7683 152 7717
rect 218 7683 252 7717
rect 518 7683 552 7717
rect 618 7683 652 7717
rect 1118 7683 1152 7717
rect 1218 7683 1252 7717
rect 1418 7683 1452 7717
rect 1512 7683 1546 7717
rect 24 7543 58 7577
rect 118 7543 152 7577
rect 218 7543 252 7577
rect 918 7543 952 7577
rect 1012 7543 1046 7577
rect 1124 7543 1158 7577
rect 1218 7543 1252 7577
rect 1312 7543 1346 7577
rect 1824 7963 1858 7997
rect 1918 7963 1952 7997
rect 2012 7963 2046 7997
rect 2724 8103 2758 8137
rect 2812 8103 2846 8137
rect 2124 7963 2158 7997
rect 2218 7963 2252 7997
rect 2318 7963 2352 7997
rect 2518 7963 2552 7997
rect 2618 7963 2652 7997
rect 2712 7963 2746 7997
rect 1724 7823 1758 7857
rect 1818 7823 1852 7857
rect 2018 7823 2052 7857
rect 2118 7823 2152 7857
rect 2318 7823 2352 7857
rect 2418 7823 2452 7857
rect 2512 7823 2546 7857
rect 1624 7683 1658 7717
rect 1712 7683 1746 7717
rect 3224 8243 3258 8277
rect 3318 8243 3352 8277
rect 3418 8243 3452 8277
rect 3512 8243 3546 8277
rect 4124 8523 4158 8557
rect 4218 8523 4252 8557
rect 4312 8523 4346 8557
rect 4424 8523 4458 8557
rect 4518 8523 4552 8557
rect 4618 8523 4652 8557
rect 4712 8523 4746 8557
rect 3924 8383 3958 8417
rect 4018 8383 4052 8417
rect 4218 8383 4252 8417
rect 4318 8383 4352 8417
rect 4518 8383 4552 8417
rect 4618 8383 4652 8417
rect 4712 8383 4746 8417
rect 5724 8893 5758 8927
rect 5818 8893 5852 8927
rect 6018 8893 6052 8927
rect 6112 8893 6146 8927
rect 5624 8753 5658 8787
rect 5718 8753 5752 8787
rect 5818 8753 5852 8787
rect 5912 8753 5946 8787
rect 4824 8523 4858 8557
rect 4918 8523 4952 8557
rect 5018 8523 5052 8557
rect 5218 8523 5252 8557
rect 5318 8523 5352 8557
rect 5418 8523 5452 8557
rect 5518 8523 5552 8557
rect 5612 8523 5646 8557
rect 4824 8383 4858 8417
rect 4912 8383 4946 8417
rect 6224 8893 6258 8927
rect 6318 8893 6352 8927
rect 6524 8908 6558 8942
rect 6618 8893 6652 8927
rect 6712 8878 6746 8912
rect 6828 8893 6862 8927
rect 6928 8893 6962 8927
rect 7028 8893 7062 8927
rect 7128 8893 7162 8927
rect 7228 8893 7262 8927
rect 7328 8893 7362 8927
rect 7428 8893 7462 8927
rect 6024 8753 6058 8787
rect 6118 8753 6152 8787
rect 6218 8753 6252 8787
rect 6318 8753 6352 8787
rect 6524 8768 6558 8802
rect 6618 8753 6652 8787
rect 6712 8738 6746 8772
rect 6828 8753 6862 8787
rect 6928 8753 6962 8787
rect 7028 8753 7062 8787
rect 7128 8753 7162 8787
rect 7228 8753 7262 8787
rect 7328 8753 7362 8787
rect 7428 8753 7462 8787
rect 5724 8523 5758 8557
rect 5818 8523 5852 8557
rect 6218 8523 6252 8557
rect 6318 8523 6352 8557
rect 6524 8538 6558 8572
rect 6618 8523 6652 8557
rect 6712 8508 6746 8542
rect 6828 8523 6862 8557
rect 6928 8523 6962 8557
rect 7028 8523 7062 8557
rect 7128 8523 7162 8557
rect 7228 8523 7262 8557
rect 7328 8523 7362 8557
rect 7428 8523 7462 8557
rect 5024 8383 5058 8417
rect 5118 8383 5152 8417
rect 5218 8383 5252 8417
rect 5318 8383 5352 8417
rect 5718 8383 5752 8417
rect 5812 8383 5846 8417
rect 5924 8383 5958 8417
rect 6018 8383 6052 8417
rect 6118 8383 6152 8417
rect 6318 8383 6352 8417
rect 6412 8383 6446 8417
rect 6524 8398 6558 8432
rect 6618 8383 6652 8417
rect 6712 8368 6746 8402
rect 6828 8383 6862 8417
rect 6928 8383 6962 8417
rect 7028 8383 7062 8417
rect 7128 8383 7162 8417
rect 7228 8383 7262 8417
rect 7328 8383 7362 8417
rect 7428 8383 7462 8417
rect 3624 8243 3658 8277
rect 3718 8243 3752 8277
rect 3818 8243 3852 8277
rect 4218 8243 4252 8277
rect 4318 8243 4352 8277
rect 4618 8243 4652 8277
rect 4718 8243 4752 8277
rect 5018 8243 5052 8277
rect 5118 8243 5152 8277
rect 5218 8243 5252 8277
rect 5518 8243 5552 8277
rect 5618 8243 5652 8277
rect 6118 8243 6152 8277
rect 6218 8243 6252 8277
rect 6318 8243 6352 8277
rect 6412 8243 6446 8277
rect 6524 8258 6558 8292
rect 6618 8243 6652 8277
rect 6712 8228 6746 8262
rect 6828 8243 6862 8277
rect 6928 8243 6962 8277
rect 7028 8243 7062 8277
rect 7128 8243 7162 8277
rect 7228 8243 7262 8277
rect 7328 8243 7362 8277
rect 7428 8243 7462 8277
rect 2924 8103 2958 8137
rect 3018 8103 3052 8137
rect 3518 8103 3552 8137
rect 3618 8103 3652 8137
rect 3712 8103 3746 8137
rect 2824 7963 2858 7997
rect 2912 7963 2946 7997
rect 3824 8103 3858 8137
rect 3918 8103 3952 8137
rect 4018 8103 4052 8137
rect 4118 8103 4152 8137
rect 4218 8103 4252 8137
rect 4318 8103 4352 8137
rect 4418 8103 4452 8137
rect 4718 8103 4752 8137
rect 4818 8103 4852 8137
rect 4918 8103 4952 8137
rect 5218 8103 5252 8137
rect 5318 8103 5352 8137
rect 5418 8103 5452 8137
rect 5518 8103 5552 8137
rect 5718 8103 5752 8137
rect 5818 8103 5852 8137
rect 5918 8103 5952 8137
rect 6018 8103 6052 8137
rect 6118 8103 6152 8137
rect 6218 8103 6252 8137
rect 6524 8118 6558 8152
rect 6618 8103 6652 8137
rect 6712 8088 6746 8122
rect 6828 8103 6862 8137
rect 6928 8103 6962 8137
rect 7028 8103 7062 8137
rect 7128 8103 7162 8137
rect 7228 8103 7262 8137
rect 7328 8103 7362 8137
rect 7428 8103 7462 8137
rect 3024 7963 3058 7997
rect 3118 7963 3152 7997
rect 3318 7963 3352 7997
rect 3418 7963 3452 7997
rect 3618 7963 3652 7997
rect 3718 7963 3752 7997
rect 3918 7963 3952 7997
rect 4018 7963 4052 7997
rect 4118 7963 4152 7997
rect 4318 7963 4352 7997
rect 4418 7963 4452 7997
rect 4518 7963 4552 7997
rect 4718 7963 4752 7997
rect 4818 7963 4852 7997
rect 4912 7963 4946 7997
rect 2624 7823 2658 7857
rect 2718 7823 2752 7857
rect 2918 7823 2952 7857
rect 3018 7823 3052 7857
rect 3218 7823 3252 7857
rect 3312 7823 3346 7857
rect 1824 7683 1858 7717
rect 1918 7683 1952 7717
rect 2018 7683 2052 7717
rect 2118 7683 2152 7717
rect 2518 7683 2552 7717
rect 2618 7683 2652 7717
rect 2712 7683 2746 7717
rect 1424 7543 1458 7577
rect 1518 7543 1552 7577
rect 1618 7543 1652 7577
rect 1718 7543 1752 7577
rect 1918 7543 1952 7577
rect 2018 7543 2052 7577
rect 2318 7543 2352 7577
rect 2418 7543 2452 7577
rect 2618 7543 2652 7577
rect 2712 7543 2746 7577
rect 218 7313 252 7347
rect 318 7313 352 7347
rect 418 7313 452 7347
rect 518 7313 552 7347
rect 818 7313 852 7347
rect 918 7313 952 7347
rect 1018 7313 1052 7347
rect 1118 7313 1152 7347
rect 1212 7313 1246 7347
rect 118 7173 152 7207
rect 218 7173 252 7207
rect 312 7173 346 7207
rect 24 7033 58 7067
rect 118 7033 152 7067
rect 218 7033 252 7067
rect 312 7033 346 7067
rect 1324 7313 1358 7347
rect 1418 7313 1452 7347
rect 1512 7313 1546 7347
rect 1624 7313 1658 7347
rect 1718 7313 1752 7347
rect 2018 7313 2052 7347
rect 2112 7313 2146 7347
rect 2224 7313 2258 7347
rect 2312 7313 2346 7347
rect 2424 7313 2458 7347
rect 2512 7313 2546 7347
rect 424 7173 458 7207
rect 518 7173 552 7207
rect 618 7173 652 7207
rect 718 7173 752 7207
rect 818 7173 852 7207
rect 918 7173 952 7207
rect 1018 7173 1052 7207
rect 1318 7173 1352 7207
rect 1418 7173 1452 7207
rect 1518 7173 1552 7207
rect 1918 7173 1952 7207
rect 2018 7173 2052 7207
rect 2118 7173 2152 7207
rect 2218 7173 2252 7207
rect 2318 7173 2352 7207
rect 2418 7173 2452 7207
rect 2512 7173 2546 7207
rect 424 7033 458 7067
rect 518 7033 552 7067
rect 618 7033 652 7067
rect 718 7033 752 7067
rect 818 7033 852 7067
rect 918 7033 952 7067
rect 1018 7033 1052 7067
rect 1118 7033 1152 7067
rect 1212 7033 1246 7067
rect 1324 7033 1358 7067
rect 1418 7033 1452 7067
rect 1518 7033 1552 7067
rect 1618 7033 1652 7067
rect 1718 7033 1752 7067
rect 2018 7033 2052 7067
rect 2118 7033 2152 7067
rect 2212 7033 2246 7067
rect 24 6893 58 6927
rect 118 6893 152 6927
rect 218 6893 252 6927
rect 618 6893 652 6927
rect 718 6893 752 6927
rect 1118 6893 1152 6927
rect 1218 6893 1252 6927
rect 1318 6893 1352 6927
rect 1412 6893 1446 6927
rect 218 6753 252 6787
rect 318 6753 352 6787
rect 518 6753 552 6787
rect 618 6753 652 6787
rect 718 6753 752 6787
rect 818 6753 852 6787
rect 918 6753 952 6787
rect 1018 6753 1052 6787
rect 1118 6753 1152 6787
rect 1218 6753 1252 6787
rect 1312 6753 1346 6787
rect 24 6613 58 6647
rect 118 6613 152 6647
rect 212 6613 246 6647
rect 324 6613 358 6647
rect 418 6613 452 6647
rect 518 6613 552 6647
rect 818 6613 852 6647
rect 918 6613 952 6647
rect 1012 6613 1046 6647
rect 118 6473 152 6507
rect 218 6473 252 6507
rect 318 6473 352 6507
rect 418 6473 452 6507
rect 512 6473 546 6507
rect 24 6333 58 6367
rect 112 6333 146 6367
rect 1124 6613 1158 6647
rect 1212 6613 1246 6647
rect 1524 6893 1558 6927
rect 1618 6893 1652 6927
rect 1718 6893 1752 6927
rect 1818 6893 1852 6927
rect 1918 6893 1952 6927
rect 2012 6893 2046 6927
rect 1424 6753 1458 6787
rect 1512 6753 1546 6787
rect 3424 7823 3458 7857
rect 3518 7823 3552 7857
rect 3618 7823 3652 7857
rect 3712 7823 3746 7857
rect 3824 7823 3858 7857
rect 3912 7823 3946 7857
rect 4024 7823 4058 7857
rect 4112 7823 4146 7857
rect 2824 7683 2858 7717
rect 2918 7683 2952 7717
rect 3018 7683 3052 7717
rect 3118 7683 3152 7717
rect 3218 7683 3252 7717
rect 3518 7683 3552 7717
rect 3618 7683 3652 7717
rect 3718 7683 3752 7717
rect 3818 7683 3852 7717
rect 4018 7683 4052 7717
rect 4112 7683 4146 7717
rect 2824 7543 2858 7577
rect 2918 7543 2952 7577
rect 3012 7543 3046 7577
rect 3124 7543 3158 7577
rect 3212 7543 3246 7577
rect 3324 7543 3358 7577
rect 3418 7543 3452 7577
rect 3818 7543 3852 7577
rect 3912 7543 3946 7577
rect 4224 7823 4258 7857
rect 4318 7823 4352 7857
rect 4418 7823 4452 7857
rect 4512 7823 4546 7857
rect 4224 7683 4258 7717
rect 4312 7683 4346 7717
rect 4624 7823 4658 7857
rect 4712 7823 4746 7857
rect 4824 7823 4858 7857
rect 4912 7823 4946 7857
rect 5024 7963 5058 7997
rect 5118 7963 5152 7997
rect 5518 7963 5552 7997
rect 5618 7963 5652 7997
rect 5718 7963 5752 7997
rect 5918 7963 5952 7997
rect 6018 7963 6052 7997
rect 6524 7978 6558 8012
rect 6618 7963 6652 7997
rect 6712 7948 6746 7982
rect 6828 7963 6862 7997
rect 6928 7963 6962 7997
rect 7028 7963 7062 7997
rect 7128 7963 7162 7997
rect 7228 7963 7262 7997
rect 7328 7963 7362 7997
rect 7428 7963 7462 7997
rect 5024 7823 5058 7857
rect 5118 7823 5152 7857
rect 5218 7823 5252 7857
rect 5318 7823 5352 7857
rect 5418 7823 5452 7857
rect 5512 7823 5546 7857
rect 4424 7683 4458 7717
rect 4518 7683 4552 7717
rect 4818 7683 4852 7717
rect 4918 7683 4952 7717
rect 5018 7683 5052 7717
rect 5118 7683 5152 7717
rect 5418 7683 5452 7717
rect 5512 7683 5546 7717
rect 4024 7543 4058 7577
rect 4118 7543 4152 7577
rect 4218 7543 4252 7577
rect 4618 7543 4652 7577
rect 4718 7543 4752 7577
rect 4818 7543 4852 7577
rect 4912 7543 4946 7577
rect 5024 7543 5058 7577
rect 5112 7543 5146 7577
rect 5624 7823 5658 7857
rect 5712 7823 5746 7857
rect 5624 7683 5658 7717
rect 5712 7683 5746 7717
rect 5824 7823 5858 7857
rect 5918 7823 5952 7857
rect 6018 7823 6052 7857
rect 6218 7823 6252 7857
rect 6318 7823 6352 7857
rect 6412 7823 6446 7857
rect 6524 7838 6558 7872
rect 6618 7823 6652 7857
rect 6712 7808 6746 7842
rect 6828 7823 6862 7857
rect 6928 7823 6962 7857
rect 7028 7823 7062 7857
rect 7128 7823 7162 7857
rect 7228 7823 7262 7857
rect 7328 7823 7362 7857
rect 7428 7823 7462 7857
rect 5824 7683 5858 7717
rect 5918 7683 5952 7717
rect 6118 7683 6152 7717
rect 6218 7683 6252 7717
rect 6318 7683 6352 7717
rect 6524 7698 6558 7732
rect 6618 7683 6652 7717
rect 6712 7668 6746 7702
rect 6828 7683 6862 7717
rect 6928 7683 6962 7717
rect 7028 7683 7062 7717
rect 7128 7683 7162 7717
rect 7228 7683 7262 7717
rect 7328 7683 7362 7717
rect 7428 7683 7462 7717
rect 5224 7543 5258 7577
rect 5318 7543 5352 7577
rect 5418 7543 5452 7577
rect 5518 7543 5552 7577
rect 5618 7543 5652 7577
rect 5718 7543 5752 7577
rect 5818 7543 5852 7577
rect 5918 7543 5952 7577
rect 6018 7543 6052 7577
rect 6118 7543 6152 7577
rect 6318 7543 6352 7577
rect 6412 7543 6446 7577
rect 6524 7558 6558 7592
rect 6618 7543 6652 7577
rect 6712 7528 6746 7562
rect 6828 7543 6862 7577
rect 6928 7543 6962 7577
rect 7028 7543 7062 7577
rect 7128 7543 7162 7577
rect 7228 7543 7262 7577
rect 7328 7543 7362 7577
rect 7428 7543 7462 7577
rect 2624 7313 2658 7347
rect 2718 7313 2752 7347
rect 2818 7313 2852 7347
rect 2918 7313 2952 7347
rect 3018 7313 3052 7347
rect 3218 7313 3252 7347
rect 3318 7313 3352 7347
rect 3418 7313 3452 7347
rect 3618 7313 3652 7347
rect 3718 7313 3752 7347
rect 3818 7313 3852 7347
rect 4018 7313 4052 7347
rect 4118 7313 4152 7347
rect 4518 7313 4552 7347
rect 4618 7313 4652 7347
rect 4718 7313 4752 7347
rect 4818 7313 4852 7347
rect 4918 7313 4952 7347
rect 5018 7313 5052 7347
rect 5218 7313 5252 7347
rect 5318 7313 5352 7347
rect 5618 7313 5652 7347
rect 5718 7313 5752 7347
rect 6524 7328 6558 7362
rect 6618 7313 6652 7347
rect 6712 7298 6746 7332
rect 6828 7313 6862 7347
rect 6928 7313 6962 7347
rect 7028 7313 7062 7347
rect 7128 7313 7162 7347
rect 7228 7313 7262 7347
rect 7328 7313 7362 7347
rect 7428 7313 7462 7347
rect 2624 7173 2658 7207
rect 2718 7173 2752 7207
rect 2818 7173 2852 7207
rect 2912 7173 2946 7207
rect 3024 7173 3058 7207
rect 3118 7173 3152 7207
rect 3212 7173 3246 7207
rect 2324 7033 2358 7067
rect 2418 7033 2452 7067
rect 2518 7033 2552 7067
rect 2618 7033 2652 7067
rect 2718 7033 2752 7067
rect 2818 7033 2852 7067
rect 2918 7033 2952 7067
rect 3012 7033 3046 7067
rect 2124 6893 2158 6927
rect 2218 6893 2252 6927
rect 2318 6893 2352 6927
rect 2718 6893 2752 6927
rect 2818 6893 2852 6927
rect 2912 6893 2946 6927
rect 1624 6753 1658 6787
rect 1718 6753 1752 6787
rect 1918 6753 1952 6787
rect 2018 6753 2052 6787
rect 2112 6753 2146 6787
rect 3324 7173 3358 7207
rect 3418 7173 3452 7207
rect 3818 7173 3852 7207
rect 3918 7173 3952 7207
rect 4018 7173 4052 7207
rect 4218 7173 4252 7207
rect 4312 7173 4346 7207
rect 3124 7033 3158 7067
rect 3218 7033 3252 7067
rect 3318 7033 3352 7067
rect 3412 7033 3446 7067
rect 3024 6893 3058 6927
rect 3112 6893 3146 6927
rect 3224 6893 3258 6927
rect 3318 6893 3352 6927
rect 3412 6893 3446 6927
rect 3524 7033 3558 7067
rect 3618 7033 3652 7067
rect 3718 7033 3752 7067
rect 3818 7033 3852 7067
rect 3918 7033 3952 7067
rect 4012 7033 4046 7067
rect 4424 7173 4458 7207
rect 4518 7173 4552 7207
rect 4612 7173 4646 7207
rect 4724 7173 4758 7207
rect 4818 7173 4852 7207
rect 4918 7173 4952 7207
rect 5012 7173 5046 7207
rect 5124 7173 5158 7207
rect 5218 7173 5252 7207
rect 5618 7173 5652 7207
rect 5718 7173 5752 7207
rect 5918 7173 5952 7207
rect 6012 7173 6046 7207
rect 4124 7033 4158 7067
rect 4218 7033 4252 7067
rect 4318 7033 4352 7067
rect 4618 7033 4652 7067
rect 4718 7033 4752 7067
rect 5018 7033 5052 7067
rect 5112 7033 5146 7067
rect 3524 6893 3558 6927
rect 3618 6893 3652 6927
rect 3918 6893 3952 6927
rect 4018 6893 4052 6927
rect 4118 6893 4152 6927
rect 4212 6893 4246 6927
rect 4324 6893 4358 6927
rect 4418 6893 4452 6927
rect 4518 6893 4552 6927
rect 4618 6893 4652 6927
rect 4718 6893 4752 6927
rect 4812 6893 4846 6927
rect 4924 6893 4958 6927
rect 5018 6893 5052 6927
rect 5112 6893 5146 6927
rect 6124 7173 6158 7207
rect 6218 7173 6252 7207
rect 6318 7173 6352 7207
rect 6412 7173 6446 7207
rect 6524 7188 6558 7222
rect 6618 7173 6652 7207
rect 6712 7158 6746 7192
rect 6828 7173 6862 7207
rect 6928 7173 6962 7207
rect 7028 7173 7062 7207
rect 7128 7173 7162 7207
rect 7228 7173 7262 7207
rect 7328 7173 7362 7207
rect 7428 7173 7462 7207
rect 5224 7033 5258 7067
rect 5318 7033 5352 7067
rect 5418 7033 5452 7067
rect 5518 7033 5552 7067
rect 5618 7033 5652 7067
rect 5718 7033 5752 7067
rect 5818 7033 5852 7067
rect 6018 7033 6052 7067
rect 6112 7033 6146 7067
rect 5224 6893 5258 6927
rect 5312 6893 5346 6927
rect 5424 6893 5458 6927
rect 5518 6893 5552 6927
rect 5718 6893 5752 6927
rect 5818 6893 5852 6927
rect 6018 6893 6052 6927
rect 6112 6893 6146 6927
rect 2224 6753 2258 6787
rect 2318 6753 2352 6787
rect 2818 6753 2852 6787
rect 2918 6753 2952 6787
rect 4018 6753 4052 6787
rect 4118 6753 4152 6787
rect 4318 6753 4352 6787
rect 4418 6753 4452 6787
rect 4518 6753 4552 6787
rect 4718 6753 4752 6787
rect 4818 6753 4852 6787
rect 4918 6753 4952 6787
rect 5018 6753 5052 6787
rect 5118 6753 5152 6787
rect 5318 6753 5352 6787
rect 5412 6753 5446 6787
rect 1324 6613 1358 6647
rect 1418 6613 1452 6647
rect 1818 6613 1852 6647
rect 1918 6613 1952 6647
rect 2018 6613 2052 6647
rect 2118 6613 2152 6647
rect 2218 6613 2252 6647
rect 2318 6613 2352 6647
rect 2518 6613 2552 6647
rect 2618 6613 2652 6647
rect 3018 6613 3052 6647
rect 3118 6613 3152 6647
rect 3318 6613 3352 6647
rect 3412 6613 3446 6647
rect 624 6473 658 6507
rect 718 6473 752 6507
rect 818 6473 852 6507
rect 918 6473 952 6507
rect 1018 6473 1052 6507
rect 1118 6473 1152 6507
rect 1218 6473 1252 6507
rect 1418 6473 1452 6507
rect 1518 6473 1552 6507
rect 1612 6473 1646 6507
rect 224 6333 258 6367
rect 318 6333 352 6367
rect 418 6333 452 6367
rect 518 6333 552 6367
rect 718 6333 752 6367
rect 812 6333 846 6367
rect 924 6333 958 6367
rect 1012 6333 1046 6367
rect 1124 6333 1158 6367
rect 1218 6333 1252 6367
rect 1318 6333 1352 6367
rect 1518 6333 1552 6367
rect 1612 6333 1646 6367
rect 3524 6613 3558 6647
rect 3612 6613 3646 6647
rect 3724 6613 3758 6647
rect 3818 6613 3852 6647
rect 3918 6613 3952 6647
rect 4218 6613 4252 6647
rect 4318 6613 4352 6647
rect 4412 6613 4446 6647
rect 1724 6473 1758 6507
rect 1818 6473 1852 6507
rect 2118 6473 2152 6507
rect 2218 6473 2252 6507
rect 3218 6473 3252 6507
rect 3318 6473 3352 6507
rect 3418 6473 3452 6507
rect 3618 6473 3652 6507
rect 3712 6473 3746 6507
rect 1724 6333 1758 6367
rect 1818 6333 1852 6367
rect 1912 6333 1946 6367
rect 2024 6333 2058 6367
rect 2118 6333 2152 6367
rect 2218 6333 2252 6367
rect 2318 6333 2352 6367
rect 2618 6333 2652 6367
rect 2718 6333 2752 6367
rect 2812 6333 2846 6367
rect 318 6103 352 6137
rect 418 6103 452 6137
rect 818 6103 852 6137
rect 918 6103 952 6137
rect 1018 6103 1052 6137
rect 1218 6103 1252 6137
rect 1318 6103 1352 6137
rect 1518 6103 1552 6137
rect 1618 6103 1652 6137
rect 1918 6103 1952 6137
rect 2018 6103 2052 6137
rect 2218 6103 2252 6137
rect 2318 6103 2352 6137
rect 2412 6103 2446 6137
rect 218 5963 252 5997
rect 318 5963 352 5997
rect 412 5963 446 5997
rect 524 5963 558 5997
rect 618 5963 652 5997
rect 818 5963 852 5997
rect 918 5963 952 5997
rect 1018 5963 1052 5997
rect 1218 5963 1252 5997
rect 1312 5963 1346 5997
rect 2924 6333 2958 6367
rect 3018 6333 3052 6367
rect 3218 6333 3252 6367
rect 3312 6333 3346 6367
rect 5524 6753 5558 6787
rect 5612 6753 5646 6787
rect 5724 6753 5758 6787
rect 5812 6753 5846 6787
rect 4524 6613 4558 6647
rect 4618 6613 4652 6647
rect 4718 6613 4752 6647
rect 4818 6613 4852 6647
rect 4918 6613 4952 6647
rect 5418 6613 5452 6647
rect 5518 6613 5552 6647
rect 5718 6613 5752 6647
rect 5812 6613 5846 6647
rect 3824 6473 3858 6507
rect 3918 6473 3952 6507
rect 4018 6473 4052 6507
rect 4118 6473 4152 6507
rect 4218 6473 4252 6507
rect 4618 6473 4652 6507
rect 4718 6473 4752 6507
rect 4818 6473 4852 6507
rect 4918 6473 4952 6507
rect 5018 6473 5052 6507
rect 5112 6473 5146 6507
rect 3424 6333 3458 6367
rect 3518 6333 3552 6367
rect 3618 6333 3652 6367
rect 3918 6333 3952 6367
rect 4018 6333 4052 6367
rect 4118 6333 4152 6367
rect 4518 6333 4552 6367
rect 4618 6333 4652 6367
rect 4818 6333 4852 6367
rect 4918 6333 4952 6367
rect 5012 6333 5046 6367
rect 2524 6103 2558 6137
rect 2618 6103 2652 6137
rect 2718 6103 2752 6137
rect 2918 6103 2952 6137
rect 3018 6103 3052 6137
rect 3218 6103 3252 6137
rect 3318 6103 3352 6137
rect 3418 6103 3452 6137
rect 3618 6103 3652 6137
rect 3712 6103 3746 6137
rect 1424 5963 1458 5997
rect 1518 5963 1552 5997
rect 1618 5963 1652 5997
rect 1718 5963 1752 5997
rect 1818 5963 1852 5997
rect 1918 5963 1952 5997
rect 2618 5963 2652 5997
rect 2718 5963 2752 5997
rect 2818 5963 2852 5997
rect 2918 5963 2952 5997
rect 3218 5963 3252 5997
rect 3312 5963 3346 5997
rect 24 5823 58 5857
rect 118 5823 152 5857
rect 218 5823 252 5857
rect 518 5823 552 5857
rect 618 5823 652 5857
rect 918 5823 952 5857
rect 1018 5823 1052 5857
rect 1118 5823 1152 5857
rect 1318 5823 1352 5857
rect 1418 5823 1452 5857
rect 1518 5823 1552 5857
rect 1618 5823 1652 5857
rect 1718 5823 1752 5857
rect 1918 5823 1952 5857
rect 2012 5823 2046 5857
rect 218 5683 252 5717
rect 312 5683 346 5717
rect 424 5683 458 5717
rect 518 5683 552 5717
rect 618 5683 652 5717
rect 718 5683 752 5717
rect 818 5683 852 5717
rect 918 5683 952 5717
rect 1012 5683 1046 5717
rect 3824 6103 3858 6137
rect 3918 6103 3952 6137
rect 4012 6103 4046 6137
rect 4124 6103 4158 6137
rect 4218 6103 4252 6137
rect 4318 6103 4352 6137
rect 4412 6103 4446 6137
rect 4524 6103 4558 6137
rect 4612 6103 4646 6137
rect 5224 6473 5258 6507
rect 5312 6473 5346 6507
rect 5124 6333 5158 6367
rect 5218 6333 5252 6367
rect 5312 6333 5346 6367
rect 6224 7033 6258 7067
rect 6318 7033 6352 7067
rect 6524 7048 6558 7082
rect 6618 7033 6652 7067
rect 6712 7018 6746 7052
rect 6828 7033 6862 7067
rect 6928 7033 6962 7067
rect 7028 7033 7062 7067
rect 7128 7033 7162 7067
rect 7228 7033 7262 7067
rect 7328 7033 7362 7067
rect 7428 7033 7462 7067
rect 6224 6893 6258 6927
rect 6318 6893 6352 6927
rect 6524 6908 6558 6942
rect 6618 6893 6652 6927
rect 6712 6878 6746 6912
rect 6828 6893 6862 6927
rect 6928 6893 6962 6927
rect 7028 6893 7062 6927
rect 7128 6893 7162 6927
rect 7228 6893 7262 6927
rect 7328 6893 7362 6927
rect 7428 6893 7462 6927
rect 5924 6753 5958 6787
rect 6018 6753 6052 6787
rect 6118 6753 6152 6787
rect 6218 6753 6252 6787
rect 6318 6753 6352 6787
rect 6524 6768 6558 6802
rect 6618 6753 6652 6787
rect 6712 6738 6746 6772
rect 6828 6753 6862 6787
rect 6928 6753 6962 6787
rect 7028 6753 7062 6787
rect 7128 6753 7162 6787
rect 7228 6753 7262 6787
rect 7328 6753 7362 6787
rect 7428 6753 7462 6787
rect 5924 6613 5958 6647
rect 6018 6613 6052 6647
rect 6118 6613 6152 6647
rect 6524 6628 6558 6662
rect 6618 6613 6652 6647
rect 6712 6598 6746 6632
rect 6828 6613 6862 6647
rect 6928 6613 6962 6647
rect 7028 6613 7062 6647
rect 7128 6613 7162 6647
rect 7228 6613 7262 6647
rect 7328 6613 7362 6647
rect 7428 6613 7462 6647
rect 5424 6473 5458 6507
rect 5518 6473 5552 6507
rect 5618 6473 5652 6507
rect 5718 6473 5752 6507
rect 5818 6473 5852 6507
rect 5918 6473 5952 6507
rect 6018 6473 6052 6507
rect 6218 6473 6252 6507
rect 6318 6473 6352 6507
rect 6524 6488 6558 6522
rect 6618 6473 6652 6507
rect 6712 6458 6746 6492
rect 6828 6473 6862 6507
rect 6928 6473 6962 6507
rect 7028 6473 7062 6507
rect 7128 6473 7162 6507
rect 7228 6473 7262 6507
rect 7328 6473 7362 6507
rect 7428 6473 7462 6507
rect 5424 6333 5458 6367
rect 5518 6333 5552 6367
rect 5818 6333 5852 6367
rect 5918 6333 5952 6367
rect 6018 6333 6052 6367
rect 6112 6333 6146 6367
rect 6224 6333 6258 6367
rect 6318 6333 6352 6367
rect 6412 6333 6446 6367
rect 6524 6348 6558 6382
rect 6618 6333 6652 6367
rect 6712 6318 6746 6352
rect 6828 6333 6862 6367
rect 6928 6333 6962 6367
rect 7028 6333 7062 6367
rect 7128 6333 7162 6367
rect 7228 6333 7262 6367
rect 7328 6333 7362 6367
rect 7428 6333 7462 6367
rect 4724 6103 4758 6137
rect 4818 6103 4852 6137
rect 4918 6103 4952 6137
rect 5418 6103 5452 6137
rect 5518 6103 5552 6137
rect 5718 6103 5752 6137
rect 5818 6103 5852 6137
rect 5918 6103 5952 6137
rect 6012 6103 6046 6137
rect 3424 5963 3458 5997
rect 3518 5963 3552 5997
rect 3618 5963 3652 5997
rect 3718 5963 3752 5997
rect 3818 5963 3852 5997
rect 3918 5963 3952 5997
rect 4218 5963 4252 5997
rect 4318 5963 4352 5997
rect 4518 5963 4552 5997
rect 4618 5963 4652 5997
rect 4918 5963 4952 5997
rect 5018 5963 5052 5997
rect 5118 5963 5152 5997
rect 5212 5963 5246 5997
rect 2124 5823 2158 5857
rect 2218 5823 2252 5857
rect 2318 5823 2352 5857
rect 2518 5823 2552 5857
rect 2618 5823 2652 5857
rect 2718 5823 2752 5857
rect 2818 5823 2852 5857
rect 2918 5823 2952 5857
rect 3118 5823 3152 5857
rect 3218 5823 3252 5857
rect 3318 5823 3352 5857
rect 3412 5823 3446 5857
rect 1124 5683 1158 5717
rect 1218 5683 1252 5717
rect 1318 5683 1352 5717
rect 1418 5683 1452 5717
rect 1518 5683 1552 5717
rect 1618 5683 1652 5717
rect 1718 5683 1752 5717
rect 1818 5683 1852 5717
rect 1918 5683 1952 5717
rect 2118 5683 2152 5717
rect 2218 5683 2252 5717
rect 2318 5683 2352 5717
rect 2718 5683 2752 5717
rect 2812 5683 2846 5717
rect 118 5543 152 5577
rect 218 5543 252 5577
rect 318 5543 352 5577
rect 418 5543 452 5577
rect 518 5543 552 5577
rect 718 5543 752 5577
rect 818 5543 852 5577
rect 1018 5543 1052 5577
rect 1112 5543 1146 5577
rect 24 5403 58 5437
rect 118 5403 152 5437
rect 218 5403 252 5437
rect 318 5403 352 5437
rect 412 5403 446 5437
rect 1224 5543 1258 5577
rect 1312 5543 1346 5577
rect 1424 5543 1458 5577
rect 1518 5543 1552 5577
rect 1618 5543 1652 5577
rect 1718 5543 1752 5577
rect 1818 5543 1852 5577
rect 1912 5543 1946 5577
rect 524 5403 558 5437
rect 618 5403 652 5437
rect 718 5403 752 5437
rect 1318 5403 1352 5437
rect 1412 5403 1446 5437
rect 1524 5403 1558 5437
rect 1618 5403 1652 5437
rect 1712 5403 1746 5437
rect 2024 5543 2058 5577
rect 2118 5543 2152 5577
rect 2212 5543 2246 5577
rect 1824 5403 1858 5437
rect 1918 5403 1952 5437
rect 2018 5403 2052 5437
rect 2118 5403 2152 5437
rect 2212 5403 2246 5437
rect 318 5263 352 5297
rect 418 5263 452 5297
rect 718 5263 752 5297
rect 818 5263 852 5297
rect 1218 5263 1252 5297
rect 1318 5263 1352 5297
rect 1418 5263 1452 5297
rect 1618 5263 1652 5297
rect 1718 5263 1752 5297
rect 2018 5263 2052 5297
rect 2112 5263 2146 5297
rect 118 5123 152 5157
rect 218 5123 252 5157
rect 318 5123 352 5157
rect 418 5123 452 5157
rect 618 5123 652 5157
rect 718 5123 752 5157
rect 818 5123 852 5157
rect 1218 5123 1252 5157
rect 1312 5123 1346 5157
rect 24 4753 58 4787
rect 118 4753 152 4787
rect 212 4753 246 4787
rect 324 4753 358 4787
rect 418 4753 452 4787
rect 618 4753 652 4787
rect 718 4753 752 4787
rect 1018 4753 1052 4787
rect 1112 4753 1146 4787
rect 1424 5123 1458 5157
rect 1518 5123 1552 5157
rect 1618 5123 1652 5157
rect 1718 5123 1752 5157
rect 2018 5123 2052 5157
rect 2112 5123 2146 5157
rect 2924 5683 2958 5717
rect 3012 5683 3046 5717
rect 3124 5683 3158 5717
rect 3212 5683 3246 5717
rect 3324 5683 3358 5717
rect 3412 5683 3446 5717
rect 3524 5823 3558 5857
rect 3618 5823 3652 5857
rect 3718 5823 3752 5857
rect 4018 5823 4052 5857
rect 4112 5823 4146 5857
rect 3524 5683 3558 5717
rect 3612 5683 3646 5717
rect 3724 5683 3758 5717
rect 3818 5683 3852 5717
rect 4018 5683 4052 5717
rect 4112 5683 4146 5717
rect 2324 5543 2358 5577
rect 2418 5543 2452 5577
rect 2518 5543 2552 5577
rect 3018 5543 3052 5577
rect 3118 5543 3152 5577
rect 3218 5543 3252 5577
rect 3318 5543 3352 5577
rect 3418 5543 3452 5577
rect 3518 5543 3552 5577
rect 3618 5543 3652 5577
rect 3818 5543 3852 5577
rect 3918 5543 3952 5577
rect 4012 5543 4046 5577
rect 2324 5403 2358 5437
rect 2418 5403 2452 5437
rect 2718 5403 2752 5437
rect 2818 5403 2852 5437
rect 3018 5403 3052 5437
rect 3118 5403 3152 5437
rect 3518 5403 3552 5437
rect 3618 5403 3652 5437
rect 3712 5403 3746 5437
rect 2224 5263 2258 5297
rect 2312 5263 2346 5297
rect 2424 5263 2458 5297
rect 2518 5263 2552 5297
rect 2612 5263 2646 5297
rect 2724 5263 2758 5297
rect 2818 5263 2852 5297
rect 2912 5263 2946 5297
rect 3024 5263 3058 5297
rect 3112 5263 3146 5297
rect 5324 5963 5358 5997
rect 5418 5963 5452 5997
rect 5518 5963 5552 5997
rect 5618 5963 5652 5997
rect 5718 5963 5752 5997
rect 5812 5963 5846 5997
rect 4224 5823 4258 5857
rect 4318 5823 4352 5857
rect 4518 5823 4552 5857
rect 4618 5823 4652 5857
rect 4718 5823 4752 5857
rect 4918 5823 4952 5857
rect 5018 5823 5052 5857
rect 5118 5823 5152 5857
rect 5218 5823 5252 5857
rect 5318 5823 5352 5857
rect 5618 5823 5652 5857
rect 5712 5823 5746 5857
rect 4224 5683 4258 5717
rect 4312 5683 4346 5717
rect 4424 5683 4458 5717
rect 4512 5683 4546 5717
rect 4624 5683 4658 5717
rect 4718 5683 4752 5717
rect 4918 5683 4952 5717
rect 5018 5683 5052 5717
rect 5218 5683 5252 5717
rect 5318 5683 5352 5717
rect 5418 5683 5452 5717
rect 5512 5683 5546 5717
rect 6124 6103 6158 6137
rect 6212 6103 6246 6137
rect 6324 6103 6358 6137
rect 6412 6103 6446 6137
rect 6524 6118 6558 6152
rect 6618 6103 6652 6137
rect 6712 6088 6746 6122
rect 6828 6103 6862 6137
rect 6928 6103 6962 6137
rect 7028 6103 7062 6137
rect 7128 6103 7162 6137
rect 7228 6103 7262 6137
rect 7328 6103 7362 6137
rect 7428 6103 7462 6137
rect 5924 5963 5958 5997
rect 6018 5963 6052 5997
rect 6318 5963 6352 5997
rect 6412 5963 6446 5997
rect 6524 5978 6558 6012
rect 6618 5963 6652 5997
rect 6712 5948 6746 5982
rect 6828 5963 6862 5997
rect 6928 5963 6962 5997
rect 7028 5963 7062 5997
rect 7128 5963 7162 5997
rect 7228 5963 7262 5997
rect 7328 5963 7362 5997
rect 7428 5963 7462 5997
rect 5824 5823 5858 5857
rect 5912 5823 5946 5857
rect 6024 5823 6058 5857
rect 6118 5823 6152 5857
rect 6218 5823 6252 5857
rect 6318 5823 6352 5857
rect 6524 5838 6558 5872
rect 6618 5823 6652 5857
rect 6712 5808 6746 5842
rect 6828 5823 6862 5857
rect 6928 5823 6962 5857
rect 7028 5823 7062 5857
rect 7128 5823 7162 5857
rect 7228 5823 7262 5857
rect 7328 5823 7362 5857
rect 7428 5823 7462 5857
rect 5624 5683 5658 5717
rect 5718 5683 5752 5717
rect 5818 5683 5852 5717
rect 6018 5683 6052 5717
rect 6118 5683 6152 5717
rect 6218 5683 6252 5717
rect 6318 5683 6352 5717
rect 6524 5698 6558 5732
rect 6618 5683 6652 5717
rect 6712 5668 6746 5702
rect 6828 5683 6862 5717
rect 6928 5683 6962 5717
rect 7028 5683 7062 5717
rect 7128 5683 7162 5717
rect 7228 5683 7262 5717
rect 7328 5683 7362 5717
rect 7428 5683 7462 5717
rect 4124 5543 4158 5577
rect 4218 5543 4252 5577
rect 4518 5543 4552 5577
rect 4618 5543 4652 5577
rect 4718 5543 4752 5577
rect 4818 5543 4852 5577
rect 5118 5543 5152 5577
rect 5218 5543 5252 5577
rect 5318 5543 5352 5577
rect 5418 5543 5452 5577
rect 5718 5543 5752 5577
rect 5818 5543 5852 5577
rect 5918 5543 5952 5577
rect 6018 5543 6052 5577
rect 6524 5558 6558 5592
rect 6618 5543 6652 5577
rect 6712 5528 6746 5562
rect 6828 5543 6862 5577
rect 6928 5543 6962 5577
rect 7028 5543 7062 5577
rect 7128 5543 7162 5577
rect 7228 5543 7262 5577
rect 7328 5543 7362 5577
rect 7428 5543 7462 5577
rect 3824 5403 3858 5437
rect 3918 5403 3952 5437
rect 4018 5403 4052 5437
rect 4118 5403 4152 5437
rect 4218 5403 4252 5437
rect 4418 5403 4452 5437
rect 4518 5403 4552 5437
rect 4618 5403 4652 5437
rect 4718 5403 4752 5437
rect 5018 5403 5052 5437
rect 5112 5403 5146 5437
rect 5224 5403 5258 5437
rect 5312 5403 5346 5437
rect 3224 5263 3258 5297
rect 3318 5263 3352 5297
rect 3518 5263 3552 5297
rect 3618 5263 3652 5297
rect 4018 5263 4052 5297
rect 4118 5263 4152 5297
rect 4218 5263 4252 5297
rect 4318 5263 4352 5297
rect 4418 5263 4452 5297
rect 4518 5263 4552 5297
rect 4718 5263 4752 5297
rect 4818 5263 4852 5297
rect 4918 5263 4952 5297
rect 5018 5263 5052 5297
rect 5118 5263 5152 5297
rect 5212 5263 5246 5297
rect 2224 5123 2258 5157
rect 2318 5123 2352 5157
rect 2418 5123 2452 5157
rect 2518 5123 2552 5157
rect 2818 5123 2852 5157
rect 2918 5123 2952 5157
rect 3018 5123 3052 5157
rect 3118 5123 3152 5157
rect 3518 5123 3552 5157
rect 3618 5123 3652 5157
rect 4018 5123 4052 5157
rect 4118 5123 4152 5157
rect 4218 5123 4252 5157
rect 4312 5123 4346 5157
rect 1224 4753 1258 4787
rect 1318 4753 1352 4787
rect 1518 4753 1552 4787
rect 1618 4753 1652 4787
rect 2018 4753 2052 4787
rect 2118 4753 2152 4787
rect 2218 4753 2252 4787
rect 2718 4753 2752 4787
rect 2812 4753 2846 4787
rect 24 4613 58 4647
rect 118 4613 152 4647
rect 318 4613 352 4647
rect 418 4613 452 4647
rect 518 4613 552 4647
rect 818 4613 852 4647
rect 918 4613 952 4647
rect 1218 4613 1252 4647
rect 1318 4613 1352 4647
rect 1518 4613 1552 4647
rect 1618 4613 1652 4647
rect 1718 4613 1752 4647
rect 1812 4613 1846 4647
rect 24 4473 58 4507
rect 112 4473 146 4507
rect 224 4473 258 4507
rect 318 4473 352 4507
rect 718 4473 752 4507
rect 818 4473 852 4507
rect 918 4473 952 4507
rect 1318 4473 1352 4507
rect 1418 4473 1452 4507
rect 1518 4473 1552 4507
rect 1612 4473 1646 4507
rect 24 4333 58 4367
rect 118 4333 152 4367
rect 218 4333 252 4367
rect 318 4333 352 4367
rect 412 4333 446 4367
rect 24 4193 58 4227
rect 112 4193 146 4227
rect 224 4193 258 4227
rect 312 4193 346 4227
rect 524 4333 558 4367
rect 618 4333 652 4367
rect 712 4333 746 4367
rect 1924 4613 1958 4647
rect 2012 4613 2046 4647
rect 4424 5123 4458 5157
rect 4518 5123 4552 5157
rect 4618 5123 4652 5157
rect 4712 5123 4746 5157
rect 5424 5403 5458 5437
rect 5512 5403 5546 5437
rect 5324 5263 5358 5297
rect 5412 5263 5446 5297
rect 5624 5403 5658 5437
rect 5712 5403 5746 5437
rect 5824 5403 5858 5437
rect 5918 5403 5952 5437
rect 6018 5403 6052 5437
rect 6524 5418 6558 5452
rect 6618 5403 6652 5437
rect 6712 5388 6746 5422
rect 6828 5403 6862 5437
rect 6928 5403 6962 5437
rect 7028 5403 7062 5437
rect 7128 5403 7162 5437
rect 7228 5403 7262 5437
rect 7328 5403 7362 5437
rect 7428 5403 7462 5437
rect 5524 5263 5558 5297
rect 5618 5263 5652 5297
rect 5818 5263 5852 5297
rect 5918 5263 5952 5297
rect 6218 5263 6252 5297
rect 6318 5263 6352 5297
rect 6412 5263 6446 5297
rect 6524 5278 6558 5312
rect 6618 5263 6652 5297
rect 6712 5248 6746 5282
rect 6828 5263 6862 5297
rect 6928 5263 6962 5297
rect 7028 5263 7062 5297
rect 7128 5263 7162 5297
rect 7228 5263 7262 5297
rect 7328 5263 7362 5297
rect 7428 5263 7462 5297
rect 4824 5123 4858 5157
rect 4918 5123 4952 5157
rect 5018 5123 5052 5157
rect 5118 5123 5152 5157
rect 5218 5123 5252 5157
rect 5518 5123 5552 5157
rect 5618 5123 5652 5157
rect 5712 5123 5746 5157
rect 2924 4753 2958 4787
rect 3018 4753 3052 4787
rect 3418 4753 3452 4787
rect 3518 4753 3552 4787
rect 3618 4753 3652 4787
rect 4218 4753 4252 4787
rect 4318 4753 4352 4787
rect 4518 4753 4552 4787
rect 4612 4753 4646 4787
rect 2124 4613 2158 4647
rect 2218 4613 2252 4647
rect 2518 4613 2552 4647
rect 2618 4613 2652 4647
rect 2818 4613 2852 4647
rect 2918 4613 2952 4647
rect 3018 4613 3052 4647
rect 3118 4613 3152 4647
rect 3212 4613 3246 4647
rect 1724 4473 1758 4507
rect 1818 4473 1852 4507
rect 2018 4473 2052 4507
rect 2118 4473 2152 4507
rect 2318 4473 2352 4507
rect 2412 4473 2446 4507
rect 824 4333 858 4367
rect 918 4333 952 4367
rect 1018 4333 1052 4367
rect 1618 4333 1652 4367
rect 1718 4333 1752 4367
rect 2018 4333 2052 4367
rect 2118 4333 2152 4367
rect 2318 4333 2352 4367
rect 2412 4333 2446 4367
rect 424 4193 458 4227
rect 518 4193 552 4227
rect 918 4193 952 4227
rect 1018 4193 1052 4227
rect 1118 4193 1152 4227
rect 1218 4193 1252 4227
rect 1318 4193 1352 4227
rect 1412 4193 1446 4227
rect 24 4053 58 4087
rect 118 4053 152 4087
rect 318 4053 352 4087
rect 412 4053 446 4087
rect 524 4053 558 4087
rect 612 4053 646 4087
rect 218 3913 252 3947
rect 318 3913 352 3947
rect 418 3913 452 3947
rect 512 3913 546 3947
rect 3324 4613 3358 4647
rect 3418 4613 3452 4647
rect 3518 4613 3552 4647
rect 3718 4613 3752 4647
rect 3818 4613 3852 4647
rect 3918 4613 3952 4647
rect 4118 4613 4152 4647
rect 4218 4613 4252 4647
rect 4318 4613 4352 4647
rect 4418 4613 4452 4647
rect 4512 4613 4546 4647
rect 2524 4473 2558 4507
rect 2618 4473 2652 4507
rect 2818 4473 2852 4507
rect 2918 4473 2952 4507
rect 3018 4473 3052 4507
rect 3218 4473 3252 4507
rect 3312 4473 3346 4507
rect 2524 4333 2558 4367
rect 2618 4333 2652 4367
rect 2718 4333 2752 4367
rect 2812 4333 2846 4367
rect 2924 4333 2958 4367
rect 3018 4333 3052 4367
rect 3118 4333 3152 4367
rect 3212 4333 3246 4367
rect 3424 4473 3458 4507
rect 3518 4473 3552 4507
rect 3718 4473 3752 4507
rect 3818 4473 3852 4507
rect 4118 4473 4152 4507
rect 4218 4473 4252 4507
rect 4312 4473 4346 4507
rect 4724 4753 4758 4787
rect 4818 4753 4852 4787
rect 5118 4753 5152 4787
rect 5218 4753 5252 4787
rect 5318 4753 5352 4787
rect 5412 4753 5446 4787
rect 5824 5123 5858 5157
rect 5918 5123 5952 5157
rect 6524 5138 6558 5172
rect 6618 5123 6652 5157
rect 6712 5108 6746 5142
rect 6828 5123 6862 5157
rect 6928 5123 6962 5157
rect 7028 5123 7062 5157
rect 7128 5123 7162 5157
rect 7228 5123 7262 5157
rect 7328 5123 7362 5157
rect 7428 5123 7462 5157
rect 5524 4753 5558 4787
rect 5618 4753 5652 4787
rect 5818 4753 5852 4787
rect 5912 4753 5946 4787
rect 6024 4753 6058 4787
rect 6112 4753 6146 4787
rect 4624 4613 4658 4647
rect 4718 4613 4752 4647
rect 5018 4613 5052 4647
rect 5118 4613 5152 4647
rect 5218 4613 5252 4647
rect 5318 4613 5352 4647
rect 5418 4613 5452 4647
rect 5718 4613 5752 4647
rect 5818 4613 5852 4647
rect 5918 4613 5952 4647
rect 6012 4613 6046 4647
rect 4424 4473 4458 4507
rect 4518 4473 4552 4507
rect 4618 4473 4652 4507
rect 5018 4473 5052 4507
rect 5118 4473 5152 4507
rect 5212 4473 5246 4507
rect 3324 4333 3358 4367
rect 3418 4333 3452 4367
rect 3518 4333 3552 4367
rect 3618 4333 3652 4367
rect 4018 4333 4052 4367
rect 4118 4333 4152 4367
rect 4218 4333 4252 4367
rect 4818 4333 4852 4367
rect 4918 4333 4952 4367
rect 5012 4333 5046 4367
rect 1524 4193 1558 4227
rect 1618 4193 1652 4227
rect 1918 4193 1952 4227
rect 2018 4193 2052 4227
rect 2118 4193 2152 4227
rect 2218 4193 2252 4227
rect 2518 4193 2552 4227
rect 2618 4193 2652 4227
rect 2818 4193 2852 4227
rect 2918 4193 2952 4227
rect 3018 4193 3052 4227
rect 3218 4193 3252 4227
rect 3318 4193 3352 4227
rect 3412 4193 3446 4227
rect 724 4053 758 4087
rect 818 4053 852 4087
rect 918 4053 952 4087
rect 1318 4053 1352 4087
rect 1418 4053 1452 4087
rect 1512 4053 1546 4087
rect 1624 4053 1658 4087
rect 1712 4053 1746 4087
rect 1824 4053 1858 4087
rect 1912 4053 1946 4087
rect 2024 4053 2058 4087
rect 2118 4053 2152 4087
rect 2212 4053 2246 4087
rect 624 3913 658 3947
rect 718 3913 752 3947
rect 1118 3913 1152 3947
rect 1218 3913 1252 3947
rect 1518 3913 1552 3947
rect 1618 3913 1652 3947
rect 1918 3913 1952 3947
rect 2018 3913 2052 3947
rect 2112 3913 2146 3947
rect 118 3773 152 3807
rect 218 3773 252 3807
rect 318 3773 352 3807
rect 418 3773 452 3807
rect 518 3773 552 3807
rect 818 3773 852 3807
rect 918 3773 952 3807
rect 1018 3773 1052 3807
rect 1118 3773 1152 3807
rect 1212 3773 1246 3807
rect 118 3543 152 3577
rect 212 3543 246 3577
rect 1324 3773 1358 3807
rect 1412 3773 1446 3807
rect 324 3543 358 3577
rect 418 3543 452 3577
rect 518 3543 552 3577
rect 618 3543 652 3577
rect 718 3543 752 3577
rect 818 3543 852 3577
rect 1018 3543 1052 3577
rect 1118 3543 1152 3577
rect 1218 3543 1252 3577
rect 1312 3543 1346 3577
rect 318 3403 352 3437
rect 418 3403 452 3437
rect 512 3403 546 3437
rect 624 3403 658 3437
rect 712 3403 746 3437
rect 1524 3773 1558 3807
rect 1618 3773 1652 3807
rect 1712 3773 1746 3807
rect 1424 3543 1458 3577
rect 1512 3543 1546 3577
rect 2324 4053 2358 4087
rect 2412 4053 2446 4087
rect 2524 4053 2558 4087
rect 2618 4053 2652 4087
rect 3118 4053 3152 4087
rect 3212 4053 3246 4087
rect 2224 3913 2258 3947
rect 2318 3913 2352 3947
rect 2418 3913 2452 3947
rect 2518 3913 2552 3947
rect 2818 3913 2852 3947
rect 2918 3913 2952 3947
rect 3118 3913 3152 3947
rect 3212 3913 3246 3947
rect 3324 4053 3358 4087
rect 3412 4053 3446 4087
rect 3524 4193 3558 4227
rect 3612 4193 3646 4227
rect 3724 4193 3758 4227
rect 3818 4193 3852 4227
rect 3918 4193 3952 4227
rect 4318 4193 4352 4227
rect 4412 4193 4446 4227
rect 4524 4193 4558 4227
rect 4618 4193 4652 4227
rect 4918 4193 4952 4227
rect 5012 4193 5046 4227
rect 3524 4053 3558 4087
rect 3618 4053 3652 4087
rect 3918 4053 3952 4087
rect 4018 4053 4052 4087
rect 4218 4053 4252 4087
rect 4318 4053 4352 4087
rect 4518 4053 4552 4087
rect 4618 4053 4652 4087
rect 4712 4053 4746 4087
rect 3324 3913 3358 3947
rect 3418 3913 3452 3947
rect 3518 3913 3552 3947
rect 4018 3913 4052 3947
rect 4112 3913 4146 3947
rect 1824 3773 1858 3807
rect 1918 3773 1952 3807
rect 2118 3773 2152 3807
rect 2218 3773 2252 3807
rect 2318 3773 2352 3807
rect 2618 3773 2652 3807
rect 2718 3773 2752 3807
rect 2818 3773 2852 3807
rect 2918 3773 2952 3807
rect 3218 3773 3252 3807
rect 3318 3773 3352 3807
rect 3412 3773 3446 3807
rect 1624 3543 1658 3577
rect 1718 3543 1752 3577
rect 1818 3543 1852 3577
rect 1918 3543 1952 3577
rect 2118 3543 2152 3577
rect 2212 3543 2246 3577
rect 824 3403 858 3437
rect 918 3403 952 3437
rect 1018 3403 1052 3437
rect 1218 3403 1252 3437
rect 1318 3403 1352 3437
rect 1518 3403 1552 3437
rect 1618 3403 1652 3437
rect 1718 3403 1752 3437
rect 1818 3403 1852 3437
rect 1912 3403 1946 3437
rect 24 3263 58 3297
rect 118 3263 152 3297
rect 218 3263 252 3297
rect 318 3263 352 3297
rect 718 3263 752 3297
rect 818 3263 852 3297
rect 918 3263 952 3297
rect 1118 3263 1152 3297
rect 1212 3263 1246 3297
rect 218 3123 252 3157
rect 318 3123 352 3157
rect 412 3123 446 3157
rect 524 3123 558 3157
rect 618 3123 652 3157
rect 718 3123 752 3157
rect 918 3123 952 3157
rect 1018 3123 1052 3157
rect 1112 3123 1146 3157
rect 4224 3913 4258 3947
rect 4318 3913 4352 3947
rect 4418 3913 4452 3947
rect 4512 3913 4546 3947
rect 5324 4473 5358 4507
rect 5418 4473 5452 4507
rect 5518 4473 5552 4507
rect 5618 4473 5652 4507
rect 5712 4473 5746 4507
rect 5124 4333 5158 4367
rect 5218 4333 5252 4367
rect 5318 4333 5352 4367
rect 5412 4333 5446 4367
rect 5124 4193 5158 4227
rect 5218 4193 5252 4227
rect 5318 4193 5352 4227
rect 5412 4193 5446 4227
rect 6224 4753 6258 4787
rect 6318 4753 6352 4787
rect 6524 4768 6558 4802
rect 6618 4753 6652 4787
rect 6712 4738 6746 4772
rect 6828 4753 6862 4787
rect 6928 4753 6962 4787
rect 7028 4753 7062 4787
rect 7128 4753 7162 4787
rect 7228 4753 7262 4787
rect 7328 4753 7362 4787
rect 7428 4753 7462 4787
rect 6124 4613 6158 4647
rect 6212 4613 6246 4647
rect 5824 4473 5858 4507
rect 5918 4473 5952 4507
rect 6118 4473 6152 4507
rect 6212 4473 6246 4507
rect 5524 4333 5558 4367
rect 5618 4333 5652 4367
rect 5918 4333 5952 4367
rect 6012 4333 6046 4367
rect 5524 4193 5558 4227
rect 5618 4193 5652 4227
rect 5718 4193 5752 4227
rect 5812 4193 5846 4227
rect 4824 4053 4858 4087
rect 4918 4053 4952 4087
rect 5018 4053 5052 4087
rect 5218 4053 5252 4087
rect 5318 4053 5352 4087
rect 5518 4053 5552 4087
rect 5612 4053 5646 4087
rect 6124 4333 6158 4367
rect 6212 4333 6246 4367
rect 6324 4613 6358 4647
rect 6412 4613 6446 4647
rect 6524 4628 6558 4662
rect 6618 4613 6652 4647
rect 6712 4598 6746 4632
rect 6828 4613 6862 4647
rect 6928 4613 6962 4647
rect 7028 4613 7062 4647
rect 7128 4613 7162 4647
rect 7228 4613 7262 4647
rect 7328 4613 7362 4647
rect 7428 4613 7462 4647
rect 6324 4473 6358 4507
rect 6412 4473 6446 4507
rect 6524 4488 6558 4522
rect 6618 4473 6652 4507
rect 6712 4458 6746 4492
rect 6828 4473 6862 4507
rect 6928 4473 6962 4507
rect 7028 4473 7062 4507
rect 7128 4473 7162 4507
rect 7228 4473 7262 4507
rect 7328 4473 7362 4507
rect 7428 4473 7462 4507
rect 6324 4333 6358 4367
rect 6412 4333 6446 4367
rect 6524 4348 6558 4382
rect 6618 4333 6652 4367
rect 6712 4318 6746 4352
rect 6828 4333 6862 4367
rect 6928 4333 6962 4367
rect 7028 4333 7062 4367
rect 7128 4333 7162 4367
rect 7228 4333 7262 4367
rect 7328 4333 7362 4367
rect 7428 4333 7462 4367
rect 5924 4193 5958 4227
rect 6018 4193 6052 4227
rect 6118 4193 6152 4227
rect 6318 4193 6352 4227
rect 6412 4193 6446 4227
rect 6524 4208 6558 4242
rect 6618 4193 6652 4227
rect 6712 4178 6746 4212
rect 6828 4193 6862 4227
rect 6928 4193 6962 4227
rect 7028 4193 7062 4227
rect 7128 4193 7162 4227
rect 7228 4193 7262 4227
rect 7328 4193 7362 4227
rect 7428 4193 7462 4227
rect 5724 4053 5758 4087
rect 5818 4053 5852 4087
rect 6118 4053 6152 4087
rect 6218 4053 6252 4087
rect 6318 4053 6352 4087
rect 6412 4053 6446 4087
rect 6524 4068 6558 4102
rect 6618 4053 6652 4087
rect 6712 4038 6746 4072
rect 6828 4053 6862 4087
rect 6928 4053 6962 4087
rect 7028 4053 7062 4087
rect 7128 4053 7162 4087
rect 7228 4053 7262 4087
rect 7328 4053 7362 4087
rect 7428 4053 7462 4087
rect 4624 3913 4658 3947
rect 4718 3913 4752 3947
rect 5018 3913 5052 3947
rect 5118 3913 5152 3947
rect 5418 3913 5452 3947
rect 5518 3913 5552 3947
rect 5718 3913 5752 3947
rect 5818 3913 5852 3947
rect 5918 3913 5952 3947
rect 6012 3913 6046 3947
rect 3524 3773 3558 3807
rect 3618 3773 3652 3807
rect 3718 3773 3752 3807
rect 4618 3773 4652 3807
rect 4712 3773 4746 3807
rect 2324 3543 2358 3577
rect 2418 3543 2452 3577
rect 2518 3543 2552 3577
rect 2618 3543 2652 3577
rect 2718 3543 2752 3577
rect 3018 3543 3052 3577
rect 3118 3543 3152 3577
rect 3418 3543 3452 3577
rect 3512 3543 3546 3577
rect 2024 3403 2058 3437
rect 2118 3403 2152 3437
rect 2218 3403 2252 3437
rect 2318 3403 2352 3437
rect 2418 3403 2452 3437
rect 2518 3403 2552 3437
rect 2618 3403 2652 3437
rect 2718 3403 2752 3437
rect 2812 3403 2846 3437
rect 1324 3263 1358 3297
rect 1418 3263 1452 3297
rect 1518 3263 1552 3297
rect 1718 3263 1752 3297
rect 1818 3263 1852 3297
rect 1918 3263 1952 3297
rect 2018 3263 2052 3297
rect 2118 3263 2152 3297
rect 2218 3263 2252 3297
rect 2318 3263 2352 3297
rect 2418 3263 2452 3297
rect 2518 3263 2552 3297
rect 2618 3263 2652 3297
rect 2712 3263 2746 3297
rect 1224 3123 1258 3157
rect 1318 3123 1352 3157
rect 1718 3123 1752 3157
rect 1818 3123 1852 3157
rect 1918 3123 1952 3157
rect 2018 3123 2052 3157
rect 2118 3123 2152 3157
rect 2318 3123 2352 3157
rect 2412 3123 2446 3157
rect 3624 3543 3658 3577
rect 3712 3543 3746 3577
rect 3824 3543 3858 3577
rect 3918 3543 3952 3577
rect 4018 3543 4052 3577
rect 4118 3543 4152 3577
rect 4212 3543 4246 3577
rect 4824 3773 4858 3807
rect 4918 3773 4952 3807
rect 5018 3773 5052 3807
rect 5418 3773 5452 3807
rect 5518 3773 5552 3807
rect 5612 3773 5646 3807
rect 4324 3543 4358 3577
rect 4418 3543 4452 3577
rect 4618 3543 4652 3577
rect 4712 3543 4746 3577
rect 4824 3543 4858 3577
rect 4918 3543 4952 3577
rect 5118 3543 5152 3577
rect 5212 3543 5246 3577
rect 6124 3913 6158 3947
rect 6218 3913 6252 3947
rect 6318 3913 6352 3947
rect 6524 3928 6558 3962
rect 6618 3913 6652 3947
rect 6712 3898 6746 3932
rect 6828 3913 6862 3947
rect 6928 3913 6962 3947
rect 7028 3913 7062 3947
rect 7128 3913 7162 3947
rect 7228 3913 7262 3947
rect 7328 3913 7362 3947
rect 7428 3913 7462 3947
rect 5724 3773 5758 3807
rect 5818 3773 5852 3807
rect 6018 3773 6052 3807
rect 6118 3773 6152 3807
rect 6218 3773 6252 3807
rect 6318 3773 6352 3807
rect 6524 3788 6558 3822
rect 6618 3773 6652 3807
rect 6712 3758 6746 3792
rect 6828 3773 6862 3807
rect 6928 3773 6962 3807
rect 7028 3773 7062 3807
rect 7128 3773 7162 3807
rect 7228 3773 7262 3807
rect 7328 3773 7362 3807
rect 7428 3773 7462 3807
rect 5324 3543 5358 3577
rect 5418 3543 5452 3577
rect 5518 3543 5552 3577
rect 5618 3543 5652 3577
rect 5718 3543 5752 3577
rect 5818 3543 5852 3577
rect 5918 3543 5952 3577
rect 6218 3543 6252 3577
rect 6318 3543 6352 3577
rect 6412 3543 6446 3577
rect 6524 3558 6558 3592
rect 6618 3543 6652 3577
rect 6712 3528 6746 3562
rect 6828 3543 6862 3577
rect 6928 3543 6962 3577
rect 7028 3543 7062 3577
rect 7128 3543 7162 3577
rect 7228 3543 7262 3577
rect 7328 3543 7362 3577
rect 7428 3543 7462 3577
rect 2924 3403 2958 3437
rect 3018 3403 3052 3437
rect 3118 3403 3152 3437
rect 3218 3403 3252 3437
rect 3318 3403 3352 3437
rect 3418 3403 3452 3437
rect 3518 3403 3552 3437
rect 3918 3403 3952 3437
rect 4018 3403 4052 3437
rect 4118 3403 4152 3437
rect 4218 3403 4252 3437
rect 4618 3403 4652 3437
rect 4718 3403 4752 3437
rect 5018 3403 5052 3437
rect 5118 3403 5152 3437
rect 5218 3403 5252 3437
rect 5318 3403 5352 3437
rect 5418 3403 5452 3437
rect 5518 3403 5552 3437
rect 5618 3403 5652 3437
rect 5818 3403 5852 3437
rect 5912 3403 5946 3437
rect 2824 3263 2858 3297
rect 2912 3263 2946 3297
rect 3024 3263 3058 3297
rect 3118 3263 3152 3297
rect 3618 3263 3652 3297
rect 3718 3263 3752 3297
rect 3818 3263 3852 3297
rect 3918 3263 3952 3297
rect 4218 3263 4252 3297
rect 4312 3263 4346 3297
rect 2524 3123 2558 3157
rect 2618 3123 2652 3157
rect 3118 3123 3152 3157
rect 3212 3123 3246 3157
rect 3324 3123 3358 3157
rect 3418 3123 3452 3157
rect 3518 3123 3552 3157
rect 3612 3123 3646 3157
rect 118 2983 152 3017
rect 218 2983 252 3017
rect 418 2983 452 3017
rect 518 2983 552 3017
rect 618 2983 652 3017
rect 718 2983 752 3017
rect 818 2983 852 3017
rect 1018 2983 1052 3017
rect 1118 2983 1152 3017
rect 1618 2983 1652 3017
rect 1718 2983 1752 3017
rect 2018 2983 2052 3017
rect 2118 2983 2152 3017
rect 2518 2983 2552 3017
rect 2618 2983 2652 3017
rect 2718 2983 2752 3017
rect 2818 2983 2852 3017
rect 3218 2983 3252 3017
rect 3312 2983 3346 3017
rect 118 2843 152 2877
rect 218 2843 252 2877
rect 312 2843 346 2877
rect 424 2843 458 2877
rect 518 2843 552 2877
rect 618 2843 652 2877
rect 712 2843 746 2877
rect 824 2843 858 2877
rect 918 2843 952 2877
rect 1018 2843 1052 2877
rect 1118 2843 1152 2877
rect 1218 2843 1252 2877
rect 1318 2843 1352 2877
rect 1412 2843 1446 2877
rect 118 2703 152 2737
rect 218 2703 252 2737
rect 318 2703 352 2737
rect 518 2703 552 2737
rect 618 2703 652 2737
rect 818 2703 852 2737
rect 918 2703 952 2737
rect 1118 2703 1152 2737
rect 1218 2703 1252 2737
rect 1312 2703 1346 2737
rect 1524 2843 1558 2877
rect 1618 2843 1652 2877
rect 1918 2843 1952 2877
rect 2018 2843 2052 2877
rect 2112 2843 2146 2877
rect 1424 2703 1458 2737
rect 1512 2703 1546 2737
rect 218 2563 252 2597
rect 318 2563 352 2597
rect 518 2563 552 2597
rect 618 2563 652 2597
rect 718 2563 752 2597
rect 1018 2563 1052 2597
rect 1118 2563 1152 2597
rect 1418 2563 1452 2597
rect 1512 2563 1546 2597
rect 1624 2703 1658 2737
rect 1718 2703 1752 2737
rect 1818 2703 1852 2737
rect 1918 2703 1952 2737
rect 2012 2703 2046 2737
rect 2224 2843 2258 2877
rect 2312 2843 2346 2877
rect 2424 2843 2458 2877
rect 2512 2843 2546 2877
rect 2624 2843 2658 2877
rect 2718 2843 2752 2877
rect 2918 2843 2952 2877
rect 3012 2843 3046 2877
rect 2124 2703 2158 2737
rect 2218 2703 2252 2737
rect 2518 2703 2552 2737
rect 2618 2703 2652 2737
rect 2718 2703 2752 2737
rect 2812 2703 2846 2737
rect 1624 2563 1658 2597
rect 1718 2563 1752 2597
rect 1818 2563 1852 2597
rect 2018 2563 2052 2597
rect 2112 2563 2146 2597
rect 2224 2563 2258 2597
rect 2318 2563 2352 2597
rect 2412 2563 2446 2597
rect 2524 2563 2558 2597
rect 2612 2563 2646 2597
rect 3724 3123 3758 3157
rect 3818 3123 3852 3157
rect 3918 3123 3952 3157
rect 4118 3123 4152 3157
rect 4212 3123 4246 3157
rect 3424 2983 3458 3017
rect 3518 2983 3552 3017
rect 3618 2983 3652 3017
rect 3718 2983 3752 3017
rect 3812 2983 3846 3017
rect 3924 2983 3958 3017
rect 4012 2983 4046 3017
rect 4424 3263 4458 3297
rect 4518 3263 4552 3297
rect 4618 3263 4652 3297
rect 4718 3263 4752 3297
rect 4812 3263 4846 3297
rect 4324 3123 4358 3157
rect 4418 3123 4452 3157
rect 4512 3123 4546 3157
rect 4124 2983 4158 3017
rect 4218 2983 4252 3017
rect 4318 2983 4352 3017
rect 4418 2983 4452 3017
rect 4512 2983 4546 3017
rect 4624 3123 4658 3157
rect 4712 3123 4746 3157
rect 4924 3263 4958 3297
rect 5018 3263 5052 3297
rect 5218 3263 5252 3297
rect 5318 3263 5352 3297
rect 5418 3263 5452 3297
rect 5512 3263 5546 3297
rect 4824 3123 4858 3157
rect 4918 3123 4952 3157
rect 5012 3123 5046 3157
rect 5124 3123 5158 3157
rect 5218 3123 5252 3157
rect 5418 3123 5452 3157
rect 5512 3123 5546 3157
rect 6024 3403 6058 3437
rect 6118 3403 6152 3437
rect 6218 3403 6252 3437
rect 6318 3403 6352 3437
rect 6524 3418 6558 3452
rect 6618 3403 6652 3437
rect 6712 3388 6746 3422
rect 6828 3403 6862 3437
rect 6928 3403 6962 3437
rect 7028 3403 7062 3437
rect 7128 3403 7162 3437
rect 7228 3403 7262 3437
rect 7328 3403 7362 3437
rect 7428 3403 7462 3437
rect 5624 3263 5658 3297
rect 5718 3263 5752 3297
rect 5918 3263 5952 3297
rect 6018 3263 6052 3297
rect 6118 3263 6152 3297
rect 6218 3263 6252 3297
rect 6318 3263 6352 3297
rect 6524 3278 6558 3312
rect 6618 3263 6652 3297
rect 6712 3248 6746 3282
rect 6828 3263 6862 3297
rect 6928 3263 6962 3297
rect 7028 3263 7062 3297
rect 7128 3263 7162 3297
rect 7228 3263 7262 3297
rect 7328 3263 7362 3297
rect 7428 3263 7462 3297
rect 5624 3123 5658 3157
rect 5712 3123 5746 3157
rect 5824 3123 5858 3157
rect 5918 3123 5952 3157
rect 6018 3123 6052 3157
rect 6118 3123 6152 3157
rect 6524 3138 6558 3172
rect 6618 3123 6652 3157
rect 6712 3108 6746 3142
rect 6828 3123 6862 3157
rect 6928 3123 6962 3157
rect 7028 3123 7062 3157
rect 7128 3123 7162 3157
rect 7228 3123 7262 3157
rect 7328 3123 7362 3157
rect 7428 3123 7462 3157
rect 4624 2983 4658 3017
rect 4718 2983 4752 3017
rect 4918 2983 4952 3017
rect 5018 2983 5052 3017
rect 5118 2983 5152 3017
rect 5318 2983 5352 3017
rect 5418 2983 5452 3017
rect 5518 2983 5552 3017
rect 5618 2983 5652 3017
rect 5818 2983 5852 3017
rect 5912 2983 5946 3017
rect 6024 2983 6058 3017
rect 6118 2983 6152 3017
rect 6218 2983 6252 3017
rect 6524 2998 6558 3032
rect 6618 2983 6652 3017
rect 6712 2968 6746 3002
rect 6828 2983 6862 3017
rect 6928 2983 6962 3017
rect 7028 2983 7062 3017
rect 7128 2983 7162 3017
rect 7228 2983 7262 3017
rect 7328 2983 7362 3017
rect 7428 2983 7462 3017
rect 3124 2843 3158 2877
rect 3218 2843 3252 2877
rect 3318 2843 3352 2877
rect 3918 2843 3952 2877
rect 4018 2843 4052 2877
rect 4418 2843 4452 2877
rect 4518 2843 4552 2877
rect 4618 2843 4652 2877
rect 4818 2843 4852 2877
rect 4918 2843 4952 2877
rect 5018 2843 5052 2877
rect 5118 2843 5152 2877
rect 5218 2843 5252 2877
rect 5518 2843 5552 2877
rect 5618 2843 5652 2877
rect 5918 2843 5952 2877
rect 6012 2843 6046 2877
rect 2924 2703 2958 2737
rect 3018 2703 3052 2737
rect 3112 2703 3146 2737
rect 3224 2703 3258 2737
rect 3318 2703 3352 2737
rect 3418 2703 3452 2737
rect 3918 2703 3952 2737
rect 4018 2703 4052 2737
rect 4118 2703 4152 2737
rect 4318 2703 4352 2737
rect 4412 2703 4446 2737
rect 2724 2563 2758 2597
rect 2818 2563 2852 2597
rect 2918 2563 2952 2597
rect 3018 2563 3052 2597
rect 3118 2563 3152 2597
rect 3212 2563 3246 2597
rect 3324 2563 3358 2597
rect 3412 2563 3446 2597
rect 4524 2703 4558 2737
rect 4612 2703 4646 2737
rect 4724 2703 4758 2737
rect 4818 2703 4852 2737
rect 5018 2703 5052 2737
rect 5118 2703 5152 2737
rect 5318 2703 5352 2737
rect 5412 2703 5446 2737
rect 6124 2843 6158 2877
rect 6218 2843 6252 2877
rect 6318 2843 6352 2877
rect 6412 2843 6446 2877
rect 6524 2858 6558 2892
rect 6618 2843 6652 2877
rect 6712 2828 6746 2862
rect 6828 2843 6862 2877
rect 6928 2843 6962 2877
rect 7028 2843 7062 2877
rect 7128 2843 7162 2877
rect 7228 2843 7262 2877
rect 7328 2843 7362 2877
rect 7428 2843 7462 2877
rect 5524 2703 5558 2737
rect 5618 2703 5652 2737
rect 5718 2703 5752 2737
rect 6118 2703 6152 2737
rect 6218 2703 6252 2737
rect 6318 2703 6352 2737
rect 6524 2718 6558 2752
rect 6618 2703 6652 2737
rect 6712 2688 6746 2722
rect 6828 2703 6862 2737
rect 6928 2703 6962 2737
rect 7028 2703 7062 2737
rect 7128 2703 7162 2737
rect 7228 2703 7262 2737
rect 7328 2703 7362 2737
rect 7428 2703 7462 2737
rect 3524 2563 3558 2597
rect 3618 2563 3652 2597
rect 3718 2563 3752 2597
rect 3818 2563 3852 2597
rect 4018 2563 4052 2597
rect 4118 2563 4152 2597
rect 4218 2563 4252 2597
rect 4418 2563 4452 2597
rect 4518 2563 4552 2597
rect 4718 2563 4752 2597
rect 4818 2563 4852 2597
rect 5018 2563 5052 2597
rect 5118 2563 5152 2597
rect 5218 2563 5252 2597
rect 5418 2563 5452 2597
rect 5512 2563 5546 2597
rect 5624 2563 5658 2597
rect 5718 2563 5752 2597
rect 5918 2563 5952 2597
rect 6018 2563 6052 2597
rect 6218 2563 6252 2597
rect 6318 2563 6352 2597
rect 6524 2578 6558 2612
rect 6618 2563 6652 2597
rect 6712 2548 6746 2582
rect 6828 2563 6862 2597
rect 6928 2563 6962 2597
rect 7028 2563 7062 2597
rect 7128 2563 7162 2597
rect 7228 2563 7262 2597
rect 7328 2563 7362 2597
rect 7428 2563 7462 2597
rect 418 2333 452 2367
rect 518 2333 552 2367
rect 818 2333 852 2367
rect 918 2333 952 2367
rect 1018 2333 1052 2367
rect 1518 2333 1552 2367
rect 1618 2333 1652 2367
rect 1818 2333 1852 2367
rect 1918 2333 1952 2367
rect 2018 2333 2052 2367
rect 2118 2333 2152 2367
rect 2318 2333 2352 2367
rect 2418 2333 2452 2367
rect 2518 2333 2552 2367
rect 2718 2333 2752 2367
rect 2818 2333 2852 2367
rect 3318 2333 3352 2367
rect 3418 2333 3452 2367
rect 4018 2333 4052 2367
rect 4118 2333 4152 2367
rect 4318 2333 4352 2367
rect 4418 2333 4452 2367
rect 4718 2333 4752 2367
rect 4818 2333 4852 2367
rect 4918 2333 4952 2367
rect 5018 2333 5052 2367
rect 5318 2333 5352 2367
rect 5412 2333 5446 2367
rect 24 2193 58 2227
rect 118 2193 152 2227
rect 212 2193 246 2227
rect 324 2193 358 2227
rect 418 2193 452 2227
rect 518 2193 552 2227
rect 618 2193 652 2227
rect 1018 2193 1052 2227
rect 1118 2193 1152 2227
rect 1218 2193 1252 2227
rect 1312 2193 1346 2227
rect 24 2053 58 2087
rect 118 2053 152 2087
rect 218 2053 252 2087
rect 312 2053 346 2087
rect 218 1913 252 1947
rect 312 1913 346 1947
rect 424 2053 458 2087
rect 518 2053 552 2087
rect 618 2053 652 2087
rect 818 2053 852 2087
rect 918 2053 952 2087
rect 1218 2053 1252 2087
rect 1312 2053 1346 2087
rect 1424 2193 1458 2227
rect 1512 2193 1546 2227
rect 1424 2053 1458 2087
rect 1512 2053 1546 2087
rect 424 1913 458 1947
rect 518 1913 552 1947
rect 718 1913 752 1947
rect 818 1913 852 1947
rect 918 1913 952 1947
rect 1018 1913 1052 1947
rect 1118 1913 1152 1947
rect 1218 1913 1252 1947
rect 1318 1913 1352 1947
rect 1412 1913 1446 1947
rect 118 1773 152 1807
rect 218 1773 252 1807
rect 718 1773 752 1807
rect 818 1773 852 1807
rect 912 1773 946 1807
rect 24 1633 58 1667
rect 112 1633 146 1667
rect 24 1493 58 1527
rect 112 1493 146 1527
rect 224 1633 258 1667
rect 318 1633 352 1667
rect 418 1633 452 1667
rect 618 1633 652 1667
rect 712 1633 746 1667
rect 224 1493 258 1527
rect 318 1493 352 1527
rect 412 1493 446 1527
rect 118 1353 152 1387
rect 212 1353 246 1387
rect 824 1633 858 1667
rect 912 1633 946 1667
rect 1624 2193 1658 2227
rect 1718 2193 1752 2227
rect 1812 2193 1846 2227
rect 1624 2053 1658 2087
rect 1718 2053 1752 2087
rect 1812 2053 1846 2087
rect 1924 2193 1958 2227
rect 2018 2193 2052 2227
rect 2118 2193 2152 2227
rect 2212 2193 2246 2227
rect 1924 2053 1958 2087
rect 2018 2053 2052 2087
rect 2118 2053 2152 2087
rect 2212 2053 2246 2087
rect 2324 2193 2358 2227
rect 2418 2193 2452 2227
rect 2618 2193 2652 2227
rect 2718 2193 2752 2227
rect 2812 2193 2846 2227
rect 2324 2053 2358 2087
rect 2412 2053 2446 2087
rect 1524 1913 1558 1947
rect 1618 1913 1652 1947
rect 1718 1913 1752 1947
rect 1818 1913 1852 1947
rect 1918 1913 1952 1947
rect 2018 1913 2052 1947
rect 2318 1913 2352 1947
rect 2412 1913 2446 1947
rect 1024 1773 1058 1807
rect 1118 1773 1152 1807
rect 1418 1773 1452 1807
rect 1518 1773 1552 1807
rect 1718 1773 1752 1807
rect 1812 1773 1846 1807
rect 1024 1633 1058 1667
rect 1118 1633 1152 1667
rect 1218 1633 1252 1667
rect 1318 1633 1352 1667
rect 1418 1633 1452 1667
rect 1512 1633 1546 1667
rect 1624 1633 1658 1667
rect 1712 1633 1746 1667
rect 524 1493 558 1527
rect 618 1493 652 1527
rect 818 1493 852 1527
rect 918 1493 952 1527
rect 1118 1493 1152 1527
rect 1218 1493 1252 1527
rect 1318 1493 1352 1527
rect 1518 1493 1552 1527
rect 1612 1493 1646 1527
rect 324 1353 358 1387
rect 418 1353 452 1387
rect 512 1353 546 1387
rect 218 1123 252 1157
rect 312 1123 346 1157
rect 624 1353 658 1387
rect 718 1353 752 1387
rect 1018 1353 1052 1387
rect 1118 1353 1152 1387
rect 1318 1353 1352 1387
rect 1418 1353 1452 1387
rect 1512 1353 1546 1387
rect 424 1123 458 1157
rect 512 1123 546 1157
rect 624 1123 658 1157
rect 712 1123 746 1157
rect 824 1123 858 1157
rect 918 1123 952 1157
rect 1018 1123 1052 1157
rect 1118 1123 1152 1157
rect 1212 1123 1246 1157
rect 118 983 152 1017
rect 218 983 252 1017
rect 518 983 552 1017
rect 618 983 652 1017
rect 818 983 852 1017
rect 912 983 946 1017
rect 1024 983 1058 1017
rect 1112 983 1146 1017
rect 918 843 952 877
rect 1012 843 1046 877
rect 24 703 58 737
rect 118 703 152 737
rect 218 703 252 737
rect 318 703 352 737
rect 618 703 652 737
rect 718 703 752 737
rect 818 703 852 737
rect 912 703 946 737
rect 218 563 252 597
rect 318 563 352 597
rect 418 563 452 597
rect 512 563 546 597
rect 118 423 152 457
rect 212 423 246 457
rect 324 423 358 457
rect 412 423 446 457
rect 2924 2193 2958 2227
rect 3018 2193 3052 2227
rect 3118 2193 3152 2227
rect 3218 2193 3252 2227
rect 3318 2193 3352 2227
rect 3418 2193 3452 2227
rect 3512 2193 3546 2227
rect 2524 2053 2558 2087
rect 2618 2053 2652 2087
rect 2718 2053 2752 2087
rect 2818 2053 2852 2087
rect 2918 2053 2952 2087
rect 3218 2053 3252 2087
rect 3312 2053 3346 2087
rect 2524 1913 2558 1947
rect 2618 1913 2652 1947
rect 2918 1913 2952 1947
rect 3012 1913 3046 1947
rect 3624 2193 3658 2227
rect 3718 2193 3752 2227
rect 3818 2193 3852 2227
rect 4018 2193 4052 2227
rect 4118 2193 4152 2227
rect 4212 2193 4246 2227
rect 3424 2053 3458 2087
rect 3518 2053 3552 2087
rect 3612 2053 3646 2087
rect 3724 2053 3758 2087
rect 3818 2053 3852 2087
rect 3912 2053 3946 2087
rect 3124 1913 3158 1947
rect 3218 1913 3252 1947
rect 3518 1913 3552 1947
rect 3618 1913 3652 1947
rect 3718 1913 3752 1947
rect 3812 1913 3846 1947
rect 1924 1773 1958 1807
rect 2018 1773 2052 1807
rect 2218 1773 2252 1807
rect 2318 1773 2352 1807
rect 2618 1773 2652 1807
rect 2718 1773 2752 1807
rect 2818 1773 2852 1807
rect 2918 1773 2952 1807
rect 3018 1773 3052 1807
rect 3318 1773 3352 1807
rect 3412 1773 3446 1807
rect 1824 1633 1858 1667
rect 1912 1633 1946 1667
rect 2024 1633 2058 1667
rect 2118 1633 2152 1667
rect 2218 1633 2252 1667
rect 2518 1633 2552 1667
rect 2612 1633 2646 1667
rect 2724 1633 2758 1667
rect 2818 1633 2852 1667
rect 2918 1633 2952 1667
rect 3018 1633 3052 1667
rect 3118 1633 3152 1667
rect 3318 1633 3352 1667
rect 3412 1633 3446 1667
rect 3524 1773 3558 1807
rect 3612 1773 3646 1807
rect 4324 2193 4358 2227
rect 4412 2193 4446 2227
rect 4024 2053 4058 2087
rect 4118 2053 4152 2087
rect 4318 2053 4352 2087
rect 4412 2053 4446 2087
rect 3924 1913 3958 1947
rect 4018 1913 4052 1947
rect 4118 1913 4152 1947
rect 4218 1913 4252 1947
rect 4318 1913 4352 1947
rect 4412 1913 4446 1947
rect 3724 1773 3758 1807
rect 3818 1773 3852 1807
rect 3912 1773 3946 1807
rect 3524 1633 3558 1667
rect 3618 1633 3652 1667
rect 3712 1633 3746 1667
rect 5524 2333 5558 2367
rect 5618 2333 5652 2367
rect 5718 2333 5752 2367
rect 5918 2333 5952 2367
rect 6018 2333 6052 2367
rect 6318 2333 6352 2367
rect 6412 2333 6446 2367
rect 6524 2348 6558 2382
rect 6618 2333 6652 2367
rect 6712 2318 6746 2352
rect 6828 2333 6862 2367
rect 6928 2333 6962 2367
rect 7028 2333 7062 2367
rect 7128 2333 7162 2367
rect 7228 2333 7262 2367
rect 7328 2333 7362 2367
rect 7428 2333 7462 2367
rect 4524 2193 4558 2227
rect 4618 2193 4652 2227
rect 4718 2193 4752 2227
rect 4918 2193 4952 2227
rect 5018 2193 5052 2227
rect 5118 2193 5152 2227
rect 5418 2193 5452 2227
rect 5518 2193 5552 2227
rect 5618 2193 5652 2227
rect 5718 2193 5752 2227
rect 5818 2193 5852 2227
rect 5918 2193 5952 2227
rect 6218 2193 6252 2227
rect 6318 2193 6352 2227
rect 6412 2193 6446 2227
rect 6524 2208 6558 2242
rect 6618 2193 6652 2227
rect 6712 2178 6746 2212
rect 6828 2193 6862 2227
rect 6928 2193 6962 2227
rect 7028 2193 7062 2227
rect 7128 2193 7162 2227
rect 7228 2193 7262 2227
rect 7328 2193 7362 2227
rect 7428 2193 7462 2227
rect 4524 2053 4558 2087
rect 4618 2053 4652 2087
rect 4718 2053 4752 2087
rect 4918 2053 4952 2087
rect 5018 2053 5052 2087
rect 5318 2053 5352 2087
rect 5418 2053 5452 2087
rect 5518 2053 5552 2087
rect 5618 2053 5652 2087
rect 5818 2053 5852 2087
rect 5918 2053 5952 2087
rect 6118 2053 6152 2087
rect 6218 2053 6252 2087
rect 6318 2053 6352 2087
rect 6524 2068 6558 2102
rect 6618 2053 6652 2087
rect 6712 2038 6746 2072
rect 6828 2053 6862 2087
rect 6928 2053 6962 2087
rect 7028 2053 7062 2087
rect 7128 2053 7162 2087
rect 7228 2053 7262 2087
rect 7328 2053 7362 2087
rect 7428 2053 7462 2087
rect 4524 1913 4558 1947
rect 4618 1913 4652 1947
rect 4718 1913 4752 1947
rect 4818 1913 4852 1947
rect 4912 1913 4946 1947
rect 4024 1773 4058 1807
rect 4118 1773 4152 1807
rect 4318 1773 4352 1807
rect 4418 1773 4452 1807
rect 4518 1773 4552 1807
rect 4718 1773 4752 1807
rect 4812 1773 4846 1807
rect 3824 1633 3858 1667
rect 3918 1633 3952 1667
rect 4018 1633 4052 1667
rect 4218 1633 4252 1667
rect 4318 1633 4352 1667
rect 4412 1633 4446 1667
rect 1724 1493 1758 1527
rect 1818 1493 1852 1527
rect 1918 1493 1952 1527
rect 2018 1493 2052 1527
rect 2118 1493 2152 1527
rect 2218 1493 2252 1527
rect 2418 1493 2452 1527
rect 2518 1493 2552 1527
rect 2618 1493 2652 1527
rect 2718 1493 2752 1527
rect 3018 1493 3052 1527
rect 3118 1493 3152 1527
rect 3218 1493 3252 1527
rect 3318 1493 3352 1527
rect 3418 1493 3452 1527
rect 3618 1493 3652 1527
rect 3718 1493 3752 1527
rect 3918 1493 3952 1527
rect 4018 1493 4052 1527
rect 4112 1493 4146 1527
rect 1624 1353 1658 1387
rect 1712 1353 1746 1387
rect 1824 1353 1858 1387
rect 1918 1353 1952 1387
rect 2218 1353 2252 1387
rect 2318 1353 2352 1387
rect 2418 1353 2452 1387
rect 2718 1353 2752 1387
rect 2818 1353 2852 1387
rect 2912 1353 2946 1387
rect 1324 1123 1358 1157
rect 1418 1123 1452 1157
rect 1618 1123 1652 1157
rect 1718 1123 1752 1157
rect 1818 1123 1852 1157
rect 1918 1123 1952 1157
rect 2118 1123 2152 1157
rect 2218 1123 2252 1157
rect 2318 1123 2352 1157
rect 2418 1123 2452 1157
rect 2512 1123 2546 1157
rect 1224 983 1258 1017
rect 1318 983 1352 1017
rect 1518 983 1552 1017
rect 1618 983 1652 1017
rect 1818 983 1852 1017
rect 1918 983 1952 1017
rect 2018 983 2052 1017
rect 2112 983 2146 1017
rect 1124 843 1158 877
rect 1218 843 1252 877
rect 1318 843 1352 877
rect 1518 843 1552 877
rect 1618 843 1652 877
rect 1712 843 1746 877
rect 2224 983 2258 1017
rect 2318 983 2352 1017
rect 2412 983 2446 1017
rect 2624 1123 2658 1157
rect 2712 1123 2746 1157
rect 3024 1353 3058 1387
rect 3118 1353 3152 1387
rect 3318 1353 3352 1387
rect 3418 1353 3452 1387
rect 3512 1353 3546 1387
rect 3624 1353 3658 1387
rect 3718 1353 3752 1387
rect 3812 1353 3846 1387
rect 4224 1493 4258 1527
rect 4318 1493 4352 1527
rect 4412 1493 4446 1527
rect 5024 1913 5058 1947
rect 5112 1913 5146 1947
rect 5224 1913 5258 1947
rect 5312 1913 5346 1947
rect 5424 1913 5458 1947
rect 5518 1913 5552 1947
rect 5618 1913 5652 1947
rect 5712 1913 5746 1947
rect 5824 1913 5858 1947
rect 5918 1913 5952 1947
rect 6012 1913 6046 1947
rect 6124 1913 6158 1947
rect 6218 1913 6252 1947
rect 6524 1928 6558 1962
rect 6618 1913 6652 1947
rect 6712 1898 6746 1932
rect 6828 1913 6862 1947
rect 6928 1913 6962 1947
rect 7028 1913 7062 1947
rect 7128 1913 7162 1947
rect 7228 1913 7262 1947
rect 7328 1913 7362 1947
rect 7428 1913 7462 1947
rect 4924 1773 4958 1807
rect 5018 1773 5052 1807
rect 5318 1773 5352 1807
rect 5418 1773 5452 1807
rect 5518 1773 5552 1807
rect 5718 1773 5752 1807
rect 5818 1773 5852 1807
rect 6118 1773 6152 1807
rect 6218 1773 6252 1807
rect 6318 1773 6352 1807
rect 6524 1788 6558 1822
rect 6618 1773 6652 1807
rect 6712 1758 6746 1792
rect 6828 1773 6862 1807
rect 6928 1773 6962 1807
rect 7028 1773 7062 1807
rect 7128 1773 7162 1807
rect 7228 1773 7262 1807
rect 7328 1773 7362 1807
rect 7428 1773 7462 1807
rect 4524 1633 4558 1667
rect 4618 1633 4652 1667
rect 4818 1633 4852 1667
rect 4918 1633 4952 1667
rect 5018 1633 5052 1667
rect 5118 1633 5152 1667
rect 5218 1633 5252 1667
rect 5312 1633 5346 1667
rect 4524 1493 4558 1527
rect 4618 1493 4652 1527
rect 4918 1493 4952 1527
rect 5012 1493 5046 1527
rect 3924 1353 3958 1387
rect 4018 1353 4052 1387
rect 4118 1353 4152 1387
rect 4218 1353 4252 1387
rect 4718 1353 4752 1387
rect 4812 1353 4846 1387
rect 2824 1123 2858 1157
rect 2918 1123 2952 1157
rect 3118 1123 3152 1157
rect 3218 1123 3252 1157
rect 3318 1123 3352 1157
rect 3618 1123 3652 1157
rect 3718 1123 3752 1157
rect 4118 1123 4152 1157
rect 4212 1123 4246 1157
rect 2524 983 2558 1017
rect 2618 983 2652 1017
rect 2718 983 2752 1017
rect 2818 983 2852 1017
rect 3018 983 3052 1017
rect 3118 983 3152 1017
rect 3218 983 3252 1017
rect 3418 983 3452 1017
rect 3518 983 3552 1017
rect 3718 983 3752 1017
rect 3818 983 3852 1017
rect 4118 983 4152 1017
rect 4212 983 4246 1017
rect 4924 1353 4958 1387
rect 5012 1353 5046 1387
rect 5124 1493 5158 1527
rect 5212 1493 5246 1527
rect 5424 1633 5458 1667
rect 5518 1633 5552 1667
rect 5618 1633 5652 1667
rect 5712 1633 5746 1667
rect 5324 1493 5358 1527
rect 5412 1493 5446 1527
rect 5524 1493 5558 1527
rect 5618 1493 5652 1527
rect 5712 1493 5746 1527
rect 5824 1633 5858 1667
rect 5912 1633 5946 1667
rect 5824 1493 5858 1527
rect 5912 1493 5946 1527
rect 6024 1633 6058 1667
rect 6118 1633 6152 1667
rect 6218 1633 6252 1667
rect 6524 1648 6558 1682
rect 6618 1633 6652 1667
rect 6712 1618 6746 1652
rect 6828 1633 6862 1667
rect 6928 1633 6962 1667
rect 7028 1633 7062 1667
rect 7128 1633 7162 1667
rect 7228 1633 7262 1667
rect 7328 1633 7362 1667
rect 7428 1633 7462 1667
rect 6024 1493 6058 1527
rect 6118 1493 6152 1527
rect 6212 1493 6246 1527
rect 5124 1353 5158 1387
rect 5218 1353 5252 1387
rect 5518 1353 5552 1387
rect 5618 1353 5652 1387
rect 5718 1353 5752 1387
rect 5918 1353 5952 1387
rect 6018 1353 6052 1387
rect 6112 1353 6146 1387
rect 4324 1123 4358 1157
rect 4418 1123 4452 1157
rect 4718 1123 4752 1157
rect 4818 1123 4852 1157
rect 4918 1123 4952 1157
rect 5118 1123 5152 1157
rect 5218 1123 5252 1157
rect 5318 1123 5352 1157
rect 5412 1123 5446 1157
rect 4324 983 4358 1017
rect 4418 983 4452 1017
rect 4518 983 4552 1017
rect 4618 983 4652 1017
rect 4718 983 4752 1017
rect 4812 983 4846 1017
rect 1824 843 1858 877
rect 1918 843 1952 877
rect 2018 843 2052 877
rect 2118 843 2152 877
rect 2218 843 2252 877
rect 2318 843 2352 877
rect 2418 843 2452 877
rect 2518 843 2552 877
rect 2818 843 2852 877
rect 2918 843 2952 877
rect 3118 843 3152 877
rect 3218 843 3252 877
rect 3318 843 3352 877
rect 3918 843 3952 877
rect 4018 843 4052 877
rect 4118 843 4152 877
rect 4218 843 4252 877
rect 4312 843 4346 877
rect 1024 703 1058 737
rect 1118 703 1152 737
rect 1818 703 1852 737
rect 1918 703 1952 737
rect 2012 703 2046 737
rect 624 563 658 597
rect 718 563 752 597
rect 918 563 952 597
rect 1012 563 1046 597
rect 2124 703 2158 737
rect 2212 703 2246 737
rect 4424 843 4458 877
rect 4512 843 4546 877
rect 2324 703 2358 737
rect 2418 703 2452 737
rect 2718 703 2752 737
rect 2818 703 2852 737
rect 2918 703 2952 737
rect 3018 703 3052 737
rect 3118 703 3152 737
rect 3218 703 3252 737
rect 3518 703 3552 737
rect 3618 703 3652 737
rect 3918 703 3952 737
rect 4018 703 4052 737
rect 4118 703 4152 737
rect 4318 703 4352 737
rect 4412 703 4446 737
rect 1124 563 1158 597
rect 1218 563 1252 597
rect 1518 563 1552 597
rect 1618 563 1652 597
rect 1818 563 1852 597
rect 1918 563 1952 597
rect 2018 563 2052 597
rect 2118 563 2152 597
rect 2518 563 2552 597
rect 2618 563 2652 597
rect 2718 563 2752 597
rect 3118 563 3152 597
rect 3218 563 3252 597
rect 3518 563 3552 597
rect 3618 563 3652 597
rect 3712 563 3746 597
rect 524 423 558 457
rect 618 423 652 457
rect 718 423 752 457
rect 818 423 852 457
rect 918 423 952 457
rect 1018 423 1052 457
rect 1218 423 1252 457
rect 1318 423 1352 457
rect 1412 423 1446 457
rect 118 283 152 317
rect 218 283 252 317
rect 418 283 452 317
rect 518 283 552 317
rect 612 283 646 317
rect 1524 423 1558 457
rect 1618 423 1652 457
rect 1818 423 1852 457
rect 1918 423 1952 457
rect 2018 423 2052 457
rect 2218 423 2252 457
rect 2318 423 2352 457
rect 2718 423 2752 457
rect 2818 423 2852 457
rect 2918 423 2952 457
rect 3012 423 3046 457
rect 724 283 758 317
rect 818 283 852 317
rect 918 283 952 317
rect 1418 283 1452 317
rect 1512 283 1546 317
rect 24 143 58 177
rect 118 143 152 177
rect 218 143 252 177
rect 318 143 352 177
rect 418 143 452 177
rect 618 143 652 177
rect 718 143 752 177
rect 812 143 846 177
rect 1624 283 1658 317
rect 1718 283 1752 317
rect 2018 283 2052 317
rect 2118 283 2152 317
rect 2212 283 2246 317
rect 924 143 958 177
rect 1018 143 1052 177
rect 1318 143 1352 177
rect 1418 143 1452 177
rect 1518 143 1552 177
rect 1718 143 1752 177
rect 1818 143 1852 177
rect 1912 143 1946 177
rect 2324 283 2358 317
rect 2412 283 2446 317
rect 2524 283 2558 317
rect 2612 283 2646 317
rect 2724 283 2758 317
rect 2812 283 2846 317
rect 3124 423 3158 457
rect 3212 423 3246 457
rect 3324 423 3358 457
rect 3418 423 3452 457
rect 3512 423 3546 457
rect 2924 283 2958 317
rect 3018 283 3052 317
rect 3118 283 3152 317
rect 3318 283 3352 317
rect 3418 283 3452 317
rect 3512 283 3546 317
rect 2024 143 2058 177
rect 2118 143 2152 177
rect 2218 143 2252 177
rect 2418 143 2452 177
rect 2518 143 2552 177
rect 2618 143 2652 177
rect 3018 143 3052 177
rect 3118 143 3152 177
rect 3218 143 3252 177
rect 3418 143 3452 177
rect 3512 143 3546 177
rect 3624 423 3658 457
rect 3712 423 3746 457
rect 3824 563 3858 597
rect 3918 563 3952 597
rect 4012 563 4046 597
rect 4124 563 4158 597
rect 4212 563 4246 597
rect 4924 983 4958 1017
rect 5012 983 5046 1017
rect 5524 1123 5558 1157
rect 5618 1123 5652 1157
rect 5718 1123 5752 1157
rect 5818 1123 5852 1157
rect 5912 1123 5946 1157
rect 6324 1493 6358 1527
rect 6412 1493 6446 1527
rect 6524 1508 6558 1542
rect 6618 1493 6652 1527
rect 6712 1478 6746 1512
rect 6828 1493 6862 1527
rect 6928 1493 6962 1527
rect 7028 1493 7062 1527
rect 7128 1493 7162 1527
rect 7228 1493 7262 1527
rect 7328 1493 7362 1527
rect 7428 1493 7462 1527
rect 6224 1353 6258 1387
rect 6318 1353 6352 1387
rect 6524 1368 6558 1402
rect 6618 1353 6652 1387
rect 6712 1338 6746 1372
rect 6828 1353 6862 1387
rect 6928 1353 6962 1387
rect 7028 1353 7062 1387
rect 7128 1353 7162 1387
rect 7228 1353 7262 1387
rect 7328 1353 7362 1387
rect 7428 1353 7462 1387
rect 6024 1123 6058 1157
rect 6118 1123 6152 1157
rect 6218 1123 6252 1157
rect 6318 1123 6352 1157
rect 6412 1123 6446 1157
rect 6524 1138 6558 1172
rect 6618 1123 6652 1157
rect 6712 1108 6746 1142
rect 6828 1123 6862 1157
rect 6928 1123 6962 1157
rect 7028 1123 7062 1157
rect 7128 1123 7162 1157
rect 7228 1123 7262 1157
rect 7328 1123 7362 1157
rect 7428 1123 7462 1157
rect 5124 983 5158 1017
rect 5218 983 5252 1017
rect 5318 983 5352 1017
rect 5418 983 5452 1017
rect 5518 983 5552 1017
rect 5718 983 5752 1017
rect 5818 983 5852 1017
rect 6118 983 6152 1017
rect 6212 983 6246 1017
rect 6324 983 6358 1017
rect 6412 983 6446 1017
rect 6524 998 6558 1032
rect 6618 983 6652 1017
rect 6712 968 6746 1002
rect 6828 983 6862 1017
rect 6928 983 6962 1017
rect 7028 983 7062 1017
rect 7128 983 7162 1017
rect 7228 983 7262 1017
rect 7328 983 7362 1017
rect 7428 983 7462 1017
rect 4624 843 4658 877
rect 4718 843 4752 877
rect 4818 843 4852 877
rect 5018 843 5052 877
rect 5118 843 5152 877
rect 5218 843 5252 877
rect 5318 843 5352 877
rect 5618 843 5652 877
rect 5718 843 5752 877
rect 6018 843 6052 877
rect 6118 843 6152 877
rect 6524 858 6558 892
rect 6618 843 6652 877
rect 6712 828 6746 862
rect 6828 843 6862 877
rect 6928 843 6962 877
rect 7028 843 7062 877
rect 7128 843 7162 877
rect 7228 843 7262 877
rect 7328 843 7362 877
rect 7428 843 7462 877
rect 4524 703 4558 737
rect 4618 703 4652 737
rect 4818 703 4852 737
rect 4918 703 4952 737
rect 5018 703 5052 737
rect 5318 703 5352 737
rect 5418 703 5452 737
rect 5512 703 5546 737
rect 4324 563 4358 597
rect 4418 563 4452 597
rect 4518 563 4552 597
rect 4612 563 4646 597
rect 4724 563 4758 597
rect 4818 563 4852 597
rect 5018 563 5052 597
rect 5118 563 5152 597
rect 5212 563 5246 597
rect 5624 703 5658 737
rect 5712 703 5746 737
rect 5824 703 5858 737
rect 5918 703 5952 737
rect 6018 703 6052 737
rect 6218 703 6252 737
rect 6318 703 6352 737
rect 6524 718 6558 752
rect 6618 703 6652 737
rect 6712 688 6746 722
rect 6828 703 6862 737
rect 6928 703 6962 737
rect 7028 703 7062 737
rect 7128 703 7162 737
rect 7228 703 7262 737
rect 7328 703 7362 737
rect 7428 703 7462 737
rect 5324 563 5358 597
rect 5418 563 5452 597
rect 5718 563 5752 597
rect 5818 563 5852 597
rect 5918 563 5952 597
rect 6012 563 6046 597
rect 3824 423 3858 457
rect 3918 423 3952 457
rect 4018 423 4052 457
rect 4318 423 4352 457
rect 4418 423 4452 457
rect 4518 423 4552 457
rect 4618 423 4652 457
rect 4818 423 4852 457
rect 4918 423 4952 457
rect 5018 423 5052 457
rect 5118 423 5152 457
rect 5218 423 5252 457
rect 5318 423 5352 457
rect 5418 423 5452 457
rect 5512 423 5546 457
rect 6124 563 6158 597
rect 6218 563 6252 597
rect 6318 563 6352 597
rect 6412 563 6446 597
rect 6524 578 6558 612
rect 6618 563 6652 597
rect 6712 548 6746 582
rect 6828 563 6862 597
rect 6928 563 6962 597
rect 7028 563 7062 597
rect 7128 563 7162 597
rect 7228 563 7262 597
rect 7328 563 7362 597
rect 7428 563 7462 597
rect 5624 423 5658 457
rect 5718 423 5752 457
rect 6018 423 6052 457
rect 6118 423 6152 457
rect 6212 423 6246 457
rect 3624 283 3658 317
rect 3718 283 3752 317
rect 3818 283 3852 317
rect 3918 283 3952 317
rect 4118 283 4152 317
rect 4218 283 4252 317
rect 4318 283 4352 317
rect 4418 283 4452 317
rect 4518 283 4552 317
rect 4618 283 4652 317
rect 4718 283 4752 317
rect 5118 283 5152 317
rect 5218 283 5252 317
rect 5518 283 5552 317
rect 5612 283 5646 317
rect 3624 143 3658 177
rect 3718 143 3752 177
rect 3918 143 3952 177
rect 4018 143 4052 177
rect 4418 143 4452 177
rect 4518 143 4552 177
rect 4618 143 4652 177
rect 4712 143 4746 177
rect 6324 423 6358 457
rect 6412 423 6446 457
rect 6524 438 6558 472
rect 6618 423 6652 457
rect 6712 408 6746 442
rect 6828 423 6862 457
rect 6928 423 6962 457
rect 7028 423 7062 457
rect 7128 423 7162 457
rect 7228 423 7262 457
rect 7328 423 7362 457
rect 7428 423 7462 457
rect 5724 283 5758 317
rect 5818 283 5852 317
rect 5918 283 5952 317
rect 6018 283 6052 317
rect 6118 283 6152 317
rect 6218 283 6252 317
rect 6318 283 6352 317
rect 6412 283 6446 317
rect 6524 298 6558 332
rect 6618 283 6652 317
rect 6712 268 6746 302
rect 6828 283 6862 317
rect 6928 283 6962 317
rect 7028 283 7062 317
rect 7128 283 7162 317
rect 7228 283 7262 317
rect 7328 283 7362 317
rect 7428 283 7462 317
rect 4824 143 4858 177
rect 4918 143 4952 177
rect 5018 143 5052 177
rect 5118 143 5152 177
rect 5218 143 5252 177
rect 5418 143 5452 177
rect 5518 143 5552 177
rect 5718 143 5752 177
rect 5818 143 5852 177
rect 6018 143 6052 177
rect 6112 143 6146 177
rect 6224 143 6258 177
rect 6318 143 6352 177
rect 6412 143 6446 177
rect 6524 158 6558 192
rect 6618 143 6652 177
rect 6712 128 6746 162
rect 6828 143 6862 177
rect 6928 143 6962 177
rect 7028 143 7062 177
rect 7128 143 7162 177
rect 7228 143 7262 177
rect 7328 143 7362 177
rect 7428 143 7462 177
rect 8162 -42 8196 -8
rect 8230 -42 8264 -8
rect 9278 -42 9312 -8
rect 9346 -42 9380 -8
rect -82 -183 -48 -149
rect 18 -183 52 -149
rect 118 -183 152 -149
rect 218 -183 252 -149
rect 318 -183 352 -149
rect 418 -183 452 -149
rect 518 -183 552 -149
rect 618 -183 652 -149
rect 718 -183 752 -149
rect 818 -183 852 -149
rect 918 -183 952 -149
rect 1018 -183 1052 -149
rect 1118 -183 1152 -149
rect 1218 -183 1252 -149
rect 1318 -183 1352 -149
rect 1418 -183 1452 -149
rect 1518 -183 1552 -149
rect 1618 -183 1652 -149
rect 1718 -183 1752 -149
rect 1818 -183 1852 -149
rect 1918 -183 1952 -149
rect 2018 -183 2052 -149
rect 2118 -183 2152 -149
rect 2218 -183 2252 -149
rect 2318 -183 2352 -149
rect 2418 -183 2452 -149
rect 2518 -183 2552 -149
rect 2618 -183 2652 -149
rect 2718 -183 2752 -149
rect 2818 -183 2852 -149
rect 2918 -183 2952 -149
rect 3018 -183 3052 -149
rect 3118 -183 3152 -149
rect 3218 -183 3252 -149
rect 3318 -183 3352 -149
rect 3418 -183 3452 -149
rect 3518 -183 3552 -149
rect 3618 -183 3652 -149
rect 3718 -183 3752 -149
rect 3818 -183 3852 -149
rect 3918 -183 3952 -149
rect 4018 -183 4052 -149
rect 4118 -183 4152 -149
rect 4218 -183 4252 -149
rect 4318 -183 4352 -149
rect 4418 -183 4452 -149
rect 4518 -183 4552 -149
rect 4618 -183 4652 -149
rect 4718 -183 4752 -149
rect 4818 -183 4852 -149
rect 4918 -183 4952 -149
rect 5018 -183 5052 -149
rect 5118 -183 5152 -149
rect 5218 -183 5252 -149
rect 5318 -183 5352 -149
rect 5418 -183 5452 -149
rect 5518 -183 5552 -149
rect 5618 -183 5652 -149
rect 5718 -183 5752 -149
rect 5818 -183 5852 -149
rect 5918 -183 5952 -149
rect 6018 -183 6052 -149
rect 6118 -183 6152 -149
rect 6218 -183 6252 -149
rect 6318 -183 6352 -149
rect 8162 -142 8196 -108
rect 8230 -142 8264 -108
rect 9278 -142 9312 -108
rect 9346 -142 9380 -108
rect 8162 -242 8196 -208
rect 8230 -242 8264 -208
rect 9278 -242 9312 -208
rect 9346 -242 9380 -208
rect 8162 -342 8196 -308
rect 8230 -342 8264 -308
rect 9278 -342 9312 -308
rect 9346 -342 9380 -308
rect 8162 -442 8196 -408
rect 8230 -442 8264 -408
rect 9278 -442 9312 -408
rect 9346 -442 9380 -408
rect 8162 -542 8196 -508
rect 8230 -542 8264 -508
rect 9278 -542 9312 -508
rect 9346 -542 9380 -508
rect 8162 -642 8196 -608
rect 8230 -642 8264 -608
rect 9278 -642 9312 -608
rect 9346 -642 9380 -608
rect 8162 -742 8196 -708
rect 8230 -742 8264 -708
rect 9278 -742 9312 -708
rect 9346 -742 9380 -708
rect 8162 -842 8196 -808
rect 8230 -842 8264 -808
rect -2 -892 32 -858
rect 66 -892 100 -858
rect 170 -892 204 -858
rect 238 -892 272 -858
rect 398 -892 432 -858
rect 466 -892 500 -858
rect 570 -892 604 -858
rect 638 -892 672 -858
rect 798 -892 832 -858
rect 866 -892 900 -858
rect -2 -992 32 -958
rect 66 -992 100 -958
rect 170 -992 204 -958
rect 238 -992 272 -958
rect 398 -992 432 -958
rect 466 -992 500 -958
rect 970 -892 1004 -858
rect 1038 -892 1072 -858
rect 1198 -892 1232 -858
rect 1266 -892 1300 -858
rect 1370 -892 1404 -858
rect 1438 -892 1472 -858
rect 1598 -892 1632 -858
rect 1666 -892 1700 -858
rect 570 -992 604 -958
rect 638 -992 672 -958
rect 798 -992 832 -958
rect 866 -992 900 -958
rect -2 -1092 32 -1058
rect 66 -1092 100 -1058
rect 170 -1092 204 -1058
rect 238 -1092 272 -1058
rect 398 -1092 432 -1058
rect 466 -1092 500 -1058
rect 970 -992 1004 -958
rect 1038 -992 1072 -958
rect 1198 -992 1232 -958
rect 1266 -992 1300 -958
rect 1770 -892 1804 -858
rect 1838 -892 1872 -858
rect 1998 -892 2032 -858
rect 2066 -892 2100 -858
rect 2170 -892 2204 -858
rect 2238 -892 2272 -858
rect 2398 -892 2432 -858
rect 2466 -892 2500 -858
rect 1370 -992 1404 -958
rect 1438 -992 1472 -958
rect 1598 -992 1632 -958
rect 1666 -992 1700 -958
rect 570 -1092 604 -1058
rect 638 -1092 672 -1058
rect 798 -1092 832 -1058
rect 866 -1092 900 -1058
rect -2 -1192 32 -1158
rect 66 -1192 100 -1158
rect 170 -1192 204 -1158
rect 238 -1192 272 -1158
rect 398 -1192 432 -1158
rect 466 -1192 500 -1158
rect 970 -1092 1004 -1058
rect 1038 -1092 1072 -1058
rect 1198 -1092 1232 -1058
rect 1266 -1092 1300 -1058
rect 1770 -992 1804 -958
rect 1838 -992 1872 -958
rect 1998 -992 2032 -958
rect 2066 -992 2100 -958
rect 2570 -892 2604 -858
rect 2638 -892 2672 -858
rect 2798 -892 2832 -858
rect 2866 -892 2900 -858
rect 2970 -892 3004 -858
rect 3038 -892 3072 -858
rect 3198 -892 3232 -858
rect 3266 -892 3300 -858
rect 2170 -992 2204 -958
rect 2238 -992 2272 -958
rect 2398 -992 2432 -958
rect 2466 -992 2500 -958
rect 1370 -1092 1404 -1058
rect 1438 -1092 1472 -1058
rect 1598 -1092 1632 -1058
rect 1666 -1092 1700 -1058
rect 570 -1192 604 -1158
rect 638 -1192 672 -1158
rect 798 -1192 832 -1158
rect 866 -1192 900 -1158
rect -2 -1292 32 -1258
rect 66 -1292 100 -1258
rect 170 -1292 204 -1258
rect 238 -1292 272 -1258
rect 398 -1292 432 -1258
rect 466 -1292 500 -1258
rect 970 -1192 1004 -1158
rect 1038 -1192 1072 -1158
rect 1198 -1192 1232 -1158
rect 1266 -1192 1300 -1158
rect 1770 -1092 1804 -1058
rect 1838 -1092 1872 -1058
rect 1998 -1092 2032 -1058
rect 2066 -1092 2100 -1058
rect 2570 -992 2604 -958
rect 2638 -992 2672 -958
rect 2798 -992 2832 -958
rect 2866 -992 2900 -958
rect 3370 -892 3404 -858
rect 3438 -892 3472 -858
rect 3598 -892 3632 -858
rect 3666 -892 3700 -858
rect 3770 -892 3804 -858
rect 3838 -892 3872 -858
rect 3998 -892 4032 -858
rect 4066 -892 4100 -858
rect 2970 -992 3004 -958
rect 3038 -992 3072 -958
rect 3198 -992 3232 -958
rect 3266 -992 3300 -958
rect 2170 -1092 2204 -1058
rect 2238 -1092 2272 -1058
rect 2398 -1092 2432 -1058
rect 2466 -1092 2500 -1058
rect 1370 -1192 1404 -1158
rect 1438 -1192 1472 -1158
rect 1598 -1192 1632 -1158
rect 1666 -1192 1700 -1158
rect 570 -1292 604 -1258
rect 638 -1292 672 -1258
rect 798 -1292 832 -1258
rect 866 -1292 900 -1258
rect -2 -1392 32 -1358
rect 66 -1392 100 -1358
rect 170 -1392 204 -1358
rect 238 -1392 272 -1358
rect 398 -1392 432 -1358
rect 466 -1392 500 -1358
rect 970 -1292 1004 -1258
rect 1038 -1292 1072 -1258
rect 1198 -1292 1232 -1258
rect 1266 -1292 1300 -1258
rect 1770 -1192 1804 -1158
rect 1838 -1192 1872 -1158
rect 1998 -1192 2032 -1158
rect 2066 -1192 2100 -1158
rect 2570 -1092 2604 -1058
rect 2638 -1092 2672 -1058
rect 2798 -1092 2832 -1058
rect 2866 -1092 2900 -1058
rect 3370 -992 3404 -958
rect 3438 -992 3472 -958
rect 3598 -992 3632 -958
rect 3666 -992 3700 -958
rect 4170 -892 4204 -858
rect 4238 -892 4272 -858
rect 4398 -892 4432 -858
rect 4466 -892 4500 -858
rect 4570 -892 4604 -858
rect 4638 -892 4672 -858
rect 4798 -892 4832 -858
rect 4866 -892 4900 -858
rect 3770 -992 3804 -958
rect 3838 -992 3872 -958
rect 3998 -992 4032 -958
rect 4066 -992 4100 -958
rect 2970 -1092 3004 -1058
rect 3038 -1092 3072 -1058
rect 3198 -1092 3232 -1058
rect 3266 -1092 3300 -1058
rect 2170 -1192 2204 -1158
rect 2238 -1192 2272 -1158
rect 2398 -1192 2432 -1158
rect 2466 -1192 2500 -1158
rect 1370 -1292 1404 -1258
rect 1438 -1292 1472 -1258
rect 1598 -1292 1632 -1258
rect 1666 -1292 1700 -1258
rect 570 -1392 604 -1358
rect 638 -1392 672 -1358
rect 798 -1392 832 -1358
rect 866 -1392 900 -1358
rect -2 -1492 32 -1458
rect 66 -1492 100 -1458
rect 170 -1492 204 -1458
rect 238 -1492 272 -1458
rect 398 -1492 432 -1458
rect 466 -1492 500 -1458
rect 970 -1392 1004 -1358
rect 1038 -1392 1072 -1358
rect 1198 -1392 1232 -1358
rect 1266 -1392 1300 -1358
rect 1770 -1292 1804 -1258
rect 1838 -1292 1872 -1258
rect 1998 -1292 2032 -1258
rect 2066 -1292 2100 -1258
rect 2570 -1192 2604 -1158
rect 2638 -1192 2672 -1158
rect 2798 -1192 2832 -1158
rect 2866 -1192 2900 -1158
rect 3370 -1092 3404 -1058
rect 3438 -1092 3472 -1058
rect 3598 -1092 3632 -1058
rect 3666 -1092 3700 -1058
rect 4170 -992 4204 -958
rect 4238 -992 4272 -958
rect 4398 -992 4432 -958
rect 4466 -992 4500 -958
rect 4970 -892 5004 -858
rect 5038 -892 5072 -858
rect 5198 -892 5232 -858
rect 5266 -892 5300 -858
rect 5370 -892 5404 -858
rect 5438 -892 5472 -858
rect 5598 -892 5632 -858
rect 5666 -892 5700 -858
rect 4570 -992 4604 -958
rect 4638 -992 4672 -958
rect 4798 -992 4832 -958
rect 4866 -992 4900 -958
rect 3770 -1092 3804 -1058
rect 3838 -1092 3872 -1058
rect 3998 -1092 4032 -1058
rect 4066 -1092 4100 -1058
rect 2970 -1192 3004 -1158
rect 3038 -1192 3072 -1158
rect 3198 -1192 3232 -1158
rect 3266 -1192 3300 -1158
rect 2170 -1292 2204 -1258
rect 2238 -1292 2272 -1258
rect 2398 -1292 2432 -1258
rect 2466 -1292 2500 -1258
rect 1370 -1392 1404 -1358
rect 1438 -1392 1472 -1358
rect 1598 -1392 1632 -1358
rect 1666 -1392 1700 -1358
rect 570 -1492 604 -1458
rect 638 -1492 672 -1458
rect 798 -1492 832 -1458
rect 866 -1492 900 -1458
rect -2 -1592 32 -1558
rect 66 -1592 100 -1558
rect 170 -1592 204 -1558
rect 238 -1592 272 -1558
rect 398 -1592 432 -1558
rect 466 -1592 500 -1558
rect 970 -1492 1004 -1458
rect 1038 -1492 1072 -1458
rect 1198 -1492 1232 -1458
rect 1266 -1492 1300 -1458
rect 1770 -1392 1804 -1358
rect 1838 -1392 1872 -1358
rect 1998 -1392 2032 -1358
rect 2066 -1392 2100 -1358
rect 2570 -1292 2604 -1258
rect 2638 -1292 2672 -1258
rect 2798 -1292 2832 -1258
rect 2866 -1292 2900 -1258
rect 3370 -1192 3404 -1158
rect 3438 -1192 3472 -1158
rect 3598 -1192 3632 -1158
rect 3666 -1192 3700 -1158
rect 4170 -1092 4204 -1058
rect 4238 -1092 4272 -1058
rect 4398 -1092 4432 -1058
rect 4466 -1092 4500 -1058
rect 4970 -992 5004 -958
rect 5038 -992 5072 -958
rect 5198 -992 5232 -958
rect 5266 -992 5300 -958
rect 5770 -892 5804 -858
rect 5838 -892 5872 -858
rect 5998 -892 6032 -858
rect 6066 -892 6100 -858
rect 6170 -892 6204 -858
rect 6238 -892 6272 -858
rect 9278 -842 9312 -808
rect 9346 -842 9380 -808
rect 5370 -992 5404 -958
rect 5438 -992 5472 -958
rect 5598 -992 5632 -958
rect 5666 -992 5700 -958
rect 4570 -1092 4604 -1058
rect 4638 -1092 4672 -1058
rect 4798 -1092 4832 -1058
rect 4866 -1092 4900 -1058
rect 3770 -1192 3804 -1158
rect 3838 -1192 3872 -1158
rect 3998 -1192 4032 -1158
rect 4066 -1192 4100 -1158
rect 2970 -1292 3004 -1258
rect 3038 -1292 3072 -1258
rect 3198 -1292 3232 -1258
rect 3266 -1292 3300 -1258
rect 2170 -1392 2204 -1358
rect 2238 -1392 2272 -1358
rect 2398 -1392 2432 -1358
rect 2466 -1392 2500 -1358
rect 1370 -1492 1404 -1458
rect 1438 -1492 1472 -1458
rect 1598 -1492 1632 -1458
rect 1666 -1492 1700 -1458
rect 570 -1592 604 -1558
rect 638 -1592 672 -1558
rect 798 -1592 832 -1558
rect 866 -1592 900 -1558
rect -2 -1692 32 -1658
rect 66 -1692 100 -1658
rect 170 -1692 204 -1658
rect 238 -1692 272 -1658
rect 398 -1692 432 -1658
rect 466 -1692 500 -1658
rect 970 -1592 1004 -1558
rect 1038 -1592 1072 -1558
rect 1198 -1592 1232 -1558
rect 1266 -1592 1300 -1558
rect 1770 -1492 1804 -1458
rect 1838 -1492 1872 -1458
rect 1998 -1492 2032 -1458
rect 2066 -1492 2100 -1458
rect 2570 -1392 2604 -1358
rect 2638 -1392 2672 -1358
rect 2798 -1392 2832 -1358
rect 2866 -1392 2900 -1358
rect 3370 -1292 3404 -1258
rect 3438 -1292 3472 -1258
rect 3598 -1292 3632 -1258
rect 3666 -1292 3700 -1258
rect 4170 -1192 4204 -1158
rect 4238 -1192 4272 -1158
rect 4398 -1192 4432 -1158
rect 4466 -1192 4500 -1158
rect 4970 -1092 5004 -1058
rect 5038 -1092 5072 -1058
rect 5198 -1092 5232 -1058
rect 5266 -1092 5300 -1058
rect 5770 -992 5804 -958
rect 5838 -992 5872 -958
rect 5998 -992 6032 -958
rect 6066 -992 6100 -958
rect 8162 -942 8196 -908
rect 8230 -942 8264 -908
rect 6170 -992 6204 -958
rect 6238 -992 6272 -958
rect 9278 -942 9312 -908
rect 9346 -942 9380 -908
rect 5370 -1092 5404 -1058
rect 5438 -1092 5472 -1058
rect 5598 -1092 5632 -1058
rect 5666 -1092 5700 -1058
rect 4570 -1192 4604 -1158
rect 4638 -1192 4672 -1158
rect 4798 -1192 4832 -1158
rect 4866 -1192 4900 -1158
rect 3770 -1292 3804 -1258
rect 3838 -1292 3872 -1258
rect 3998 -1292 4032 -1258
rect 4066 -1292 4100 -1258
rect 2970 -1392 3004 -1358
rect 3038 -1392 3072 -1358
rect 3198 -1392 3232 -1358
rect 3266 -1392 3300 -1358
rect 2170 -1492 2204 -1458
rect 2238 -1492 2272 -1458
rect 2398 -1492 2432 -1458
rect 2466 -1492 2500 -1458
rect 1370 -1592 1404 -1558
rect 1438 -1592 1472 -1558
rect 1598 -1592 1632 -1558
rect 1666 -1592 1700 -1558
rect 570 -1692 604 -1658
rect 638 -1692 672 -1658
rect 798 -1692 832 -1658
rect 866 -1692 900 -1658
rect -2 -1792 32 -1758
rect 66 -1792 100 -1758
rect 170 -1792 204 -1758
rect 238 -1792 272 -1758
rect 398 -1792 432 -1758
rect 466 -1792 500 -1758
rect 970 -1692 1004 -1658
rect 1038 -1692 1072 -1658
rect 1198 -1692 1232 -1658
rect 1266 -1692 1300 -1658
rect 1770 -1592 1804 -1558
rect 1838 -1592 1872 -1558
rect 1998 -1592 2032 -1558
rect 2066 -1592 2100 -1558
rect 2570 -1492 2604 -1458
rect 2638 -1492 2672 -1458
rect 2798 -1492 2832 -1458
rect 2866 -1492 2900 -1458
rect 3370 -1392 3404 -1358
rect 3438 -1392 3472 -1358
rect 3598 -1392 3632 -1358
rect 3666 -1392 3700 -1358
rect 4170 -1292 4204 -1258
rect 4238 -1292 4272 -1258
rect 4398 -1292 4432 -1258
rect 4466 -1292 4500 -1258
rect 4970 -1192 5004 -1158
rect 5038 -1192 5072 -1158
rect 5198 -1192 5232 -1158
rect 5266 -1192 5300 -1158
rect 5770 -1092 5804 -1058
rect 5838 -1092 5872 -1058
rect 5998 -1092 6032 -1058
rect 6066 -1092 6100 -1058
rect 8162 -1042 8196 -1008
rect 8230 -1042 8264 -1008
rect 6170 -1092 6204 -1058
rect 6238 -1092 6272 -1058
rect 9278 -1042 9312 -1008
rect 9346 -1042 9380 -1008
rect 5370 -1192 5404 -1158
rect 5438 -1192 5472 -1158
rect 5598 -1192 5632 -1158
rect 5666 -1192 5700 -1158
rect 4570 -1292 4604 -1258
rect 4638 -1292 4672 -1258
rect 4798 -1292 4832 -1258
rect 4866 -1292 4900 -1258
rect 3770 -1392 3804 -1358
rect 3838 -1392 3872 -1358
rect 3998 -1392 4032 -1358
rect 4066 -1392 4100 -1358
rect 2970 -1492 3004 -1458
rect 3038 -1492 3072 -1458
rect 3198 -1492 3232 -1458
rect 3266 -1492 3300 -1458
rect 2170 -1592 2204 -1558
rect 2238 -1592 2272 -1558
rect 2398 -1592 2432 -1558
rect 2466 -1592 2500 -1558
rect 1370 -1692 1404 -1658
rect 1438 -1692 1472 -1658
rect 1598 -1692 1632 -1658
rect 1666 -1692 1700 -1658
rect 570 -1792 604 -1758
rect 638 -1792 672 -1758
rect 798 -1792 832 -1758
rect 866 -1792 900 -1758
rect -2 -1892 32 -1858
rect 66 -1892 100 -1858
rect 170 -1892 204 -1858
rect 238 -1892 272 -1858
rect 398 -1892 432 -1858
rect 466 -1892 500 -1858
rect 970 -1792 1004 -1758
rect 1038 -1792 1072 -1758
rect 1198 -1792 1232 -1758
rect 1266 -1792 1300 -1758
rect 1770 -1692 1804 -1658
rect 1838 -1692 1872 -1658
rect 1998 -1692 2032 -1658
rect 2066 -1692 2100 -1658
rect 2570 -1592 2604 -1558
rect 2638 -1592 2672 -1558
rect 2798 -1592 2832 -1558
rect 2866 -1592 2900 -1558
rect 3370 -1492 3404 -1458
rect 3438 -1492 3472 -1458
rect 3598 -1492 3632 -1458
rect 3666 -1492 3700 -1458
rect 4170 -1392 4204 -1358
rect 4238 -1392 4272 -1358
rect 4398 -1392 4432 -1358
rect 4466 -1392 4500 -1358
rect 4970 -1292 5004 -1258
rect 5038 -1292 5072 -1258
rect 5198 -1292 5232 -1258
rect 5266 -1292 5300 -1258
rect 5770 -1192 5804 -1158
rect 5838 -1192 5872 -1158
rect 5998 -1192 6032 -1158
rect 6066 -1192 6100 -1158
rect 8162 -1142 8196 -1108
rect 8230 -1142 8264 -1108
rect 6170 -1192 6204 -1158
rect 6238 -1192 6272 -1158
rect 9278 -1142 9312 -1108
rect 9346 -1142 9380 -1108
rect 5370 -1292 5404 -1258
rect 5438 -1292 5472 -1258
rect 5598 -1292 5632 -1258
rect 5666 -1292 5700 -1258
rect 4570 -1392 4604 -1358
rect 4638 -1392 4672 -1358
rect 4798 -1392 4832 -1358
rect 4866 -1392 4900 -1358
rect 3770 -1492 3804 -1458
rect 3838 -1492 3872 -1458
rect 3998 -1492 4032 -1458
rect 4066 -1492 4100 -1458
rect 2970 -1592 3004 -1558
rect 3038 -1592 3072 -1558
rect 3198 -1592 3232 -1558
rect 3266 -1592 3300 -1558
rect 2170 -1692 2204 -1658
rect 2238 -1692 2272 -1658
rect 2398 -1692 2432 -1658
rect 2466 -1692 2500 -1658
rect 1370 -1792 1404 -1758
rect 1438 -1792 1472 -1758
rect 1598 -1792 1632 -1758
rect 1666 -1792 1700 -1758
rect 570 -1892 604 -1858
rect 638 -1892 672 -1858
rect 798 -1892 832 -1858
rect 866 -1892 900 -1858
rect 970 -1892 1004 -1858
rect 1038 -1892 1072 -1858
rect 1198 -1892 1232 -1858
rect 1266 -1892 1300 -1858
rect 1770 -1792 1804 -1758
rect 1838 -1792 1872 -1758
rect 1998 -1792 2032 -1758
rect 2066 -1792 2100 -1758
rect 2570 -1692 2604 -1658
rect 2638 -1692 2672 -1658
rect 2798 -1692 2832 -1658
rect 2866 -1692 2900 -1658
rect 3370 -1592 3404 -1558
rect 3438 -1592 3472 -1558
rect 3598 -1592 3632 -1558
rect 3666 -1592 3700 -1558
rect 4170 -1492 4204 -1458
rect 4238 -1492 4272 -1458
rect 4398 -1492 4432 -1458
rect 4466 -1492 4500 -1458
rect 4970 -1392 5004 -1358
rect 5038 -1392 5072 -1358
rect 5198 -1392 5232 -1358
rect 5266 -1392 5300 -1358
rect 5770 -1292 5804 -1258
rect 5838 -1292 5872 -1258
rect 5998 -1292 6032 -1258
rect 6066 -1292 6100 -1258
rect 8162 -1242 8196 -1208
rect 8230 -1242 8264 -1208
rect 6170 -1292 6204 -1258
rect 6238 -1292 6272 -1258
rect 9278 -1242 9312 -1208
rect 9346 -1242 9380 -1208
rect 5370 -1392 5404 -1358
rect 5438 -1392 5472 -1358
rect 5598 -1392 5632 -1358
rect 5666 -1392 5700 -1358
rect 4570 -1492 4604 -1458
rect 4638 -1492 4672 -1458
rect 4798 -1492 4832 -1458
rect 4866 -1492 4900 -1458
rect 3770 -1592 3804 -1558
rect 3838 -1592 3872 -1558
rect 3998 -1592 4032 -1558
rect 4066 -1592 4100 -1558
rect 2970 -1692 3004 -1658
rect 3038 -1692 3072 -1658
rect 3198 -1692 3232 -1658
rect 3266 -1692 3300 -1658
rect 2170 -1792 2204 -1758
rect 2238 -1792 2272 -1758
rect 2398 -1792 2432 -1758
rect 2466 -1792 2500 -1758
rect 1370 -1892 1404 -1858
rect 1438 -1892 1472 -1858
rect 1598 -1892 1632 -1858
rect 1666 -1892 1700 -1858
rect 1770 -1892 1804 -1858
rect 1838 -1892 1872 -1858
rect 1998 -1892 2032 -1858
rect 2066 -1892 2100 -1858
rect 2570 -1792 2604 -1758
rect 2638 -1792 2672 -1758
rect 2798 -1792 2832 -1758
rect 2866 -1792 2900 -1758
rect 3370 -1692 3404 -1658
rect 3438 -1692 3472 -1658
rect 3598 -1692 3632 -1658
rect 3666 -1692 3700 -1658
rect 4170 -1592 4204 -1558
rect 4238 -1592 4272 -1558
rect 4398 -1592 4432 -1558
rect 4466 -1592 4500 -1558
rect 4970 -1492 5004 -1458
rect 5038 -1492 5072 -1458
rect 5198 -1492 5232 -1458
rect 5266 -1492 5300 -1458
rect 5770 -1392 5804 -1358
rect 5838 -1392 5872 -1358
rect 5998 -1392 6032 -1358
rect 6066 -1392 6100 -1358
rect 8162 -1342 8196 -1308
rect 8230 -1342 8264 -1308
rect 6170 -1392 6204 -1358
rect 6238 -1392 6272 -1358
rect 9278 -1342 9312 -1308
rect 9346 -1342 9380 -1308
rect 5370 -1492 5404 -1458
rect 5438 -1492 5472 -1458
rect 5598 -1492 5632 -1458
rect 5666 -1492 5700 -1458
rect 4570 -1592 4604 -1558
rect 4638 -1592 4672 -1558
rect 4798 -1592 4832 -1558
rect 4866 -1592 4900 -1558
rect 3770 -1692 3804 -1658
rect 3838 -1692 3872 -1658
rect 3998 -1692 4032 -1658
rect 4066 -1692 4100 -1658
rect 2970 -1792 3004 -1758
rect 3038 -1792 3072 -1758
rect 3198 -1792 3232 -1758
rect 3266 -1792 3300 -1758
rect 2170 -1892 2204 -1858
rect 2238 -1892 2272 -1858
rect 2398 -1892 2432 -1858
rect 2466 -1892 2500 -1858
rect 2570 -1892 2604 -1858
rect 2638 -1892 2672 -1858
rect 2798 -1892 2832 -1858
rect 2866 -1892 2900 -1858
rect 3370 -1792 3404 -1758
rect 3438 -1792 3472 -1758
rect 3598 -1792 3632 -1758
rect 3666 -1792 3700 -1758
rect 4170 -1692 4204 -1658
rect 4238 -1692 4272 -1658
rect 4398 -1692 4432 -1658
rect 4466 -1692 4500 -1658
rect 4970 -1592 5004 -1558
rect 5038 -1592 5072 -1558
rect 5198 -1592 5232 -1558
rect 5266 -1592 5300 -1558
rect 5770 -1492 5804 -1458
rect 5838 -1492 5872 -1458
rect 5998 -1492 6032 -1458
rect 6066 -1492 6100 -1458
rect 8162 -1442 8196 -1408
rect 8230 -1442 8264 -1408
rect 6170 -1492 6204 -1458
rect 6238 -1492 6272 -1458
rect 9278 -1442 9312 -1408
rect 9346 -1442 9380 -1408
rect 5370 -1592 5404 -1558
rect 5438 -1592 5472 -1558
rect 5598 -1592 5632 -1558
rect 5666 -1592 5700 -1558
rect 4570 -1692 4604 -1658
rect 4638 -1692 4672 -1658
rect 4798 -1692 4832 -1658
rect 4866 -1692 4900 -1658
rect 3770 -1792 3804 -1758
rect 3838 -1792 3872 -1758
rect 3998 -1792 4032 -1758
rect 4066 -1792 4100 -1758
rect 2970 -1892 3004 -1858
rect 3038 -1892 3072 -1858
rect 3198 -1892 3232 -1858
rect 3266 -1892 3300 -1858
rect 3370 -1892 3404 -1858
rect 3438 -1892 3472 -1858
rect 3598 -1892 3632 -1858
rect 3666 -1892 3700 -1858
rect 4170 -1792 4204 -1758
rect 4238 -1792 4272 -1758
rect 4398 -1792 4432 -1758
rect 4466 -1792 4500 -1758
rect 4970 -1692 5004 -1658
rect 5038 -1692 5072 -1658
rect 5198 -1692 5232 -1658
rect 5266 -1692 5300 -1658
rect 5770 -1592 5804 -1558
rect 5838 -1592 5872 -1558
rect 5998 -1592 6032 -1558
rect 6066 -1592 6100 -1558
rect 8162 -1542 8196 -1508
rect 8230 -1542 8264 -1508
rect 6170 -1592 6204 -1558
rect 6238 -1592 6272 -1558
rect 9278 -1542 9312 -1508
rect 9346 -1542 9380 -1508
rect 5370 -1692 5404 -1658
rect 5438 -1692 5472 -1658
rect 5598 -1692 5632 -1658
rect 5666 -1692 5700 -1658
rect 4570 -1792 4604 -1758
rect 4638 -1792 4672 -1758
rect 4798 -1792 4832 -1758
rect 4866 -1792 4900 -1758
rect 3770 -1892 3804 -1858
rect 3838 -1892 3872 -1858
rect 3998 -1892 4032 -1858
rect 4066 -1892 4100 -1858
rect 4170 -1892 4204 -1858
rect 4238 -1892 4272 -1858
rect 4398 -1892 4432 -1858
rect 4466 -1892 4500 -1858
rect 4970 -1792 5004 -1758
rect 5038 -1792 5072 -1758
rect 5198 -1792 5232 -1758
rect 5266 -1792 5300 -1758
rect 5770 -1692 5804 -1658
rect 5838 -1692 5872 -1658
rect 5998 -1692 6032 -1658
rect 6066 -1692 6100 -1658
rect 8162 -1642 8196 -1608
rect 8230 -1642 8264 -1608
rect 6170 -1692 6204 -1658
rect 6238 -1692 6272 -1658
rect 9278 -1642 9312 -1608
rect 9346 -1642 9380 -1608
rect 5370 -1792 5404 -1758
rect 5438 -1792 5472 -1758
rect 5598 -1792 5632 -1758
rect 5666 -1792 5700 -1758
rect 4570 -1892 4604 -1858
rect 4638 -1892 4672 -1858
rect 4798 -1892 4832 -1858
rect 4866 -1892 4900 -1858
rect 4970 -1892 5004 -1858
rect 5038 -1892 5072 -1858
rect 5198 -1892 5232 -1858
rect 5266 -1892 5300 -1858
rect 5770 -1792 5804 -1758
rect 5838 -1792 5872 -1758
rect 5998 -1792 6032 -1758
rect 6066 -1792 6100 -1758
rect 8162 -1742 8196 -1708
rect 8230 -1742 8264 -1708
rect 6170 -1792 6204 -1758
rect 6238 -1792 6272 -1758
rect 9278 -1742 9312 -1708
rect 9346 -1742 9380 -1708
rect 5370 -1892 5404 -1858
rect 5438 -1892 5472 -1858
rect 5598 -1892 5632 -1858
rect 5666 -1892 5700 -1858
rect 5770 -1892 5804 -1858
rect 5838 -1892 5872 -1858
rect 5998 -1892 6032 -1858
rect 6066 -1892 6100 -1858
rect 8162 -1842 8196 -1808
rect 8230 -1842 8264 -1808
rect 6170 -1892 6204 -1858
rect 6238 -1892 6272 -1858
rect 9278 -1842 9312 -1808
rect 9346 -1842 9380 -1808
<< pdiffc >>
rect 8447 -42 8481 -8
rect 8515 -42 8549 -8
rect 8583 -42 8617 -8
rect 8651 -42 8685 -8
rect 8857 -42 8891 -8
rect 8925 -42 8959 -8
rect 8993 -42 9027 -8
rect 9061 -42 9095 -8
rect 8447 -142 8481 -108
rect 8515 -142 8549 -108
rect 8583 -142 8617 -108
rect 8651 -142 8685 -108
rect 8857 -142 8891 -108
rect 8925 -142 8959 -108
rect 8993 -142 9027 -108
rect 9061 -142 9095 -108
rect 8447 -242 8481 -208
rect 8515 -242 8549 -208
rect 8583 -242 8617 -208
rect 8651 -242 8685 -208
rect 8857 -242 8891 -208
rect 8925 -242 8959 -208
rect 8993 -242 9027 -208
rect 9061 -242 9095 -208
rect -82 -397 -48 -363
rect -82 -465 -48 -431
rect 18 -397 52 -363
rect 18 -465 52 -431
rect 118 -397 152 -363
rect 118 -465 152 -431
rect 218 -397 252 -363
rect 218 -465 252 -431
rect 318 -397 352 -363
rect 318 -465 352 -431
rect 418 -397 452 -363
rect 418 -465 452 -431
rect 518 -397 552 -363
rect 518 -465 552 -431
rect 618 -397 652 -363
rect 618 -465 652 -431
rect 718 -397 752 -363
rect 718 -465 752 -431
rect 818 -397 852 -363
rect 818 -465 852 -431
rect 918 -397 952 -363
rect 918 -465 952 -431
rect 1018 -397 1052 -363
rect 1018 -465 1052 -431
rect 1118 -397 1152 -363
rect 1118 -465 1152 -431
rect 1218 -397 1252 -363
rect 1218 -465 1252 -431
rect 1318 -397 1352 -363
rect 1318 -465 1352 -431
rect 1418 -397 1452 -363
rect 1418 -465 1452 -431
rect 1518 -397 1552 -363
rect 1518 -465 1552 -431
rect 1618 -397 1652 -363
rect 1618 -465 1652 -431
rect 1718 -397 1752 -363
rect 1718 -465 1752 -431
rect 1818 -397 1852 -363
rect 1818 -465 1852 -431
rect 1918 -397 1952 -363
rect 1918 -465 1952 -431
rect 2018 -397 2052 -363
rect 2018 -465 2052 -431
rect 2118 -397 2152 -363
rect 2118 -465 2152 -431
rect 2218 -397 2252 -363
rect 2218 -465 2252 -431
rect 2318 -397 2352 -363
rect 2318 -465 2352 -431
rect 2418 -397 2452 -363
rect 2418 -465 2452 -431
rect 2518 -397 2552 -363
rect 2518 -465 2552 -431
rect 2618 -397 2652 -363
rect 2618 -465 2652 -431
rect 2718 -397 2752 -363
rect 2718 -465 2752 -431
rect 2818 -397 2852 -363
rect 2818 -465 2852 -431
rect 2918 -397 2952 -363
rect 2918 -465 2952 -431
rect 3018 -397 3052 -363
rect 3018 -465 3052 -431
rect 3118 -397 3152 -363
rect 3118 -465 3152 -431
rect 3218 -397 3252 -363
rect 3218 -465 3252 -431
rect 3318 -397 3352 -363
rect 3318 -465 3352 -431
rect 3418 -397 3452 -363
rect 3418 -465 3452 -431
rect 3518 -397 3552 -363
rect 3518 -465 3552 -431
rect 3618 -397 3652 -363
rect 3618 -465 3652 -431
rect 3718 -397 3752 -363
rect 3718 -465 3752 -431
rect 3818 -397 3852 -363
rect 3818 -465 3852 -431
rect 3918 -397 3952 -363
rect 3918 -465 3952 -431
rect 4018 -397 4052 -363
rect 4018 -465 4052 -431
rect 4118 -397 4152 -363
rect 4118 -465 4152 -431
rect 4218 -397 4252 -363
rect 4218 -465 4252 -431
rect 4318 -397 4352 -363
rect 4318 -465 4352 -431
rect 4418 -397 4452 -363
rect 4418 -465 4452 -431
rect 4518 -397 4552 -363
rect 4518 -465 4552 -431
rect 4618 -397 4652 -363
rect 4618 -465 4652 -431
rect 4718 -397 4752 -363
rect 4718 -465 4752 -431
rect 4818 -397 4852 -363
rect 4818 -465 4852 -431
rect 4918 -397 4952 -363
rect 4918 -465 4952 -431
rect 5018 -397 5052 -363
rect 5018 -465 5052 -431
rect 5118 -397 5152 -363
rect 5118 -465 5152 -431
rect 5218 -397 5252 -363
rect 5218 -465 5252 -431
rect 5318 -397 5352 -363
rect 5318 -465 5352 -431
rect 5418 -397 5452 -363
rect 5418 -465 5452 -431
rect 5518 -397 5552 -363
rect 5518 -465 5552 -431
rect 5618 -397 5652 -363
rect 5618 -465 5652 -431
rect 5718 -397 5752 -363
rect 5718 -465 5752 -431
rect 5818 -397 5852 -363
rect 5818 -465 5852 -431
rect 5918 -397 5952 -363
rect 5918 -465 5952 -431
rect 6018 -397 6052 -363
rect 6018 -465 6052 -431
rect 6118 -397 6152 -363
rect 6118 -465 6152 -431
rect 6218 -397 6252 -363
rect 6218 -465 6252 -431
rect 8447 -342 8481 -308
rect 8515 -342 8549 -308
rect 8583 -342 8617 -308
rect 8651 -342 8685 -308
rect 8857 -342 8891 -308
rect 8925 -342 8959 -308
rect 8993 -342 9027 -308
rect 9061 -342 9095 -308
rect 6318 -397 6352 -363
rect 6318 -465 6352 -431
rect 8447 -442 8481 -408
rect 8515 -442 8549 -408
rect 8583 -442 8617 -408
rect 8651 -442 8685 -408
rect 8857 -442 8891 -408
rect 8925 -442 8959 -408
rect 8993 -442 9027 -408
rect 9061 -442 9095 -408
rect 8447 -542 8481 -508
rect 8515 -542 8549 -508
rect 8583 -542 8617 -508
rect 8651 -542 8685 -508
rect 8857 -542 8891 -508
rect 8925 -542 8959 -508
rect 8993 -542 9027 -508
rect 9061 -542 9095 -508
rect -30 -717 4 -683
rect 118 -717 152 -683
rect 266 -717 300 -683
rect 370 -717 404 -683
rect 518 -717 552 -683
rect 666 -717 700 -683
rect 770 -717 804 -683
rect 918 -717 952 -683
rect 1066 -717 1100 -683
rect 1170 -717 1204 -683
rect 1318 -717 1352 -683
rect 1466 -717 1500 -683
rect 1570 -717 1604 -683
rect 1718 -717 1752 -683
rect 1866 -717 1900 -683
rect 1970 -717 2004 -683
rect 2118 -717 2152 -683
rect 2266 -717 2300 -683
rect 2370 -717 2404 -683
rect 2518 -717 2552 -683
rect 2666 -717 2700 -683
rect 2770 -717 2804 -683
rect 2918 -717 2952 -683
rect 3066 -717 3100 -683
rect 3170 -717 3204 -683
rect 3318 -717 3352 -683
rect 3466 -717 3500 -683
rect 3570 -717 3604 -683
rect 3718 -717 3752 -683
rect 3866 -717 3900 -683
rect 3970 -717 4004 -683
rect 4118 -717 4152 -683
rect 4266 -717 4300 -683
rect 4370 -717 4404 -683
rect 4518 -717 4552 -683
rect 4666 -717 4700 -683
rect 4770 -717 4804 -683
rect 4918 -717 4952 -683
rect 5066 -717 5100 -683
rect 5170 -717 5204 -683
rect 5318 -717 5352 -683
rect 5466 -717 5500 -683
rect 5570 -717 5604 -683
rect 5718 -717 5752 -683
rect 5866 -717 5900 -683
rect 5970 -717 6004 -683
rect 6118 -717 6152 -683
rect 8447 -642 8481 -608
rect 8515 -642 8549 -608
rect 8583 -642 8617 -608
rect 8651 -642 8685 -608
rect 8857 -642 8891 -608
rect 8925 -642 8959 -608
rect 8993 -642 9027 -608
rect 9061 -642 9095 -608
rect 6266 -717 6300 -683
rect 8447 -742 8481 -708
rect 8515 -742 8549 -708
rect 8583 -742 8617 -708
rect 8651 -742 8685 -708
rect 8857 -742 8891 -708
rect 8925 -742 8959 -708
rect 8993 -742 9027 -708
rect 9061 -742 9095 -708
rect 8447 -842 8481 -808
rect 8515 -842 8549 -808
rect 8583 -842 8617 -808
rect 8651 -842 8685 -808
rect 8857 -842 8891 -808
rect 8925 -842 8959 -808
rect 8993 -842 9027 -808
rect 9061 -842 9095 -808
rect 8447 -942 8481 -908
rect 8515 -942 8549 -908
rect 8583 -942 8617 -908
rect 8651 -942 8685 -908
rect 8857 -942 8891 -908
rect 8925 -942 8959 -908
rect 8993 -942 9027 -908
rect 9061 -942 9095 -908
rect 8447 -1042 8481 -1008
rect 8515 -1042 8549 -1008
rect 8583 -1042 8617 -1008
rect 8651 -1042 8685 -1008
rect 8857 -1042 8891 -1008
rect 8925 -1042 8959 -1008
rect 8993 -1042 9027 -1008
rect 9061 -1042 9095 -1008
rect 8447 -1142 8481 -1108
rect 8515 -1142 8549 -1108
rect 8583 -1142 8617 -1108
rect 8651 -1142 8685 -1108
rect 8857 -1142 8891 -1108
rect 8925 -1142 8959 -1108
rect 8993 -1142 9027 -1108
rect 9061 -1142 9095 -1108
rect 8447 -1242 8481 -1208
rect 8515 -1242 8549 -1208
rect 8583 -1242 8617 -1208
rect 8651 -1242 8685 -1208
rect 8857 -1242 8891 -1208
rect 8925 -1242 8959 -1208
rect 8993 -1242 9027 -1208
rect 9061 -1242 9095 -1208
rect 8447 -1342 8481 -1308
rect 8515 -1342 8549 -1308
rect 8583 -1342 8617 -1308
rect 8651 -1342 8685 -1308
rect 8857 -1342 8891 -1308
rect 8925 -1342 8959 -1308
rect 8993 -1342 9027 -1308
rect 9061 -1342 9095 -1308
rect 8447 -1442 8481 -1408
rect 8515 -1442 8549 -1408
rect 8583 -1442 8617 -1408
rect 8651 -1442 8685 -1408
rect 8857 -1442 8891 -1408
rect 8925 -1442 8959 -1408
rect 8993 -1442 9027 -1408
rect 9061 -1442 9095 -1408
rect 8447 -1542 8481 -1508
rect 8515 -1542 8549 -1508
rect 8583 -1542 8617 -1508
rect 8651 -1542 8685 -1508
rect 8857 -1542 8891 -1508
rect 8925 -1542 8959 -1508
rect 8993 -1542 9027 -1508
rect 9061 -1542 9095 -1508
rect 8447 -1642 8481 -1608
rect 8515 -1642 8549 -1608
rect 8583 -1642 8617 -1608
rect 8651 -1642 8685 -1608
rect 8857 -1642 8891 -1608
rect 8925 -1642 8959 -1608
rect 8993 -1642 9027 -1608
rect 9061 -1642 9095 -1608
rect 8447 -1742 8481 -1708
rect 8515 -1742 8549 -1708
rect 8583 -1742 8617 -1708
rect 8651 -1742 8685 -1708
rect 8857 -1742 8891 -1708
rect 8925 -1742 8959 -1708
rect 8993 -1742 9027 -1708
rect 9061 -1742 9095 -1708
rect 8447 -1842 8481 -1808
rect 8515 -1842 8549 -1808
rect 8583 -1842 8617 -1808
rect 8651 -1842 8685 -1808
rect 8857 -1842 8891 -1808
rect 8925 -1842 8959 -1808
rect 8993 -1842 9027 -1808
rect 9061 -1842 9095 -1808
<< psubdiff >>
rect 116 9997 154 10021
rect 116 9963 118 9997
rect 152 9963 154 9997
rect 116 9939 154 9963
rect 316 9997 354 10021
rect 316 9963 318 9997
rect 352 9963 354 9997
rect 316 9939 354 9963
rect 516 9997 554 10021
rect 516 9963 518 9997
rect 552 9963 554 9997
rect 516 9939 554 9963
rect 716 9997 754 10021
rect 716 9963 718 9997
rect 752 9963 754 9997
rect 716 9939 754 9963
rect 916 9997 954 10021
rect 916 9963 918 9997
rect 952 9963 954 9997
rect 916 9939 954 9963
rect 1116 9997 1154 10021
rect 1116 9963 1118 9997
rect 1152 9963 1154 9997
rect 1116 9939 1154 9963
rect 1316 9997 1354 10021
rect 1316 9963 1318 9997
rect 1352 9963 1354 9997
rect 1316 9939 1354 9963
rect 1516 9997 1554 10021
rect 1516 9963 1518 9997
rect 1552 9963 1554 9997
rect 1516 9939 1554 9963
rect 1716 9997 1754 10021
rect 1716 9963 1718 9997
rect 1752 9963 1754 9997
rect 1716 9939 1754 9963
rect 1916 9997 1954 10021
rect 1916 9963 1918 9997
rect 1952 9963 1954 9997
rect 1916 9939 1954 9963
rect 2116 9997 2154 10021
rect 2116 9963 2118 9997
rect 2152 9963 2154 9997
rect 2116 9939 2154 9963
rect 2316 9997 2354 10021
rect 2316 9963 2318 9997
rect 2352 9963 2354 9997
rect 2316 9939 2354 9963
rect 2516 9997 2554 10021
rect 2516 9963 2518 9997
rect 2552 9963 2554 9997
rect 2516 9939 2554 9963
rect 2716 9997 2754 10021
rect 2716 9963 2718 9997
rect 2752 9963 2754 9997
rect 2716 9939 2754 9963
rect 2916 9997 2954 10021
rect 2916 9963 2918 9997
rect 2952 9963 2954 9997
rect 2916 9939 2954 9963
rect 3116 9997 3154 10021
rect 3116 9963 3118 9997
rect 3152 9963 3154 9997
rect 3116 9939 3154 9963
rect 3316 9997 3354 10021
rect 3316 9963 3318 9997
rect 3352 9963 3354 9997
rect 3316 9939 3354 9963
rect 3516 9997 3554 10021
rect 3516 9963 3518 9997
rect 3552 9963 3554 9997
rect 3516 9939 3554 9963
rect 3716 9997 3754 10021
rect 3716 9963 3718 9997
rect 3752 9963 3754 9997
rect 3716 9939 3754 9963
rect 3916 9997 3954 10021
rect 3916 9963 3918 9997
rect 3952 9963 3954 9997
rect 3916 9939 3954 9963
rect 4116 9997 4154 10021
rect 4116 9963 4118 9997
rect 4152 9963 4154 9997
rect 4116 9939 4154 9963
rect 4316 9997 4354 10021
rect 4316 9963 4318 9997
rect 4352 9963 4354 9997
rect 4316 9939 4354 9963
rect 4516 9997 4554 10021
rect 4516 9963 4518 9997
rect 4552 9963 4554 9997
rect 4516 9939 4554 9963
rect 4716 9997 4754 10021
rect 4716 9963 4718 9997
rect 4752 9963 4754 9997
rect 4716 9939 4754 9963
rect 4916 9997 4954 10021
rect 4916 9963 4918 9997
rect 4952 9963 4954 9997
rect 4916 9939 4954 9963
rect 5116 9997 5154 10021
rect 5116 9963 5118 9997
rect 5152 9963 5154 9997
rect 5116 9939 5154 9963
rect 5316 9997 5354 10021
rect 5316 9963 5318 9997
rect 5352 9963 5354 9997
rect 5316 9939 5354 9963
rect 5516 9997 5554 10021
rect 5516 9963 5518 9997
rect 5552 9963 5554 9997
rect 5516 9939 5554 9963
rect 5716 9997 5754 10021
rect 5716 9963 5718 9997
rect 5752 9963 5754 9997
rect 5716 9939 5754 9963
rect 5916 9997 5954 10021
rect 5916 9963 5918 9997
rect 5952 9963 5954 9997
rect 5916 9939 5954 9963
rect 6116 9997 6154 10021
rect 6116 9963 6118 9997
rect 6152 9963 6154 9997
rect 6116 9939 6154 9963
rect 6316 9997 6354 10021
rect 6316 9963 6318 9997
rect 6352 9963 6354 9997
rect 6316 9939 6354 9963
rect 116 5017 154 5041
rect 116 4983 118 5017
rect 152 4983 154 5017
rect 116 4959 154 4983
rect 316 5017 354 5041
rect 316 4983 318 5017
rect 352 4983 354 5017
rect 316 4959 354 4983
rect 516 5017 554 5041
rect 516 4983 518 5017
rect 552 4983 554 5017
rect 516 4959 554 4983
rect 716 5017 754 5041
rect 716 4983 718 5017
rect 752 4983 754 5017
rect 716 4959 754 4983
rect 916 5017 954 5041
rect 916 4983 918 5017
rect 952 4983 954 5017
rect 916 4959 954 4983
rect 1116 5017 1154 5041
rect 1116 4983 1118 5017
rect 1152 4983 1154 5017
rect 1116 4959 1154 4983
rect 1316 5017 1354 5041
rect 1316 4983 1318 5017
rect 1352 4983 1354 5017
rect 1316 4959 1354 4983
rect 1516 5017 1554 5041
rect 1516 4983 1518 5017
rect 1552 4983 1554 5017
rect 1516 4959 1554 4983
rect 1716 5017 1754 5041
rect 1716 4983 1718 5017
rect 1752 4983 1754 5017
rect 1716 4959 1754 4983
rect 1916 5017 1954 5041
rect 1916 4983 1918 5017
rect 1952 4983 1954 5017
rect 1916 4959 1954 4983
rect 2116 5017 2154 5041
rect 2116 4983 2118 5017
rect 2152 4983 2154 5017
rect 2116 4959 2154 4983
rect 2316 5017 2354 5041
rect 2316 4983 2318 5017
rect 2352 4983 2354 5017
rect 2316 4959 2354 4983
rect 2516 5017 2554 5041
rect 2516 4983 2518 5017
rect 2552 4983 2554 5017
rect 2516 4959 2554 4983
rect 2716 5017 2754 5041
rect 2716 4983 2718 5017
rect 2752 4983 2754 5017
rect 2716 4959 2754 4983
rect 2916 5017 2954 5041
rect 2916 4983 2918 5017
rect 2952 4983 2954 5017
rect 2916 4959 2954 4983
rect 3116 5017 3154 5041
rect 3116 4983 3118 5017
rect 3152 4983 3154 5017
rect 3116 4959 3154 4983
rect 3316 5017 3354 5041
rect 3316 4983 3318 5017
rect 3352 4983 3354 5017
rect 3316 4959 3354 4983
rect 3516 5017 3554 5041
rect 3516 4983 3518 5017
rect 3552 4983 3554 5017
rect 3516 4959 3554 4983
rect 3716 5017 3754 5041
rect 3716 4983 3718 5017
rect 3752 4983 3754 5017
rect 3716 4959 3754 4983
rect 3916 5017 3954 5041
rect 3916 4983 3918 5017
rect 3952 4983 3954 5017
rect 3916 4959 3954 4983
rect 4116 5017 4154 5041
rect 4116 4983 4118 5017
rect 4152 4983 4154 5017
rect 4116 4959 4154 4983
rect 4316 5017 4354 5041
rect 4316 4983 4318 5017
rect 4352 4983 4354 5017
rect 4316 4959 4354 4983
rect 4516 5017 4554 5041
rect 4516 4983 4518 5017
rect 4552 4983 4554 5017
rect 4516 4959 4554 4983
rect 4716 5017 4754 5041
rect 4716 4983 4718 5017
rect 4752 4983 4754 5017
rect 4716 4959 4754 4983
rect 4916 5017 4954 5041
rect 4916 4983 4918 5017
rect 4952 4983 4954 5017
rect 4916 4959 4954 4983
rect 5116 5017 5154 5041
rect 5116 4983 5118 5017
rect 5152 4983 5154 5017
rect 5116 4959 5154 4983
rect 5316 5017 5354 5041
rect 5316 4983 5318 5017
rect 5352 4983 5354 5017
rect 5316 4959 5354 4983
rect 5516 5017 5554 5041
rect 5516 4983 5518 5017
rect 5552 4983 5554 5017
rect 5516 4959 5554 4983
rect 5716 5017 5754 5041
rect 5716 4983 5718 5017
rect 5752 4983 5754 5017
rect 5716 4959 5754 4983
rect 5916 5017 5954 5041
rect 5916 4983 5918 5017
rect 5952 4983 5954 5017
rect 5916 4959 5954 4983
rect 6116 5017 6154 5041
rect 6116 4983 6118 5017
rect 6152 4983 6154 5017
rect 6116 4959 6154 4983
rect 6316 5017 6354 5041
rect 6316 4983 6318 5017
rect 6352 4983 6354 5017
rect 6316 4959 6354 4983
rect 8140 85 8290 87
rect 8140 51 8164 85
rect 8198 51 8232 85
rect 8266 51 8290 85
rect 8140 29 8290 51
rect -140 -61 -116 -27
rect -82 -61 -48 -27
rect -14 -61 84 -27
rect 118 -61 152 -27
rect 186 -61 284 -27
rect 318 -61 352 -27
rect 386 -61 484 -27
rect 518 -61 552 -27
rect 586 -61 684 -27
rect 718 -61 752 -27
rect 786 -61 884 -27
rect 918 -61 952 -27
rect 986 -61 1084 -27
rect 1118 -61 1152 -27
rect 1186 -61 1284 -27
rect 1318 -61 1352 -27
rect 1386 -61 1484 -27
rect 1518 -61 1552 -27
rect 1586 -61 1684 -27
rect 1718 -61 1752 -27
rect 1786 -61 1884 -27
rect 1918 -61 1952 -27
rect 1986 -61 2084 -27
rect 2118 -61 2152 -27
rect 2186 -61 2284 -27
rect 2318 -61 2352 -27
rect 2386 -61 2484 -27
rect 2518 -61 2552 -27
rect 2586 -61 2684 -27
rect 2718 -61 2752 -27
rect 2786 -61 2884 -27
rect 2918 -61 2952 -27
rect 2986 -61 3084 -27
rect 3118 -61 3152 -27
rect 3186 -61 3284 -27
rect 3318 -61 3352 -27
rect 3386 -61 3484 -27
rect 3518 -61 3552 -27
rect 3586 -61 3684 -27
rect 3718 -61 3752 -27
rect 3786 -61 3884 -27
rect 3918 -61 3952 -27
rect 3986 -61 4084 -27
rect 4118 -61 4152 -27
rect 4186 -61 4284 -27
rect 4318 -61 4352 -27
rect 4386 -61 4484 -27
rect 4518 -61 4552 -27
rect 4586 -61 4684 -27
rect 4718 -61 4752 -27
rect 4786 -61 4884 -27
rect 4918 -61 4952 -27
rect 4986 -61 5084 -27
rect 5118 -61 5152 -27
rect 5186 -61 5284 -27
rect 5318 -61 5352 -27
rect 5386 -61 5484 -27
rect 5518 -61 5552 -27
rect 5586 -61 5684 -27
rect 5718 -61 5752 -27
rect 5786 -61 5884 -27
rect 5918 -61 5952 -27
rect 5986 -61 6084 -27
rect 6118 -61 6152 -27
rect 6186 -61 6284 -27
rect 6318 -61 6352 -27
rect 6386 -61 6410 -27
rect 9252 85 9402 87
rect 9252 51 9276 85
rect 9310 51 9344 85
rect 9378 51 9402 85
rect 9252 29 9402 51
rect -10 -1951 108 -1929
rect -10 -1985 32 -1951
rect 66 -1985 108 -1951
rect -10 -1987 108 -1985
rect 162 -1951 280 -1929
rect 162 -1985 204 -1951
rect 238 -1985 280 -1951
rect 162 -1987 280 -1985
rect 390 -1951 508 -1929
rect 390 -1985 432 -1951
rect 466 -1985 508 -1951
rect 390 -1987 508 -1985
rect 562 -1951 680 -1929
rect 562 -1985 604 -1951
rect 638 -1985 680 -1951
rect 562 -1987 680 -1985
rect 790 -1951 908 -1929
rect 790 -1985 832 -1951
rect 866 -1985 908 -1951
rect 790 -1987 908 -1985
rect 962 -1951 1080 -1929
rect 962 -1985 1004 -1951
rect 1038 -1985 1080 -1951
rect 962 -1987 1080 -1985
rect 1190 -1951 1308 -1929
rect 1190 -1985 1232 -1951
rect 1266 -1985 1308 -1951
rect 1190 -1987 1308 -1985
rect 1362 -1951 1480 -1929
rect 1362 -1985 1404 -1951
rect 1438 -1985 1480 -1951
rect 1362 -1987 1480 -1985
rect 1590 -1951 1708 -1929
rect 1590 -1985 1632 -1951
rect 1666 -1985 1708 -1951
rect 1590 -1987 1708 -1985
rect 1762 -1951 1880 -1929
rect 1762 -1985 1804 -1951
rect 1838 -1985 1880 -1951
rect 1762 -1987 1880 -1985
rect 1990 -1951 2108 -1929
rect 1990 -1985 2032 -1951
rect 2066 -1985 2108 -1951
rect 1990 -1987 2108 -1985
rect 2162 -1951 2280 -1929
rect 2162 -1985 2204 -1951
rect 2238 -1985 2280 -1951
rect 2162 -1987 2280 -1985
rect 2390 -1951 2508 -1929
rect 2390 -1985 2432 -1951
rect 2466 -1985 2508 -1951
rect 2390 -1987 2508 -1985
rect 2562 -1951 2680 -1929
rect 2562 -1985 2604 -1951
rect 2638 -1985 2680 -1951
rect 2562 -1987 2680 -1985
rect 2790 -1951 2908 -1929
rect 2790 -1985 2832 -1951
rect 2866 -1985 2908 -1951
rect 2790 -1987 2908 -1985
rect 2962 -1951 3080 -1929
rect 2962 -1985 3004 -1951
rect 3038 -1985 3080 -1951
rect 2962 -1987 3080 -1985
rect 3190 -1951 3308 -1929
rect 3190 -1985 3232 -1951
rect 3266 -1985 3308 -1951
rect 3190 -1987 3308 -1985
rect 3362 -1951 3480 -1929
rect 3362 -1985 3404 -1951
rect 3438 -1985 3480 -1951
rect 3362 -1987 3480 -1985
rect 3590 -1951 3708 -1929
rect 3590 -1985 3632 -1951
rect 3666 -1985 3708 -1951
rect 3590 -1987 3708 -1985
rect 3762 -1951 3880 -1929
rect 3762 -1985 3804 -1951
rect 3838 -1985 3880 -1951
rect 3762 -1987 3880 -1985
rect 3990 -1951 4108 -1929
rect 3990 -1985 4032 -1951
rect 4066 -1985 4108 -1951
rect 3990 -1987 4108 -1985
rect 4162 -1951 4280 -1929
rect 4162 -1985 4204 -1951
rect 4238 -1985 4280 -1951
rect 4162 -1987 4280 -1985
rect 4390 -1951 4508 -1929
rect 4390 -1985 4432 -1951
rect 4466 -1985 4508 -1951
rect 4390 -1987 4508 -1985
rect 4562 -1951 4680 -1929
rect 4562 -1985 4604 -1951
rect 4638 -1985 4680 -1951
rect 4562 -1987 4680 -1985
rect 4790 -1951 4908 -1929
rect 4790 -1985 4832 -1951
rect 4866 -1985 4908 -1951
rect 4790 -1987 4908 -1985
rect 4962 -1951 5080 -1929
rect 4962 -1985 5004 -1951
rect 5038 -1985 5080 -1951
rect 4962 -1987 5080 -1985
rect 5190 -1951 5308 -1929
rect 5190 -1985 5232 -1951
rect 5266 -1985 5308 -1951
rect 5190 -1987 5308 -1985
rect 5362 -1951 5480 -1929
rect 5362 -1985 5404 -1951
rect 5438 -1985 5480 -1951
rect 5362 -1987 5480 -1985
rect 5590 -1951 5708 -1929
rect 5590 -1985 5632 -1951
rect 5666 -1985 5708 -1951
rect 5590 -1987 5708 -1985
rect 5762 -1951 5880 -1929
rect 5762 -1985 5804 -1951
rect 5838 -1985 5880 -1951
rect 5762 -1987 5880 -1985
rect 5990 -1951 6108 -1929
rect 5990 -1985 6032 -1951
rect 6066 -1985 6108 -1951
rect 5990 -1987 6108 -1985
rect 6162 -1951 6280 -1929
rect 8140 -1901 8290 -1879
rect 8140 -1935 8164 -1901
rect 8198 -1935 8232 -1901
rect 8266 -1935 8290 -1901
rect 8140 -1937 8290 -1935
rect 9252 -1901 9402 -1879
rect 9252 -1935 9276 -1901
rect 9310 -1935 9344 -1901
rect 9378 -1935 9402 -1901
rect 9252 -1937 9402 -1935
rect 6162 -1985 6204 -1951
rect 6238 -1985 6280 -1951
rect 6162 -1987 6280 -1985
<< nsubdiff >>
rect 8416 85 8716 87
rect 8416 51 8447 85
rect 8481 51 8515 85
rect 8549 51 8583 85
rect 8617 51 8651 85
rect 8685 51 8716 85
rect 8416 29 8716 51
rect 8826 85 9126 87
rect 8826 51 8857 85
rect 8891 51 8925 85
rect 8959 51 8993 85
rect 9027 51 9061 85
rect 9095 51 9126 85
rect 8826 29 9126 51
rect -133 -595 -82 -561
rect -48 -595 3 -561
rect 267 -595 318 -561
rect 352 -595 403 -561
rect 667 -595 718 -561
rect 752 -595 803 -561
rect 1067 -595 1118 -561
rect 1152 -595 1203 -561
rect 1467 -595 1518 -561
rect 1552 -595 1603 -561
rect 1867 -595 1918 -561
rect 1952 -595 2003 -561
rect 2267 -595 2318 -561
rect 2352 -595 2403 -561
rect 2667 -595 2718 -561
rect 2752 -595 2803 -561
rect 3067 -595 3118 -561
rect 3152 -595 3203 -561
rect 3467 -595 3518 -561
rect 3552 -595 3603 -561
rect 3867 -595 3918 -561
rect 3952 -595 4003 -561
rect 4267 -595 4318 -561
rect 4352 -595 4403 -561
rect 4667 -595 4718 -561
rect 4752 -595 4803 -561
rect 5067 -595 5118 -561
rect 5152 -595 5203 -561
rect 5467 -595 5518 -561
rect 5552 -595 5603 -561
rect 5867 -595 5918 -561
rect 5952 -595 6003 -561
rect 6267 -595 6318 -561
rect 6352 -595 6403 -561
rect 8416 -1901 8716 -1879
rect 8416 -1935 8447 -1901
rect 8481 -1935 8515 -1901
rect 8549 -1935 8583 -1901
rect 8617 -1935 8651 -1901
rect 8685 -1935 8716 -1901
rect 8416 -1937 8716 -1935
rect 8826 -1901 9126 -1879
rect 8826 -1935 8857 -1901
rect 8891 -1935 8925 -1901
rect 8959 -1935 8993 -1901
rect 9027 -1935 9061 -1901
rect 9095 -1935 9126 -1901
rect 8826 -1937 9126 -1935
<< psubdiffcont >>
rect 118 9963 152 9997
rect 318 9963 352 9997
rect 518 9963 552 9997
rect 718 9963 752 9997
rect 918 9963 952 9997
rect 1118 9963 1152 9997
rect 1318 9963 1352 9997
rect 1518 9963 1552 9997
rect 1718 9963 1752 9997
rect 1918 9963 1952 9997
rect 2118 9963 2152 9997
rect 2318 9963 2352 9997
rect 2518 9963 2552 9997
rect 2718 9963 2752 9997
rect 2918 9963 2952 9997
rect 3118 9963 3152 9997
rect 3318 9963 3352 9997
rect 3518 9963 3552 9997
rect 3718 9963 3752 9997
rect 3918 9963 3952 9997
rect 4118 9963 4152 9997
rect 4318 9963 4352 9997
rect 4518 9963 4552 9997
rect 4718 9963 4752 9997
rect 4918 9963 4952 9997
rect 5118 9963 5152 9997
rect 5318 9963 5352 9997
rect 5518 9963 5552 9997
rect 5718 9963 5752 9997
rect 5918 9963 5952 9997
rect 6118 9963 6152 9997
rect 6318 9963 6352 9997
rect 118 4983 152 5017
rect 318 4983 352 5017
rect 518 4983 552 5017
rect 718 4983 752 5017
rect 918 4983 952 5017
rect 1118 4983 1152 5017
rect 1318 4983 1352 5017
rect 1518 4983 1552 5017
rect 1718 4983 1752 5017
rect 1918 4983 1952 5017
rect 2118 4983 2152 5017
rect 2318 4983 2352 5017
rect 2518 4983 2552 5017
rect 2718 4983 2752 5017
rect 2918 4983 2952 5017
rect 3118 4983 3152 5017
rect 3318 4983 3352 5017
rect 3518 4983 3552 5017
rect 3718 4983 3752 5017
rect 3918 4983 3952 5017
rect 4118 4983 4152 5017
rect 4318 4983 4352 5017
rect 4518 4983 4552 5017
rect 4718 4983 4752 5017
rect 4918 4983 4952 5017
rect 5118 4983 5152 5017
rect 5318 4983 5352 5017
rect 5518 4983 5552 5017
rect 5718 4983 5752 5017
rect 5918 4983 5952 5017
rect 6118 4983 6152 5017
rect 6318 4983 6352 5017
rect 8164 51 8198 85
rect 8232 51 8266 85
rect -116 -61 -82 -27
rect -48 -61 -14 -27
rect 84 -61 118 -27
rect 152 -61 186 -27
rect 284 -61 318 -27
rect 352 -61 386 -27
rect 484 -61 518 -27
rect 552 -61 586 -27
rect 684 -61 718 -27
rect 752 -61 786 -27
rect 884 -61 918 -27
rect 952 -61 986 -27
rect 1084 -61 1118 -27
rect 1152 -61 1186 -27
rect 1284 -61 1318 -27
rect 1352 -61 1386 -27
rect 1484 -61 1518 -27
rect 1552 -61 1586 -27
rect 1684 -61 1718 -27
rect 1752 -61 1786 -27
rect 1884 -61 1918 -27
rect 1952 -61 1986 -27
rect 2084 -61 2118 -27
rect 2152 -61 2186 -27
rect 2284 -61 2318 -27
rect 2352 -61 2386 -27
rect 2484 -61 2518 -27
rect 2552 -61 2586 -27
rect 2684 -61 2718 -27
rect 2752 -61 2786 -27
rect 2884 -61 2918 -27
rect 2952 -61 2986 -27
rect 3084 -61 3118 -27
rect 3152 -61 3186 -27
rect 3284 -61 3318 -27
rect 3352 -61 3386 -27
rect 3484 -61 3518 -27
rect 3552 -61 3586 -27
rect 3684 -61 3718 -27
rect 3752 -61 3786 -27
rect 3884 -61 3918 -27
rect 3952 -61 3986 -27
rect 4084 -61 4118 -27
rect 4152 -61 4186 -27
rect 4284 -61 4318 -27
rect 4352 -61 4386 -27
rect 4484 -61 4518 -27
rect 4552 -61 4586 -27
rect 4684 -61 4718 -27
rect 4752 -61 4786 -27
rect 4884 -61 4918 -27
rect 4952 -61 4986 -27
rect 5084 -61 5118 -27
rect 5152 -61 5186 -27
rect 5284 -61 5318 -27
rect 5352 -61 5386 -27
rect 5484 -61 5518 -27
rect 5552 -61 5586 -27
rect 5684 -61 5718 -27
rect 5752 -61 5786 -27
rect 5884 -61 5918 -27
rect 5952 -61 5986 -27
rect 6084 -61 6118 -27
rect 6152 -61 6186 -27
rect 6284 -61 6318 -27
rect 6352 -61 6386 -27
rect 9276 51 9310 85
rect 9344 51 9378 85
rect 32 -1985 66 -1951
rect 204 -1985 238 -1951
rect 432 -1985 466 -1951
rect 604 -1985 638 -1951
rect 832 -1985 866 -1951
rect 1004 -1985 1038 -1951
rect 1232 -1985 1266 -1951
rect 1404 -1985 1438 -1951
rect 1632 -1985 1666 -1951
rect 1804 -1985 1838 -1951
rect 2032 -1985 2066 -1951
rect 2204 -1985 2238 -1951
rect 2432 -1985 2466 -1951
rect 2604 -1985 2638 -1951
rect 2832 -1985 2866 -1951
rect 3004 -1985 3038 -1951
rect 3232 -1985 3266 -1951
rect 3404 -1985 3438 -1951
rect 3632 -1985 3666 -1951
rect 3804 -1985 3838 -1951
rect 4032 -1985 4066 -1951
rect 4204 -1985 4238 -1951
rect 4432 -1985 4466 -1951
rect 4604 -1985 4638 -1951
rect 4832 -1985 4866 -1951
rect 5004 -1985 5038 -1951
rect 5232 -1985 5266 -1951
rect 5404 -1985 5438 -1951
rect 5632 -1985 5666 -1951
rect 5804 -1985 5838 -1951
rect 6032 -1985 6066 -1951
rect 8164 -1935 8198 -1901
rect 8232 -1935 8266 -1901
rect 9276 -1935 9310 -1901
rect 9344 -1935 9378 -1901
rect 6204 -1985 6238 -1951
<< nsubdiffcont >>
rect 8447 51 8481 85
rect 8515 51 8549 85
rect 8583 51 8617 85
rect 8651 51 8685 85
rect 8857 51 8891 85
rect 8925 51 8959 85
rect 8993 51 9027 85
rect 9061 51 9095 85
rect -82 -595 -48 -561
rect 318 -595 352 -561
rect 718 -595 752 -561
rect 1118 -595 1152 -561
rect 1518 -595 1552 -561
rect 1918 -595 1952 -561
rect 2318 -595 2352 -561
rect 2718 -595 2752 -561
rect 3118 -595 3152 -561
rect 3518 -595 3552 -561
rect 3918 -595 3952 -561
rect 4318 -595 4352 -561
rect 4718 -595 4752 -561
rect 5118 -595 5152 -561
rect 5518 -595 5552 -561
rect 5918 -595 5952 -561
rect 6318 -595 6352 -561
rect 8447 -1935 8481 -1901
rect 8515 -1935 8549 -1901
rect 8583 -1935 8617 -1901
rect 8651 -1935 8685 -1901
rect 8857 -1935 8891 -1901
rect 8925 -1935 8959 -1901
rect 8993 -1935 9027 -1901
rect 9061 -1935 9095 -1901
<< poly >>
rect 70 9884 100 10050
rect 170 9884 200 10050
rect 70 9874 200 9884
rect 70 9840 118 9874
rect 152 9840 200 9874
rect 70 9830 200 9840
rect 70 9793 100 9830
rect 170 9793 200 9830
rect 270 9900 300 10050
rect 370 9900 400 10050
rect 270 9890 400 9900
rect 270 9856 318 9890
rect 352 9856 400 9890
rect 270 9846 400 9856
rect 270 9793 300 9846
rect 370 9793 400 9846
rect 470 9884 500 10050
rect 570 9884 600 10050
rect 470 9874 600 9884
rect 470 9840 518 9874
rect 552 9840 600 9874
rect 470 9830 600 9840
rect 470 9793 500 9830
rect 570 9793 600 9830
rect 670 9900 700 10050
rect 770 9900 800 10050
rect 670 9890 800 9900
rect 670 9856 718 9890
rect 752 9856 800 9890
rect 670 9846 800 9856
rect 670 9793 700 9846
rect 770 9793 800 9846
rect 870 9884 900 10050
rect 970 9884 1000 10050
rect 870 9874 1000 9884
rect 870 9840 918 9874
rect 952 9840 1000 9874
rect 870 9830 1000 9840
rect 870 9793 900 9830
rect 970 9793 1000 9830
rect 1070 9900 1100 10050
rect 1170 9900 1200 10050
rect 1070 9890 1200 9900
rect 1070 9856 1118 9890
rect 1152 9856 1200 9890
rect 1070 9846 1200 9856
rect 1070 9793 1100 9846
rect 1170 9793 1200 9846
rect 1270 9884 1300 10050
rect 1370 9884 1400 10050
rect 1270 9874 1400 9884
rect 1270 9840 1318 9874
rect 1352 9840 1400 9874
rect 1270 9830 1400 9840
rect 1270 9793 1300 9830
rect 1370 9793 1400 9830
rect 1470 9900 1500 10050
rect 1570 9900 1600 10050
rect 1470 9890 1600 9900
rect 1470 9856 1518 9890
rect 1552 9856 1600 9890
rect 1470 9846 1600 9856
rect 1470 9793 1500 9846
rect 70 9653 100 9707
rect 170 9653 200 9707
rect 270 9653 300 9707
rect 370 9653 400 9707
rect 470 9653 500 9707
rect 570 9653 600 9707
rect 70 9513 100 9567
rect 170 9513 200 9567
rect 270 9513 300 9567
rect 370 9513 400 9567
rect 70 9373 100 9427
rect 170 9373 200 9427
rect 270 9373 300 9427
rect 370 9373 400 9427
rect 470 9373 500 9567
rect 570 9513 600 9567
rect 670 9513 700 9707
rect 770 9653 800 9707
rect 870 9653 900 9707
rect 970 9653 1000 9707
rect 1070 9653 1100 9707
rect 1170 9653 1200 9707
rect 1270 9653 1300 9707
rect 1370 9653 1400 9707
rect 1470 9653 1500 9707
rect 1570 9653 1600 9846
rect 1670 9884 1700 10050
rect 1770 9884 1800 10050
rect 1670 9874 1800 9884
rect 1670 9840 1718 9874
rect 1752 9840 1800 9874
rect 1670 9830 1800 9840
rect 1670 9793 1700 9830
rect 1770 9793 1800 9830
rect 1870 9900 1900 10050
rect 1970 9900 2000 10050
rect 1870 9890 2000 9900
rect 1870 9856 1918 9890
rect 1952 9856 2000 9890
rect 1870 9846 2000 9856
rect 1870 9793 1900 9846
rect 1970 9793 2000 9846
rect 2070 9884 2100 10050
rect 2170 9884 2200 10050
rect 2070 9874 2200 9884
rect 2070 9840 2118 9874
rect 2152 9840 2200 9874
rect 2070 9830 2200 9840
rect 2070 9793 2100 9830
rect 1670 9653 1700 9707
rect 1770 9653 1800 9707
rect 1870 9653 1900 9707
rect 1970 9653 2000 9707
rect 2070 9653 2100 9707
rect 770 9513 800 9567
rect 870 9513 900 9567
rect 570 9373 600 9427
rect 670 9373 700 9427
rect 770 9373 800 9427
rect 870 9373 900 9427
rect 970 9373 1000 9567
rect 1070 9513 1100 9567
rect 1070 9373 1100 9427
rect 1170 9373 1200 9567
rect 1270 9513 1300 9567
rect 1370 9513 1400 9567
rect 1470 9513 1500 9567
rect 1570 9513 1600 9567
rect 1670 9513 1700 9567
rect 1270 9373 1300 9427
rect 1370 9373 1400 9427
rect 1470 9373 1500 9427
rect 1570 9373 1600 9427
rect 1670 9373 1700 9427
rect 70 9233 100 9287
rect 170 9233 200 9287
rect 270 9233 300 9287
rect 370 9233 400 9287
rect 470 9233 500 9287
rect 570 9233 600 9287
rect 670 9233 700 9287
rect 770 9233 800 9287
rect 870 9233 900 9287
rect 970 9233 1000 9287
rect 1070 9233 1100 9287
rect 1170 9233 1200 9287
rect 1270 9233 1300 9287
rect 1370 9233 1400 9287
rect 1470 9233 1500 9287
rect 70 9093 100 9147
rect 170 9093 200 9147
rect 270 9093 300 9147
rect 370 9093 400 9147
rect 470 9093 500 9147
rect 570 9093 600 9147
rect 70 8953 100 9007
rect 170 8953 200 9007
rect 270 8953 300 9007
rect 370 8953 400 9007
rect 470 8953 500 9007
rect 570 8953 600 9007
rect 670 8953 700 9147
rect 770 9093 800 9147
rect 870 9093 900 9147
rect 970 9093 1000 9147
rect 1070 9093 1100 9147
rect 1170 9093 1200 9147
rect 1270 9093 1300 9147
rect 1370 9093 1400 9147
rect 1470 9093 1500 9147
rect 1570 9093 1600 9287
rect 1670 9233 1700 9287
rect 1770 9233 1800 9567
rect 1870 9513 1900 9567
rect 1970 9513 2000 9567
rect 1870 9373 1900 9427
rect 1970 9373 2000 9427
rect 2070 9373 2100 9567
rect 2170 9513 2200 9830
rect 2270 9900 2300 10050
rect 2370 9900 2400 10050
rect 2270 9890 2400 9900
rect 2270 9856 2318 9890
rect 2352 9856 2400 9890
rect 2270 9846 2400 9856
rect 2270 9793 2300 9846
rect 2370 9793 2400 9846
rect 2470 9884 2500 10050
rect 2570 9884 2600 10050
rect 2470 9874 2600 9884
rect 2470 9840 2518 9874
rect 2552 9840 2600 9874
rect 2470 9830 2600 9840
rect 2470 9793 2500 9830
rect 2570 9793 2600 9830
rect 2670 9900 2700 10050
rect 2770 9900 2800 10050
rect 2670 9890 2800 9900
rect 2670 9856 2718 9890
rect 2752 9856 2800 9890
rect 2670 9846 2800 9856
rect 2670 9793 2700 9846
rect 2270 9653 2300 9707
rect 2270 9513 2300 9567
rect 2170 9373 2200 9427
rect 2270 9373 2300 9427
rect 2370 9373 2400 9707
rect 2470 9653 2500 9707
rect 2570 9653 2600 9707
rect 2670 9653 2700 9707
rect 2770 9653 2800 9846
rect 2870 9884 2900 10050
rect 2970 9884 3000 10050
rect 2870 9874 3000 9884
rect 2870 9840 2918 9874
rect 2952 9840 3000 9874
rect 2870 9830 3000 9840
rect 2870 9793 2900 9830
rect 2970 9793 3000 9830
rect 3070 9900 3100 10050
rect 3170 9900 3200 10050
rect 3070 9890 3200 9900
rect 3070 9856 3118 9890
rect 3152 9856 3200 9890
rect 3070 9846 3200 9856
rect 3070 9793 3100 9846
rect 3170 9793 3200 9846
rect 3270 9884 3300 10050
rect 3370 9884 3400 10050
rect 3270 9874 3400 9884
rect 3270 9840 3318 9874
rect 3352 9840 3400 9874
rect 3270 9830 3400 9840
rect 2870 9653 2900 9707
rect 2470 9513 2500 9567
rect 2470 9373 2500 9427
rect 2570 9373 2600 9567
rect 2670 9513 2700 9567
rect 2670 9373 2700 9427
rect 2770 9373 2800 9567
rect 2870 9513 2900 9567
rect 2970 9513 3000 9707
rect 3070 9653 3100 9707
rect 3170 9653 3200 9707
rect 3270 9653 3300 9830
rect 3370 9793 3400 9830
rect 3470 9900 3500 10050
rect 3570 9900 3600 10050
rect 3470 9890 3600 9900
rect 3470 9856 3518 9890
rect 3552 9856 3600 9890
rect 3470 9846 3600 9856
rect 3470 9793 3500 9846
rect 3370 9653 3400 9707
rect 3470 9653 3500 9707
rect 3570 9653 3600 9846
rect 3670 9884 3700 10050
rect 3770 9884 3800 10050
rect 3670 9874 3800 9884
rect 3670 9840 3718 9874
rect 3752 9840 3800 9874
rect 3670 9830 3800 9840
rect 3670 9793 3700 9830
rect 3770 9793 3800 9830
rect 3870 9900 3900 10050
rect 3970 9900 4000 10050
rect 3870 9890 4000 9900
rect 3870 9856 3918 9890
rect 3952 9856 4000 9890
rect 3870 9846 4000 9856
rect 3870 9793 3900 9846
rect 3970 9793 4000 9846
rect 4070 9884 4100 10050
rect 4170 9884 4200 10050
rect 4070 9874 4200 9884
rect 4070 9840 4118 9874
rect 4152 9840 4200 9874
rect 4070 9830 4200 9840
rect 4070 9793 4100 9830
rect 4170 9793 4200 9830
rect 4270 9900 4300 10050
rect 4370 9900 4400 10050
rect 4270 9890 4400 9900
rect 4270 9856 4318 9890
rect 4352 9856 4400 9890
rect 4270 9846 4400 9856
rect 4270 9793 4300 9846
rect 4370 9793 4400 9846
rect 4470 9884 4500 10050
rect 4570 9884 4600 10050
rect 4470 9874 4600 9884
rect 4470 9840 4518 9874
rect 4552 9840 4600 9874
rect 4470 9830 4600 9840
rect 4470 9793 4500 9830
rect 4570 9793 4600 9830
rect 4670 9900 4700 10050
rect 4770 9900 4800 10050
rect 4670 9890 4800 9900
rect 4670 9856 4718 9890
rect 4752 9856 4800 9890
rect 4670 9846 4800 9856
rect 4670 9793 4700 9846
rect 4770 9793 4800 9846
rect 4870 9884 4900 10050
rect 4970 9884 5000 10050
rect 4870 9874 5000 9884
rect 4870 9840 4918 9874
rect 4952 9840 5000 9874
rect 4870 9830 5000 9840
rect 4870 9793 4900 9830
rect 4970 9793 5000 9830
rect 5070 9900 5100 10050
rect 5170 9900 5200 10050
rect 5070 9890 5200 9900
rect 5070 9856 5118 9890
rect 5152 9856 5200 9890
rect 5070 9846 5200 9856
rect 5070 9793 5100 9846
rect 5170 9793 5200 9846
rect 5270 9884 5300 10050
rect 5370 9884 5400 10050
rect 5270 9874 5400 9884
rect 5270 9840 5318 9874
rect 5352 9840 5400 9874
rect 5270 9830 5400 9840
rect 5270 9793 5300 9830
rect 5370 9793 5400 9830
rect 5470 9900 5500 10050
rect 5570 9900 5600 10050
rect 5470 9890 5600 9900
rect 5470 9856 5518 9890
rect 5552 9856 5600 9890
rect 5470 9846 5600 9856
rect 3670 9653 3700 9707
rect 3770 9653 3800 9707
rect 3870 9653 3900 9707
rect 3970 9653 4000 9707
rect 3070 9513 3100 9567
rect 3170 9513 3200 9567
rect 3270 9513 3300 9567
rect 3370 9513 3400 9567
rect 3470 9513 3500 9567
rect 3570 9513 3600 9567
rect 3670 9513 3700 9567
rect 3770 9513 3800 9567
rect 3870 9513 3900 9567
rect 3970 9513 4000 9567
rect 2870 9373 2900 9427
rect 2970 9373 3000 9427
rect 3070 9373 3100 9427
rect 3170 9373 3200 9427
rect 3270 9373 3300 9427
rect 3370 9373 3400 9427
rect 3470 9373 3500 9427
rect 3570 9373 3600 9427
rect 3670 9373 3700 9427
rect 3770 9373 3800 9427
rect 3870 9373 3900 9427
rect 3970 9373 4000 9427
rect 4070 9373 4100 9707
rect 4170 9653 4200 9707
rect 4270 9653 4300 9707
rect 4370 9653 4400 9707
rect 4470 9653 4500 9707
rect 4570 9653 4600 9707
rect 4670 9653 4700 9707
rect 4770 9653 4800 9707
rect 4870 9653 4900 9707
rect 4970 9653 5000 9707
rect 5070 9653 5100 9707
rect 5170 9653 5200 9707
rect 5270 9653 5300 9707
rect 5370 9653 5400 9707
rect 5470 9653 5500 9846
rect 5570 9793 5600 9846
rect 5670 9884 5700 10050
rect 5770 9884 5800 10050
rect 5670 9874 5800 9884
rect 5670 9840 5718 9874
rect 5752 9840 5800 9874
rect 5670 9830 5800 9840
rect 5670 9793 5700 9830
rect 5570 9653 5600 9707
rect 5670 9653 5700 9707
rect 5770 9653 5800 9830
rect 5870 9900 5900 10050
rect 5970 9900 6000 10050
rect 5870 9890 6000 9900
rect 5870 9856 5918 9890
rect 5952 9856 6000 9890
rect 5870 9846 6000 9856
rect 5870 9793 5900 9846
rect 5870 9653 5900 9707
rect 4170 9513 4200 9567
rect 4270 9513 4300 9567
rect 4370 9513 4400 9567
rect 4470 9513 4500 9567
rect 1870 9233 1900 9287
rect 1970 9233 2000 9287
rect 2070 9233 2100 9287
rect 2170 9233 2200 9287
rect 2270 9233 2300 9287
rect 2370 9233 2400 9287
rect 1670 9093 1700 9147
rect 770 8953 800 9007
rect 870 8953 900 9007
rect 970 8953 1000 9007
rect 1070 8953 1100 9007
rect 1170 8953 1200 9007
rect 1270 8953 1300 9007
rect 1370 8953 1400 9007
rect 1470 8953 1500 9007
rect 1570 8953 1600 9007
rect 1670 8953 1700 9007
rect 1770 8953 1800 9147
rect 1870 9093 1900 9147
rect 1870 8953 1900 9007
rect 1970 8953 2000 9147
rect 2070 9093 2100 9147
rect 2170 9093 2200 9147
rect 2270 9093 2300 9147
rect 2370 9093 2400 9147
rect 2470 9093 2500 9287
rect 2570 9233 2600 9287
rect 2670 9233 2700 9287
rect 2770 9233 2800 9287
rect 2870 9233 2900 9287
rect 2970 9233 3000 9287
rect 3070 9233 3100 9287
rect 3170 9233 3200 9287
rect 3270 9233 3300 9287
rect 3370 9233 3400 9287
rect 3470 9233 3500 9287
rect 3570 9233 3600 9287
rect 3670 9233 3700 9287
rect 3770 9233 3800 9287
rect 3870 9233 3900 9287
rect 3970 9233 4000 9287
rect 2570 9093 2600 9147
rect 2070 8953 2100 9007
rect 2170 8953 2200 9007
rect 2270 8953 2300 9007
rect 2370 8953 2400 9007
rect 2470 8953 2500 9007
rect 2570 8953 2600 9007
rect 70 8813 100 8867
rect 170 8813 200 8867
rect 70 8674 100 8727
rect 170 8674 200 8727
rect 70 8664 200 8674
rect 70 8630 118 8664
rect 152 8630 200 8664
rect 70 8620 200 8630
rect 70 8583 100 8620
rect 170 8583 200 8620
rect 270 8690 300 8867
rect 370 8813 400 8867
rect 470 8813 500 8867
rect 570 8813 600 8867
rect 670 8813 700 8867
rect 770 8813 800 8867
rect 870 8813 900 8867
rect 970 8813 1000 8867
rect 1070 8813 1100 8867
rect 1170 8813 1200 8867
rect 1270 8813 1300 8867
rect 1370 8813 1400 8867
rect 1470 8813 1500 8867
rect 1570 8813 1600 8867
rect 1670 8813 1700 8867
rect 1770 8813 1800 8867
rect 1870 8813 1900 8867
rect 1970 8813 2000 8867
rect 2070 8813 2100 8867
rect 2170 8813 2200 8867
rect 2270 8813 2300 8867
rect 2370 8813 2400 8867
rect 2470 8813 2500 8867
rect 2570 8813 2600 8867
rect 370 8690 400 8727
rect 270 8680 400 8690
rect 270 8646 318 8680
rect 352 8646 400 8680
rect 270 8636 400 8646
rect 270 8583 300 8636
rect 370 8583 400 8636
rect 470 8674 500 8727
rect 570 8674 600 8727
rect 470 8664 600 8674
rect 470 8630 518 8664
rect 552 8630 600 8664
rect 470 8620 600 8630
rect 470 8583 500 8620
rect 570 8583 600 8620
rect 670 8690 700 8727
rect 770 8690 800 8727
rect 670 8680 800 8690
rect 670 8646 718 8680
rect 752 8646 800 8680
rect 670 8636 800 8646
rect 670 8583 700 8636
rect 770 8583 800 8636
rect 870 8674 900 8727
rect 970 8674 1000 8727
rect 870 8664 1000 8674
rect 870 8630 918 8664
rect 952 8630 1000 8664
rect 870 8620 1000 8630
rect 70 8443 100 8497
rect 170 8443 200 8497
rect 270 8443 300 8497
rect 370 8443 400 8497
rect 470 8443 500 8497
rect 570 8443 600 8497
rect 670 8443 700 8497
rect 770 8443 800 8497
rect 870 8443 900 8620
rect 970 8583 1000 8620
rect 1070 8690 1100 8727
rect 1170 8690 1200 8727
rect 1070 8680 1200 8690
rect 1070 8646 1118 8680
rect 1152 8646 1200 8680
rect 1070 8636 1200 8646
rect 970 8443 1000 8497
rect 1070 8443 1100 8636
rect 1170 8583 1200 8636
rect 1270 8674 1300 8727
rect 1370 8674 1400 8727
rect 1270 8664 1400 8674
rect 1270 8630 1318 8664
rect 1352 8630 1400 8664
rect 1270 8620 1400 8630
rect 1270 8583 1300 8620
rect 1370 8583 1400 8620
rect 1470 8690 1500 8727
rect 1570 8690 1600 8727
rect 1470 8680 1600 8690
rect 1470 8646 1518 8680
rect 1552 8646 1600 8680
rect 1470 8636 1600 8646
rect 1470 8583 1500 8636
rect 1570 8583 1600 8636
rect 1670 8674 1700 8727
rect 1770 8674 1800 8727
rect 1670 8664 1800 8674
rect 1670 8630 1718 8664
rect 1752 8630 1800 8664
rect 1670 8620 1800 8630
rect 1670 8583 1700 8620
rect 1770 8583 1800 8620
rect 1870 8690 1900 8727
rect 1970 8690 2000 8727
rect 1870 8680 2000 8690
rect 1870 8646 1918 8680
rect 1952 8646 2000 8680
rect 1870 8636 2000 8646
rect 1870 8583 1900 8636
rect 1970 8583 2000 8636
rect 2070 8674 2100 8727
rect 2170 8674 2200 8727
rect 2070 8664 2200 8674
rect 2070 8630 2118 8664
rect 2152 8630 2200 8664
rect 2070 8620 2200 8630
rect 2070 8583 2100 8620
rect 2170 8583 2200 8620
rect 2270 8690 2300 8727
rect 2370 8690 2400 8727
rect 2270 8680 2400 8690
rect 2270 8646 2318 8680
rect 2352 8646 2400 8680
rect 2270 8636 2400 8646
rect 2270 8583 2300 8636
rect 2370 8583 2400 8636
rect 2470 8674 2500 8727
rect 2570 8674 2600 8727
rect 2470 8664 2600 8674
rect 2470 8630 2518 8664
rect 2552 8630 2600 8664
rect 2470 8620 2600 8630
rect 2470 8583 2500 8620
rect 2570 8583 2600 8620
rect 2670 8690 2700 9147
rect 2770 9093 2800 9147
rect 2770 8953 2800 9007
rect 2870 8953 2900 9147
rect 2970 9093 3000 9147
rect 3070 9093 3100 9147
rect 3170 9093 3200 9147
rect 2970 8953 3000 9007
rect 3070 8953 3100 9007
rect 3170 8953 3200 9007
rect 3270 8953 3300 9147
rect 3370 9093 3400 9147
rect 3470 9093 3500 9147
rect 3570 9093 3600 9147
rect 3670 9093 3700 9147
rect 3770 9093 3800 9147
rect 3870 9093 3900 9147
rect 3970 9093 4000 9147
rect 4070 9093 4100 9287
rect 4170 9233 4200 9427
rect 4270 9373 4300 9427
rect 4370 9373 4400 9427
rect 4470 9373 4500 9427
rect 4570 9373 4600 9567
rect 4670 9513 4700 9567
rect 4770 9513 4800 9567
rect 4670 9373 4700 9427
rect 4770 9373 4800 9427
rect 4870 9373 4900 9567
rect 4970 9513 5000 9567
rect 4970 9373 5000 9427
rect 5070 9373 5100 9567
rect 5170 9513 5200 9567
rect 5170 9373 5200 9427
rect 5270 9373 5300 9567
rect 5370 9513 5400 9567
rect 5470 9513 5500 9567
rect 5570 9513 5600 9567
rect 5370 9373 5400 9427
rect 5470 9373 5500 9427
rect 5570 9373 5600 9427
rect 5670 9373 5700 9567
rect 5770 9513 5800 9567
rect 5770 9373 5800 9427
rect 5870 9373 5900 9567
rect 5970 9513 6000 9846
rect 6070 9884 6100 10050
rect 6170 9884 6200 10050
rect 6070 9874 6200 9884
rect 6070 9840 6118 9874
rect 6152 9840 6200 9874
rect 6070 9830 6200 9840
rect 6070 9793 6100 9830
rect 6170 9793 6200 9830
rect 6270 9900 6300 10050
rect 6370 9900 6400 10050
rect 6570 9904 6600 10050
rect 6670 9904 6700 10050
rect 6880 9904 6910 10050
rect 6980 9904 7010 10050
rect 7080 9904 7110 10050
rect 7180 9904 7210 10050
rect 7280 9904 7310 10050
rect 7380 9904 7410 10050
rect 6270 9890 6400 9900
rect 6270 9856 6318 9890
rect 6352 9856 6400 9890
rect 6270 9846 6400 9856
rect 6270 9793 6300 9846
rect 6370 9793 6400 9846
rect 6558 9888 6612 9904
rect 6558 9854 6568 9888
rect 6602 9854 6612 9888
rect 6558 9838 6612 9854
rect 6658 9888 6712 9904
rect 6658 9854 6668 9888
rect 6702 9854 6712 9888
rect 6658 9838 6712 9854
rect 6868 9888 6922 9904
rect 6868 9854 6878 9888
rect 6912 9854 6922 9888
rect 6868 9838 6922 9854
rect 6968 9888 7022 9904
rect 6968 9854 6978 9888
rect 7012 9854 7022 9888
rect 6968 9838 7022 9854
rect 7068 9888 7122 9904
rect 7068 9854 7078 9888
rect 7112 9854 7122 9888
rect 7068 9838 7122 9854
rect 7168 9888 7222 9904
rect 7168 9854 7178 9888
rect 7212 9854 7222 9888
rect 7168 9838 7222 9854
rect 7268 9888 7322 9904
rect 7268 9854 7278 9888
rect 7312 9854 7322 9888
rect 7268 9838 7322 9854
rect 7368 9888 7422 9904
rect 7368 9854 7378 9888
rect 7412 9854 7422 9888
rect 7368 9838 7422 9854
rect 6570 9793 6600 9838
rect 6670 9793 6700 9838
rect 6880 9793 6910 9838
rect 6980 9793 7010 9838
rect 7080 9793 7110 9838
rect 7180 9793 7210 9838
rect 7280 9793 7310 9838
rect 7380 9793 7410 9838
rect 6070 9653 6100 9707
rect 6170 9653 6200 9707
rect 6270 9653 6300 9707
rect 6370 9653 6400 9707
rect 6570 9653 6600 9707
rect 6670 9653 6700 9707
rect 6880 9653 6910 9707
rect 6980 9653 7010 9707
rect 7080 9653 7110 9707
rect 7180 9653 7210 9707
rect 7280 9653 7310 9707
rect 7380 9653 7410 9707
rect 6070 9513 6100 9567
rect 5970 9373 6000 9427
rect 6070 9373 6100 9427
rect 6170 9373 6200 9567
rect 6270 9513 6300 9567
rect 6370 9513 6400 9567
rect 6570 9513 6600 9567
rect 6670 9513 6700 9567
rect 6880 9513 6910 9567
rect 6980 9513 7010 9567
rect 7080 9513 7110 9567
rect 7180 9513 7210 9567
rect 7280 9513 7310 9567
rect 7380 9513 7410 9567
rect 6270 9373 6300 9427
rect 6370 9373 6400 9427
rect 6570 9373 6600 9427
rect 6670 9373 6700 9427
rect 6880 9373 6910 9427
rect 6980 9373 7010 9427
rect 7080 9373 7110 9427
rect 7180 9373 7210 9427
rect 7280 9373 7310 9427
rect 7380 9373 7410 9427
rect 4270 9233 4300 9287
rect 4370 9233 4400 9287
rect 4470 9233 4500 9287
rect 4570 9233 4600 9287
rect 4670 9233 4700 9287
rect 4770 9233 4800 9287
rect 4870 9233 4900 9287
rect 4970 9233 5000 9287
rect 4170 9093 4200 9147
rect 4270 9093 4300 9147
rect 4370 9093 4400 9147
rect 4470 9093 4500 9147
rect 3370 8953 3400 9007
rect 3470 8953 3500 9007
rect 3570 8953 3600 9007
rect 3670 8953 3700 9007
rect 3770 8953 3800 9007
rect 3870 8953 3900 9007
rect 3970 8953 4000 9007
rect 4070 8953 4100 9007
rect 4170 8953 4200 9007
rect 4270 8953 4300 9007
rect 4370 8953 4400 9007
rect 2770 8813 2800 8867
rect 2870 8813 2900 8867
rect 2970 8813 3000 8867
rect 3070 8813 3100 8867
rect 2770 8690 2800 8727
rect 2670 8680 2800 8690
rect 2670 8646 2718 8680
rect 2752 8646 2800 8680
rect 2670 8636 2800 8646
rect 2670 8583 2700 8636
rect 1170 8443 1200 8497
rect 1270 8443 1300 8497
rect 70 8303 100 8357
rect 170 8303 200 8357
rect 270 8303 300 8357
rect 370 8303 400 8357
rect 470 8303 500 8357
rect 570 8303 600 8357
rect 70 8163 100 8217
rect 170 8163 200 8217
rect 270 8163 300 8217
rect 370 8163 400 8217
rect 470 8163 500 8217
rect 570 8163 600 8217
rect 670 8163 700 8357
rect 770 8303 800 8357
rect 770 8163 800 8217
rect 870 8163 900 8357
rect 970 8303 1000 8357
rect 1070 8303 1100 8357
rect 1170 8303 1200 8357
rect 1270 8303 1300 8357
rect 1370 8303 1400 8497
rect 1470 8443 1500 8497
rect 1570 8443 1600 8497
rect 1670 8443 1700 8497
rect 1770 8443 1800 8497
rect 1470 8303 1500 8357
rect 1570 8303 1600 8357
rect 1670 8303 1700 8357
rect 1770 8303 1800 8357
rect 1870 8303 1900 8497
rect 1970 8443 2000 8497
rect 970 8163 1000 8217
rect 1070 8163 1100 8217
rect 1170 8163 1200 8217
rect 70 8023 100 8077
rect 170 8023 200 8077
rect 70 7883 100 7937
rect 170 7883 200 7937
rect 270 7883 300 8077
rect 370 8023 400 8077
rect 470 8023 500 8077
rect 570 8023 600 8077
rect 670 8023 700 8077
rect 770 8023 800 8077
rect 870 8023 900 8077
rect 970 8023 1000 8077
rect 370 7883 400 7937
rect 470 7883 500 7937
rect 570 7883 600 7937
rect 70 7743 100 7797
rect 170 7743 200 7797
rect 270 7743 300 7797
rect 370 7743 400 7797
rect 470 7743 500 7797
rect 570 7743 600 7797
rect 670 7743 700 7937
rect 770 7883 800 7937
rect 770 7743 800 7797
rect 870 7743 900 7937
rect 970 7883 1000 7937
rect 1070 7883 1100 8077
rect 1170 8023 1200 8077
rect 1270 8023 1300 8217
rect 1370 8163 1400 8217
rect 1470 8163 1500 8217
rect 1570 8163 1600 8217
rect 1670 8163 1700 8217
rect 1770 8163 1800 8217
rect 1870 8163 1900 8217
rect 1970 8163 2000 8357
rect 2070 8303 2100 8497
rect 2170 8443 2200 8497
rect 2270 8443 2300 8497
rect 2170 8303 2200 8357
rect 2270 8303 2300 8357
rect 2070 8163 2100 8217
rect 2170 8163 2200 8217
rect 2270 8163 2300 8217
rect 2370 8163 2400 8497
rect 2470 8443 2500 8497
rect 2570 8443 2600 8497
rect 2670 8443 2700 8497
rect 2770 8443 2800 8636
rect 2870 8674 2900 8727
rect 2970 8674 3000 8727
rect 2870 8664 3000 8674
rect 2870 8630 2918 8664
rect 2952 8630 3000 8664
rect 2870 8620 3000 8630
rect 2870 8583 2900 8620
rect 2970 8583 3000 8620
rect 3070 8690 3100 8727
rect 3170 8690 3200 8867
rect 3270 8813 3300 8867
rect 3370 8813 3400 8867
rect 3470 8813 3500 8867
rect 3570 8813 3600 8867
rect 3670 8813 3700 8867
rect 3770 8813 3800 8867
rect 3870 8813 3900 8867
rect 3970 8813 4000 8867
rect 4070 8813 4100 8867
rect 4170 8813 4200 8867
rect 4270 8813 4300 8867
rect 4370 8813 4400 8867
rect 4470 8813 4500 9007
rect 4570 8953 4600 9147
rect 4670 9093 4700 9147
rect 4570 8813 4600 8867
rect 4670 8813 4700 9007
rect 4770 8953 4800 9147
rect 4870 9093 4900 9147
rect 4970 9093 5000 9147
rect 5070 9093 5100 9287
rect 5170 9233 5200 9287
rect 5270 9233 5300 9287
rect 5370 9233 5400 9287
rect 5170 9093 5200 9147
rect 4770 8813 4800 8867
rect 4870 8813 4900 9007
rect 4970 8953 5000 9007
rect 5070 8953 5100 9007
rect 5170 8953 5200 9007
rect 5270 8953 5300 9147
rect 5370 9093 5400 9147
rect 5470 9093 5500 9287
rect 5570 9233 5600 9287
rect 5670 9233 5700 9287
rect 5570 9093 5600 9147
rect 5670 9093 5700 9147
rect 5770 9093 5800 9287
rect 5870 9233 5900 9287
rect 5970 9233 6000 9287
rect 6070 9233 6100 9287
rect 6170 9233 6200 9287
rect 6270 9233 6300 9287
rect 6370 9233 6400 9287
rect 6570 9233 6600 9287
rect 6670 9233 6700 9287
rect 6880 9233 6910 9287
rect 6980 9233 7010 9287
rect 7080 9233 7110 9287
rect 7180 9233 7210 9287
rect 7280 9233 7310 9287
rect 7380 9233 7410 9287
rect 5870 9093 5900 9147
rect 5970 9093 6000 9147
rect 6070 9093 6100 9147
rect 6170 9093 6200 9147
rect 6270 9093 6300 9147
rect 6370 9093 6400 9147
rect 6570 9093 6600 9147
rect 6670 9093 6700 9147
rect 6880 9093 6910 9147
rect 6980 9093 7010 9147
rect 7080 9093 7110 9147
rect 7180 9093 7210 9147
rect 7280 9093 7310 9147
rect 7380 9093 7410 9147
rect 5370 8953 5400 9007
rect 5470 8953 5500 9007
rect 5570 8953 5600 9007
rect 4970 8813 5000 8867
rect 5070 8813 5100 8867
rect 5170 8813 5200 8867
rect 5270 8813 5300 8867
rect 5370 8813 5400 8867
rect 5470 8813 5500 8867
rect 3070 8680 3200 8690
rect 3070 8646 3118 8680
rect 3152 8646 3200 8680
rect 3070 8636 3200 8646
rect 3070 8583 3100 8636
rect 3170 8583 3200 8636
rect 3270 8674 3300 8727
rect 3370 8674 3400 8727
rect 3270 8664 3400 8674
rect 3270 8630 3318 8664
rect 3352 8630 3400 8664
rect 3270 8620 3400 8630
rect 3270 8583 3300 8620
rect 2870 8443 2900 8497
rect 2970 8443 3000 8497
rect 3070 8443 3100 8497
rect 3170 8443 3200 8497
rect 3270 8443 3300 8497
rect 3370 8443 3400 8620
rect 3470 8690 3500 8727
rect 3570 8690 3600 8727
rect 3470 8680 3600 8690
rect 3470 8646 3518 8680
rect 3552 8646 3600 8680
rect 3470 8636 3600 8646
rect 3470 8583 3500 8636
rect 3470 8443 3500 8497
rect 3570 8443 3600 8636
rect 3670 8674 3700 8727
rect 3770 8674 3800 8727
rect 3670 8664 3800 8674
rect 3670 8630 3718 8664
rect 3752 8630 3800 8664
rect 3670 8620 3800 8630
rect 3670 8583 3700 8620
rect 3770 8583 3800 8620
rect 3870 8690 3900 8727
rect 3970 8690 4000 8727
rect 3870 8680 4000 8690
rect 3870 8646 3918 8680
rect 3952 8646 4000 8680
rect 3870 8636 4000 8646
rect 3870 8583 3900 8636
rect 3970 8583 4000 8636
rect 4070 8674 4100 8727
rect 4170 8674 4200 8727
rect 4070 8664 4200 8674
rect 4070 8630 4118 8664
rect 4152 8630 4200 8664
rect 4070 8620 4200 8630
rect 3670 8443 3700 8497
rect 3770 8443 3800 8497
rect 2470 8303 2500 8357
rect 2470 8163 2500 8217
rect 2570 8163 2600 8357
rect 2670 8303 2700 8357
rect 2770 8303 2800 8357
rect 2870 8303 2900 8357
rect 2970 8303 3000 8357
rect 3070 8303 3100 8357
rect 1170 7883 1200 7937
rect 1270 7883 1300 7937
rect 1370 7883 1400 8077
rect 1470 8023 1500 8077
rect 1570 8023 1600 8077
rect 1670 8023 1700 8077
rect 970 7743 1000 7797
rect 1070 7743 1100 7797
rect 1170 7743 1200 7797
rect 1270 7743 1300 7797
rect 1370 7743 1400 7797
rect 1470 7743 1500 7937
rect 1570 7883 1600 7937
rect 70 7603 100 7657
rect 170 7603 200 7657
rect 270 7603 300 7657
rect 370 7603 400 7657
rect 470 7603 500 7657
rect 570 7603 600 7657
rect 670 7603 700 7657
rect 770 7603 800 7657
rect 870 7603 900 7657
rect 970 7603 1000 7657
rect 70 7464 100 7517
rect 170 7464 200 7517
rect 70 7454 200 7464
rect 70 7420 118 7454
rect 152 7420 200 7454
rect 70 7410 200 7420
rect 70 7373 100 7410
rect 170 7373 200 7410
rect 270 7480 300 7517
rect 370 7480 400 7517
rect 270 7470 400 7480
rect 270 7436 318 7470
rect 352 7436 400 7470
rect 270 7426 400 7436
rect 270 7373 300 7426
rect 370 7373 400 7426
rect 470 7464 500 7517
rect 570 7464 600 7517
rect 470 7454 600 7464
rect 470 7420 518 7454
rect 552 7420 600 7454
rect 470 7410 600 7420
rect 470 7373 500 7410
rect 570 7373 600 7410
rect 670 7480 700 7517
rect 770 7480 800 7517
rect 670 7470 800 7480
rect 670 7436 718 7470
rect 752 7436 800 7470
rect 670 7426 800 7436
rect 670 7373 700 7426
rect 770 7373 800 7426
rect 870 7464 900 7517
rect 970 7464 1000 7517
rect 870 7454 1000 7464
rect 870 7420 918 7454
rect 952 7420 1000 7454
rect 870 7410 1000 7420
rect 870 7373 900 7410
rect 970 7373 1000 7410
rect 1070 7480 1100 7657
rect 1170 7603 1200 7657
rect 1270 7603 1300 7657
rect 1170 7480 1200 7517
rect 1070 7470 1200 7480
rect 1070 7436 1118 7470
rect 1152 7436 1200 7470
rect 1070 7426 1200 7436
rect 1070 7373 1100 7426
rect 1170 7373 1200 7426
rect 1270 7464 1300 7517
rect 1370 7464 1400 7657
rect 1470 7603 1500 7657
rect 1570 7603 1600 7797
rect 1670 7743 1700 7937
rect 1770 7883 1800 8077
rect 1870 8023 1900 8077
rect 1970 8023 2000 8077
rect 1870 7883 1900 7937
rect 1970 7883 2000 7937
rect 2070 7883 2100 8077
rect 2170 8023 2200 8077
rect 2270 8023 2300 8077
rect 2370 8023 2400 8077
rect 2470 8023 2500 8077
rect 2570 8023 2600 8077
rect 2670 8023 2700 8217
rect 2770 8163 2800 8217
rect 2170 7883 2200 7937
rect 2270 7883 2300 7937
rect 2370 7883 2400 7937
rect 2470 7883 2500 7937
rect 1670 7603 1700 7657
rect 1770 7603 1800 7797
rect 1870 7743 1900 7797
rect 1970 7743 2000 7797
rect 2070 7743 2100 7797
rect 2170 7743 2200 7797
rect 2270 7743 2300 7797
rect 2370 7743 2400 7797
rect 2470 7743 2500 7797
rect 2570 7743 2600 7937
rect 2670 7883 2700 7937
rect 2770 7883 2800 8077
rect 2870 8023 2900 8217
rect 2970 8163 3000 8217
rect 3070 8163 3100 8217
rect 3170 8163 3200 8357
rect 3270 8303 3300 8357
rect 3370 8303 3400 8357
rect 3470 8303 3500 8357
rect 3270 8163 3300 8217
rect 3370 8163 3400 8217
rect 3470 8163 3500 8217
rect 3570 8163 3600 8357
rect 3670 8303 3700 8357
rect 3770 8303 3800 8357
rect 3870 8303 3900 8497
rect 3970 8443 4000 8497
rect 4070 8443 4100 8620
rect 4170 8583 4200 8620
rect 4270 8690 4300 8727
rect 4370 8690 4400 8727
rect 4270 8680 4400 8690
rect 4270 8646 4318 8680
rect 4352 8646 4400 8680
rect 4270 8636 4400 8646
rect 4270 8583 4300 8636
rect 4170 8443 4200 8497
rect 4270 8443 4300 8497
rect 4370 8443 4400 8636
rect 4470 8674 4500 8727
rect 4570 8674 4600 8727
rect 4470 8664 4600 8674
rect 4470 8630 4518 8664
rect 4552 8630 4600 8664
rect 4470 8620 4600 8630
rect 4470 8583 4500 8620
rect 4570 8583 4600 8620
rect 4670 8690 4700 8727
rect 4770 8690 4800 8727
rect 4670 8680 4800 8690
rect 4670 8646 4718 8680
rect 4752 8646 4800 8680
rect 4670 8636 4800 8646
rect 4670 8583 4700 8636
rect 4470 8443 4500 8497
rect 4570 8443 4600 8497
rect 4670 8443 4700 8497
rect 3970 8303 4000 8357
rect 4070 8303 4100 8357
rect 4170 8303 4200 8357
rect 4270 8303 4300 8357
rect 4370 8303 4400 8357
rect 4470 8303 4500 8357
rect 4570 8303 4600 8357
rect 4670 8303 4700 8357
rect 4770 8303 4800 8636
rect 4870 8674 4900 8727
rect 4970 8674 5000 8727
rect 4870 8664 5000 8674
rect 4870 8630 4918 8664
rect 4952 8630 5000 8664
rect 4870 8620 5000 8630
rect 4870 8583 4900 8620
rect 4970 8583 5000 8620
rect 5070 8690 5100 8727
rect 5170 8690 5200 8727
rect 5070 8680 5200 8690
rect 5070 8646 5118 8680
rect 5152 8646 5200 8680
rect 5070 8636 5200 8646
rect 5070 8583 5100 8636
rect 5170 8583 5200 8636
rect 5270 8674 5300 8727
rect 5370 8674 5400 8727
rect 5270 8664 5400 8674
rect 5270 8630 5318 8664
rect 5352 8630 5400 8664
rect 5270 8620 5400 8630
rect 5270 8583 5300 8620
rect 5370 8583 5400 8620
rect 5470 8690 5500 8727
rect 5570 8690 5600 8867
rect 5670 8813 5700 9007
rect 5770 8953 5800 9007
rect 5870 8953 5900 9007
rect 5970 8953 6000 9007
rect 6070 8953 6100 9007
rect 5770 8813 5800 8867
rect 5870 8813 5900 8867
rect 5470 8680 5600 8690
rect 5470 8646 5518 8680
rect 5552 8646 5600 8680
rect 5470 8636 5600 8646
rect 5470 8583 5500 8636
rect 5570 8583 5600 8636
rect 5670 8674 5700 8727
rect 5770 8674 5800 8727
rect 5670 8664 5800 8674
rect 5670 8630 5718 8664
rect 5752 8630 5800 8664
rect 5670 8620 5800 8630
rect 4870 8443 4900 8497
rect 4870 8303 4900 8357
rect 4970 8303 5000 8497
rect 5070 8443 5100 8497
rect 5170 8443 5200 8497
rect 5270 8443 5300 8497
rect 5370 8443 5400 8497
rect 5470 8443 5500 8497
rect 5570 8443 5600 8497
rect 5670 8443 5700 8620
rect 5770 8583 5800 8620
rect 5870 8690 5900 8727
rect 5970 8690 6000 8867
rect 6070 8813 6100 8867
rect 6170 8813 6200 9007
rect 6270 8953 6300 9007
rect 6370 8953 6400 9007
rect 6570 8953 6600 9007
rect 6670 8953 6700 9007
rect 6880 8953 6910 9007
rect 6980 8953 7010 9007
rect 7080 8953 7110 9007
rect 7180 8953 7210 9007
rect 7280 8953 7310 9007
rect 7380 8953 7410 9007
rect 6270 8813 6300 8867
rect 6370 8813 6400 8867
rect 6570 8813 6600 8867
rect 6670 8813 6700 8867
rect 6880 8813 6910 8867
rect 6980 8813 7010 8867
rect 7080 8813 7110 8867
rect 7180 8813 7210 8867
rect 7280 8813 7310 8867
rect 7380 8813 7410 8867
rect 5870 8680 6000 8690
rect 5870 8646 5918 8680
rect 5952 8646 6000 8680
rect 5870 8636 6000 8646
rect 5870 8583 5900 8636
rect 5970 8583 6000 8636
rect 6070 8674 6100 8727
rect 6170 8674 6200 8727
rect 6070 8664 6200 8674
rect 6070 8630 6118 8664
rect 6152 8630 6200 8664
rect 6070 8620 6200 8630
rect 6070 8583 6100 8620
rect 6170 8583 6200 8620
rect 6270 8690 6300 8727
rect 6370 8690 6400 8727
rect 6570 8694 6600 8727
rect 6670 8694 6700 8727
rect 6880 8694 6910 8727
rect 6980 8694 7010 8727
rect 7080 8694 7110 8727
rect 7180 8694 7210 8727
rect 7280 8694 7310 8727
rect 7380 8694 7410 8727
rect 6270 8680 6400 8690
rect 6270 8646 6318 8680
rect 6352 8646 6400 8680
rect 6270 8636 6400 8646
rect 6270 8583 6300 8636
rect 6370 8583 6400 8636
rect 6558 8678 6612 8694
rect 6558 8644 6568 8678
rect 6602 8644 6612 8678
rect 6558 8628 6612 8644
rect 6658 8678 6712 8694
rect 6658 8644 6668 8678
rect 6702 8644 6712 8678
rect 6658 8628 6712 8644
rect 6868 8678 6922 8694
rect 6868 8644 6878 8678
rect 6912 8644 6922 8678
rect 6868 8628 6922 8644
rect 6968 8678 7022 8694
rect 6968 8644 6978 8678
rect 7012 8644 7022 8678
rect 6968 8628 7022 8644
rect 7068 8678 7122 8694
rect 7068 8644 7078 8678
rect 7112 8644 7122 8678
rect 7068 8628 7122 8644
rect 7168 8678 7222 8694
rect 7168 8644 7178 8678
rect 7212 8644 7222 8678
rect 7168 8628 7222 8644
rect 7268 8678 7322 8694
rect 7268 8644 7278 8678
rect 7312 8644 7322 8678
rect 7268 8628 7322 8644
rect 7368 8678 7422 8694
rect 7368 8644 7378 8678
rect 7412 8644 7422 8678
rect 7368 8628 7422 8644
rect 6570 8583 6600 8628
rect 6670 8583 6700 8628
rect 6880 8583 6910 8628
rect 6980 8583 7010 8628
rect 7080 8583 7110 8628
rect 7180 8583 7210 8628
rect 7280 8583 7310 8628
rect 7380 8583 7410 8628
rect 5770 8443 5800 8497
rect 5070 8303 5100 8357
rect 5170 8303 5200 8357
rect 5270 8303 5300 8357
rect 5370 8303 5400 8357
rect 5470 8303 5500 8357
rect 5570 8303 5600 8357
rect 5670 8303 5700 8357
rect 5770 8303 5800 8357
rect 5870 8303 5900 8497
rect 5970 8443 6000 8497
rect 6070 8443 6100 8497
rect 6170 8443 6200 8497
rect 6270 8443 6300 8497
rect 6370 8443 6400 8497
rect 6570 8443 6600 8497
rect 6670 8443 6700 8497
rect 6880 8443 6910 8497
rect 6980 8443 7010 8497
rect 7080 8443 7110 8497
rect 7180 8443 7210 8497
rect 7280 8443 7310 8497
rect 7380 8443 7410 8497
rect 5970 8303 6000 8357
rect 6070 8303 6100 8357
rect 6170 8303 6200 8357
rect 6270 8303 6300 8357
rect 6370 8303 6400 8357
rect 6570 8303 6600 8357
rect 6670 8303 6700 8357
rect 6880 8303 6910 8357
rect 6980 8303 7010 8357
rect 7080 8303 7110 8357
rect 7180 8303 7210 8357
rect 7280 8303 7310 8357
rect 7380 8303 7410 8357
rect 3670 8163 3700 8217
rect 2870 7883 2900 7937
rect 2970 7883 3000 8077
rect 3070 8023 3100 8077
rect 3170 8023 3200 8077
rect 3270 8023 3300 8077
rect 3370 8023 3400 8077
rect 3470 8023 3500 8077
rect 3570 8023 3600 8077
rect 3670 8023 3700 8077
rect 3770 8023 3800 8217
rect 3870 8163 3900 8217
rect 3970 8163 4000 8217
rect 4070 8163 4100 8217
rect 4170 8163 4200 8217
rect 4270 8163 4300 8217
rect 4370 8163 4400 8217
rect 4470 8163 4500 8217
rect 4570 8163 4600 8217
rect 4670 8163 4700 8217
rect 4770 8163 4800 8217
rect 4870 8163 4900 8217
rect 4970 8163 5000 8217
rect 5070 8163 5100 8217
rect 5170 8163 5200 8217
rect 5270 8163 5300 8217
rect 5370 8163 5400 8217
rect 5470 8163 5500 8217
rect 5570 8163 5600 8217
rect 5670 8163 5700 8217
rect 5770 8163 5800 8217
rect 5870 8163 5900 8217
rect 5970 8163 6000 8217
rect 6070 8163 6100 8217
rect 6170 8163 6200 8217
rect 6270 8163 6300 8217
rect 6370 8163 6400 8217
rect 6570 8163 6600 8217
rect 6670 8163 6700 8217
rect 6880 8163 6910 8217
rect 6980 8163 7010 8217
rect 7080 8163 7110 8217
rect 7180 8163 7210 8217
rect 7280 8163 7310 8217
rect 7380 8163 7410 8217
rect 3870 8023 3900 8077
rect 3970 8023 4000 8077
rect 4070 8023 4100 8077
rect 4170 8023 4200 8077
rect 4270 8023 4300 8077
rect 4370 8023 4400 8077
rect 4470 8023 4500 8077
rect 4570 8023 4600 8077
rect 4670 8023 4700 8077
rect 4770 8023 4800 8077
rect 4870 8023 4900 8077
rect 3070 7883 3100 7937
rect 3170 7883 3200 7937
rect 3270 7883 3300 7937
rect 2670 7743 2700 7797
rect 1870 7603 1900 7657
rect 1970 7603 2000 7657
rect 2070 7603 2100 7657
rect 2170 7603 2200 7657
rect 2270 7603 2300 7657
rect 2370 7603 2400 7657
rect 2470 7603 2500 7657
rect 2570 7603 2600 7657
rect 2670 7603 2700 7657
rect 1270 7454 1400 7464
rect 1270 7420 1318 7454
rect 1352 7420 1400 7454
rect 1270 7410 1400 7420
rect 70 7233 100 7287
rect 170 7233 200 7287
rect 270 7233 300 7287
rect 70 7093 100 7147
rect 170 7093 200 7147
rect 270 7093 300 7147
rect 70 6953 100 7007
rect 170 6953 200 7007
rect 270 6953 300 7007
rect 370 6953 400 7287
rect 470 7233 500 7287
rect 570 7233 600 7287
rect 670 7233 700 7287
rect 770 7233 800 7287
rect 870 7233 900 7287
rect 970 7233 1000 7287
rect 1070 7233 1100 7287
rect 1170 7233 1200 7287
rect 1270 7233 1300 7410
rect 1370 7373 1400 7410
rect 1470 7480 1500 7517
rect 1570 7480 1600 7517
rect 1470 7470 1600 7480
rect 1470 7436 1518 7470
rect 1552 7436 1600 7470
rect 1470 7426 1600 7436
rect 1470 7373 1500 7426
rect 1370 7233 1400 7287
rect 1470 7233 1500 7287
rect 1570 7233 1600 7426
rect 1670 7464 1700 7517
rect 1770 7464 1800 7517
rect 1670 7454 1800 7464
rect 1670 7420 1718 7454
rect 1752 7420 1800 7454
rect 1670 7410 1800 7420
rect 1670 7373 1700 7410
rect 1770 7373 1800 7410
rect 1870 7480 1900 7517
rect 1970 7480 2000 7517
rect 1870 7470 2000 7480
rect 1870 7436 1918 7470
rect 1952 7436 2000 7470
rect 1870 7426 2000 7436
rect 1870 7373 1900 7426
rect 1970 7373 2000 7426
rect 2070 7464 2100 7517
rect 2170 7464 2200 7517
rect 2070 7454 2200 7464
rect 2070 7420 2118 7454
rect 2152 7420 2200 7454
rect 2070 7410 2200 7420
rect 2070 7373 2100 7410
rect 1670 7233 1700 7287
rect 1770 7233 1800 7287
rect 1870 7233 1900 7287
rect 1970 7233 2000 7287
rect 2070 7233 2100 7287
rect 2170 7233 2200 7410
rect 2270 7480 2300 7517
rect 2370 7480 2400 7517
rect 2270 7470 2400 7480
rect 2270 7436 2318 7470
rect 2352 7436 2400 7470
rect 2270 7426 2400 7436
rect 2270 7373 2300 7426
rect 2270 7233 2300 7287
rect 2370 7233 2400 7426
rect 2470 7464 2500 7517
rect 2570 7464 2600 7517
rect 2470 7454 2600 7464
rect 2470 7420 2518 7454
rect 2552 7420 2600 7454
rect 2470 7410 2600 7420
rect 2470 7373 2500 7410
rect 2470 7233 2500 7287
rect 470 7093 500 7147
rect 570 7093 600 7147
rect 670 7093 700 7147
rect 770 7093 800 7147
rect 870 7093 900 7147
rect 970 7093 1000 7147
rect 1070 7093 1100 7147
rect 1170 7093 1200 7147
rect 470 6953 500 7007
rect 570 6953 600 7007
rect 670 6953 700 7007
rect 770 6953 800 7007
rect 870 6953 900 7007
rect 970 6953 1000 7007
rect 1070 6953 1100 7007
rect 1170 6953 1200 7007
rect 1270 6953 1300 7147
rect 1370 7093 1400 7147
rect 1470 7093 1500 7147
rect 1570 7093 1600 7147
rect 1670 7093 1700 7147
rect 1770 7093 1800 7147
rect 1870 7093 1900 7147
rect 1970 7093 2000 7147
rect 2070 7093 2100 7147
rect 2170 7093 2200 7147
rect 1370 6953 1400 7007
rect 70 6813 100 6867
rect 170 6813 200 6867
rect 270 6813 300 6867
rect 370 6813 400 6867
rect 470 6813 500 6867
rect 570 6813 600 6867
rect 670 6813 700 6867
rect 770 6813 800 6867
rect 870 6813 900 6867
rect 970 6813 1000 6867
rect 1070 6813 1100 6867
rect 1170 6813 1200 6867
rect 1270 6813 1300 6867
rect 70 6673 100 6727
rect 170 6673 200 6727
rect 70 6533 100 6587
rect 170 6533 200 6587
rect 270 6533 300 6727
rect 370 6673 400 6727
rect 470 6673 500 6727
rect 570 6673 600 6727
rect 670 6673 700 6727
rect 770 6673 800 6727
rect 870 6673 900 6727
rect 970 6673 1000 6727
rect 370 6533 400 6587
rect 470 6533 500 6587
rect 70 6393 100 6447
rect 70 6254 100 6307
rect 170 6254 200 6447
rect 270 6393 300 6447
rect 370 6393 400 6447
rect 470 6393 500 6447
rect 570 6393 600 6587
rect 670 6533 700 6587
rect 770 6533 800 6587
rect 870 6533 900 6587
rect 970 6533 1000 6587
rect 1070 6533 1100 6727
rect 1170 6673 1200 6727
rect 1170 6533 1200 6587
rect 1270 6533 1300 6727
rect 1370 6673 1400 6867
rect 1470 6813 1500 7007
rect 1570 6953 1600 7007
rect 1670 6953 1700 7007
rect 1770 6953 1800 7007
rect 1870 6953 1900 7007
rect 1970 6953 2000 7007
rect 1470 6673 1500 6727
rect 1570 6673 1600 6867
rect 1670 6813 1700 6867
rect 1770 6813 1800 6867
rect 1870 6813 1900 6867
rect 1970 6813 2000 6867
rect 2070 6813 2100 7007
rect 2170 6953 2200 7007
rect 2270 6953 2300 7147
rect 2370 7093 2400 7147
rect 2470 7093 2500 7147
rect 2570 7093 2600 7410
rect 2670 7480 2700 7517
rect 2770 7480 2800 7797
rect 2870 7743 2900 7797
rect 2970 7743 3000 7797
rect 3070 7743 3100 7797
rect 3170 7743 3200 7797
rect 3270 7743 3300 7797
rect 3370 7743 3400 7937
rect 3470 7883 3500 7937
rect 3570 7883 3600 7937
rect 3670 7883 3700 7937
rect 3470 7743 3500 7797
rect 3570 7743 3600 7797
rect 3670 7743 3700 7797
rect 3770 7743 3800 7937
rect 3870 7883 3900 7937
rect 3870 7743 3900 7797
rect 3970 7743 4000 7937
rect 4070 7883 4100 7937
rect 4070 7743 4100 7797
rect 2870 7603 2900 7657
rect 2970 7603 3000 7657
rect 2670 7470 2800 7480
rect 2670 7436 2718 7470
rect 2752 7436 2800 7470
rect 2670 7426 2800 7436
rect 2670 7373 2700 7426
rect 2770 7373 2800 7426
rect 2870 7464 2900 7517
rect 2970 7464 3000 7517
rect 2870 7454 3000 7464
rect 2870 7420 2918 7454
rect 2952 7420 3000 7454
rect 2870 7410 3000 7420
rect 2870 7373 2900 7410
rect 2970 7373 3000 7410
rect 3070 7480 3100 7657
rect 3170 7603 3200 7657
rect 3170 7480 3200 7517
rect 3070 7470 3200 7480
rect 3070 7436 3118 7470
rect 3152 7436 3200 7470
rect 3070 7426 3200 7436
rect 3070 7373 3100 7426
rect 3170 7373 3200 7426
rect 3270 7464 3300 7657
rect 3370 7603 3400 7657
rect 3470 7603 3500 7657
rect 3570 7603 3600 7657
rect 3670 7603 3700 7657
rect 3770 7603 3800 7657
rect 3870 7603 3900 7657
rect 3370 7464 3400 7517
rect 3270 7454 3400 7464
rect 3270 7420 3318 7454
rect 3352 7420 3400 7454
rect 3270 7410 3400 7420
rect 3270 7373 3300 7410
rect 3370 7373 3400 7410
rect 3470 7480 3500 7517
rect 3570 7480 3600 7517
rect 3470 7470 3600 7480
rect 3470 7436 3518 7470
rect 3552 7436 3600 7470
rect 3470 7426 3600 7436
rect 3470 7373 3500 7426
rect 3570 7373 3600 7426
rect 3670 7464 3700 7517
rect 3770 7464 3800 7517
rect 3670 7454 3800 7464
rect 3670 7420 3718 7454
rect 3752 7420 3800 7454
rect 3670 7410 3800 7420
rect 3670 7373 3700 7410
rect 3770 7373 3800 7410
rect 3870 7480 3900 7517
rect 3970 7480 4000 7657
rect 4070 7603 4100 7657
rect 4170 7603 4200 7937
rect 4270 7883 4300 7937
rect 4370 7883 4400 7937
rect 4470 7883 4500 7937
rect 4270 7743 4300 7797
rect 4270 7603 4300 7657
rect 4370 7603 4400 7797
rect 4470 7743 4500 7797
rect 4570 7743 4600 7937
rect 4670 7883 4700 7937
rect 4670 7743 4700 7797
rect 4770 7743 4800 7937
rect 4870 7883 4900 7937
rect 4870 7743 4900 7797
rect 4970 7743 5000 8077
rect 5070 8023 5100 8077
rect 5170 8023 5200 8077
rect 5270 8023 5300 8077
rect 5370 8023 5400 8077
rect 5470 8023 5500 8077
rect 5570 8023 5600 8077
rect 5670 8023 5700 8077
rect 5770 8023 5800 8077
rect 5870 8023 5900 8077
rect 5970 8023 6000 8077
rect 6070 8023 6100 8077
rect 6170 8023 6200 8077
rect 6270 8023 6300 8077
rect 6370 8023 6400 8077
rect 6570 8023 6600 8077
rect 6670 8023 6700 8077
rect 6880 8023 6910 8077
rect 6980 8023 7010 8077
rect 7080 8023 7110 8077
rect 7180 8023 7210 8077
rect 7280 8023 7310 8077
rect 7380 8023 7410 8077
rect 5070 7883 5100 7937
rect 5170 7883 5200 7937
rect 5270 7883 5300 7937
rect 5370 7883 5400 7937
rect 5470 7883 5500 7937
rect 5070 7743 5100 7797
rect 5170 7743 5200 7797
rect 5270 7743 5300 7797
rect 5370 7743 5400 7797
rect 5470 7743 5500 7797
rect 4470 7603 4500 7657
rect 4570 7603 4600 7657
rect 4670 7603 4700 7657
rect 4770 7603 4800 7657
rect 4870 7603 4900 7657
rect 3870 7470 4000 7480
rect 3870 7436 3918 7470
rect 3952 7436 4000 7470
rect 3870 7426 4000 7436
rect 3870 7373 3900 7426
rect 3970 7373 4000 7426
rect 4070 7464 4100 7517
rect 4170 7464 4200 7517
rect 4070 7454 4200 7464
rect 4070 7420 4118 7454
rect 4152 7420 4200 7454
rect 4070 7410 4200 7420
rect 4070 7373 4100 7410
rect 4170 7373 4200 7410
rect 4270 7480 4300 7517
rect 4370 7480 4400 7517
rect 4270 7470 4400 7480
rect 4270 7436 4318 7470
rect 4352 7436 4400 7470
rect 4270 7426 4400 7436
rect 4270 7373 4300 7426
rect 4370 7373 4400 7426
rect 4470 7464 4500 7517
rect 4570 7464 4600 7517
rect 4470 7454 4600 7464
rect 4470 7420 4518 7454
rect 4552 7420 4600 7454
rect 4470 7410 4600 7420
rect 4470 7373 4500 7410
rect 4570 7373 4600 7410
rect 4670 7480 4700 7517
rect 4770 7480 4800 7517
rect 4670 7470 4800 7480
rect 4670 7436 4718 7470
rect 4752 7436 4800 7470
rect 4670 7426 4800 7436
rect 4670 7373 4700 7426
rect 4770 7373 4800 7426
rect 4870 7464 4900 7517
rect 4970 7464 5000 7657
rect 5070 7603 5100 7657
rect 4870 7454 5000 7464
rect 4870 7420 4918 7454
rect 4952 7420 5000 7454
rect 4870 7410 5000 7420
rect 4870 7373 4900 7410
rect 4970 7373 5000 7410
rect 5070 7480 5100 7517
rect 5170 7480 5200 7657
rect 5270 7603 5300 7657
rect 5370 7603 5400 7657
rect 5470 7603 5500 7657
rect 5570 7603 5600 7937
rect 5670 7883 5700 7937
rect 5670 7743 5700 7797
rect 5670 7603 5700 7657
rect 5770 7603 5800 7937
rect 5870 7883 5900 7937
rect 5970 7883 6000 7937
rect 6070 7883 6100 7937
rect 6170 7883 6200 7937
rect 6270 7883 6300 7937
rect 6370 7883 6400 7937
rect 6570 7883 6600 7937
rect 6670 7883 6700 7937
rect 6880 7883 6910 7937
rect 6980 7883 7010 7937
rect 7080 7883 7110 7937
rect 7180 7883 7210 7937
rect 7280 7883 7310 7937
rect 7380 7883 7410 7937
rect 5870 7743 5900 7797
rect 5970 7743 6000 7797
rect 6070 7743 6100 7797
rect 6170 7743 6200 7797
rect 6270 7743 6300 7797
rect 6370 7743 6400 7797
rect 6570 7743 6600 7797
rect 6670 7743 6700 7797
rect 6880 7743 6910 7797
rect 6980 7743 7010 7797
rect 7080 7743 7110 7797
rect 7180 7743 7210 7797
rect 7280 7743 7310 7797
rect 7380 7743 7410 7797
rect 5870 7603 5900 7657
rect 5970 7603 6000 7657
rect 6070 7603 6100 7657
rect 6170 7603 6200 7657
rect 6270 7603 6300 7657
rect 6370 7603 6400 7657
rect 6570 7603 6600 7657
rect 6670 7603 6700 7657
rect 6880 7603 6910 7657
rect 6980 7603 7010 7657
rect 7080 7603 7110 7657
rect 7180 7603 7210 7657
rect 7280 7603 7310 7657
rect 7380 7603 7410 7657
rect 5070 7470 5200 7480
rect 5070 7436 5118 7470
rect 5152 7436 5200 7470
rect 5070 7426 5200 7436
rect 5070 7373 5100 7426
rect 5170 7373 5200 7426
rect 5270 7464 5300 7517
rect 5370 7464 5400 7517
rect 5270 7454 5400 7464
rect 5270 7420 5318 7454
rect 5352 7420 5400 7454
rect 5270 7410 5400 7420
rect 5270 7373 5300 7410
rect 5370 7373 5400 7410
rect 5470 7480 5500 7517
rect 5570 7480 5600 7517
rect 5470 7470 5600 7480
rect 5470 7436 5518 7470
rect 5552 7436 5600 7470
rect 5470 7426 5600 7436
rect 5470 7373 5500 7426
rect 5570 7373 5600 7426
rect 5670 7464 5700 7517
rect 5770 7464 5800 7517
rect 5670 7454 5800 7464
rect 5670 7420 5718 7454
rect 5752 7420 5800 7454
rect 5670 7410 5800 7420
rect 5670 7373 5700 7410
rect 5770 7373 5800 7410
rect 5870 7480 5900 7517
rect 5970 7480 6000 7517
rect 5870 7470 6000 7480
rect 5870 7436 5918 7470
rect 5952 7436 6000 7470
rect 5870 7426 6000 7436
rect 5870 7373 5900 7426
rect 5970 7373 6000 7426
rect 6070 7464 6100 7517
rect 6170 7464 6200 7517
rect 6070 7454 6200 7464
rect 6070 7420 6118 7454
rect 6152 7420 6200 7454
rect 6070 7410 6200 7420
rect 6070 7373 6100 7410
rect 6170 7373 6200 7410
rect 6270 7480 6300 7517
rect 6370 7480 6400 7517
rect 6570 7484 6600 7517
rect 6670 7484 6700 7517
rect 6880 7484 6910 7517
rect 6980 7484 7010 7517
rect 7080 7484 7110 7517
rect 7180 7484 7210 7517
rect 7280 7484 7310 7517
rect 7380 7484 7410 7517
rect 6270 7470 6400 7480
rect 6270 7436 6318 7470
rect 6352 7436 6400 7470
rect 6270 7426 6400 7436
rect 6270 7373 6300 7426
rect 6370 7373 6400 7426
rect 6558 7468 6612 7484
rect 6558 7434 6568 7468
rect 6602 7434 6612 7468
rect 6558 7418 6612 7434
rect 6658 7468 6712 7484
rect 6658 7434 6668 7468
rect 6702 7434 6712 7468
rect 6658 7418 6712 7434
rect 6868 7468 6922 7484
rect 6868 7434 6878 7468
rect 6912 7434 6922 7468
rect 6868 7418 6922 7434
rect 6968 7468 7022 7484
rect 6968 7434 6978 7468
rect 7012 7434 7022 7468
rect 6968 7418 7022 7434
rect 7068 7468 7122 7484
rect 7068 7434 7078 7468
rect 7112 7434 7122 7468
rect 7068 7418 7122 7434
rect 7168 7468 7222 7484
rect 7168 7434 7178 7468
rect 7212 7434 7222 7468
rect 7168 7418 7222 7434
rect 7268 7468 7322 7484
rect 7268 7434 7278 7468
rect 7312 7434 7322 7468
rect 7268 7418 7322 7434
rect 7368 7468 7422 7484
rect 7368 7434 7378 7468
rect 7412 7434 7422 7468
rect 7368 7418 7422 7434
rect 6570 7373 6600 7418
rect 6670 7373 6700 7418
rect 6880 7373 6910 7418
rect 6980 7373 7010 7418
rect 7080 7373 7110 7418
rect 7180 7373 7210 7418
rect 7280 7373 7310 7418
rect 7380 7373 7410 7418
rect 2670 7233 2700 7287
rect 2770 7233 2800 7287
rect 2870 7233 2900 7287
rect 2670 7093 2700 7147
rect 2770 7093 2800 7147
rect 2870 7093 2900 7147
rect 2970 7093 3000 7287
rect 3070 7233 3100 7287
rect 3170 7233 3200 7287
rect 2370 6953 2400 7007
rect 2470 6953 2500 7007
rect 2570 6953 2600 7007
rect 2670 6953 2700 7007
rect 2770 6953 2800 7007
rect 2870 6953 2900 7007
rect 1670 6673 1700 6727
rect 1770 6673 1800 6727
rect 1870 6673 1900 6727
rect 1970 6673 2000 6727
rect 2070 6673 2100 6727
rect 2170 6673 2200 6867
rect 2270 6813 2300 6867
rect 2370 6813 2400 6867
rect 2470 6813 2500 6867
rect 2570 6813 2600 6867
rect 2670 6813 2700 6867
rect 2770 6813 2800 6867
rect 2870 6813 2900 6867
rect 2970 6813 3000 7007
rect 3070 6953 3100 7147
rect 3170 7093 3200 7147
rect 3270 7093 3300 7287
rect 3370 7233 3400 7287
rect 3470 7233 3500 7287
rect 3570 7233 3600 7287
rect 3670 7233 3700 7287
rect 3770 7233 3800 7287
rect 3870 7233 3900 7287
rect 3970 7233 4000 7287
rect 4070 7233 4100 7287
rect 4170 7233 4200 7287
rect 4270 7233 4300 7287
rect 3370 7093 3400 7147
rect 3070 6813 3100 6867
rect 3170 6813 3200 7007
rect 3270 6953 3300 7007
rect 3370 6953 3400 7007
rect 3270 6813 3300 6867
rect 3370 6813 3400 6867
rect 3470 6813 3500 7147
rect 3570 7093 3600 7147
rect 3670 7093 3700 7147
rect 3770 7093 3800 7147
rect 3870 7093 3900 7147
rect 3970 7093 4000 7147
rect 3570 6953 3600 7007
rect 3670 6953 3700 7007
rect 3770 6953 3800 7007
rect 3870 6953 3900 7007
rect 3970 6953 4000 7007
rect 4070 6953 4100 7147
rect 4170 7093 4200 7147
rect 4270 7093 4300 7147
rect 4370 7093 4400 7287
rect 4470 7233 4500 7287
rect 4570 7233 4600 7287
rect 4470 7093 4500 7147
rect 4570 7093 4600 7147
rect 4670 7093 4700 7287
rect 4770 7233 4800 7287
rect 4870 7233 4900 7287
rect 4970 7233 5000 7287
rect 4770 7093 4800 7147
rect 4870 7093 4900 7147
rect 4970 7093 5000 7147
rect 5070 7093 5100 7287
rect 5170 7233 5200 7287
rect 5270 7233 5300 7287
rect 5370 7233 5400 7287
rect 5470 7233 5500 7287
rect 5570 7233 5600 7287
rect 5670 7233 5700 7287
rect 5770 7233 5800 7287
rect 5870 7233 5900 7287
rect 5970 7233 6000 7287
rect 4170 6953 4200 7007
rect 3570 6813 3600 6867
rect 3670 6813 3700 6867
rect 3770 6813 3800 6867
rect 3870 6813 3900 6867
rect 3970 6813 4000 6867
rect 4070 6813 4100 6867
rect 4170 6813 4200 6867
rect 4270 6813 4300 7007
rect 4370 6953 4400 7007
rect 4470 6953 4500 7007
rect 4570 6953 4600 7007
rect 4670 6953 4700 7007
rect 4770 6953 4800 7007
rect 4370 6813 4400 6867
rect 4470 6813 4500 6867
rect 4570 6813 4600 6867
rect 4670 6813 4700 6867
rect 4770 6813 4800 6867
rect 4870 6813 4900 7007
rect 4970 6953 5000 7007
rect 5070 6953 5100 7007
rect 4970 6813 5000 6867
rect 5070 6813 5100 6867
rect 5170 6813 5200 7147
rect 5270 7093 5300 7147
rect 5370 7093 5400 7147
rect 5470 7093 5500 7147
rect 5570 7093 5600 7147
rect 5670 7093 5700 7147
rect 5770 7093 5800 7147
rect 5870 7093 5900 7147
rect 5970 7093 6000 7147
rect 6070 7093 6100 7287
rect 6170 7233 6200 7287
rect 6270 7233 6300 7287
rect 6370 7233 6400 7287
rect 6570 7233 6600 7287
rect 6670 7233 6700 7287
rect 6880 7233 6910 7287
rect 6980 7233 7010 7287
rect 7080 7233 7110 7287
rect 7180 7233 7210 7287
rect 7280 7233 7310 7287
rect 7380 7233 7410 7287
rect 5270 6953 5300 7007
rect 5270 6813 5300 6867
rect 5370 6813 5400 7007
rect 5470 6953 5500 7007
rect 5570 6953 5600 7007
rect 5670 6953 5700 7007
rect 5770 6953 5800 7007
rect 5870 6953 5900 7007
rect 5970 6953 6000 7007
rect 6070 6953 6100 7007
rect 2270 6673 2300 6727
rect 2370 6673 2400 6727
rect 2470 6673 2500 6727
rect 2570 6673 2600 6727
rect 2670 6673 2700 6727
rect 2770 6673 2800 6727
rect 2870 6673 2900 6727
rect 2970 6673 3000 6727
rect 3070 6673 3100 6727
rect 3170 6673 3200 6727
rect 3270 6673 3300 6727
rect 3370 6673 3400 6727
rect 1370 6533 1400 6587
rect 1470 6533 1500 6587
rect 1570 6533 1600 6587
rect 670 6393 700 6447
rect 770 6393 800 6447
rect 70 6244 200 6254
rect 70 6210 118 6244
rect 152 6210 200 6244
rect 70 6200 200 6210
rect 70 6163 100 6200
rect 170 6163 200 6200
rect 270 6270 300 6307
rect 370 6270 400 6307
rect 270 6260 400 6270
rect 270 6226 318 6260
rect 352 6226 400 6260
rect 270 6216 400 6226
rect 270 6163 300 6216
rect 370 6163 400 6216
rect 470 6254 500 6307
rect 570 6254 600 6307
rect 470 6244 600 6254
rect 470 6210 518 6244
rect 552 6210 600 6244
rect 470 6200 600 6210
rect 470 6163 500 6200
rect 570 6163 600 6200
rect 670 6270 700 6307
rect 770 6270 800 6307
rect 670 6260 800 6270
rect 670 6226 718 6260
rect 752 6226 800 6260
rect 670 6216 800 6226
rect 670 6163 700 6216
rect 770 6163 800 6216
rect 870 6254 900 6447
rect 970 6393 1000 6447
rect 970 6254 1000 6307
rect 870 6244 1000 6254
rect 870 6210 918 6244
rect 952 6210 1000 6244
rect 870 6200 1000 6210
rect 870 6163 900 6200
rect 970 6163 1000 6200
rect 1070 6270 1100 6447
rect 1170 6393 1200 6447
rect 1270 6393 1300 6447
rect 1370 6393 1400 6447
rect 1470 6393 1500 6447
rect 1570 6393 1600 6447
rect 1170 6270 1200 6307
rect 1070 6260 1200 6270
rect 1070 6226 1118 6260
rect 1152 6226 1200 6260
rect 1070 6216 1200 6226
rect 1070 6163 1100 6216
rect 1170 6163 1200 6216
rect 1270 6254 1300 6307
rect 1370 6254 1400 6307
rect 1270 6244 1400 6254
rect 1270 6210 1318 6244
rect 1352 6210 1400 6244
rect 1270 6200 1400 6210
rect 1270 6163 1300 6200
rect 1370 6163 1400 6200
rect 1470 6270 1500 6307
rect 1570 6270 1600 6307
rect 1470 6260 1600 6270
rect 1470 6226 1518 6260
rect 1552 6226 1600 6260
rect 1470 6216 1600 6226
rect 1470 6163 1500 6216
rect 1570 6163 1600 6216
rect 1670 6254 1700 6587
rect 1770 6533 1800 6587
rect 1870 6533 1900 6587
rect 1970 6533 2000 6587
rect 2070 6533 2100 6587
rect 2170 6533 2200 6587
rect 2270 6533 2300 6587
rect 2370 6533 2400 6587
rect 2470 6533 2500 6587
rect 2570 6533 2600 6587
rect 2670 6533 2700 6587
rect 2770 6533 2800 6587
rect 2870 6533 2900 6587
rect 2970 6533 3000 6587
rect 3070 6533 3100 6587
rect 3170 6533 3200 6587
rect 3270 6533 3300 6587
rect 3370 6533 3400 6587
rect 3470 6533 3500 6727
rect 3570 6673 3600 6727
rect 3570 6533 3600 6587
rect 3670 6533 3700 6727
rect 3770 6673 3800 6727
rect 3870 6673 3900 6727
rect 3970 6673 4000 6727
rect 4070 6673 4100 6727
rect 4170 6673 4200 6727
rect 4270 6673 4300 6727
rect 4370 6673 4400 6727
rect 1770 6393 1800 6447
rect 1870 6393 1900 6447
rect 1770 6254 1800 6307
rect 1670 6244 1800 6254
rect 1670 6210 1718 6244
rect 1752 6210 1800 6244
rect 1670 6200 1800 6210
rect 1670 6163 1700 6200
rect 1770 6163 1800 6200
rect 1870 6270 1900 6307
rect 1970 6270 2000 6447
rect 2070 6393 2100 6447
rect 2170 6393 2200 6447
rect 2270 6393 2300 6447
rect 2370 6393 2400 6447
rect 2470 6393 2500 6447
rect 2570 6393 2600 6447
rect 2670 6393 2700 6447
rect 2770 6393 2800 6447
rect 1870 6260 2000 6270
rect 1870 6226 1918 6260
rect 1952 6226 2000 6260
rect 1870 6216 2000 6226
rect 1870 6163 1900 6216
rect 1970 6163 2000 6216
rect 2070 6254 2100 6307
rect 2170 6254 2200 6307
rect 2070 6244 2200 6254
rect 2070 6210 2118 6244
rect 2152 6210 2200 6244
rect 2070 6200 2200 6210
rect 2070 6163 2100 6200
rect 2170 6163 2200 6200
rect 2270 6270 2300 6307
rect 2370 6270 2400 6307
rect 2270 6260 2400 6270
rect 2270 6226 2318 6260
rect 2352 6226 2400 6260
rect 2270 6216 2400 6226
rect 2270 6163 2300 6216
rect 2370 6163 2400 6216
rect 2470 6254 2500 6307
rect 2570 6254 2600 6307
rect 2470 6244 2600 6254
rect 2470 6210 2518 6244
rect 2552 6210 2600 6244
rect 2470 6200 2600 6210
rect 70 6023 100 6077
rect 170 6023 200 6077
rect 270 6023 300 6077
rect 370 6023 400 6077
rect 70 5883 100 5937
rect 170 5883 200 5937
rect 270 5883 300 5937
rect 370 5883 400 5937
rect 470 5883 500 6077
rect 570 6023 600 6077
rect 670 6023 700 6077
rect 770 6023 800 6077
rect 870 6023 900 6077
rect 970 6023 1000 6077
rect 1070 6023 1100 6077
rect 1170 6023 1200 6077
rect 1270 6023 1300 6077
rect 570 5883 600 5937
rect 670 5883 700 5937
rect 770 5883 800 5937
rect 870 5883 900 5937
rect 970 5883 1000 5937
rect 1070 5883 1100 5937
rect 1170 5883 1200 5937
rect 1270 5883 1300 5937
rect 1370 5883 1400 6077
rect 1470 6023 1500 6077
rect 1570 6023 1600 6077
rect 1670 6023 1700 6077
rect 1770 6023 1800 6077
rect 1870 6023 1900 6077
rect 1970 6023 2000 6077
rect 2070 6023 2100 6077
rect 2170 6023 2200 6077
rect 2270 6023 2300 6077
rect 2370 6023 2400 6077
rect 2470 6023 2500 6200
rect 2570 6163 2600 6200
rect 2670 6270 2700 6307
rect 2770 6270 2800 6307
rect 2670 6260 2800 6270
rect 2670 6226 2718 6260
rect 2752 6226 2800 6260
rect 2670 6216 2800 6226
rect 2670 6163 2700 6216
rect 2770 6163 2800 6216
rect 2870 6254 2900 6447
rect 2970 6393 3000 6447
rect 3070 6393 3100 6447
rect 3170 6393 3200 6447
rect 3270 6393 3300 6447
rect 2970 6254 3000 6307
rect 2870 6244 3000 6254
rect 2870 6210 2918 6244
rect 2952 6210 3000 6244
rect 2870 6200 3000 6210
rect 2870 6163 2900 6200
rect 2970 6163 3000 6200
rect 3070 6270 3100 6307
rect 3170 6270 3200 6307
rect 3070 6260 3200 6270
rect 3070 6226 3118 6260
rect 3152 6226 3200 6260
rect 3070 6216 3200 6226
rect 3070 6163 3100 6216
rect 3170 6163 3200 6216
rect 3270 6254 3300 6307
rect 3370 6254 3400 6447
rect 3470 6393 3500 6447
rect 3570 6393 3600 6447
rect 3670 6393 3700 6447
rect 3770 6393 3800 6587
rect 3870 6533 3900 6587
rect 3970 6533 4000 6587
rect 4070 6533 4100 6587
rect 4170 6533 4200 6587
rect 4270 6533 4300 6587
rect 4370 6533 4400 6587
rect 4470 6533 4500 6727
rect 4570 6673 4600 6727
rect 4670 6673 4700 6727
rect 4770 6673 4800 6727
rect 4870 6673 4900 6727
rect 4970 6673 5000 6727
rect 5070 6673 5100 6727
rect 5170 6673 5200 6727
rect 5270 6673 5300 6727
rect 5370 6673 5400 6727
rect 5470 6673 5500 6867
rect 5570 6813 5600 6867
rect 5570 6673 5600 6727
rect 5670 6673 5700 6867
rect 5770 6813 5800 6867
rect 5770 6673 5800 6727
rect 4570 6533 4600 6587
rect 4670 6533 4700 6587
rect 4770 6533 4800 6587
rect 4870 6533 4900 6587
rect 4970 6533 5000 6587
rect 5070 6533 5100 6587
rect 3870 6393 3900 6447
rect 3970 6393 4000 6447
rect 4070 6393 4100 6447
rect 4170 6393 4200 6447
rect 4270 6393 4300 6447
rect 4370 6393 4400 6447
rect 4470 6393 4500 6447
rect 4570 6393 4600 6447
rect 4670 6393 4700 6447
rect 4770 6393 4800 6447
rect 4870 6393 4900 6447
rect 4970 6393 5000 6447
rect 3270 6244 3400 6254
rect 3270 6210 3318 6244
rect 3352 6210 3400 6244
rect 3270 6200 3400 6210
rect 3270 6163 3300 6200
rect 3370 6163 3400 6200
rect 3470 6270 3500 6307
rect 3570 6270 3600 6307
rect 3470 6260 3600 6270
rect 3470 6226 3518 6260
rect 3552 6226 3600 6260
rect 3470 6216 3600 6226
rect 3470 6163 3500 6216
rect 3570 6163 3600 6216
rect 3670 6254 3700 6307
rect 3770 6254 3800 6307
rect 3670 6244 3800 6254
rect 3670 6210 3718 6244
rect 3752 6210 3800 6244
rect 3670 6200 3800 6210
rect 3670 6163 3700 6200
rect 2570 6023 2600 6077
rect 2670 6023 2700 6077
rect 2770 6023 2800 6077
rect 2870 6023 2900 6077
rect 2970 6023 3000 6077
rect 3070 6023 3100 6077
rect 3170 6023 3200 6077
rect 3270 6023 3300 6077
rect 1470 5883 1500 5937
rect 1570 5883 1600 5937
rect 1670 5883 1700 5937
rect 1770 5883 1800 5937
rect 1870 5883 1900 5937
rect 1970 5883 2000 5937
rect 70 5743 100 5797
rect 170 5743 200 5797
rect 270 5743 300 5797
rect 70 5603 100 5657
rect 170 5603 200 5657
rect 270 5603 300 5657
rect 370 5603 400 5797
rect 470 5743 500 5797
rect 570 5743 600 5797
rect 670 5743 700 5797
rect 770 5743 800 5797
rect 870 5743 900 5797
rect 970 5743 1000 5797
rect 470 5603 500 5657
rect 570 5603 600 5657
rect 670 5603 700 5657
rect 770 5603 800 5657
rect 870 5603 900 5657
rect 970 5603 1000 5657
rect 1070 5603 1100 5797
rect 1170 5743 1200 5797
rect 1270 5743 1300 5797
rect 1370 5743 1400 5797
rect 1470 5743 1500 5797
rect 1570 5743 1600 5797
rect 1670 5743 1700 5797
rect 1770 5743 1800 5797
rect 1870 5743 1900 5797
rect 1970 5743 2000 5797
rect 2070 5743 2100 5937
rect 2170 5883 2200 5937
rect 2270 5883 2300 5937
rect 2370 5883 2400 5937
rect 2470 5883 2500 5937
rect 2570 5883 2600 5937
rect 2670 5883 2700 5937
rect 2770 5883 2800 5937
rect 2870 5883 2900 5937
rect 2970 5883 3000 5937
rect 3070 5883 3100 5937
rect 3170 5883 3200 5937
rect 3270 5883 3300 5937
rect 3370 5883 3400 6077
rect 3470 6023 3500 6077
rect 3570 6023 3600 6077
rect 3670 6023 3700 6077
rect 3770 6023 3800 6200
rect 3870 6270 3900 6307
rect 3970 6270 4000 6307
rect 3870 6260 4000 6270
rect 3870 6226 3918 6260
rect 3952 6226 4000 6260
rect 3870 6216 4000 6226
rect 3870 6163 3900 6216
rect 3970 6163 4000 6216
rect 4070 6254 4100 6307
rect 4170 6254 4200 6307
rect 4070 6244 4200 6254
rect 4070 6210 4118 6244
rect 4152 6210 4200 6244
rect 4070 6200 4200 6210
rect 3870 6023 3900 6077
rect 3970 6023 4000 6077
rect 4070 6023 4100 6200
rect 4170 6163 4200 6200
rect 4270 6270 4300 6307
rect 4370 6270 4400 6307
rect 4270 6260 4400 6270
rect 4270 6226 4318 6260
rect 4352 6226 4400 6260
rect 4270 6216 4400 6226
rect 4270 6163 4300 6216
rect 4370 6163 4400 6216
rect 4470 6254 4500 6307
rect 4570 6254 4600 6307
rect 4470 6244 4600 6254
rect 4470 6210 4518 6244
rect 4552 6210 4600 6244
rect 4470 6200 4600 6210
rect 4170 6023 4200 6077
rect 4270 6023 4300 6077
rect 4370 6023 4400 6077
rect 4470 6023 4500 6200
rect 4570 6163 4600 6200
rect 4670 6270 4700 6307
rect 4770 6270 4800 6307
rect 4670 6260 4800 6270
rect 4670 6226 4718 6260
rect 4752 6226 4800 6260
rect 4670 6216 4800 6226
rect 4570 6023 4600 6077
rect 4670 6023 4700 6216
rect 4770 6163 4800 6216
rect 4870 6254 4900 6307
rect 4970 6254 5000 6307
rect 4870 6244 5000 6254
rect 4870 6210 4918 6244
rect 4952 6210 5000 6244
rect 4870 6200 5000 6210
rect 4870 6163 4900 6200
rect 4970 6163 5000 6200
rect 5070 6270 5100 6447
rect 5170 6393 5200 6587
rect 5270 6533 5300 6587
rect 5270 6393 5300 6447
rect 5170 6270 5200 6307
rect 5070 6260 5200 6270
rect 5070 6226 5118 6260
rect 5152 6226 5200 6260
rect 5070 6216 5200 6226
rect 5070 6163 5100 6216
rect 5170 6163 5200 6216
rect 5270 6254 5300 6307
rect 5370 6254 5400 6587
rect 5470 6533 5500 6587
rect 5570 6533 5600 6587
rect 5670 6533 5700 6587
rect 5770 6533 5800 6587
rect 5870 6533 5900 6867
rect 5970 6813 6000 6867
rect 6070 6813 6100 6867
rect 6170 6813 6200 7147
rect 6270 7093 6300 7147
rect 6370 7093 6400 7147
rect 6570 7093 6600 7147
rect 6670 7093 6700 7147
rect 6880 7093 6910 7147
rect 6980 7093 7010 7147
rect 7080 7093 7110 7147
rect 7180 7093 7210 7147
rect 7280 7093 7310 7147
rect 7380 7093 7410 7147
rect 6270 6953 6300 7007
rect 6370 6953 6400 7007
rect 6570 6953 6600 7007
rect 6670 6953 6700 7007
rect 6880 6953 6910 7007
rect 6980 6953 7010 7007
rect 7080 6953 7110 7007
rect 7180 6953 7210 7007
rect 7280 6953 7310 7007
rect 7380 6953 7410 7007
rect 6270 6813 6300 6867
rect 6370 6813 6400 6867
rect 6570 6813 6600 6867
rect 6670 6813 6700 6867
rect 6880 6813 6910 6867
rect 6980 6813 7010 6867
rect 7080 6813 7110 6867
rect 7180 6813 7210 6867
rect 7280 6813 7310 6867
rect 7380 6813 7410 6867
rect 5970 6673 6000 6727
rect 6070 6673 6100 6727
rect 6170 6673 6200 6727
rect 6270 6673 6300 6727
rect 6370 6673 6400 6727
rect 6570 6673 6600 6727
rect 6670 6673 6700 6727
rect 6880 6673 6910 6727
rect 6980 6673 7010 6727
rect 7080 6673 7110 6727
rect 7180 6673 7210 6727
rect 7280 6673 7310 6727
rect 7380 6673 7410 6727
rect 5970 6533 6000 6587
rect 6070 6533 6100 6587
rect 6170 6533 6200 6587
rect 6270 6533 6300 6587
rect 6370 6533 6400 6587
rect 6570 6533 6600 6587
rect 6670 6533 6700 6587
rect 6880 6533 6910 6587
rect 6980 6533 7010 6587
rect 7080 6533 7110 6587
rect 7180 6533 7210 6587
rect 7280 6533 7310 6587
rect 7380 6533 7410 6587
rect 5470 6393 5500 6447
rect 5570 6393 5600 6447
rect 5670 6393 5700 6447
rect 5770 6393 5800 6447
rect 5870 6393 5900 6447
rect 5970 6393 6000 6447
rect 6070 6393 6100 6447
rect 5270 6244 5400 6254
rect 5270 6210 5318 6244
rect 5352 6210 5400 6244
rect 5270 6200 5400 6210
rect 5270 6163 5300 6200
rect 5370 6163 5400 6200
rect 5470 6270 5500 6307
rect 5570 6270 5600 6307
rect 5470 6260 5600 6270
rect 5470 6226 5518 6260
rect 5552 6226 5600 6260
rect 5470 6216 5600 6226
rect 5470 6163 5500 6216
rect 5570 6163 5600 6216
rect 5670 6254 5700 6307
rect 5770 6254 5800 6307
rect 5670 6244 5800 6254
rect 5670 6210 5718 6244
rect 5752 6210 5800 6244
rect 5670 6200 5800 6210
rect 5670 6163 5700 6200
rect 5770 6163 5800 6200
rect 5870 6270 5900 6307
rect 5970 6270 6000 6307
rect 5870 6260 6000 6270
rect 5870 6226 5918 6260
rect 5952 6226 6000 6260
rect 5870 6216 6000 6226
rect 5870 6163 5900 6216
rect 5970 6163 6000 6216
rect 6070 6254 6100 6307
rect 6170 6254 6200 6447
rect 6270 6393 6300 6447
rect 6370 6393 6400 6447
rect 6570 6393 6600 6447
rect 6670 6393 6700 6447
rect 6880 6393 6910 6447
rect 6980 6393 7010 6447
rect 7080 6393 7110 6447
rect 7180 6393 7210 6447
rect 7280 6393 7310 6447
rect 7380 6393 7410 6447
rect 6070 6244 6200 6254
rect 6070 6210 6118 6244
rect 6152 6210 6200 6244
rect 6070 6200 6200 6210
rect 4770 6023 4800 6077
rect 4870 6023 4900 6077
rect 4970 6023 5000 6077
rect 5070 6023 5100 6077
rect 5170 6023 5200 6077
rect 2170 5743 2200 5797
rect 2270 5743 2300 5797
rect 2370 5743 2400 5797
rect 2470 5743 2500 5797
rect 2570 5743 2600 5797
rect 2670 5743 2700 5797
rect 2770 5743 2800 5797
rect 70 5463 100 5517
rect 170 5463 200 5517
rect 270 5463 300 5517
rect 370 5463 400 5517
rect 70 5323 100 5377
rect 170 5323 200 5377
rect 270 5323 300 5377
rect 370 5323 400 5377
rect 470 5323 500 5517
rect 570 5463 600 5517
rect 670 5463 700 5517
rect 770 5463 800 5517
rect 870 5463 900 5517
rect 970 5463 1000 5517
rect 1070 5463 1100 5517
rect 1170 5463 1200 5657
rect 1270 5603 1300 5657
rect 1270 5463 1300 5517
rect 1370 5463 1400 5657
rect 1470 5603 1500 5657
rect 1570 5603 1600 5657
rect 1670 5603 1700 5657
rect 1770 5603 1800 5657
rect 1870 5603 1900 5657
rect 570 5323 600 5377
rect 670 5323 700 5377
rect 770 5323 800 5377
rect 870 5323 900 5377
rect 970 5323 1000 5377
rect 1070 5323 1100 5377
rect 1170 5323 1200 5377
rect 1270 5323 1300 5377
rect 1370 5323 1400 5377
rect 1470 5323 1500 5517
rect 1570 5463 1600 5517
rect 1670 5463 1700 5517
rect 1570 5323 1600 5377
rect 1670 5323 1700 5377
rect 1770 5323 1800 5517
rect 1870 5463 1900 5517
rect 1970 5463 2000 5657
rect 2070 5603 2100 5657
rect 2170 5603 2200 5657
rect 2070 5463 2100 5517
rect 2170 5463 2200 5517
rect 1870 5323 1900 5377
rect 1970 5323 2000 5377
rect 2070 5323 2100 5377
rect 70 5183 100 5237
rect 170 5183 200 5237
rect 270 5183 300 5237
rect 370 5183 400 5237
rect 470 5183 500 5237
rect 570 5183 600 5237
rect 670 5183 700 5237
rect 770 5183 800 5237
rect 870 5183 900 5237
rect 970 5183 1000 5237
rect 1070 5183 1100 5237
rect 1170 5183 1200 5237
rect 1270 5183 1300 5237
rect 70 4904 100 5097
rect 170 4904 200 5097
rect 70 4894 200 4904
rect 70 4860 118 4894
rect 152 4860 200 4894
rect 70 4850 200 4860
rect 70 4813 100 4850
rect 170 4813 200 4850
rect 270 4920 300 5097
rect 370 4920 400 5097
rect 270 4910 400 4920
rect 270 4876 318 4910
rect 352 4876 400 4910
rect 270 4866 400 4876
rect 70 4673 100 4727
rect 170 4673 200 4727
rect 270 4673 300 4866
rect 370 4813 400 4866
rect 470 4904 500 5097
rect 570 4904 600 5097
rect 470 4894 600 4904
rect 470 4860 518 4894
rect 552 4860 600 4894
rect 470 4850 600 4860
rect 470 4813 500 4850
rect 570 4813 600 4850
rect 670 4920 700 5097
rect 770 4920 800 5097
rect 670 4910 800 4920
rect 670 4876 718 4910
rect 752 4876 800 4910
rect 670 4866 800 4876
rect 670 4813 700 4866
rect 770 4813 800 4866
rect 870 4904 900 5097
rect 970 4904 1000 5097
rect 870 4894 1000 4904
rect 870 4860 918 4894
rect 952 4860 1000 4894
rect 870 4850 1000 4860
rect 870 4813 900 4850
rect 970 4813 1000 4850
rect 1070 4920 1100 5097
rect 1170 4920 1200 5097
rect 1070 4910 1200 4920
rect 1070 4876 1118 4910
rect 1152 4876 1200 4910
rect 1070 4866 1200 4876
rect 1070 4813 1100 4866
rect 370 4673 400 4727
rect 470 4673 500 4727
rect 570 4673 600 4727
rect 670 4673 700 4727
rect 770 4673 800 4727
rect 870 4673 900 4727
rect 970 4673 1000 4727
rect 1070 4673 1100 4727
rect 1170 4673 1200 4866
rect 1270 4904 1300 5097
rect 1370 4904 1400 5237
rect 1470 5183 1500 5237
rect 1570 5183 1600 5237
rect 1670 5183 1700 5237
rect 1770 5183 1800 5237
rect 1870 5183 1900 5237
rect 1970 5183 2000 5237
rect 2070 5183 2100 5237
rect 1270 4894 1400 4904
rect 1270 4860 1318 4894
rect 1352 4860 1400 4894
rect 1270 4850 1400 4860
rect 1270 4813 1300 4850
rect 1370 4813 1400 4850
rect 1470 4920 1500 5097
rect 1570 4920 1600 5097
rect 1470 4910 1600 4920
rect 1470 4876 1518 4910
rect 1552 4876 1600 4910
rect 1470 4866 1600 4876
rect 1470 4813 1500 4866
rect 1570 4813 1600 4866
rect 1670 4904 1700 5097
rect 1770 4904 1800 5097
rect 1670 4894 1800 4904
rect 1670 4860 1718 4894
rect 1752 4860 1800 4894
rect 1670 4850 1800 4860
rect 1670 4813 1700 4850
rect 1770 4813 1800 4850
rect 1870 4920 1900 5097
rect 1970 4920 2000 5097
rect 1870 4910 2000 4920
rect 1870 4876 1918 4910
rect 1952 4876 2000 4910
rect 1870 4866 2000 4876
rect 1870 4813 1900 4866
rect 1970 4813 2000 4866
rect 2070 4904 2100 5097
rect 2170 4904 2200 5377
rect 2270 5323 2300 5657
rect 2370 5603 2400 5657
rect 2470 5603 2500 5657
rect 2570 5603 2600 5657
rect 2670 5603 2700 5657
rect 2770 5603 2800 5657
rect 2870 5603 2900 5797
rect 2970 5743 3000 5797
rect 2970 5603 3000 5657
rect 3070 5603 3100 5797
rect 3170 5743 3200 5797
rect 3170 5603 3200 5657
rect 3270 5603 3300 5797
rect 3370 5743 3400 5797
rect 3370 5603 3400 5657
rect 3470 5603 3500 5937
rect 3570 5883 3600 5937
rect 3670 5883 3700 5937
rect 3770 5883 3800 5937
rect 3870 5883 3900 5937
rect 3970 5883 4000 5937
rect 4070 5883 4100 5937
rect 3570 5743 3600 5797
rect 3570 5603 3600 5657
rect 3670 5603 3700 5797
rect 3770 5743 3800 5797
rect 3870 5743 3900 5797
rect 3970 5743 4000 5797
rect 4070 5743 4100 5797
rect 3770 5603 3800 5657
rect 3870 5603 3900 5657
rect 3970 5603 4000 5657
rect 2370 5463 2400 5517
rect 2470 5463 2500 5517
rect 2570 5463 2600 5517
rect 2670 5463 2700 5517
rect 2770 5463 2800 5517
rect 2870 5463 2900 5517
rect 2970 5463 3000 5517
rect 3070 5463 3100 5517
rect 3170 5463 3200 5517
rect 3270 5463 3300 5517
rect 3370 5463 3400 5517
rect 3470 5463 3500 5517
rect 3570 5463 3600 5517
rect 3670 5463 3700 5517
rect 2270 5183 2300 5237
rect 2370 5183 2400 5377
rect 2470 5323 2500 5377
rect 2570 5323 2600 5377
rect 2470 5183 2500 5237
rect 2570 5183 2600 5237
rect 2670 5183 2700 5377
rect 2770 5323 2800 5377
rect 2870 5323 2900 5377
rect 2770 5183 2800 5237
rect 2870 5183 2900 5237
rect 2970 5183 3000 5377
rect 3070 5323 3100 5377
rect 3070 5183 3100 5237
rect 3170 5183 3200 5377
rect 3270 5323 3300 5377
rect 3370 5323 3400 5377
rect 3470 5323 3500 5377
rect 3570 5323 3600 5377
rect 3670 5323 3700 5377
rect 3770 5323 3800 5517
rect 3870 5463 3900 5517
rect 3970 5463 4000 5517
rect 4070 5463 4100 5657
rect 4170 5603 4200 5937
rect 4270 5883 4300 5937
rect 4370 5883 4400 5937
rect 4470 5883 4500 5937
rect 4570 5883 4600 5937
rect 4670 5883 4700 5937
rect 4770 5883 4800 5937
rect 4870 5883 4900 5937
rect 4970 5883 5000 5937
rect 5070 5883 5100 5937
rect 5170 5883 5200 5937
rect 5270 5883 5300 6077
rect 5370 6023 5400 6077
rect 5470 6023 5500 6077
rect 5570 6023 5600 6077
rect 5670 6023 5700 6077
rect 5770 6023 5800 6077
rect 5370 5883 5400 5937
rect 5470 5883 5500 5937
rect 5570 5883 5600 5937
rect 5670 5883 5700 5937
rect 4270 5743 4300 5797
rect 4270 5603 4300 5657
rect 4370 5603 4400 5797
rect 4470 5743 4500 5797
rect 4470 5603 4500 5657
rect 4570 5603 4600 5797
rect 4670 5743 4700 5797
rect 4770 5743 4800 5797
rect 4870 5743 4900 5797
rect 4970 5743 5000 5797
rect 5070 5743 5100 5797
rect 5170 5743 5200 5797
rect 5270 5743 5300 5797
rect 5370 5743 5400 5797
rect 5470 5743 5500 5797
rect 4670 5603 4700 5657
rect 4770 5603 4800 5657
rect 4870 5603 4900 5657
rect 4970 5603 5000 5657
rect 5070 5603 5100 5657
rect 5170 5603 5200 5657
rect 5270 5603 5300 5657
rect 5370 5603 5400 5657
rect 5470 5603 5500 5657
rect 5570 5603 5600 5797
rect 5670 5743 5700 5797
rect 5770 5743 5800 5937
rect 5870 5883 5900 6077
rect 5970 6023 6000 6077
rect 6070 6023 6100 6200
rect 6170 6163 6200 6200
rect 6270 6270 6300 6307
rect 6370 6270 6400 6307
rect 6570 6274 6600 6307
rect 6670 6274 6700 6307
rect 6880 6274 6910 6307
rect 6980 6274 7010 6307
rect 7080 6274 7110 6307
rect 7180 6274 7210 6307
rect 7280 6274 7310 6307
rect 7380 6274 7410 6307
rect 6270 6260 6400 6270
rect 6270 6226 6318 6260
rect 6352 6226 6400 6260
rect 6270 6216 6400 6226
rect 6170 6023 6200 6077
rect 6270 6023 6300 6216
rect 6370 6163 6400 6216
rect 6558 6258 6612 6274
rect 6558 6224 6568 6258
rect 6602 6224 6612 6258
rect 6558 6208 6612 6224
rect 6658 6258 6712 6274
rect 6658 6224 6668 6258
rect 6702 6224 6712 6258
rect 6658 6208 6712 6224
rect 6868 6258 6922 6274
rect 6868 6224 6878 6258
rect 6912 6224 6922 6258
rect 6868 6208 6922 6224
rect 6968 6258 7022 6274
rect 6968 6224 6978 6258
rect 7012 6224 7022 6258
rect 6968 6208 7022 6224
rect 7068 6258 7122 6274
rect 7068 6224 7078 6258
rect 7112 6224 7122 6258
rect 7068 6208 7122 6224
rect 7168 6258 7222 6274
rect 7168 6224 7178 6258
rect 7212 6224 7222 6258
rect 7168 6208 7222 6224
rect 7268 6258 7322 6274
rect 7268 6224 7278 6258
rect 7312 6224 7322 6258
rect 7268 6208 7322 6224
rect 7368 6258 7422 6274
rect 7368 6224 7378 6258
rect 7412 6224 7422 6258
rect 7368 6208 7422 6224
rect 6570 6163 6600 6208
rect 6670 6163 6700 6208
rect 6880 6163 6910 6208
rect 6980 6163 7010 6208
rect 7080 6163 7110 6208
rect 7180 6163 7210 6208
rect 7280 6163 7310 6208
rect 7380 6163 7410 6208
rect 6370 6023 6400 6077
rect 6570 6023 6600 6077
rect 6670 6023 6700 6077
rect 6880 6023 6910 6077
rect 6980 6023 7010 6077
rect 7080 6023 7110 6077
rect 7180 6023 7210 6077
rect 7280 6023 7310 6077
rect 7380 6023 7410 6077
rect 5870 5743 5900 5797
rect 5970 5743 6000 5937
rect 6070 5883 6100 5937
rect 6170 5883 6200 5937
rect 6270 5883 6300 5937
rect 6370 5883 6400 5937
rect 6570 5883 6600 5937
rect 6670 5883 6700 5937
rect 6880 5883 6910 5937
rect 6980 5883 7010 5937
rect 7080 5883 7110 5937
rect 7180 5883 7210 5937
rect 7280 5883 7310 5937
rect 7380 5883 7410 5937
rect 6070 5743 6100 5797
rect 6170 5743 6200 5797
rect 6270 5743 6300 5797
rect 6370 5743 6400 5797
rect 6570 5743 6600 5797
rect 6670 5743 6700 5797
rect 6880 5743 6910 5797
rect 6980 5743 7010 5797
rect 7080 5743 7110 5797
rect 7180 5743 7210 5797
rect 7280 5743 7310 5797
rect 7380 5743 7410 5797
rect 5670 5603 5700 5657
rect 5770 5603 5800 5657
rect 5870 5603 5900 5657
rect 5970 5603 6000 5657
rect 6070 5603 6100 5657
rect 6170 5603 6200 5657
rect 6270 5603 6300 5657
rect 6370 5603 6400 5657
rect 6570 5603 6600 5657
rect 6670 5603 6700 5657
rect 6880 5603 6910 5657
rect 6980 5603 7010 5657
rect 7080 5603 7110 5657
rect 7180 5603 7210 5657
rect 7280 5603 7310 5657
rect 7380 5603 7410 5657
rect 4170 5463 4200 5517
rect 4270 5463 4300 5517
rect 4370 5463 4400 5517
rect 4470 5463 4500 5517
rect 4570 5463 4600 5517
rect 4670 5463 4700 5517
rect 4770 5463 4800 5517
rect 4870 5463 4900 5517
rect 4970 5463 5000 5517
rect 5070 5463 5100 5517
rect 3870 5323 3900 5377
rect 3970 5323 4000 5377
rect 4070 5323 4100 5377
rect 4170 5323 4200 5377
rect 4270 5323 4300 5377
rect 4370 5323 4400 5377
rect 4470 5323 4500 5377
rect 4570 5323 4600 5377
rect 4670 5323 4700 5377
rect 4770 5323 4800 5377
rect 4870 5323 4900 5377
rect 4970 5323 5000 5377
rect 5070 5323 5100 5377
rect 5170 5323 5200 5517
rect 5270 5463 5300 5517
rect 3270 5183 3300 5237
rect 3370 5183 3400 5237
rect 3470 5183 3500 5237
rect 3570 5183 3600 5237
rect 3670 5183 3700 5237
rect 3770 5183 3800 5237
rect 3870 5183 3900 5237
rect 3970 5183 4000 5237
rect 4070 5183 4100 5237
rect 4170 5183 4200 5237
rect 4270 5183 4300 5237
rect 2070 4894 2200 4904
rect 2070 4860 2118 4894
rect 2152 4860 2200 4894
rect 2070 4850 2200 4860
rect 2070 4813 2100 4850
rect 2170 4813 2200 4850
rect 2270 4920 2300 5097
rect 2370 4920 2400 5097
rect 2270 4910 2400 4920
rect 2270 4876 2318 4910
rect 2352 4876 2400 4910
rect 2270 4866 2400 4876
rect 2270 4813 2300 4866
rect 2370 4813 2400 4866
rect 2470 4904 2500 5097
rect 2570 4904 2600 5097
rect 2470 4894 2600 4904
rect 2470 4860 2518 4894
rect 2552 4860 2600 4894
rect 2470 4850 2600 4860
rect 2470 4813 2500 4850
rect 2570 4813 2600 4850
rect 2670 4920 2700 5097
rect 2770 4920 2800 5097
rect 2670 4910 2800 4920
rect 2670 4876 2718 4910
rect 2752 4876 2800 4910
rect 2670 4866 2800 4876
rect 2670 4813 2700 4866
rect 2770 4813 2800 4866
rect 2870 4904 2900 5097
rect 2970 4904 3000 5097
rect 2870 4894 3000 4904
rect 2870 4860 2918 4894
rect 2952 4860 3000 4894
rect 2870 4850 3000 4860
rect 1270 4673 1300 4727
rect 1370 4673 1400 4727
rect 1470 4673 1500 4727
rect 1570 4673 1600 4727
rect 1670 4673 1700 4727
rect 1770 4673 1800 4727
rect 70 4533 100 4587
rect 70 4393 100 4447
rect 170 4393 200 4587
rect 270 4533 300 4587
rect 370 4533 400 4587
rect 470 4533 500 4587
rect 570 4533 600 4587
rect 670 4533 700 4587
rect 770 4533 800 4587
rect 870 4533 900 4587
rect 970 4533 1000 4587
rect 1070 4533 1100 4587
rect 1170 4533 1200 4587
rect 1270 4533 1300 4587
rect 1370 4533 1400 4587
rect 1470 4533 1500 4587
rect 1570 4533 1600 4587
rect 270 4393 300 4447
rect 370 4393 400 4447
rect 70 4253 100 4307
rect 70 4113 100 4167
rect 170 4113 200 4307
rect 270 4253 300 4307
rect 270 4113 300 4167
rect 370 4113 400 4307
rect 470 4253 500 4447
rect 570 4393 600 4447
rect 670 4393 700 4447
rect 570 4253 600 4307
rect 670 4253 700 4307
rect 770 4253 800 4447
rect 870 4393 900 4447
rect 970 4393 1000 4447
rect 1070 4393 1100 4447
rect 1170 4393 1200 4447
rect 1270 4393 1300 4447
rect 1370 4393 1400 4447
rect 1470 4393 1500 4447
rect 1570 4393 1600 4447
rect 1670 4393 1700 4587
rect 1770 4533 1800 4587
rect 1870 4533 1900 4727
rect 1970 4673 2000 4727
rect 1970 4533 2000 4587
rect 2070 4533 2100 4727
rect 2170 4673 2200 4727
rect 2270 4673 2300 4727
rect 2370 4673 2400 4727
rect 2470 4673 2500 4727
rect 2570 4673 2600 4727
rect 2670 4673 2700 4727
rect 2770 4673 2800 4727
rect 2870 4673 2900 4850
rect 2970 4813 3000 4850
rect 3070 4920 3100 5097
rect 3170 4920 3200 5097
rect 3070 4910 3200 4920
rect 3070 4876 3118 4910
rect 3152 4876 3200 4910
rect 3070 4866 3200 4876
rect 3070 4813 3100 4866
rect 3170 4813 3200 4866
rect 3270 4904 3300 5097
rect 3370 4904 3400 5097
rect 3270 4894 3400 4904
rect 3270 4860 3318 4894
rect 3352 4860 3400 4894
rect 3270 4850 3400 4860
rect 3270 4813 3300 4850
rect 3370 4813 3400 4850
rect 3470 4920 3500 5097
rect 3570 4920 3600 5097
rect 3470 4910 3600 4920
rect 3470 4876 3518 4910
rect 3552 4876 3600 4910
rect 3470 4866 3600 4876
rect 3470 4813 3500 4866
rect 3570 4813 3600 4866
rect 3670 4904 3700 5097
rect 3770 4904 3800 5097
rect 3670 4894 3800 4904
rect 3670 4860 3718 4894
rect 3752 4860 3800 4894
rect 3670 4850 3800 4860
rect 3670 4813 3700 4850
rect 3770 4813 3800 4850
rect 3870 4920 3900 5097
rect 3970 4920 4000 5097
rect 3870 4910 4000 4920
rect 3870 4876 3918 4910
rect 3952 4876 4000 4910
rect 3870 4866 4000 4876
rect 3870 4813 3900 4866
rect 3970 4813 4000 4866
rect 4070 4904 4100 5097
rect 4170 4904 4200 5097
rect 4070 4894 4200 4904
rect 4070 4860 4118 4894
rect 4152 4860 4200 4894
rect 4070 4850 4200 4860
rect 4070 4813 4100 4850
rect 4170 4813 4200 4850
rect 4270 4920 4300 5097
rect 4370 4920 4400 5237
rect 4470 5183 4500 5237
rect 4570 5183 4600 5237
rect 4670 5183 4700 5237
rect 4270 4910 4400 4920
rect 4270 4876 4318 4910
rect 4352 4876 4400 4910
rect 4270 4866 4400 4876
rect 4270 4813 4300 4866
rect 4370 4813 4400 4866
rect 4470 4904 4500 5097
rect 4570 4904 4600 5097
rect 4470 4894 4600 4904
rect 4470 4860 4518 4894
rect 4552 4860 4600 4894
rect 4470 4850 4600 4860
rect 4470 4813 4500 4850
rect 4570 4813 4600 4850
rect 4670 4920 4700 5097
rect 4770 4920 4800 5237
rect 4870 5183 4900 5237
rect 4970 5183 5000 5237
rect 5070 5183 5100 5237
rect 5170 5183 5200 5237
rect 5270 5183 5300 5377
rect 5370 5323 5400 5517
rect 5470 5463 5500 5517
rect 5370 5183 5400 5237
rect 5470 5183 5500 5377
rect 5570 5323 5600 5517
rect 5670 5463 5700 5517
rect 5670 5323 5700 5377
rect 5770 5323 5800 5517
rect 5870 5463 5900 5517
rect 5970 5463 6000 5517
rect 6070 5463 6100 5517
rect 6170 5463 6200 5517
rect 6270 5463 6300 5517
rect 6370 5463 6400 5517
rect 6570 5463 6600 5517
rect 6670 5463 6700 5517
rect 6880 5463 6910 5517
rect 6980 5463 7010 5517
rect 7080 5463 7110 5517
rect 7180 5463 7210 5517
rect 7280 5463 7310 5517
rect 7380 5463 7410 5517
rect 5870 5323 5900 5377
rect 5970 5323 6000 5377
rect 6070 5323 6100 5377
rect 6170 5323 6200 5377
rect 6270 5323 6300 5377
rect 6370 5323 6400 5377
rect 6570 5323 6600 5377
rect 6670 5323 6700 5377
rect 6880 5323 6910 5377
rect 6980 5323 7010 5377
rect 7080 5323 7110 5377
rect 7180 5323 7210 5377
rect 7280 5323 7310 5377
rect 7380 5323 7410 5377
rect 5570 5183 5600 5237
rect 5670 5183 5700 5237
rect 4670 4910 4800 4920
rect 4670 4876 4718 4910
rect 4752 4876 4800 4910
rect 4670 4866 4800 4876
rect 2970 4673 3000 4727
rect 3070 4673 3100 4727
rect 3170 4673 3200 4727
rect 2170 4533 2200 4587
rect 2270 4533 2300 4587
rect 2370 4533 2400 4587
rect 1770 4393 1800 4447
rect 1870 4393 1900 4447
rect 1970 4393 2000 4447
rect 2070 4393 2100 4447
rect 2170 4393 2200 4447
rect 2270 4393 2300 4447
rect 2370 4393 2400 4447
rect 870 4253 900 4307
rect 970 4253 1000 4307
rect 1070 4253 1100 4307
rect 1170 4253 1200 4307
rect 1270 4253 1300 4307
rect 1370 4253 1400 4307
rect 70 3973 100 4027
rect 170 3973 200 4027
rect 270 3973 300 4027
rect 370 3973 400 4027
rect 470 3973 500 4167
rect 570 4113 600 4167
rect 70 3833 100 3887
rect 170 3833 200 3887
rect 270 3833 300 3887
rect 370 3833 400 3887
rect 470 3833 500 3887
rect 570 3833 600 4027
rect 670 3973 700 4167
rect 770 4113 800 4167
rect 870 4113 900 4167
rect 970 4113 1000 4167
rect 1070 4113 1100 4167
rect 1170 4113 1200 4167
rect 1270 4113 1300 4167
rect 1370 4113 1400 4167
rect 1470 4113 1500 4307
rect 1570 4253 1600 4307
rect 1670 4253 1700 4307
rect 1770 4253 1800 4307
rect 1870 4253 1900 4307
rect 1970 4253 2000 4307
rect 2070 4253 2100 4307
rect 2170 4253 2200 4307
rect 2270 4253 2300 4307
rect 2370 4253 2400 4307
rect 2470 4253 2500 4587
rect 2570 4533 2600 4587
rect 2670 4533 2700 4587
rect 2770 4533 2800 4587
rect 2870 4533 2900 4587
rect 2970 4533 3000 4587
rect 3070 4533 3100 4587
rect 3170 4533 3200 4587
rect 3270 4533 3300 4727
rect 3370 4673 3400 4727
rect 3470 4673 3500 4727
rect 3570 4673 3600 4727
rect 3670 4673 3700 4727
rect 3770 4673 3800 4727
rect 3870 4673 3900 4727
rect 3970 4673 4000 4727
rect 4070 4673 4100 4727
rect 4170 4673 4200 4727
rect 4270 4673 4300 4727
rect 4370 4673 4400 4727
rect 4470 4673 4500 4727
rect 2570 4393 2600 4447
rect 2670 4393 2700 4447
rect 2770 4393 2800 4447
rect 2570 4253 2600 4307
rect 2670 4253 2700 4307
rect 2770 4253 2800 4307
rect 2870 4253 2900 4447
rect 2970 4393 3000 4447
rect 3070 4393 3100 4447
rect 3170 4393 3200 4447
rect 2970 4253 3000 4307
rect 3070 4253 3100 4307
rect 3170 4253 3200 4307
rect 3270 4253 3300 4447
rect 3370 4393 3400 4587
rect 3470 4533 3500 4587
rect 3570 4533 3600 4587
rect 3670 4533 3700 4587
rect 3770 4533 3800 4587
rect 3870 4533 3900 4587
rect 3970 4533 4000 4587
rect 4070 4533 4100 4587
rect 4170 4533 4200 4587
rect 4270 4533 4300 4587
rect 3470 4393 3500 4447
rect 3570 4393 3600 4447
rect 3670 4393 3700 4447
rect 3770 4393 3800 4447
rect 3870 4393 3900 4447
rect 3970 4393 4000 4447
rect 4070 4393 4100 4447
rect 4170 4393 4200 4447
rect 4270 4393 4300 4447
rect 4370 4393 4400 4587
rect 4470 4533 4500 4587
rect 4570 4533 4600 4727
rect 4670 4673 4700 4866
rect 4770 4813 4800 4866
rect 4870 4904 4900 5097
rect 4970 4904 5000 5097
rect 4870 4894 5000 4904
rect 4870 4860 4918 4894
rect 4952 4860 5000 4894
rect 4870 4850 5000 4860
rect 4870 4813 4900 4850
rect 4970 4813 5000 4850
rect 5070 4920 5100 5097
rect 5170 4920 5200 5097
rect 5070 4910 5200 4920
rect 5070 4876 5118 4910
rect 5152 4876 5200 4910
rect 5070 4866 5200 4876
rect 5070 4813 5100 4866
rect 5170 4813 5200 4866
rect 5270 4904 5300 5097
rect 5370 4904 5400 5097
rect 5270 4894 5400 4904
rect 5270 4860 5318 4894
rect 5352 4860 5400 4894
rect 5270 4850 5400 4860
rect 5270 4813 5300 4850
rect 5370 4813 5400 4850
rect 5470 4920 5500 5097
rect 5570 4920 5600 5097
rect 5470 4910 5600 4920
rect 5470 4876 5518 4910
rect 5552 4876 5600 4910
rect 5470 4866 5600 4876
rect 4770 4673 4800 4727
rect 4870 4673 4900 4727
rect 4970 4673 5000 4727
rect 5070 4673 5100 4727
rect 5170 4673 5200 4727
rect 5270 4673 5300 4727
rect 5370 4673 5400 4727
rect 5470 4673 5500 4866
rect 5570 4813 5600 4866
rect 5670 4904 5700 5097
rect 5770 4904 5800 5237
rect 5870 5183 5900 5237
rect 5970 5183 6000 5237
rect 6070 5183 6100 5237
rect 6170 5183 6200 5237
rect 6270 5183 6300 5237
rect 6370 5183 6400 5237
rect 6570 5183 6600 5237
rect 6670 5183 6700 5237
rect 6880 5183 6910 5237
rect 6980 5183 7010 5237
rect 7080 5183 7110 5237
rect 7180 5183 7210 5237
rect 7280 5183 7310 5237
rect 7380 5183 7410 5237
rect 5670 4894 5800 4904
rect 5670 4860 5718 4894
rect 5752 4860 5800 4894
rect 5670 4850 5800 4860
rect 5670 4813 5700 4850
rect 5770 4813 5800 4850
rect 5870 4920 5900 5097
rect 5970 4920 6000 5097
rect 5870 4910 6000 4920
rect 5870 4876 5918 4910
rect 5952 4876 6000 4910
rect 5870 4866 6000 4876
rect 5870 4813 5900 4866
rect 5570 4673 5600 4727
rect 5670 4673 5700 4727
rect 5770 4673 5800 4727
rect 5870 4673 5900 4727
rect 5970 4673 6000 4866
rect 6070 4904 6100 5097
rect 6170 4904 6200 5097
rect 6070 4894 6200 4904
rect 6070 4860 6118 4894
rect 6152 4860 6200 4894
rect 6070 4850 6200 4860
rect 6070 4813 6100 4850
rect 4670 4533 4700 4587
rect 4770 4533 4800 4587
rect 4870 4533 4900 4587
rect 4970 4533 5000 4587
rect 5070 4533 5100 4587
rect 5170 4533 5200 4587
rect 4470 4393 4500 4447
rect 4570 4393 4600 4447
rect 4670 4393 4700 4447
rect 4770 4393 4800 4447
rect 4870 4393 4900 4447
rect 4970 4393 5000 4447
rect 3370 4253 3400 4307
rect 770 3973 800 4027
rect 870 3973 900 4027
rect 970 3973 1000 4027
rect 1070 3973 1100 4027
rect 1170 3973 1200 4027
rect 1270 3973 1300 4027
rect 1370 3973 1400 4027
rect 1470 3973 1500 4027
rect 1570 3973 1600 4167
rect 1670 4113 1700 4167
rect 1670 3973 1700 4027
rect 1770 3973 1800 4167
rect 1870 4113 1900 4167
rect 1870 3973 1900 4027
rect 1970 3973 2000 4167
rect 2070 4113 2100 4167
rect 2170 4113 2200 4167
rect 2070 3973 2100 4027
rect 670 3833 700 3887
rect 770 3833 800 3887
rect 870 3833 900 3887
rect 970 3833 1000 3887
rect 1070 3833 1100 3887
rect 1170 3833 1200 3887
rect 70 3694 100 3747
rect 170 3694 200 3747
rect 70 3684 200 3694
rect 70 3650 118 3684
rect 152 3650 200 3684
rect 70 3640 200 3650
rect 70 3603 100 3640
rect 170 3603 200 3640
rect 270 3710 300 3747
rect 370 3710 400 3747
rect 270 3700 400 3710
rect 270 3666 318 3700
rect 352 3666 400 3700
rect 270 3656 400 3666
rect 70 3463 100 3517
rect 170 3463 200 3517
rect 270 3463 300 3656
rect 370 3603 400 3656
rect 470 3694 500 3747
rect 570 3694 600 3747
rect 470 3684 600 3694
rect 470 3650 518 3684
rect 552 3650 600 3684
rect 470 3640 600 3650
rect 470 3603 500 3640
rect 570 3603 600 3640
rect 670 3710 700 3747
rect 770 3710 800 3747
rect 670 3700 800 3710
rect 670 3666 718 3700
rect 752 3666 800 3700
rect 670 3656 800 3666
rect 670 3603 700 3656
rect 770 3603 800 3656
rect 870 3694 900 3747
rect 970 3694 1000 3747
rect 870 3684 1000 3694
rect 870 3650 918 3684
rect 952 3650 1000 3684
rect 870 3640 1000 3650
rect 870 3603 900 3640
rect 970 3603 1000 3640
rect 1070 3710 1100 3747
rect 1170 3710 1200 3747
rect 1070 3700 1200 3710
rect 1070 3666 1118 3700
rect 1152 3666 1200 3700
rect 1070 3656 1200 3666
rect 1070 3603 1100 3656
rect 1170 3603 1200 3656
rect 1270 3694 1300 3887
rect 1370 3833 1400 3887
rect 1370 3694 1400 3747
rect 1270 3684 1400 3694
rect 1270 3650 1318 3684
rect 1352 3650 1400 3684
rect 1270 3640 1400 3650
rect 1270 3603 1300 3640
rect 370 3463 400 3517
rect 470 3463 500 3517
rect 70 3323 100 3377
rect 170 3323 200 3377
rect 270 3323 300 3377
rect 370 3323 400 3377
rect 470 3323 500 3377
rect 570 3323 600 3517
rect 670 3463 700 3517
rect 670 3323 700 3377
rect 770 3323 800 3517
rect 870 3463 900 3517
rect 970 3463 1000 3517
rect 1070 3463 1100 3517
rect 1170 3463 1200 3517
rect 1270 3463 1300 3517
rect 1370 3463 1400 3640
rect 1470 3710 1500 3887
rect 1570 3833 1600 3887
rect 1670 3833 1700 3887
rect 1570 3710 1600 3747
rect 1470 3700 1600 3710
rect 1470 3666 1518 3700
rect 1552 3666 1600 3700
rect 1470 3656 1600 3666
rect 1470 3603 1500 3656
rect 1470 3463 1500 3517
rect 1570 3463 1600 3656
rect 1670 3694 1700 3747
rect 1770 3694 1800 3887
rect 1870 3833 1900 3887
rect 1970 3833 2000 3887
rect 2070 3833 2100 3887
rect 2170 3833 2200 4027
rect 2270 3973 2300 4167
rect 2370 4113 2400 4167
rect 2370 3973 2400 4027
rect 2470 3973 2500 4167
rect 2570 4113 2600 4167
rect 2670 4113 2700 4167
rect 2770 4113 2800 4167
rect 2870 4113 2900 4167
rect 2970 4113 3000 4167
rect 3070 4113 3100 4167
rect 3170 4113 3200 4167
rect 2570 3973 2600 4027
rect 2670 3973 2700 4027
rect 2770 3973 2800 4027
rect 2870 3973 2900 4027
rect 2970 3973 3000 4027
rect 3070 3973 3100 4027
rect 3170 3973 3200 4027
rect 2270 3833 2300 3887
rect 2370 3833 2400 3887
rect 2470 3833 2500 3887
rect 2570 3833 2600 3887
rect 2670 3833 2700 3887
rect 2770 3833 2800 3887
rect 2870 3833 2900 3887
rect 2970 3833 3000 3887
rect 3070 3833 3100 3887
rect 3170 3833 3200 3887
rect 3270 3833 3300 4167
rect 3370 4113 3400 4167
rect 3370 3973 3400 4027
rect 3470 3973 3500 4307
rect 3570 4253 3600 4307
rect 3570 4113 3600 4167
rect 3670 4113 3700 4307
rect 3770 4253 3800 4307
rect 3870 4253 3900 4307
rect 3970 4253 4000 4307
rect 4070 4253 4100 4307
rect 4170 4253 4200 4307
rect 4270 4253 4300 4307
rect 4370 4253 4400 4307
rect 3770 4113 3800 4167
rect 3870 4113 3900 4167
rect 3970 4113 4000 4167
rect 4070 4113 4100 4167
rect 4170 4113 4200 4167
rect 4270 4113 4300 4167
rect 4370 4113 4400 4167
rect 4470 4113 4500 4307
rect 4570 4253 4600 4307
rect 4670 4253 4700 4307
rect 4770 4253 4800 4307
rect 4870 4253 4900 4307
rect 4970 4253 5000 4307
rect 4570 4113 4600 4167
rect 4670 4113 4700 4167
rect 3570 3973 3600 4027
rect 3670 3973 3700 4027
rect 3770 3973 3800 4027
rect 3870 3973 3900 4027
rect 3970 3973 4000 4027
rect 4070 3973 4100 4027
rect 3370 3833 3400 3887
rect 1670 3684 1800 3694
rect 1670 3650 1718 3684
rect 1752 3650 1800 3684
rect 1670 3640 1800 3650
rect 1670 3603 1700 3640
rect 1770 3603 1800 3640
rect 1870 3710 1900 3747
rect 1970 3710 2000 3747
rect 1870 3700 2000 3710
rect 1870 3666 1918 3700
rect 1952 3666 2000 3700
rect 1870 3656 2000 3666
rect 1870 3603 1900 3656
rect 1970 3603 2000 3656
rect 2070 3694 2100 3747
rect 2170 3694 2200 3747
rect 2070 3684 2200 3694
rect 2070 3650 2118 3684
rect 2152 3650 2200 3684
rect 2070 3640 2200 3650
rect 2070 3603 2100 3640
rect 2170 3603 2200 3640
rect 2270 3710 2300 3747
rect 2370 3710 2400 3747
rect 2270 3700 2400 3710
rect 2270 3666 2318 3700
rect 2352 3666 2400 3700
rect 2270 3656 2400 3666
rect 1670 3463 1700 3517
rect 1770 3463 1800 3517
rect 1870 3463 1900 3517
rect 870 3323 900 3377
rect 970 3323 1000 3377
rect 1070 3323 1100 3377
rect 1170 3323 1200 3377
rect 70 3183 100 3237
rect 170 3183 200 3237
rect 270 3183 300 3237
rect 370 3183 400 3237
rect 70 3043 100 3097
rect 170 3043 200 3097
rect 270 3043 300 3097
rect 370 3043 400 3097
rect 470 3043 500 3237
rect 570 3183 600 3237
rect 670 3183 700 3237
rect 770 3183 800 3237
rect 870 3183 900 3237
rect 970 3183 1000 3237
rect 1070 3183 1100 3237
rect 570 3043 600 3097
rect 670 3043 700 3097
rect 770 3043 800 3097
rect 870 3043 900 3097
rect 970 3043 1000 3097
rect 1070 3043 1100 3097
rect 1170 3043 1200 3237
rect 1270 3183 1300 3377
rect 1370 3323 1400 3377
rect 1470 3323 1500 3377
rect 1570 3323 1600 3377
rect 1670 3323 1700 3377
rect 1770 3323 1800 3377
rect 1870 3323 1900 3377
rect 1970 3323 2000 3517
rect 2070 3463 2100 3517
rect 2170 3463 2200 3517
rect 2270 3463 2300 3656
rect 2370 3603 2400 3656
rect 2470 3694 2500 3747
rect 2570 3694 2600 3747
rect 2470 3684 2600 3694
rect 2470 3650 2518 3684
rect 2552 3650 2600 3684
rect 2470 3640 2600 3650
rect 2470 3603 2500 3640
rect 2570 3603 2600 3640
rect 2670 3710 2700 3747
rect 2770 3710 2800 3747
rect 2670 3700 2800 3710
rect 2670 3666 2718 3700
rect 2752 3666 2800 3700
rect 2670 3656 2800 3666
rect 2670 3603 2700 3656
rect 2770 3603 2800 3656
rect 2870 3694 2900 3747
rect 2970 3694 3000 3747
rect 2870 3684 3000 3694
rect 2870 3650 2918 3684
rect 2952 3650 3000 3684
rect 2870 3640 3000 3650
rect 2870 3603 2900 3640
rect 2970 3603 3000 3640
rect 3070 3710 3100 3747
rect 3170 3710 3200 3747
rect 3070 3700 3200 3710
rect 3070 3666 3118 3700
rect 3152 3666 3200 3700
rect 3070 3656 3200 3666
rect 3070 3603 3100 3656
rect 3170 3603 3200 3656
rect 3270 3694 3300 3747
rect 3370 3694 3400 3747
rect 3270 3684 3400 3694
rect 3270 3650 3318 3684
rect 3352 3650 3400 3684
rect 3270 3640 3400 3650
rect 3270 3603 3300 3640
rect 3370 3603 3400 3640
rect 3470 3710 3500 3887
rect 3570 3833 3600 3887
rect 3670 3833 3700 3887
rect 3770 3833 3800 3887
rect 3870 3833 3900 3887
rect 3970 3833 4000 3887
rect 4070 3833 4100 3887
rect 4170 3833 4200 4027
rect 4270 3973 4300 4027
rect 4370 3973 4400 4027
rect 4470 3973 4500 4027
rect 4270 3833 4300 3887
rect 4370 3833 4400 3887
rect 4470 3833 4500 3887
rect 4570 3833 4600 4027
rect 4670 3973 4700 4027
rect 4770 3973 4800 4167
rect 4870 4113 4900 4167
rect 4970 4113 5000 4167
rect 5070 4113 5100 4447
rect 5170 4393 5200 4447
rect 5270 4393 5300 4587
rect 5370 4533 5400 4587
rect 5470 4533 5500 4587
rect 5570 4533 5600 4587
rect 5670 4533 5700 4587
rect 5370 4393 5400 4447
rect 5170 4253 5200 4307
rect 5270 4253 5300 4307
rect 5370 4253 5400 4307
rect 5170 4113 5200 4167
rect 5270 4113 5300 4167
rect 5370 4113 5400 4167
rect 5470 4113 5500 4447
rect 5570 4393 5600 4447
rect 5670 4393 5700 4447
rect 5770 4393 5800 4587
rect 5870 4533 5900 4587
rect 5970 4533 6000 4587
rect 6070 4533 6100 4727
rect 6170 4673 6200 4850
rect 6270 4920 6300 5097
rect 6370 4920 6400 5097
rect 6570 4924 6600 5097
rect 6670 4924 6700 5097
rect 6880 4924 6910 5097
rect 6980 4924 7010 5097
rect 7080 4924 7110 5097
rect 7180 4924 7210 5097
rect 7280 4924 7310 5097
rect 7380 4924 7410 5097
rect 6270 4910 6400 4920
rect 6270 4876 6318 4910
rect 6352 4876 6400 4910
rect 6270 4866 6400 4876
rect 6270 4813 6300 4866
rect 6370 4813 6400 4866
rect 6558 4908 6612 4924
rect 6558 4874 6568 4908
rect 6602 4874 6612 4908
rect 6558 4858 6612 4874
rect 6658 4908 6712 4924
rect 6658 4874 6668 4908
rect 6702 4874 6712 4908
rect 6658 4858 6712 4874
rect 6868 4908 6922 4924
rect 6868 4874 6878 4908
rect 6912 4874 6922 4908
rect 6868 4858 6922 4874
rect 6968 4908 7022 4924
rect 6968 4874 6978 4908
rect 7012 4874 7022 4908
rect 6968 4858 7022 4874
rect 7068 4908 7122 4924
rect 7068 4874 7078 4908
rect 7112 4874 7122 4908
rect 7068 4858 7122 4874
rect 7168 4908 7222 4924
rect 7168 4874 7178 4908
rect 7212 4874 7222 4908
rect 7168 4858 7222 4874
rect 7268 4908 7322 4924
rect 7268 4874 7278 4908
rect 7312 4874 7322 4908
rect 7268 4858 7322 4874
rect 7368 4908 7422 4924
rect 7368 4874 7378 4908
rect 7412 4874 7422 4908
rect 7368 4858 7422 4874
rect 6570 4813 6600 4858
rect 6670 4813 6700 4858
rect 6880 4813 6910 4858
rect 6980 4813 7010 4858
rect 7080 4813 7110 4858
rect 7180 4813 7210 4858
rect 7280 4813 7310 4858
rect 7380 4813 7410 4858
rect 6170 4533 6200 4587
rect 5870 4393 5900 4447
rect 5970 4393 6000 4447
rect 5570 4253 5600 4307
rect 5670 4253 5700 4307
rect 5770 4253 5800 4307
rect 5570 4113 5600 4167
rect 4870 3973 4900 4027
rect 4970 3973 5000 4027
rect 5070 3973 5100 4027
rect 5170 3973 5200 4027
rect 5270 3973 5300 4027
rect 5370 3973 5400 4027
rect 5470 3973 5500 4027
rect 5570 3973 5600 4027
rect 5670 3973 5700 4167
rect 5770 4113 5800 4167
rect 5870 4113 5900 4307
rect 5970 4253 6000 4307
rect 6070 4253 6100 4447
rect 6170 4393 6200 4447
rect 6170 4253 6200 4307
rect 6270 4253 6300 4727
rect 6370 4673 6400 4727
rect 6570 4673 6600 4727
rect 6670 4673 6700 4727
rect 6880 4673 6910 4727
rect 6980 4673 7010 4727
rect 7080 4673 7110 4727
rect 7180 4673 7210 4727
rect 7280 4673 7310 4727
rect 7380 4673 7410 4727
rect 6370 4533 6400 4587
rect 6570 4533 6600 4587
rect 6670 4533 6700 4587
rect 6880 4533 6910 4587
rect 6980 4533 7010 4587
rect 7080 4533 7110 4587
rect 7180 4533 7210 4587
rect 7280 4533 7310 4587
rect 7380 4533 7410 4587
rect 6370 4393 6400 4447
rect 6570 4393 6600 4447
rect 6670 4393 6700 4447
rect 6880 4393 6910 4447
rect 6980 4393 7010 4447
rect 7080 4393 7110 4447
rect 7180 4393 7210 4447
rect 7280 4393 7310 4447
rect 7380 4393 7410 4447
rect 6370 4253 6400 4307
rect 6570 4253 6600 4307
rect 6670 4253 6700 4307
rect 6880 4253 6910 4307
rect 6980 4253 7010 4307
rect 7080 4253 7110 4307
rect 7180 4253 7210 4307
rect 7280 4253 7310 4307
rect 7380 4253 7410 4307
rect 5970 4113 6000 4167
rect 6070 4113 6100 4167
rect 6170 4113 6200 4167
rect 6270 4113 6300 4167
rect 6370 4113 6400 4167
rect 6570 4113 6600 4167
rect 6670 4113 6700 4167
rect 6880 4113 6910 4167
rect 6980 4113 7010 4167
rect 7080 4113 7110 4167
rect 7180 4113 7210 4167
rect 7280 4113 7310 4167
rect 7380 4113 7410 4167
rect 5770 3973 5800 4027
rect 5870 3973 5900 4027
rect 5970 3973 6000 4027
rect 4670 3833 4700 3887
rect 3570 3710 3600 3747
rect 3470 3700 3600 3710
rect 3470 3666 3518 3700
rect 3552 3666 3600 3700
rect 3470 3656 3600 3666
rect 3470 3603 3500 3656
rect 2370 3463 2400 3517
rect 2470 3463 2500 3517
rect 2570 3463 2600 3517
rect 2670 3463 2700 3517
rect 2770 3463 2800 3517
rect 2070 3323 2100 3377
rect 2170 3323 2200 3377
rect 2270 3323 2300 3377
rect 2370 3323 2400 3377
rect 2470 3323 2500 3377
rect 2570 3323 2600 3377
rect 2670 3323 2700 3377
rect 1370 3183 1400 3237
rect 1470 3183 1500 3237
rect 1570 3183 1600 3237
rect 1670 3183 1700 3237
rect 1770 3183 1800 3237
rect 1870 3183 1900 3237
rect 1970 3183 2000 3237
rect 2070 3183 2100 3237
rect 2170 3183 2200 3237
rect 2270 3183 2300 3237
rect 2370 3183 2400 3237
rect 1270 3043 1300 3097
rect 1370 3043 1400 3097
rect 1470 3043 1500 3097
rect 1570 3043 1600 3097
rect 1670 3043 1700 3097
rect 1770 3043 1800 3097
rect 1870 3043 1900 3097
rect 1970 3043 2000 3097
rect 2070 3043 2100 3097
rect 2170 3043 2200 3097
rect 2270 3043 2300 3097
rect 2370 3043 2400 3097
rect 2470 3043 2500 3237
rect 2570 3183 2600 3237
rect 2670 3183 2700 3237
rect 2770 3183 2800 3377
rect 2870 3323 2900 3517
rect 2970 3463 3000 3517
rect 3070 3463 3100 3517
rect 3170 3463 3200 3517
rect 3270 3463 3300 3517
rect 3370 3463 3400 3517
rect 3470 3463 3500 3517
rect 3570 3463 3600 3656
rect 3670 3694 3700 3747
rect 3770 3694 3800 3747
rect 3670 3684 3800 3694
rect 3670 3650 3718 3684
rect 3752 3650 3800 3684
rect 3670 3640 3800 3650
rect 3670 3603 3700 3640
rect 3670 3463 3700 3517
rect 3770 3463 3800 3640
rect 3870 3710 3900 3747
rect 3970 3710 4000 3747
rect 3870 3700 4000 3710
rect 3870 3666 3918 3700
rect 3952 3666 4000 3700
rect 3870 3656 4000 3666
rect 3870 3603 3900 3656
rect 3970 3603 4000 3656
rect 4070 3694 4100 3747
rect 4170 3694 4200 3747
rect 4070 3684 4200 3694
rect 4070 3650 4118 3684
rect 4152 3650 4200 3684
rect 4070 3640 4200 3650
rect 4070 3603 4100 3640
rect 4170 3603 4200 3640
rect 4270 3710 4300 3747
rect 4370 3710 4400 3747
rect 4270 3700 4400 3710
rect 4270 3666 4318 3700
rect 4352 3666 4400 3700
rect 4270 3656 4400 3666
rect 3870 3463 3900 3517
rect 3970 3463 4000 3517
rect 4070 3463 4100 3517
rect 4170 3463 4200 3517
rect 4270 3463 4300 3656
rect 4370 3603 4400 3656
rect 4470 3694 4500 3747
rect 4570 3694 4600 3747
rect 4470 3684 4600 3694
rect 4470 3650 4518 3684
rect 4552 3650 4600 3684
rect 4470 3640 4600 3650
rect 4470 3603 4500 3640
rect 4570 3603 4600 3640
rect 4670 3710 4700 3747
rect 4770 3710 4800 3887
rect 4870 3833 4900 3887
rect 4970 3833 5000 3887
rect 5070 3833 5100 3887
rect 5170 3833 5200 3887
rect 5270 3833 5300 3887
rect 5370 3833 5400 3887
rect 5470 3833 5500 3887
rect 5570 3833 5600 3887
rect 4670 3700 4800 3710
rect 4670 3666 4718 3700
rect 4752 3666 4800 3700
rect 4670 3656 4800 3666
rect 4670 3603 4700 3656
rect 4370 3463 4400 3517
rect 4470 3463 4500 3517
rect 4570 3463 4600 3517
rect 4670 3463 4700 3517
rect 4770 3463 4800 3656
rect 4870 3694 4900 3747
rect 4970 3694 5000 3747
rect 4870 3684 5000 3694
rect 4870 3650 4918 3684
rect 4952 3650 5000 3684
rect 4870 3640 5000 3650
rect 4870 3603 4900 3640
rect 4970 3603 5000 3640
rect 5070 3710 5100 3747
rect 5170 3710 5200 3747
rect 5070 3700 5200 3710
rect 5070 3666 5118 3700
rect 5152 3666 5200 3700
rect 5070 3656 5200 3666
rect 5070 3603 5100 3656
rect 5170 3603 5200 3656
rect 5270 3694 5300 3747
rect 5370 3694 5400 3747
rect 5270 3684 5400 3694
rect 5270 3650 5318 3684
rect 5352 3650 5400 3684
rect 5270 3640 5400 3650
rect 4870 3463 4900 3517
rect 4970 3463 5000 3517
rect 5070 3463 5100 3517
rect 5170 3463 5200 3517
rect 5270 3463 5300 3640
rect 5370 3603 5400 3640
rect 5470 3710 5500 3747
rect 5570 3710 5600 3747
rect 5470 3700 5600 3710
rect 5470 3666 5518 3700
rect 5552 3666 5600 3700
rect 5470 3656 5600 3666
rect 5470 3603 5500 3656
rect 5570 3603 5600 3656
rect 5670 3694 5700 3887
rect 5770 3833 5800 3887
rect 5870 3833 5900 3887
rect 5970 3833 6000 3887
rect 6070 3833 6100 4027
rect 6170 3973 6200 4027
rect 6270 3973 6300 4027
rect 6370 3973 6400 4027
rect 6570 3973 6600 4027
rect 6670 3973 6700 4027
rect 6880 3973 6910 4027
rect 6980 3973 7010 4027
rect 7080 3973 7110 4027
rect 7180 3973 7210 4027
rect 7280 3973 7310 4027
rect 7380 3973 7410 4027
rect 6170 3833 6200 3887
rect 6270 3833 6300 3887
rect 6370 3833 6400 3887
rect 6570 3833 6600 3887
rect 6670 3833 6700 3887
rect 6880 3833 6910 3887
rect 6980 3833 7010 3887
rect 7080 3833 7110 3887
rect 7180 3833 7210 3887
rect 7280 3833 7310 3887
rect 7380 3833 7410 3887
rect 5770 3694 5800 3747
rect 5670 3684 5800 3694
rect 5670 3650 5718 3684
rect 5752 3650 5800 3684
rect 5670 3640 5800 3650
rect 5670 3603 5700 3640
rect 5770 3603 5800 3640
rect 5870 3710 5900 3747
rect 5970 3710 6000 3747
rect 5870 3700 6000 3710
rect 5870 3666 5918 3700
rect 5952 3666 6000 3700
rect 5870 3656 6000 3666
rect 5870 3603 5900 3656
rect 5970 3603 6000 3656
rect 6070 3694 6100 3747
rect 6170 3694 6200 3747
rect 6070 3684 6200 3694
rect 6070 3650 6118 3684
rect 6152 3650 6200 3684
rect 6070 3640 6200 3650
rect 6070 3603 6100 3640
rect 6170 3603 6200 3640
rect 6270 3710 6300 3747
rect 6370 3710 6400 3747
rect 6570 3714 6600 3747
rect 6670 3714 6700 3747
rect 6880 3714 6910 3747
rect 6980 3714 7010 3747
rect 7080 3714 7110 3747
rect 7180 3714 7210 3747
rect 7280 3714 7310 3747
rect 7380 3714 7410 3747
rect 6270 3700 6400 3710
rect 6270 3666 6318 3700
rect 6352 3666 6400 3700
rect 6270 3656 6400 3666
rect 6270 3603 6300 3656
rect 6370 3603 6400 3656
rect 6558 3698 6612 3714
rect 6558 3664 6568 3698
rect 6602 3664 6612 3698
rect 6558 3648 6612 3664
rect 6658 3698 6712 3714
rect 6658 3664 6668 3698
rect 6702 3664 6712 3698
rect 6658 3648 6712 3664
rect 6868 3698 6922 3714
rect 6868 3664 6878 3698
rect 6912 3664 6922 3698
rect 6868 3648 6922 3664
rect 6968 3698 7022 3714
rect 6968 3664 6978 3698
rect 7012 3664 7022 3698
rect 6968 3648 7022 3664
rect 7068 3698 7122 3714
rect 7068 3664 7078 3698
rect 7112 3664 7122 3698
rect 7068 3648 7122 3664
rect 7168 3698 7222 3714
rect 7168 3664 7178 3698
rect 7212 3664 7222 3698
rect 7168 3648 7222 3664
rect 7268 3698 7322 3714
rect 7268 3664 7278 3698
rect 7312 3664 7322 3698
rect 7268 3648 7322 3664
rect 7368 3698 7422 3714
rect 7368 3664 7378 3698
rect 7412 3664 7422 3698
rect 7368 3648 7422 3664
rect 6570 3603 6600 3648
rect 6670 3603 6700 3648
rect 6880 3603 6910 3648
rect 6980 3603 7010 3648
rect 7080 3603 7110 3648
rect 7180 3603 7210 3648
rect 7280 3603 7310 3648
rect 7380 3603 7410 3648
rect 5370 3463 5400 3517
rect 5470 3463 5500 3517
rect 5570 3463 5600 3517
rect 5670 3463 5700 3517
rect 5770 3463 5800 3517
rect 5870 3463 5900 3517
rect 2870 3183 2900 3237
rect 2970 3183 3000 3377
rect 3070 3323 3100 3377
rect 3170 3323 3200 3377
rect 3270 3323 3300 3377
rect 3370 3323 3400 3377
rect 3470 3323 3500 3377
rect 3570 3323 3600 3377
rect 3670 3323 3700 3377
rect 3770 3323 3800 3377
rect 3870 3323 3900 3377
rect 3970 3323 4000 3377
rect 4070 3323 4100 3377
rect 4170 3323 4200 3377
rect 4270 3323 4300 3377
rect 3070 3183 3100 3237
rect 3170 3183 3200 3237
rect 2570 3043 2600 3097
rect 2670 3043 2700 3097
rect 2770 3043 2800 3097
rect 2870 3043 2900 3097
rect 2970 3043 3000 3097
rect 3070 3043 3100 3097
rect 3170 3043 3200 3097
rect 3270 3043 3300 3237
rect 3370 3183 3400 3237
rect 3470 3183 3500 3237
rect 3570 3183 3600 3237
rect 70 2903 100 2957
rect 170 2903 200 2957
rect 270 2903 300 2957
rect 70 2763 100 2817
rect 170 2763 200 2817
rect 270 2763 300 2817
rect 370 2763 400 2957
rect 470 2903 500 2957
rect 570 2903 600 2957
rect 670 2903 700 2957
rect 470 2763 500 2817
rect 570 2763 600 2817
rect 670 2763 700 2817
rect 770 2763 800 2957
rect 870 2903 900 2957
rect 970 2903 1000 2957
rect 1070 2903 1100 2957
rect 1170 2903 1200 2957
rect 1270 2903 1300 2957
rect 1370 2903 1400 2957
rect 870 2763 900 2817
rect 970 2763 1000 2817
rect 1070 2763 1100 2817
rect 1170 2763 1200 2817
rect 1270 2763 1300 2817
rect 70 2623 100 2677
rect 170 2623 200 2677
rect 270 2623 300 2677
rect 370 2623 400 2677
rect 470 2623 500 2677
rect 570 2623 600 2677
rect 670 2623 700 2677
rect 770 2623 800 2677
rect 870 2623 900 2677
rect 970 2623 1000 2677
rect 1070 2623 1100 2677
rect 1170 2623 1200 2677
rect 1270 2623 1300 2677
rect 1370 2623 1400 2817
rect 1470 2763 1500 2957
rect 1570 2903 1600 2957
rect 1670 2903 1700 2957
rect 1770 2903 1800 2957
rect 1870 2903 1900 2957
rect 1970 2903 2000 2957
rect 2070 2903 2100 2957
rect 1470 2623 1500 2677
rect 70 2484 100 2537
rect 170 2484 200 2537
rect 70 2474 200 2484
rect 70 2440 118 2474
rect 152 2440 200 2474
rect 70 2430 200 2440
rect 70 2393 100 2430
rect 170 2393 200 2430
rect 270 2500 300 2537
rect 370 2500 400 2537
rect 270 2490 400 2500
rect 270 2456 318 2490
rect 352 2456 400 2490
rect 270 2446 400 2456
rect 270 2393 300 2446
rect 370 2393 400 2446
rect 470 2484 500 2537
rect 570 2484 600 2537
rect 470 2474 600 2484
rect 470 2440 518 2474
rect 552 2440 600 2474
rect 470 2430 600 2440
rect 470 2393 500 2430
rect 570 2393 600 2430
rect 670 2500 700 2537
rect 770 2500 800 2537
rect 670 2490 800 2500
rect 670 2456 718 2490
rect 752 2456 800 2490
rect 670 2446 800 2456
rect 670 2393 700 2446
rect 770 2393 800 2446
rect 870 2484 900 2537
rect 970 2484 1000 2537
rect 870 2474 1000 2484
rect 870 2440 918 2474
rect 952 2440 1000 2474
rect 870 2430 1000 2440
rect 870 2393 900 2430
rect 970 2393 1000 2430
rect 1070 2500 1100 2537
rect 1170 2500 1200 2537
rect 1070 2490 1200 2500
rect 1070 2456 1118 2490
rect 1152 2456 1200 2490
rect 1070 2446 1200 2456
rect 1070 2393 1100 2446
rect 1170 2393 1200 2446
rect 1270 2484 1300 2537
rect 1370 2484 1400 2537
rect 1270 2474 1400 2484
rect 1270 2440 1318 2474
rect 1352 2440 1400 2474
rect 1270 2430 1400 2440
rect 1270 2393 1300 2430
rect 1370 2393 1400 2430
rect 1470 2500 1500 2537
rect 1570 2500 1600 2817
rect 1670 2763 1700 2817
rect 1770 2763 1800 2817
rect 1870 2763 1900 2817
rect 1970 2763 2000 2817
rect 1670 2623 1700 2677
rect 1770 2623 1800 2677
rect 1870 2623 1900 2677
rect 1970 2623 2000 2677
rect 2070 2623 2100 2817
rect 2170 2763 2200 2957
rect 2270 2903 2300 2957
rect 2270 2763 2300 2817
rect 2370 2763 2400 2957
rect 2470 2903 2500 2957
rect 2470 2763 2500 2817
rect 2570 2763 2600 2957
rect 2670 2903 2700 2957
rect 2770 2903 2800 2957
rect 2870 2903 2900 2957
rect 2970 2903 3000 2957
rect 2670 2763 2700 2817
rect 2770 2763 2800 2817
rect 1470 2490 1600 2500
rect 1470 2456 1518 2490
rect 1552 2456 1600 2490
rect 1470 2446 1600 2456
rect 1470 2393 1500 2446
rect 1570 2393 1600 2446
rect 1670 2484 1700 2537
rect 1770 2484 1800 2537
rect 1670 2474 1800 2484
rect 1670 2440 1718 2474
rect 1752 2440 1800 2474
rect 1670 2430 1800 2440
rect 1670 2393 1700 2430
rect 1770 2393 1800 2430
rect 1870 2500 1900 2537
rect 1970 2500 2000 2537
rect 1870 2490 2000 2500
rect 1870 2456 1918 2490
rect 1952 2456 2000 2490
rect 1870 2446 2000 2456
rect 1870 2393 1900 2446
rect 1970 2393 2000 2446
rect 2070 2484 2100 2537
rect 2170 2484 2200 2677
rect 2270 2623 2300 2677
rect 2370 2623 2400 2677
rect 2070 2474 2200 2484
rect 2070 2440 2118 2474
rect 2152 2440 2200 2474
rect 2070 2430 2200 2440
rect 2070 2393 2100 2430
rect 2170 2393 2200 2430
rect 2270 2500 2300 2537
rect 2370 2500 2400 2537
rect 2270 2490 2400 2500
rect 2270 2456 2318 2490
rect 2352 2456 2400 2490
rect 2270 2446 2400 2456
rect 2270 2393 2300 2446
rect 2370 2393 2400 2446
rect 2470 2484 2500 2677
rect 2570 2623 2600 2677
rect 2570 2484 2600 2537
rect 2470 2474 2600 2484
rect 2470 2440 2518 2474
rect 2552 2440 2600 2474
rect 2470 2430 2600 2440
rect 2470 2393 2500 2430
rect 2570 2393 2600 2430
rect 2670 2500 2700 2677
rect 2770 2623 2800 2677
rect 2870 2623 2900 2817
rect 2970 2763 3000 2817
rect 3070 2763 3100 2957
rect 3170 2903 3200 2957
rect 3270 2903 3300 2957
rect 3370 2903 3400 3097
rect 3470 3043 3500 3097
rect 3570 3043 3600 3097
rect 3670 3043 3700 3237
rect 3770 3183 3800 3237
rect 3870 3183 3900 3237
rect 3970 3183 4000 3237
rect 4070 3183 4100 3237
rect 4170 3183 4200 3237
rect 3770 3043 3800 3097
rect 3470 2903 3500 2957
rect 3570 2903 3600 2957
rect 3670 2903 3700 2957
rect 3770 2903 3800 2957
rect 3870 2903 3900 3097
rect 3970 3043 4000 3097
rect 3970 2903 4000 2957
rect 4070 2903 4100 3097
rect 4170 3043 4200 3097
rect 4270 3043 4300 3237
rect 4370 3183 4400 3377
rect 4470 3323 4500 3377
rect 4570 3323 4600 3377
rect 4670 3323 4700 3377
rect 4770 3323 4800 3377
rect 4470 3183 4500 3237
rect 4370 3043 4400 3097
rect 4470 3043 4500 3097
rect 4170 2903 4200 2957
rect 4270 2903 4300 2957
rect 4370 2903 4400 2957
rect 4470 2903 4500 2957
rect 4570 2903 4600 3237
rect 4670 3183 4700 3237
rect 4670 3043 4700 3097
rect 4770 3043 4800 3237
rect 4870 3183 4900 3377
rect 4970 3323 5000 3377
rect 5070 3323 5100 3377
rect 5170 3323 5200 3377
rect 5270 3323 5300 3377
rect 5370 3323 5400 3377
rect 5470 3323 5500 3377
rect 4970 3183 5000 3237
rect 4870 3043 4900 3097
rect 4970 3043 5000 3097
rect 5070 3043 5100 3237
rect 5170 3183 5200 3237
rect 5270 3183 5300 3237
rect 5370 3183 5400 3237
rect 5470 3183 5500 3237
rect 5170 3043 5200 3097
rect 5270 3043 5300 3097
rect 5370 3043 5400 3097
rect 5470 3043 5500 3097
rect 5570 3043 5600 3377
rect 5670 3323 5700 3377
rect 5770 3323 5800 3377
rect 5870 3323 5900 3377
rect 5970 3323 6000 3517
rect 6070 3463 6100 3517
rect 6170 3463 6200 3517
rect 6270 3463 6300 3517
rect 6370 3463 6400 3517
rect 6570 3463 6600 3517
rect 6670 3463 6700 3517
rect 6880 3463 6910 3517
rect 6980 3463 7010 3517
rect 7080 3463 7110 3517
rect 7180 3463 7210 3517
rect 7280 3463 7310 3517
rect 7380 3463 7410 3517
rect 6070 3323 6100 3377
rect 6170 3323 6200 3377
rect 6270 3323 6300 3377
rect 6370 3323 6400 3377
rect 6570 3323 6600 3377
rect 6670 3323 6700 3377
rect 6880 3323 6910 3377
rect 6980 3323 7010 3377
rect 7080 3323 7110 3377
rect 7180 3323 7210 3377
rect 7280 3323 7310 3377
rect 7380 3323 7410 3377
rect 5670 3183 5700 3237
rect 5670 3043 5700 3097
rect 5770 3043 5800 3237
rect 5870 3183 5900 3237
rect 5970 3183 6000 3237
rect 6070 3183 6100 3237
rect 6170 3183 6200 3237
rect 6270 3183 6300 3237
rect 6370 3183 6400 3237
rect 6570 3183 6600 3237
rect 6670 3183 6700 3237
rect 6880 3183 6910 3237
rect 6980 3183 7010 3237
rect 7080 3183 7110 3237
rect 7180 3183 7210 3237
rect 7280 3183 7310 3237
rect 7380 3183 7410 3237
rect 5870 3043 5900 3097
rect 4670 2903 4700 2957
rect 4770 2903 4800 2957
rect 4870 2903 4900 2957
rect 4970 2903 5000 2957
rect 5070 2903 5100 2957
rect 5170 2903 5200 2957
rect 5270 2903 5300 2957
rect 5370 2903 5400 2957
rect 5470 2903 5500 2957
rect 5570 2903 5600 2957
rect 5670 2903 5700 2957
rect 5770 2903 5800 2957
rect 5870 2903 5900 2957
rect 5970 2903 6000 3097
rect 6070 3043 6100 3097
rect 6170 3043 6200 3097
rect 6270 3043 6300 3097
rect 6370 3043 6400 3097
rect 6570 3043 6600 3097
rect 6670 3043 6700 3097
rect 6880 3043 6910 3097
rect 6980 3043 7010 3097
rect 7080 3043 7110 3097
rect 7180 3043 7210 3097
rect 7280 3043 7310 3097
rect 7380 3043 7410 3097
rect 2970 2623 3000 2677
rect 3070 2623 3100 2677
rect 3170 2623 3200 2817
rect 3270 2763 3300 2817
rect 3370 2763 3400 2817
rect 3470 2763 3500 2817
rect 3570 2763 3600 2817
rect 3670 2763 3700 2817
rect 3770 2763 3800 2817
rect 3870 2763 3900 2817
rect 3970 2763 4000 2817
rect 4070 2763 4100 2817
rect 4170 2763 4200 2817
rect 4270 2763 4300 2817
rect 4370 2763 4400 2817
rect 2770 2500 2800 2537
rect 2670 2490 2800 2500
rect 2670 2456 2718 2490
rect 2752 2456 2800 2490
rect 2670 2446 2800 2456
rect 2670 2393 2700 2446
rect 2770 2393 2800 2446
rect 2870 2484 2900 2537
rect 2970 2484 3000 2537
rect 2870 2474 3000 2484
rect 2870 2440 2918 2474
rect 2952 2440 3000 2474
rect 2870 2430 3000 2440
rect 2870 2393 2900 2430
rect 2970 2393 3000 2430
rect 3070 2500 3100 2537
rect 3170 2500 3200 2537
rect 3070 2490 3200 2500
rect 3070 2456 3118 2490
rect 3152 2456 3200 2490
rect 3070 2446 3200 2456
rect 3070 2393 3100 2446
rect 3170 2393 3200 2446
rect 3270 2484 3300 2677
rect 3370 2623 3400 2677
rect 3370 2484 3400 2537
rect 3270 2474 3400 2484
rect 3270 2440 3318 2474
rect 3352 2440 3400 2474
rect 3270 2430 3400 2440
rect 3270 2393 3300 2430
rect 3370 2393 3400 2430
rect 3470 2500 3500 2677
rect 3570 2623 3600 2677
rect 3670 2623 3700 2677
rect 3770 2623 3800 2677
rect 3870 2623 3900 2677
rect 3970 2623 4000 2677
rect 4070 2623 4100 2677
rect 4170 2623 4200 2677
rect 4270 2623 4300 2677
rect 4370 2623 4400 2677
rect 4470 2623 4500 2817
rect 4570 2763 4600 2817
rect 4570 2623 4600 2677
rect 4670 2623 4700 2817
rect 4770 2763 4800 2817
rect 4870 2763 4900 2817
rect 4970 2763 5000 2817
rect 5070 2763 5100 2817
rect 5170 2763 5200 2817
rect 5270 2763 5300 2817
rect 5370 2763 5400 2817
rect 4770 2623 4800 2677
rect 4870 2623 4900 2677
rect 4970 2623 5000 2677
rect 5070 2623 5100 2677
rect 5170 2623 5200 2677
rect 5270 2623 5300 2677
rect 5370 2623 5400 2677
rect 5470 2623 5500 2817
rect 5570 2763 5600 2817
rect 5670 2763 5700 2817
rect 5770 2763 5800 2817
rect 5870 2763 5900 2817
rect 5970 2763 6000 2817
rect 6070 2763 6100 2957
rect 6170 2903 6200 2957
rect 6270 2903 6300 2957
rect 6370 2903 6400 2957
rect 6570 2903 6600 2957
rect 6670 2903 6700 2957
rect 6880 2903 6910 2957
rect 6980 2903 7010 2957
rect 7080 2903 7110 2957
rect 7180 2903 7210 2957
rect 7280 2903 7310 2957
rect 7380 2903 7410 2957
rect 6170 2763 6200 2817
rect 6270 2763 6300 2817
rect 6370 2763 6400 2817
rect 6570 2763 6600 2817
rect 6670 2763 6700 2817
rect 6880 2763 6910 2817
rect 6980 2763 7010 2817
rect 7080 2763 7110 2817
rect 7180 2763 7210 2817
rect 7280 2763 7310 2817
rect 7380 2763 7410 2817
rect 3570 2500 3600 2537
rect 3470 2490 3600 2500
rect 3470 2456 3518 2490
rect 3552 2456 3600 2490
rect 3470 2446 3600 2456
rect 3470 2393 3500 2446
rect 3570 2393 3600 2446
rect 3670 2484 3700 2537
rect 3770 2484 3800 2537
rect 3670 2474 3800 2484
rect 3670 2440 3718 2474
rect 3752 2440 3800 2474
rect 3670 2430 3800 2440
rect 3670 2393 3700 2430
rect 3770 2393 3800 2430
rect 3870 2500 3900 2537
rect 3970 2500 4000 2537
rect 3870 2490 4000 2500
rect 3870 2456 3918 2490
rect 3952 2456 4000 2490
rect 3870 2446 4000 2456
rect 3870 2393 3900 2446
rect 3970 2393 4000 2446
rect 4070 2484 4100 2537
rect 4170 2484 4200 2537
rect 4070 2474 4200 2484
rect 4070 2440 4118 2474
rect 4152 2440 4200 2474
rect 4070 2430 4200 2440
rect 4070 2393 4100 2430
rect 4170 2393 4200 2430
rect 4270 2500 4300 2537
rect 4370 2500 4400 2537
rect 4270 2490 4400 2500
rect 4270 2456 4318 2490
rect 4352 2456 4400 2490
rect 4270 2446 4400 2456
rect 4270 2393 4300 2446
rect 4370 2393 4400 2446
rect 4470 2484 4500 2537
rect 4570 2484 4600 2537
rect 4470 2474 4600 2484
rect 4470 2440 4518 2474
rect 4552 2440 4600 2474
rect 4470 2430 4600 2440
rect 4470 2393 4500 2430
rect 4570 2393 4600 2430
rect 4670 2500 4700 2537
rect 4770 2500 4800 2537
rect 4670 2490 4800 2500
rect 4670 2456 4718 2490
rect 4752 2456 4800 2490
rect 4670 2446 4800 2456
rect 4670 2393 4700 2446
rect 4770 2393 4800 2446
rect 4870 2484 4900 2537
rect 4970 2484 5000 2537
rect 4870 2474 5000 2484
rect 4870 2440 4918 2474
rect 4952 2440 5000 2474
rect 4870 2430 5000 2440
rect 4870 2393 4900 2430
rect 4970 2393 5000 2430
rect 5070 2500 5100 2537
rect 5170 2500 5200 2537
rect 5070 2490 5200 2500
rect 5070 2456 5118 2490
rect 5152 2456 5200 2490
rect 5070 2446 5200 2456
rect 5070 2393 5100 2446
rect 5170 2393 5200 2446
rect 5270 2484 5300 2537
rect 5370 2484 5400 2537
rect 5270 2474 5400 2484
rect 5270 2440 5318 2474
rect 5352 2440 5400 2474
rect 5270 2430 5400 2440
rect 5270 2393 5300 2430
rect 5370 2393 5400 2430
rect 5470 2500 5500 2537
rect 5570 2500 5600 2677
rect 5670 2623 5700 2677
rect 5770 2623 5800 2677
rect 5870 2623 5900 2677
rect 5970 2623 6000 2677
rect 6070 2623 6100 2677
rect 6170 2623 6200 2677
rect 6270 2623 6300 2677
rect 6370 2623 6400 2677
rect 6570 2623 6600 2677
rect 6670 2623 6700 2677
rect 6880 2623 6910 2677
rect 6980 2623 7010 2677
rect 7080 2623 7110 2677
rect 7180 2623 7210 2677
rect 7280 2623 7310 2677
rect 7380 2623 7410 2677
rect 5470 2490 5600 2500
rect 5470 2456 5518 2490
rect 5552 2456 5600 2490
rect 5470 2446 5600 2456
rect 70 2253 100 2307
rect 170 2253 200 2307
rect 70 2113 100 2167
rect 170 2113 200 2167
rect 270 2113 300 2307
rect 370 2253 400 2307
rect 470 2253 500 2307
rect 570 2253 600 2307
rect 670 2253 700 2307
rect 770 2253 800 2307
rect 870 2253 900 2307
rect 970 2253 1000 2307
rect 1070 2253 1100 2307
rect 1170 2253 1200 2307
rect 1270 2253 1300 2307
rect 70 1973 100 2027
rect 170 1973 200 2027
rect 270 1973 300 2027
rect 70 1833 100 1887
rect 170 1833 200 1887
rect 270 1833 300 1887
rect 370 1833 400 2167
rect 470 2113 500 2167
rect 570 2113 600 2167
rect 670 2113 700 2167
rect 770 2113 800 2167
rect 870 2113 900 2167
rect 970 2113 1000 2167
rect 1070 2113 1100 2167
rect 1170 2113 1200 2167
rect 1270 2113 1300 2167
rect 470 1973 500 2027
rect 570 1973 600 2027
rect 670 1973 700 2027
rect 770 1973 800 2027
rect 870 1973 900 2027
rect 970 1973 1000 2027
rect 1070 1973 1100 2027
rect 1170 1973 1200 2027
rect 1270 1973 1300 2027
rect 1370 1973 1400 2307
rect 1470 2253 1500 2307
rect 1470 2113 1500 2167
rect 470 1833 500 1887
rect 570 1833 600 1887
rect 670 1833 700 1887
rect 770 1833 800 1887
rect 870 1833 900 1887
rect 70 1693 100 1747
rect 70 1553 100 1607
rect 70 1413 100 1467
rect 170 1413 200 1747
rect 270 1693 300 1747
rect 370 1693 400 1747
rect 470 1693 500 1747
rect 570 1693 600 1747
rect 670 1693 700 1747
rect 270 1553 300 1607
rect 370 1553 400 1607
rect 70 1274 100 1327
rect 170 1274 200 1327
rect 70 1264 200 1274
rect 70 1230 118 1264
rect 152 1230 200 1264
rect 70 1220 200 1230
rect 70 1183 100 1220
rect 170 1183 200 1220
rect 270 1290 300 1467
rect 370 1413 400 1467
rect 470 1413 500 1607
rect 570 1553 600 1607
rect 670 1553 700 1607
rect 770 1553 800 1747
rect 870 1693 900 1747
rect 870 1553 900 1607
rect 970 1553 1000 1887
rect 1070 1833 1100 1887
rect 1170 1833 1200 1887
rect 1270 1833 1300 1887
rect 1370 1833 1400 1887
rect 1470 1833 1500 2027
rect 1570 1973 1600 2307
rect 1670 2253 1700 2307
rect 1770 2253 1800 2307
rect 1670 2113 1700 2167
rect 1770 2113 1800 2167
rect 1670 1973 1700 2027
rect 1770 1973 1800 2027
rect 1870 1973 1900 2307
rect 1970 2253 2000 2307
rect 2070 2253 2100 2307
rect 2170 2253 2200 2307
rect 1970 2113 2000 2167
rect 2070 2113 2100 2167
rect 2170 2113 2200 2167
rect 1970 1973 2000 2027
rect 2070 1973 2100 2027
rect 2170 1973 2200 2027
rect 2270 1973 2300 2307
rect 2370 2253 2400 2307
rect 2470 2253 2500 2307
rect 2570 2253 2600 2307
rect 2670 2253 2700 2307
rect 2770 2253 2800 2307
rect 2370 2113 2400 2167
rect 2370 1973 2400 2027
rect 1570 1833 1600 1887
rect 1670 1833 1700 1887
rect 1770 1833 1800 1887
rect 1070 1693 1100 1747
rect 1170 1693 1200 1747
rect 1270 1693 1300 1747
rect 1370 1693 1400 1747
rect 1470 1693 1500 1747
rect 1070 1553 1100 1607
rect 1170 1553 1200 1607
rect 1270 1553 1300 1607
rect 1370 1553 1400 1607
rect 1470 1553 1500 1607
rect 1570 1553 1600 1747
rect 1670 1693 1700 1747
rect 370 1290 400 1327
rect 270 1280 400 1290
rect 270 1246 318 1280
rect 352 1246 400 1280
rect 270 1236 400 1246
rect 270 1183 300 1236
rect 70 1043 100 1097
rect 170 1043 200 1097
rect 270 1043 300 1097
rect 370 1043 400 1236
rect 470 1274 500 1327
rect 570 1274 600 1467
rect 670 1413 700 1467
rect 770 1413 800 1467
rect 870 1413 900 1467
rect 970 1413 1000 1467
rect 1070 1413 1100 1467
rect 1170 1413 1200 1467
rect 1270 1413 1300 1467
rect 1370 1413 1400 1467
rect 1470 1413 1500 1467
rect 470 1264 600 1274
rect 470 1230 518 1264
rect 552 1230 600 1264
rect 470 1220 600 1230
rect 470 1183 500 1220
rect 470 1043 500 1097
rect 570 1043 600 1220
rect 670 1290 700 1327
rect 770 1290 800 1327
rect 670 1280 800 1290
rect 670 1246 718 1280
rect 752 1246 800 1280
rect 670 1236 800 1246
rect 670 1183 700 1236
rect 670 1043 700 1097
rect 770 1043 800 1236
rect 870 1274 900 1327
rect 970 1274 1000 1327
rect 870 1264 1000 1274
rect 870 1230 918 1264
rect 952 1230 1000 1264
rect 870 1220 1000 1230
rect 870 1183 900 1220
rect 970 1183 1000 1220
rect 1070 1290 1100 1327
rect 1170 1290 1200 1327
rect 1070 1280 1200 1290
rect 1070 1246 1118 1280
rect 1152 1246 1200 1280
rect 1070 1236 1200 1246
rect 1070 1183 1100 1236
rect 1170 1183 1200 1236
rect 1270 1274 1300 1327
rect 1370 1274 1400 1327
rect 1270 1264 1400 1274
rect 1270 1230 1318 1264
rect 1352 1230 1400 1264
rect 1270 1220 1400 1230
rect 870 1043 900 1097
rect 70 903 100 957
rect 170 903 200 957
rect 270 903 300 957
rect 370 903 400 957
rect 470 903 500 957
rect 570 903 600 957
rect 670 903 700 957
rect 770 903 800 957
rect 870 903 900 957
rect 970 903 1000 1097
rect 1070 1043 1100 1097
rect 70 763 100 817
rect 170 763 200 817
rect 270 763 300 817
rect 370 763 400 817
rect 470 763 500 817
rect 570 763 600 817
rect 670 763 700 817
rect 770 763 800 817
rect 870 763 900 817
rect 70 623 100 677
rect 170 623 200 677
rect 270 623 300 677
rect 370 623 400 677
rect 470 623 500 677
rect 70 483 100 537
rect 170 483 200 537
rect 70 343 100 397
rect 170 343 200 397
rect 270 343 300 537
rect 370 483 400 537
rect 370 343 400 397
rect 470 343 500 537
rect 570 483 600 677
rect 670 623 700 677
rect 770 623 800 677
rect 870 623 900 677
rect 970 623 1000 817
rect 1070 763 1100 957
rect 1170 903 1200 1097
rect 1270 1043 1300 1220
rect 1370 1183 1400 1220
rect 1470 1290 1500 1327
rect 1570 1290 1600 1467
rect 1670 1413 1700 1607
rect 1770 1553 1800 1747
rect 1870 1693 1900 1887
rect 1970 1833 2000 1887
rect 2070 1833 2100 1887
rect 2170 1833 2200 1887
rect 2270 1833 2300 1887
rect 2370 1833 2400 1887
rect 2470 1833 2500 2167
rect 2570 2113 2600 2167
rect 2670 2113 2700 2167
rect 2770 2113 2800 2167
rect 2870 2113 2900 2307
rect 2970 2253 3000 2307
rect 3070 2253 3100 2307
rect 3170 2253 3200 2307
rect 3270 2253 3300 2307
rect 3370 2253 3400 2307
rect 3470 2253 3500 2307
rect 2970 2113 3000 2167
rect 3070 2113 3100 2167
rect 3170 2113 3200 2167
rect 3270 2113 3300 2167
rect 2570 1973 2600 2027
rect 2670 1973 2700 2027
rect 2770 1973 2800 2027
rect 2870 1973 2900 2027
rect 2970 1973 3000 2027
rect 2570 1833 2600 1887
rect 2670 1833 2700 1887
rect 2770 1833 2800 1887
rect 2870 1833 2900 1887
rect 2970 1833 3000 1887
rect 3070 1833 3100 2027
rect 3170 1973 3200 2027
rect 3270 1973 3300 2027
rect 3370 1973 3400 2167
rect 3470 2113 3500 2167
rect 3570 2113 3600 2307
rect 3670 2253 3700 2307
rect 3770 2253 3800 2307
rect 3870 2253 3900 2307
rect 3970 2253 4000 2307
rect 4070 2253 4100 2307
rect 4170 2253 4200 2307
rect 3470 1973 3500 2027
rect 3570 1973 3600 2027
rect 3670 1973 3700 2167
rect 3770 2113 3800 2167
rect 3870 2113 3900 2167
rect 3770 1973 3800 2027
rect 3170 1833 3200 1887
rect 3270 1833 3300 1887
rect 3370 1833 3400 1887
rect 1870 1553 1900 1607
rect 1970 1553 2000 1747
rect 2070 1693 2100 1747
rect 2170 1693 2200 1747
rect 2270 1693 2300 1747
rect 2370 1693 2400 1747
rect 2470 1693 2500 1747
rect 2570 1693 2600 1747
rect 2070 1553 2100 1607
rect 2170 1553 2200 1607
rect 2270 1553 2300 1607
rect 2370 1553 2400 1607
rect 2470 1553 2500 1607
rect 2570 1553 2600 1607
rect 2670 1553 2700 1747
rect 2770 1693 2800 1747
rect 2870 1693 2900 1747
rect 2970 1693 3000 1747
rect 3070 1693 3100 1747
rect 3170 1693 3200 1747
rect 3270 1693 3300 1747
rect 3370 1693 3400 1747
rect 2770 1553 2800 1607
rect 2870 1553 2900 1607
rect 2970 1553 3000 1607
rect 3070 1553 3100 1607
rect 3170 1553 3200 1607
rect 3270 1553 3300 1607
rect 3370 1553 3400 1607
rect 3470 1553 3500 1887
rect 3570 1833 3600 1887
rect 3570 1693 3600 1747
rect 3670 1693 3700 1887
rect 3770 1833 3800 1887
rect 3870 1833 3900 2027
rect 3970 1973 4000 2167
rect 4070 2113 4100 2167
rect 4170 2113 4200 2167
rect 4270 2113 4300 2307
rect 4370 2253 4400 2307
rect 4370 2113 4400 2167
rect 4070 1973 4100 2027
rect 4170 1973 4200 2027
rect 4270 1973 4300 2027
rect 4370 1973 4400 2027
rect 3570 1553 3600 1607
rect 3670 1553 3700 1607
rect 3770 1553 3800 1747
rect 3870 1693 3900 1747
rect 3970 1693 4000 1887
rect 4070 1833 4100 1887
rect 4170 1833 4200 1887
rect 4270 1833 4300 1887
rect 4370 1833 4400 1887
rect 4470 1833 4500 2307
rect 4570 2253 4600 2307
rect 4670 2253 4700 2307
rect 4770 2253 4800 2307
rect 4870 2253 4900 2307
rect 4970 2253 5000 2307
rect 5070 2253 5100 2307
rect 5170 2253 5200 2307
rect 5270 2253 5300 2307
rect 5370 2253 5400 2307
rect 5470 2253 5500 2446
rect 5570 2393 5600 2446
rect 5670 2484 5700 2537
rect 5770 2484 5800 2537
rect 5670 2474 5800 2484
rect 5670 2440 5718 2474
rect 5752 2440 5800 2474
rect 5670 2430 5800 2440
rect 5670 2393 5700 2430
rect 5770 2393 5800 2430
rect 5870 2500 5900 2537
rect 5970 2500 6000 2537
rect 5870 2490 6000 2500
rect 5870 2456 5918 2490
rect 5952 2456 6000 2490
rect 5870 2446 6000 2456
rect 5870 2393 5900 2446
rect 5970 2393 6000 2446
rect 6070 2484 6100 2537
rect 6170 2484 6200 2537
rect 6070 2474 6200 2484
rect 6070 2440 6118 2474
rect 6152 2440 6200 2474
rect 6070 2430 6200 2440
rect 6070 2393 6100 2430
rect 6170 2393 6200 2430
rect 6270 2500 6300 2537
rect 6370 2500 6400 2537
rect 6570 2504 6600 2537
rect 6670 2504 6700 2537
rect 6880 2504 6910 2537
rect 6980 2504 7010 2537
rect 7080 2504 7110 2537
rect 7180 2504 7210 2537
rect 7280 2504 7310 2537
rect 7380 2504 7410 2537
rect 6270 2490 6400 2500
rect 6270 2456 6318 2490
rect 6352 2456 6400 2490
rect 6270 2446 6400 2456
rect 6270 2393 6300 2446
rect 6370 2393 6400 2446
rect 6558 2488 6612 2504
rect 6558 2454 6568 2488
rect 6602 2454 6612 2488
rect 6558 2438 6612 2454
rect 6658 2488 6712 2504
rect 6658 2454 6668 2488
rect 6702 2454 6712 2488
rect 6658 2438 6712 2454
rect 6868 2488 6922 2504
rect 6868 2454 6878 2488
rect 6912 2454 6922 2488
rect 6868 2438 6922 2454
rect 6968 2488 7022 2504
rect 6968 2454 6978 2488
rect 7012 2454 7022 2488
rect 6968 2438 7022 2454
rect 7068 2488 7122 2504
rect 7068 2454 7078 2488
rect 7112 2454 7122 2488
rect 7068 2438 7122 2454
rect 7168 2488 7222 2504
rect 7168 2454 7178 2488
rect 7212 2454 7222 2488
rect 7168 2438 7222 2454
rect 7268 2488 7322 2504
rect 7268 2454 7278 2488
rect 7312 2454 7322 2488
rect 7268 2438 7322 2454
rect 7368 2488 7422 2504
rect 7368 2454 7378 2488
rect 7412 2454 7422 2488
rect 7368 2438 7422 2454
rect 6570 2393 6600 2438
rect 6670 2393 6700 2438
rect 6880 2393 6910 2438
rect 6980 2393 7010 2438
rect 7080 2393 7110 2438
rect 7180 2393 7210 2438
rect 7280 2393 7310 2438
rect 7380 2393 7410 2438
rect 5570 2253 5600 2307
rect 5670 2253 5700 2307
rect 5770 2253 5800 2307
rect 5870 2253 5900 2307
rect 5970 2253 6000 2307
rect 6070 2253 6100 2307
rect 6170 2253 6200 2307
rect 6270 2253 6300 2307
rect 6370 2253 6400 2307
rect 6570 2253 6600 2307
rect 6670 2253 6700 2307
rect 6880 2253 6910 2307
rect 6980 2253 7010 2307
rect 7080 2253 7110 2307
rect 7180 2253 7210 2307
rect 7280 2253 7310 2307
rect 7380 2253 7410 2307
rect 4570 2113 4600 2167
rect 4670 2113 4700 2167
rect 4770 2113 4800 2167
rect 4870 2113 4900 2167
rect 4970 2113 5000 2167
rect 5070 2113 5100 2167
rect 5170 2113 5200 2167
rect 5270 2113 5300 2167
rect 5370 2113 5400 2167
rect 5470 2113 5500 2167
rect 5570 2113 5600 2167
rect 5670 2113 5700 2167
rect 5770 2113 5800 2167
rect 5870 2113 5900 2167
rect 5970 2113 6000 2167
rect 6070 2113 6100 2167
rect 6170 2113 6200 2167
rect 6270 2113 6300 2167
rect 6370 2113 6400 2167
rect 6570 2113 6600 2167
rect 6670 2113 6700 2167
rect 6880 2113 6910 2167
rect 6980 2113 7010 2167
rect 7080 2113 7110 2167
rect 7180 2113 7210 2167
rect 7280 2113 7310 2167
rect 7380 2113 7410 2167
rect 4570 1973 4600 2027
rect 4670 1973 4700 2027
rect 4770 1973 4800 2027
rect 4870 1973 4900 2027
rect 4570 1833 4600 1887
rect 4670 1833 4700 1887
rect 4770 1833 4800 1887
rect 4070 1693 4100 1747
rect 4170 1693 4200 1747
rect 4270 1693 4300 1747
rect 4370 1693 4400 1747
rect 3870 1553 3900 1607
rect 3970 1553 4000 1607
rect 4070 1553 4100 1607
rect 1470 1280 1600 1290
rect 1470 1246 1518 1280
rect 1552 1246 1600 1280
rect 1470 1236 1600 1246
rect 1470 1183 1500 1236
rect 1570 1183 1600 1236
rect 1670 1274 1700 1327
rect 1770 1274 1800 1467
rect 1870 1413 1900 1467
rect 1970 1413 2000 1467
rect 2070 1413 2100 1467
rect 2170 1413 2200 1467
rect 2270 1413 2300 1467
rect 2370 1413 2400 1467
rect 2470 1413 2500 1467
rect 2570 1413 2600 1467
rect 2670 1413 2700 1467
rect 2770 1413 2800 1467
rect 2870 1413 2900 1467
rect 1670 1264 1800 1274
rect 1670 1230 1718 1264
rect 1752 1230 1800 1264
rect 1670 1220 1800 1230
rect 1670 1183 1700 1220
rect 1770 1183 1800 1220
rect 1870 1290 1900 1327
rect 1970 1290 2000 1327
rect 1870 1280 2000 1290
rect 1870 1246 1918 1280
rect 1952 1246 2000 1280
rect 1870 1236 2000 1246
rect 1870 1183 1900 1236
rect 1970 1183 2000 1236
rect 2070 1274 2100 1327
rect 2170 1274 2200 1327
rect 2070 1264 2200 1274
rect 2070 1230 2118 1264
rect 2152 1230 2200 1264
rect 2070 1220 2200 1230
rect 2070 1183 2100 1220
rect 2170 1183 2200 1220
rect 2270 1290 2300 1327
rect 2370 1290 2400 1327
rect 2270 1280 2400 1290
rect 2270 1246 2318 1280
rect 2352 1246 2400 1280
rect 2270 1236 2400 1246
rect 2270 1183 2300 1236
rect 2370 1183 2400 1236
rect 2470 1274 2500 1327
rect 2570 1274 2600 1327
rect 2470 1264 2600 1274
rect 2470 1230 2518 1264
rect 2552 1230 2600 1264
rect 2470 1220 2600 1230
rect 2470 1183 2500 1220
rect 1370 1043 1400 1097
rect 1470 1043 1500 1097
rect 1570 1043 1600 1097
rect 1670 1043 1700 1097
rect 1770 1043 1800 1097
rect 1870 1043 1900 1097
rect 1970 1043 2000 1097
rect 2070 1043 2100 1097
rect 1270 903 1300 957
rect 1370 903 1400 957
rect 1470 903 1500 957
rect 1570 903 1600 957
rect 1670 903 1700 957
rect 1170 763 1200 817
rect 1270 763 1300 817
rect 1370 763 1400 817
rect 1470 763 1500 817
rect 1570 763 1600 817
rect 1670 763 1700 817
rect 1770 763 1800 957
rect 1870 903 1900 957
rect 1970 903 2000 957
rect 2070 903 2100 957
rect 2170 903 2200 1097
rect 2270 1043 2300 1097
rect 2370 1043 2400 1097
rect 2270 903 2300 957
rect 2370 903 2400 957
rect 2470 903 2500 1097
rect 2570 1043 2600 1220
rect 2670 1290 2700 1327
rect 2770 1290 2800 1327
rect 2670 1280 2800 1290
rect 2670 1246 2718 1280
rect 2752 1246 2800 1280
rect 2670 1236 2800 1246
rect 2670 1183 2700 1236
rect 2670 1043 2700 1097
rect 2770 1043 2800 1236
rect 2870 1274 2900 1327
rect 2970 1274 3000 1467
rect 3070 1413 3100 1467
rect 3170 1413 3200 1467
rect 3270 1413 3300 1467
rect 3370 1413 3400 1467
rect 3470 1413 3500 1467
rect 2870 1264 3000 1274
rect 2870 1230 2918 1264
rect 2952 1230 3000 1264
rect 2870 1220 3000 1230
rect 2870 1183 2900 1220
rect 2970 1183 3000 1220
rect 3070 1290 3100 1327
rect 3170 1290 3200 1327
rect 3070 1280 3200 1290
rect 3070 1246 3118 1280
rect 3152 1246 3200 1280
rect 3070 1236 3200 1246
rect 3070 1183 3100 1236
rect 3170 1183 3200 1236
rect 3270 1274 3300 1327
rect 3370 1274 3400 1327
rect 3270 1264 3400 1274
rect 3270 1230 3318 1264
rect 3352 1230 3400 1264
rect 3270 1220 3400 1230
rect 3270 1183 3300 1220
rect 3370 1183 3400 1220
rect 3470 1290 3500 1327
rect 3570 1290 3600 1467
rect 3670 1413 3700 1467
rect 3770 1413 3800 1467
rect 3470 1280 3600 1290
rect 3470 1246 3518 1280
rect 3552 1246 3600 1280
rect 3470 1236 3600 1246
rect 3470 1183 3500 1236
rect 3570 1183 3600 1236
rect 3670 1274 3700 1327
rect 3770 1274 3800 1327
rect 3670 1264 3800 1274
rect 3670 1230 3718 1264
rect 3752 1230 3800 1264
rect 3670 1220 3800 1230
rect 3670 1183 3700 1220
rect 3770 1183 3800 1220
rect 3870 1290 3900 1467
rect 3970 1413 4000 1467
rect 4070 1413 4100 1467
rect 4170 1413 4200 1607
rect 4270 1553 4300 1607
rect 4370 1553 4400 1607
rect 4270 1413 4300 1467
rect 4370 1413 4400 1467
rect 4470 1413 4500 1747
rect 4570 1693 4600 1747
rect 4670 1693 4700 1747
rect 4770 1693 4800 1747
rect 4870 1693 4900 1887
rect 4970 1833 5000 2027
rect 5070 1973 5100 2027
rect 5070 1833 5100 1887
rect 5170 1833 5200 2027
rect 5270 1973 5300 2027
rect 5270 1833 5300 1887
rect 5370 1833 5400 2027
rect 5470 1973 5500 2027
rect 5570 1973 5600 2027
rect 5670 1973 5700 2027
rect 5470 1833 5500 1887
rect 5570 1833 5600 1887
rect 5670 1833 5700 1887
rect 5770 1833 5800 2027
rect 5870 1973 5900 2027
rect 5970 1973 6000 2027
rect 5870 1833 5900 1887
rect 5970 1833 6000 1887
rect 6070 1833 6100 2027
rect 6170 1973 6200 2027
rect 6270 1973 6300 2027
rect 6370 1973 6400 2027
rect 6570 1973 6600 2027
rect 6670 1973 6700 2027
rect 6880 1973 6910 2027
rect 6980 1973 7010 2027
rect 7080 1973 7110 2027
rect 7180 1973 7210 2027
rect 7280 1973 7310 2027
rect 7380 1973 7410 2027
rect 6170 1833 6200 1887
rect 6270 1833 6300 1887
rect 6370 1833 6400 1887
rect 6570 1833 6600 1887
rect 6670 1833 6700 1887
rect 6880 1833 6910 1887
rect 6980 1833 7010 1887
rect 7080 1833 7110 1887
rect 7180 1833 7210 1887
rect 7280 1833 7310 1887
rect 7380 1833 7410 1887
rect 4970 1693 5000 1747
rect 5070 1693 5100 1747
rect 5170 1693 5200 1747
rect 5270 1693 5300 1747
rect 4570 1553 4600 1607
rect 4670 1553 4700 1607
rect 4770 1553 4800 1607
rect 4870 1553 4900 1607
rect 4970 1553 5000 1607
rect 4570 1413 4600 1467
rect 4670 1413 4700 1467
rect 4770 1413 4800 1467
rect 3970 1290 4000 1327
rect 3870 1280 4000 1290
rect 3870 1246 3918 1280
rect 3952 1246 4000 1280
rect 3870 1236 4000 1246
rect 3870 1183 3900 1236
rect 3970 1183 4000 1236
rect 4070 1274 4100 1327
rect 4170 1274 4200 1327
rect 4070 1264 4200 1274
rect 4070 1230 4118 1264
rect 4152 1230 4200 1264
rect 4070 1220 4200 1230
rect 4070 1183 4100 1220
rect 4170 1183 4200 1220
rect 4270 1290 4300 1327
rect 4370 1290 4400 1327
rect 4270 1280 4400 1290
rect 4270 1246 4318 1280
rect 4352 1246 4400 1280
rect 4270 1236 4400 1246
rect 2870 1043 2900 1097
rect 2970 1043 3000 1097
rect 3070 1043 3100 1097
rect 3170 1043 3200 1097
rect 3270 1043 3300 1097
rect 3370 1043 3400 1097
rect 3470 1043 3500 1097
rect 3570 1043 3600 1097
rect 3670 1043 3700 1097
rect 3770 1043 3800 1097
rect 3870 1043 3900 1097
rect 3970 1043 4000 1097
rect 4070 1043 4100 1097
rect 4170 1043 4200 1097
rect 2570 903 2600 957
rect 2670 903 2700 957
rect 2770 903 2800 957
rect 2870 903 2900 957
rect 2970 903 3000 957
rect 3070 903 3100 957
rect 3170 903 3200 957
rect 3270 903 3300 957
rect 3370 903 3400 957
rect 3470 903 3500 957
rect 3570 903 3600 957
rect 3670 903 3700 957
rect 3770 903 3800 957
rect 3870 903 3900 957
rect 3970 903 4000 957
rect 4070 903 4100 957
rect 4170 903 4200 957
rect 4270 903 4300 1236
rect 4370 1183 4400 1236
rect 4470 1274 4500 1327
rect 4570 1274 4600 1327
rect 4470 1264 4600 1274
rect 4470 1230 4518 1264
rect 4552 1230 4600 1264
rect 4470 1220 4600 1230
rect 4470 1183 4500 1220
rect 4570 1183 4600 1220
rect 4670 1290 4700 1327
rect 4770 1290 4800 1327
rect 4670 1280 4800 1290
rect 4670 1246 4718 1280
rect 4752 1246 4800 1280
rect 4670 1236 4800 1246
rect 4670 1183 4700 1236
rect 4770 1183 4800 1236
rect 4870 1274 4900 1467
rect 4970 1413 5000 1467
rect 4970 1274 5000 1327
rect 4870 1264 5000 1274
rect 4870 1230 4918 1264
rect 4952 1230 5000 1264
rect 4870 1220 5000 1230
rect 4870 1183 4900 1220
rect 4970 1183 5000 1220
rect 5070 1290 5100 1607
rect 5170 1553 5200 1607
rect 5170 1413 5200 1467
rect 5270 1413 5300 1607
rect 5370 1553 5400 1747
rect 5470 1693 5500 1747
rect 5570 1693 5600 1747
rect 5670 1693 5700 1747
rect 5370 1413 5400 1467
rect 5470 1413 5500 1607
rect 5570 1553 5600 1607
rect 5670 1553 5700 1607
rect 5570 1413 5600 1467
rect 5670 1413 5700 1467
rect 5770 1413 5800 1747
rect 5870 1693 5900 1747
rect 5870 1553 5900 1607
rect 5870 1413 5900 1467
rect 5970 1413 6000 1747
rect 6070 1693 6100 1747
rect 6170 1693 6200 1747
rect 6270 1693 6300 1747
rect 6370 1693 6400 1747
rect 6570 1693 6600 1747
rect 6670 1693 6700 1747
rect 6880 1693 6910 1747
rect 6980 1693 7010 1747
rect 7080 1693 7110 1747
rect 7180 1693 7210 1747
rect 7280 1693 7310 1747
rect 7380 1693 7410 1747
rect 6070 1553 6100 1607
rect 6170 1553 6200 1607
rect 6070 1413 6100 1467
rect 5170 1290 5200 1327
rect 5070 1280 5200 1290
rect 5070 1246 5118 1280
rect 5152 1246 5200 1280
rect 5070 1236 5200 1246
rect 5070 1183 5100 1236
rect 5170 1183 5200 1236
rect 5270 1274 5300 1327
rect 5370 1274 5400 1327
rect 5270 1264 5400 1274
rect 5270 1230 5318 1264
rect 5352 1230 5400 1264
rect 5270 1220 5400 1230
rect 5270 1183 5300 1220
rect 5370 1183 5400 1220
rect 5470 1290 5500 1327
rect 5570 1290 5600 1327
rect 5470 1280 5600 1290
rect 5470 1246 5518 1280
rect 5552 1246 5600 1280
rect 5470 1236 5600 1246
rect 4370 1043 4400 1097
rect 4470 1043 4500 1097
rect 4570 1043 4600 1097
rect 4670 1043 4700 1097
rect 4770 1043 4800 1097
rect 1870 763 1900 817
rect 1970 763 2000 817
rect 670 483 700 537
rect 770 483 800 537
rect 870 483 900 537
rect 970 483 1000 537
rect 1070 483 1100 677
rect 1170 623 1200 677
rect 1270 623 1300 677
rect 1370 623 1400 677
rect 1470 623 1500 677
rect 1570 623 1600 677
rect 1670 623 1700 677
rect 1770 623 1800 677
rect 1870 623 1900 677
rect 1970 623 2000 677
rect 2070 623 2100 817
rect 2170 763 2200 817
rect 2170 623 2200 677
rect 2270 623 2300 817
rect 2370 763 2400 817
rect 2470 763 2500 817
rect 2570 763 2600 817
rect 2670 763 2700 817
rect 2770 763 2800 817
rect 2870 763 2900 817
rect 2970 763 3000 817
rect 3070 763 3100 817
rect 3170 763 3200 817
rect 3270 763 3300 817
rect 3370 763 3400 817
rect 3470 763 3500 817
rect 3570 763 3600 817
rect 3670 763 3700 817
rect 3770 763 3800 817
rect 3870 763 3900 817
rect 3970 763 4000 817
rect 4070 763 4100 817
rect 4170 763 4200 817
rect 4270 763 4300 817
rect 4370 763 4400 957
rect 4470 903 4500 957
rect 2370 623 2400 677
rect 2470 623 2500 677
rect 2570 623 2600 677
rect 2670 623 2700 677
rect 2770 623 2800 677
rect 2870 623 2900 677
rect 2970 623 3000 677
rect 3070 623 3100 677
rect 3170 623 3200 677
rect 3270 623 3300 677
rect 3370 623 3400 677
rect 3470 623 3500 677
rect 3570 623 3600 677
rect 3670 623 3700 677
rect 1170 483 1200 537
rect 1270 483 1300 537
rect 1370 483 1400 537
rect 570 343 600 397
rect 70 203 100 257
rect 170 203 200 257
rect 270 203 300 257
rect 370 203 400 257
rect 470 203 500 257
rect 570 203 600 257
rect 670 203 700 397
rect 770 343 800 397
rect 870 343 900 397
rect 970 343 1000 397
rect 1070 343 1100 397
rect 1170 343 1200 397
rect 1270 343 1300 397
rect 1370 343 1400 397
rect 1470 343 1500 537
rect 1570 483 1600 537
rect 1670 483 1700 537
rect 1770 483 1800 537
rect 1870 483 1900 537
rect 1970 483 2000 537
rect 2070 483 2100 537
rect 2170 483 2200 537
rect 2270 483 2300 537
rect 2370 483 2400 537
rect 2470 483 2500 537
rect 2570 483 2600 537
rect 2670 483 2700 537
rect 2770 483 2800 537
rect 2870 483 2900 537
rect 2970 483 3000 537
rect 770 203 800 257
rect 70 64 100 117
rect 170 64 200 117
rect 70 54 200 64
rect 70 20 118 54
rect 152 20 200 54
rect 70 10 200 20
rect 70 0 100 10
rect 170 0 200 10
rect 270 80 300 117
rect 370 80 400 117
rect 270 70 400 80
rect 270 36 318 70
rect 352 36 400 70
rect 270 26 400 36
rect 270 0 300 26
rect 370 0 400 26
rect 470 64 500 117
rect 570 64 600 117
rect 470 54 600 64
rect 470 20 518 54
rect 552 20 600 54
rect 470 10 600 20
rect 470 0 500 10
rect 570 0 600 10
rect 670 80 700 117
rect 770 80 800 117
rect 670 70 800 80
rect 670 36 718 70
rect 752 36 800 70
rect 670 26 800 36
rect 670 0 700 26
rect 770 0 800 26
rect 870 64 900 257
rect 970 203 1000 257
rect 1070 203 1100 257
rect 1170 203 1200 257
rect 1270 203 1300 257
rect 1370 203 1400 257
rect 1470 203 1500 257
rect 1570 203 1600 397
rect 1670 343 1700 397
rect 1770 343 1800 397
rect 1870 343 1900 397
rect 1970 343 2000 397
rect 2070 343 2100 397
rect 2170 343 2200 397
rect 1670 203 1700 257
rect 1770 203 1800 257
rect 1870 203 1900 257
rect 970 64 1000 117
rect 870 54 1000 64
rect 870 20 918 54
rect 952 20 1000 54
rect 870 10 1000 20
rect 870 0 900 10
rect 970 0 1000 10
rect 1070 80 1100 117
rect 1170 80 1200 117
rect 1070 70 1200 80
rect 1070 36 1118 70
rect 1152 36 1200 70
rect 1070 26 1200 36
rect 1070 0 1100 26
rect 1170 0 1200 26
rect 1270 64 1300 117
rect 1370 64 1400 117
rect 1270 54 1400 64
rect 1270 20 1318 54
rect 1352 20 1400 54
rect 1270 10 1400 20
rect 1270 0 1300 10
rect 1370 0 1400 10
rect 1470 80 1500 117
rect 1570 80 1600 117
rect 1470 70 1600 80
rect 1470 36 1518 70
rect 1552 36 1600 70
rect 1470 26 1600 36
rect 1470 0 1500 26
rect 1570 0 1600 26
rect 1670 64 1700 117
rect 1770 64 1800 117
rect 1670 54 1800 64
rect 1670 20 1718 54
rect 1752 20 1800 54
rect 1670 10 1800 20
rect 1670 0 1700 10
rect 1770 0 1800 10
rect 1870 80 1900 117
rect 1970 80 2000 257
rect 2070 203 2100 257
rect 2170 203 2200 257
rect 2270 203 2300 397
rect 2370 343 2400 397
rect 2370 203 2400 257
rect 2470 203 2500 397
rect 2570 343 2600 397
rect 2570 203 2600 257
rect 2670 203 2700 397
rect 2770 343 2800 397
rect 2770 203 2800 257
rect 2870 203 2900 397
rect 2970 343 3000 397
rect 3070 343 3100 537
rect 3170 483 3200 537
rect 3170 343 3200 397
rect 3270 343 3300 537
rect 3370 483 3400 537
rect 3470 483 3500 537
rect 3370 343 3400 397
rect 3470 343 3500 397
rect 2970 203 3000 257
rect 3070 203 3100 257
rect 3170 203 3200 257
rect 3270 203 3300 257
rect 3370 203 3400 257
rect 3470 203 3500 257
rect 1870 70 2000 80
rect 1870 36 1918 70
rect 1952 36 2000 70
rect 1870 26 2000 36
rect 1870 0 1900 26
rect 1970 0 2000 26
rect 2070 64 2100 117
rect 2170 64 2200 117
rect 2070 54 2200 64
rect 2070 20 2118 54
rect 2152 20 2200 54
rect 2070 10 2200 20
rect 2070 0 2100 10
rect 2170 0 2200 10
rect 2270 80 2300 117
rect 2370 80 2400 117
rect 2270 70 2400 80
rect 2270 36 2318 70
rect 2352 36 2400 70
rect 2270 26 2400 36
rect 2270 0 2300 26
rect 2370 0 2400 26
rect 2470 64 2500 117
rect 2570 64 2600 117
rect 2470 54 2600 64
rect 2470 20 2518 54
rect 2552 20 2600 54
rect 2470 10 2600 20
rect 2470 0 2500 10
rect 2570 0 2600 10
rect 2670 80 2700 117
rect 2770 80 2800 117
rect 2670 70 2800 80
rect 2670 36 2718 70
rect 2752 36 2800 70
rect 2670 26 2800 36
rect 2670 0 2700 26
rect 2770 0 2800 26
rect 2870 64 2900 117
rect 2970 64 3000 117
rect 2870 54 3000 64
rect 2870 20 2918 54
rect 2952 20 3000 54
rect 2870 10 3000 20
rect 2870 0 2900 10
rect 2970 0 3000 10
rect 3070 80 3100 117
rect 3170 80 3200 117
rect 3070 70 3200 80
rect 3070 36 3118 70
rect 3152 36 3200 70
rect 3070 26 3200 36
rect 3070 0 3100 26
rect 3170 0 3200 26
rect 3270 64 3300 117
rect 3370 64 3400 117
rect 3270 54 3400 64
rect 3270 20 3318 54
rect 3352 20 3400 54
rect 3270 10 3400 20
rect 3270 0 3300 10
rect 3370 0 3400 10
rect 3470 80 3500 117
rect 3570 80 3600 537
rect 3670 483 3700 537
rect 3670 343 3700 397
rect 3770 343 3800 677
rect 3870 623 3900 677
rect 3970 623 4000 677
rect 3870 483 3900 537
rect 3970 483 4000 537
rect 4070 483 4100 677
rect 4170 623 4200 677
rect 4170 483 4200 537
rect 4270 483 4300 677
rect 4370 623 4400 677
rect 4470 623 4500 817
rect 4570 763 4600 957
rect 4670 903 4700 957
rect 4770 903 4800 957
rect 4870 903 4900 1097
rect 4970 1043 5000 1097
rect 4970 903 5000 957
rect 5070 903 5100 1097
rect 5170 1043 5200 1097
rect 5270 1043 5300 1097
rect 5370 1043 5400 1097
rect 5470 1043 5500 1236
rect 5570 1183 5600 1236
rect 5670 1274 5700 1327
rect 5770 1274 5800 1327
rect 5670 1264 5800 1274
rect 5670 1230 5718 1264
rect 5752 1230 5800 1264
rect 5670 1220 5800 1230
rect 5670 1183 5700 1220
rect 5770 1183 5800 1220
rect 5870 1290 5900 1327
rect 5970 1290 6000 1327
rect 5870 1280 6000 1290
rect 5870 1246 5918 1280
rect 5952 1246 6000 1280
rect 5870 1236 6000 1246
rect 5870 1183 5900 1236
rect 5570 1043 5600 1097
rect 5670 1043 5700 1097
rect 5770 1043 5800 1097
rect 5870 1043 5900 1097
rect 5970 1043 6000 1236
rect 6070 1274 6100 1327
rect 6170 1274 6200 1467
rect 6270 1413 6300 1607
rect 6370 1553 6400 1607
rect 6570 1553 6600 1607
rect 6670 1553 6700 1607
rect 6880 1553 6910 1607
rect 6980 1553 7010 1607
rect 7080 1553 7110 1607
rect 7180 1553 7210 1607
rect 7280 1553 7310 1607
rect 7380 1553 7410 1607
rect 6370 1413 6400 1467
rect 6570 1413 6600 1467
rect 6670 1413 6700 1467
rect 6880 1413 6910 1467
rect 6980 1413 7010 1467
rect 7080 1413 7110 1467
rect 7180 1413 7210 1467
rect 7280 1413 7310 1467
rect 7380 1413 7410 1467
rect 6070 1264 6200 1274
rect 6070 1230 6118 1264
rect 6152 1230 6200 1264
rect 6070 1220 6200 1230
rect 6070 1183 6100 1220
rect 6170 1183 6200 1220
rect 6270 1290 6300 1327
rect 6370 1290 6400 1327
rect 6570 1294 6600 1327
rect 6670 1294 6700 1327
rect 6880 1294 6910 1327
rect 6980 1294 7010 1327
rect 7080 1294 7110 1327
rect 7180 1294 7210 1327
rect 7280 1294 7310 1327
rect 7380 1294 7410 1327
rect 6270 1280 6400 1290
rect 6270 1246 6318 1280
rect 6352 1246 6400 1280
rect 6270 1236 6400 1246
rect 6270 1183 6300 1236
rect 6370 1183 6400 1236
rect 6558 1278 6612 1294
rect 6558 1244 6568 1278
rect 6602 1244 6612 1278
rect 6558 1228 6612 1244
rect 6658 1278 6712 1294
rect 6658 1244 6668 1278
rect 6702 1244 6712 1278
rect 6658 1228 6712 1244
rect 6868 1278 6922 1294
rect 6868 1244 6878 1278
rect 6912 1244 6922 1278
rect 6868 1228 6922 1244
rect 6968 1278 7022 1294
rect 6968 1244 6978 1278
rect 7012 1244 7022 1278
rect 6968 1228 7022 1244
rect 7068 1278 7122 1294
rect 7068 1244 7078 1278
rect 7112 1244 7122 1278
rect 7068 1228 7122 1244
rect 7168 1278 7222 1294
rect 7168 1244 7178 1278
rect 7212 1244 7222 1278
rect 7168 1228 7222 1244
rect 7268 1278 7322 1294
rect 7268 1244 7278 1278
rect 7312 1244 7322 1278
rect 7268 1228 7322 1244
rect 7368 1278 7422 1294
rect 7368 1244 7378 1278
rect 7412 1244 7422 1278
rect 7368 1228 7422 1244
rect 6570 1183 6600 1228
rect 6670 1183 6700 1228
rect 6880 1183 6910 1228
rect 6980 1183 7010 1228
rect 7080 1183 7110 1228
rect 7180 1183 7210 1228
rect 7280 1183 7310 1228
rect 7380 1183 7410 1228
rect 6070 1043 6100 1097
rect 6170 1043 6200 1097
rect 5170 903 5200 957
rect 5270 903 5300 957
rect 5370 903 5400 957
rect 5470 903 5500 957
rect 5570 903 5600 957
rect 5670 903 5700 957
rect 5770 903 5800 957
rect 5870 903 5900 957
rect 5970 903 6000 957
rect 6070 903 6100 957
rect 6170 903 6200 957
rect 6270 903 6300 1097
rect 6370 1043 6400 1097
rect 6570 1043 6600 1097
rect 6670 1043 6700 1097
rect 6880 1043 6910 1097
rect 6980 1043 7010 1097
rect 7080 1043 7110 1097
rect 7180 1043 7210 1097
rect 7280 1043 7310 1097
rect 7380 1043 7410 1097
rect 6370 903 6400 957
rect 6570 903 6600 957
rect 6670 903 6700 957
rect 6880 903 6910 957
rect 6980 903 7010 957
rect 7080 903 7110 957
rect 7180 903 7210 957
rect 7280 903 7310 957
rect 7380 903 7410 957
rect 4670 763 4700 817
rect 4770 763 4800 817
rect 4870 763 4900 817
rect 4970 763 5000 817
rect 5070 763 5100 817
rect 5170 763 5200 817
rect 5270 763 5300 817
rect 5370 763 5400 817
rect 5470 763 5500 817
rect 4570 623 4600 677
rect 4370 483 4400 537
rect 4470 483 4500 537
rect 4570 483 4600 537
rect 4670 483 4700 677
rect 4770 623 4800 677
rect 4870 623 4900 677
rect 4970 623 5000 677
rect 5070 623 5100 677
rect 5170 623 5200 677
rect 4770 483 4800 537
rect 4870 483 4900 537
rect 4970 483 5000 537
rect 5070 483 5100 537
rect 5170 483 5200 537
rect 5270 483 5300 677
rect 5370 623 5400 677
rect 5470 623 5500 677
rect 5570 623 5600 817
rect 5670 763 5700 817
rect 5670 623 5700 677
rect 5770 623 5800 817
rect 5870 763 5900 817
rect 5970 763 6000 817
rect 6070 763 6100 817
rect 6170 763 6200 817
rect 6270 763 6300 817
rect 6370 763 6400 817
rect 6570 763 6600 817
rect 6670 763 6700 817
rect 6880 763 6910 817
rect 6980 763 7010 817
rect 7080 763 7110 817
rect 7180 763 7210 817
rect 7280 763 7310 817
rect 7380 763 7410 817
rect 5870 623 5900 677
rect 5970 623 6000 677
rect 5370 483 5400 537
rect 5470 483 5500 537
rect 3870 343 3900 397
rect 3970 343 4000 397
rect 4070 343 4100 397
rect 4170 343 4200 397
rect 4270 343 4300 397
rect 4370 343 4400 397
rect 4470 343 4500 397
rect 4570 343 4600 397
rect 4670 343 4700 397
rect 4770 343 4800 397
rect 4870 343 4900 397
rect 4970 343 5000 397
rect 5070 343 5100 397
rect 5170 343 5200 397
rect 5270 343 5300 397
rect 5370 343 5400 397
rect 5470 343 5500 397
rect 5570 343 5600 537
rect 5670 483 5700 537
rect 5770 483 5800 537
rect 5870 483 5900 537
rect 5970 483 6000 537
rect 6070 483 6100 677
rect 6170 623 6200 677
rect 6270 623 6300 677
rect 6370 623 6400 677
rect 6570 623 6600 677
rect 6670 623 6700 677
rect 6880 623 6910 677
rect 6980 623 7010 677
rect 7080 623 7110 677
rect 7180 623 7210 677
rect 7280 623 7310 677
rect 7380 623 7410 677
rect 6170 483 6200 537
rect 3670 203 3700 257
rect 3770 203 3800 257
rect 3870 203 3900 257
rect 3970 203 4000 257
rect 4070 203 4100 257
rect 4170 203 4200 257
rect 4270 203 4300 257
rect 4370 203 4400 257
rect 4470 203 4500 257
rect 4570 203 4600 257
rect 4670 203 4700 257
rect 3470 70 3600 80
rect 3470 36 3518 70
rect 3552 36 3600 70
rect 3470 26 3600 36
rect 3470 0 3500 26
rect 3570 0 3600 26
rect 3670 64 3700 117
rect 3770 64 3800 117
rect 3670 54 3800 64
rect 3670 20 3718 54
rect 3752 20 3800 54
rect 3670 10 3800 20
rect 3670 0 3700 10
rect 3770 0 3800 10
rect 3870 80 3900 117
rect 3970 80 4000 117
rect 3870 70 4000 80
rect 3870 36 3918 70
rect 3952 36 4000 70
rect 3870 26 4000 36
rect 3870 0 3900 26
rect 3970 0 4000 26
rect 4070 64 4100 117
rect 4170 64 4200 117
rect 4070 54 4200 64
rect 4070 20 4118 54
rect 4152 20 4200 54
rect 4070 10 4200 20
rect 4070 0 4100 10
rect 4170 0 4200 10
rect 4270 80 4300 117
rect 4370 80 4400 117
rect 4270 70 4400 80
rect 4270 36 4318 70
rect 4352 36 4400 70
rect 4270 26 4400 36
rect 4270 0 4300 26
rect 4370 0 4400 26
rect 4470 64 4500 117
rect 4570 64 4600 117
rect 4470 54 4600 64
rect 4470 20 4518 54
rect 4552 20 4600 54
rect 4470 10 4600 20
rect 4470 0 4500 10
rect 4570 0 4600 10
rect 4670 80 4700 117
rect 4770 80 4800 257
rect 4870 203 4900 257
rect 4970 203 5000 257
rect 5070 203 5100 257
rect 5170 203 5200 257
rect 5270 203 5300 257
rect 5370 203 5400 257
rect 5470 203 5500 257
rect 5570 203 5600 257
rect 5670 203 5700 397
rect 5770 343 5800 397
rect 5870 343 5900 397
rect 5970 343 6000 397
rect 6070 343 6100 397
rect 6170 343 6200 397
rect 6270 343 6300 537
rect 6370 483 6400 537
rect 6570 483 6600 537
rect 6670 483 6700 537
rect 6880 483 6910 537
rect 6980 483 7010 537
rect 7080 483 7110 537
rect 7180 483 7210 537
rect 7280 483 7310 537
rect 7380 483 7410 537
rect 6370 343 6400 397
rect 6570 343 6600 397
rect 6670 343 6700 397
rect 6880 343 6910 397
rect 6980 343 7010 397
rect 7080 343 7110 397
rect 7180 343 7210 397
rect 7280 343 7310 397
rect 7380 343 7410 397
rect 5770 203 5800 257
rect 5870 203 5900 257
rect 5970 203 6000 257
rect 6070 203 6100 257
rect 4670 70 4800 80
rect 4670 36 4718 70
rect 4752 36 4800 70
rect 4670 26 4800 36
rect 4670 0 4700 26
rect 4770 0 4800 26
rect 4870 64 4900 117
rect 4970 64 5000 117
rect 4870 54 5000 64
rect 4870 20 4918 54
rect 4952 20 5000 54
rect 4870 10 5000 20
rect 4870 0 4900 10
rect 4970 0 5000 10
rect 5070 80 5100 117
rect 5170 80 5200 117
rect 5070 70 5200 80
rect 5070 36 5118 70
rect 5152 36 5200 70
rect 5070 26 5200 36
rect 5070 0 5100 26
rect 5170 0 5200 26
rect 5270 64 5300 117
rect 5370 64 5400 117
rect 5270 54 5400 64
rect 5270 20 5318 54
rect 5352 20 5400 54
rect 5270 10 5400 20
rect 5270 0 5300 10
rect 5370 0 5400 10
rect 5470 80 5500 117
rect 5570 80 5600 117
rect 5470 70 5600 80
rect 5470 36 5518 70
rect 5552 36 5600 70
rect 5470 26 5600 36
rect 5470 0 5500 26
rect 5570 0 5600 26
rect 5670 64 5700 117
rect 5770 64 5800 117
rect 5670 54 5800 64
rect 5670 20 5718 54
rect 5752 20 5800 54
rect 5670 10 5800 20
rect 5670 0 5700 10
rect 5770 0 5800 10
rect 5870 80 5900 117
rect 5970 80 6000 117
rect 5870 70 6000 80
rect 5870 36 5918 70
rect 5952 36 6000 70
rect 5870 26 6000 36
rect 5870 0 5900 26
rect 5970 0 6000 26
rect 6070 64 6100 117
rect 6170 64 6200 257
rect 6270 203 6300 257
rect 6370 203 6400 257
rect 6570 203 6600 257
rect 6670 203 6700 257
rect 6880 203 6910 257
rect 6980 203 7010 257
rect 7080 203 7110 257
rect 7180 203 7210 257
rect 7280 203 7310 257
rect 7380 203 7410 257
rect 6070 54 6200 64
rect 6070 20 6118 54
rect 6152 20 6200 54
rect 6070 10 6200 20
rect 6070 0 6100 10
rect 6170 0 6200 10
rect 6270 80 6300 117
rect 6370 80 6400 117
rect 6570 84 6600 117
rect 6670 84 6700 117
rect 6880 84 6910 117
rect 6980 84 7010 117
rect 7080 84 7110 117
rect 7180 84 7210 117
rect 7280 84 7310 117
rect 7380 84 7410 117
rect 6270 70 6400 80
rect 6270 36 6318 70
rect 6352 36 6400 70
rect 6270 26 6400 36
rect 6270 0 6300 26
rect 6370 0 6400 26
rect 6558 68 6612 84
rect 6558 34 6568 68
rect 6602 34 6612 68
rect 6558 18 6612 34
rect 6658 68 6712 84
rect 6658 34 6668 68
rect 6702 34 6712 68
rect 6658 18 6712 34
rect 6868 68 6922 84
rect 6868 34 6878 68
rect 6912 34 6922 68
rect 6868 18 6922 34
rect 6968 68 7022 84
rect 6968 34 6978 68
rect 7012 34 7022 68
rect 6968 18 7022 34
rect 7068 68 7122 84
rect 7068 34 7078 68
rect 7112 34 7122 68
rect 7068 18 7122 34
rect 7168 68 7222 84
rect 7168 34 7178 68
rect 7212 34 7222 68
rect 7168 18 7222 34
rect 7268 68 7322 84
rect 7268 34 7278 68
rect 7312 34 7322 68
rect 7268 18 7322 34
rect 7368 68 7422 84
rect 7368 34 7378 68
rect 7412 34 7422 68
rect 7368 18 7422 34
rect 6570 0 6600 18
rect 6670 0 6700 18
rect 6880 0 6910 18
rect 6980 0 7010 18
rect 7080 0 7110 18
rect 7180 0 7210 18
rect 7280 0 7310 18
rect 7380 0 7410 18
rect 8114 -90 8140 -60
rect 8290 -90 8416 -60
rect 8716 -90 8742 -60
rect 8800 -90 8826 -60
rect 9126 -90 9252 -60
rect 9402 -90 9428 -60
rect -30 -126 0 -100
rect 70 -126 100 -100
rect 170 -126 200 -100
rect 270 -126 300 -100
rect 370 -126 400 -100
rect 470 -126 500 -100
rect 570 -126 600 -100
rect 670 -126 700 -100
rect 770 -126 800 -100
rect 870 -126 900 -100
rect 970 -126 1000 -100
rect 1070 -126 1100 -100
rect 1170 -126 1200 -100
rect 1270 -126 1300 -100
rect 1370 -126 1400 -100
rect 1470 -126 1500 -100
rect 1570 -126 1600 -100
rect 1670 -126 1700 -100
rect 1770 -126 1800 -100
rect 1870 -126 1900 -100
rect 1970 -126 2000 -100
rect 2070 -126 2100 -100
rect 2170 -126 2200 -100
rect 2270 -126 2300 -100
rect 2370 -126 2400 -100
rect 2470 -126 2500 -100
rect 2570 -126 2600 -100
rect 2670 -126 2700 -100
rect 2770 -126 2800 -100
rect 2870 -126 2900 -100
rect 2970 -126 3000 -100
rect 3070 -126 3100 -100
rect 3170 -126 3200 -100
rect 3270 -126 3300 -100
rect 3370 -126 3400 -100
rect 3470 -126 3500 -100
rect 3570 -126 3600 -100
rect 3670 -126 3700 -100
rect 3770 -126 3800 -100
rect 3870 -126 3900 -100
rect 3970 -126 4000 -100
rect 4070 -126 4100 -100
rect 4170 -126 4200 -100
rect 4270 -126 4300 -100
rect 4370 -126 4400 -100
rect 4470 -126 4500 -100
rect 4570 -126 4600 -100
rect 4670 -126 4700 -100
rect 4770 -126 4800 -100
rect 4870 -126 4900 -100
rect 4970 -126 5000 -100
rect 5070 -126 5100 -100
rect 5170 -126 5200 -100
rect 5270 -126 5300 -100
rect 5370 -126 5400 -100
rect 5470 -126 5500 -100
rect 5570 -126 5600 -100
rect 5670 -126 5700 -100
rect 5770 -126 5800 -100
rect 5870 -126 5900 -100
rect 5970 -126 6000 -100
rect 6070 -126 6100 -100
rect 6170 -126 6200 -100
rect 6270 -126 6300 -100
rect 8306 -109 8400 -90
rect 8306 -143 8334 -109
rect 8368 -143 8400 -109
rect 8306 -160 8400 -143
rect 9142 -109 9236 -90
rect 9142 -143 9174 -109
rect 9208 -143 9236 -109
rect 9142 -160 9236 -143
rect 8114 -190 8140 -160
rect 8290 -190 8416 -160
rect 8716 -190 8742 -160
rect 8800 -190 8826 -160
rect 9126 -190 9252 -160
rect 9402 -190 9428 -160
rect -30 -226 0 -210
rect 70 -226 100 -210
rect -30 -248 100 -226
rect -30 -282 18 -248
rect 52 -282 100 -248
rect -30 -314 100 -282
rect -30 -330 0 -314
rect 70 -330 100 -314
rect 170 -226 200 -210
rect 270 -226 300 -210
rect 170 -248 300 -226
rect 170 -282 218 -248
rect 252 -282 300 -248
rect 170 -314 300 -282
rect 170 -330 200 -314
rect 270 -330 300 -314
rect 370 -226 400 -210
rect 470 -226 500 -210
rect 370 -248 500 -226
rect 370 -282 418 -248
rect 452 -282 500 -248
rect 370 -314 500 -282
rect 370 -330 400 -314
rect 470 -330 500 -314
rect 570 -226 600 -210
rect 670 -226 700 -210
rect 570 -248 700 -226
rect 570 -282 618 -248
rect 652 -282 700 -248
rect 570 -314 700 -282
rect 570 -330 600 -314
rect 670 -330 700 -314
rect 770 -226 800 -210
rect 870 -226 900 -210
rect 770 -248 900 -226
rect 770 -282 818 -248
rect 852 -282 900 -248
rect 770 -314 900 -282
rect 770 -330 800 -314
rect 870 -330 900 -314
rect 970 -226 1000 -210
rect 1070 -226 1100 -210
rect 970 -248 1100 -226
rect 970 -282 1018 -248
rect 1052 -282 1100 -248
rect 970 -314 1100 -282
rect 970 -330 1000 -314
rect 1070 -330 1100 -314
rect 1170 -226 1200 -210
rect 1270 -226 1300 -210
rect 1170 -248 1300 -226
rect 1170 -282 1218 -248
rect 1252 -282 1300 -248
rect 1170 -314 1300 -282
rect 1170 -330 1200 -314
rect 1270 -330 1300 -314
rect 1370 -226 1400 -210
rect 1470 -226 1500 -210
rect 1370 -248 1500 -226
rect 1370 -282 1418 -248
rect 1452 -282 1500 -248
rect 1370 -314 1500 -282
rect 1370 -330 1400 -314
rect 1470 -330 1500 -314
rect 1570 -226 1600 -210
rect 1670 -226 1700 -210
rect 1570 -248 1700 -226
rect 1570 -282 1618 -248
rect 1652 -282 1700 -248
rect 1570 -314 1700 -282
rect 1570 -330 1600 -314
rect 1670 -330 1700 -314
rect 1770 -226 1800 -210
rect 1870 -226 1900 -210
rect 1770 -248 1900 -226
rect 1770 -282 1818 -248
rect 1852 -282 1900 -248
rect 1770 -314 1900 -282
rect 1770 -330 1800 -314
rect 1870 -330 1900 -314
rect 1970 -226 2000 -210
rect 2070 -226 2100 -210
rect 1970 -248 2100 -226
rect 1970 -282 2018 -248
rect 2052 -282 2100 -248
rect 1970 -314 2100 -282
rect 1970 -330 2000 -314
rect 2070 -330 2100 -314
rect 2170 -226 2200 -210
rect 2270 -226 2300 -210
rect 2170 -248 2300 -226
rect 2170 -282 2218 -248
rect 2252 -282 2300 -248
rect 2170 -314 2300 -282
rect 2170 -330 2200 -314
rect 2270 -330 2300 -314
rect 2370 -226 2400 -210
rect 2470 -226 2500 -210
rect 2370 -248 2500 -226
rect 2370 -282 2418 -248
rect 2452 -282 2500 -248
rect 2370 -314 2500 -282
rect 2370 -330 2400 -314
rect 2470 -330 2500 -314
rect 2570 -226 2600 -210
rect 2670 -226 2700 -210
rect 2570 -248 2700 -226
rect 2570 -282 2618 -248
rect 2652 -282 2700 -248
rect 2570 -314 2700 -282
rect 2570 -330 2600 -314
rect 2670 -330 2700 -314
rect 2770 -226 2800 -210
rect 2870 -226 2900 -210
rect 2770 -248 2900 -226
rect 2770 -282 2818 -248
rect 2852 -282 2900 -248
rect 2770 -314 2900 -282
rect 2770 -330 2800 -314
rect 2870 -330 2900 -314
rect 2970 -226 3000 -210
rect 3070 -226 3100 -210
rect 2970 -248 3100 -226
rect 2970 -282 3018 -248
rect 3052 -282 3100 -248
rect 2970 -314 3100 -282
rect 2970 -330 3000 -314
rect 3070 -330 3100 -314
rect 3170 -226 3200 -210
rect 3270 -226 3300 -210
rect 3170 -248 3300 -226
rect 3170 -282 3218 -248
rect 3252 -282 3300 -248
rect 3170 -314 3300 -282
rect 3170 -330 3200 -314
rect 3270 -330 3300 -314
rect 3370 -226 3400 -210
rect 3470 -226 3500 -210
rect 3370 -248 3500 -226
rect 3370 -282 3418 -248
rect 3452 -282 3500 -248
rect 3370 -314 3500 -282
rect 3370 -330 3400 -314
rect 3470 -330 3500 -314
rect 3570 -226 3600 -210
rect 3670 -226 3700 -210
rect 3570 -248 3700 -226
rect 3570 -282 3618 -248
rect 3652 -282 3700 -248
rect 3570 -314 3700 -282
rect 3570 -330 3600 -314
rect 3670 -330 3700 -314
rect 3770 -226 3800 -210
rect 3870 -226 3900 -210
rect 3770 -248 3900 -226
rect 3770 -282 3818 -248
rect 3852 -282 3900 -248
rect 3770 -314 3900 -282
rect 3770 -330 3800 -314
rect 3870 -330 3900 -314
rect 3970 -226 4000 -210
rect 4070 -226 4100 -210
rect 3970 -248 4100 -226
rect 3970 -282 4018 -248
rect 4052 -282 4100 -248
rect 3970 -314 4100 -282
rect 3970 -330 4000 -314
rect 4070 -330 4100 -314
rect 4170 -226 4200 -210
rect 4270 -226 4300 -210
rect 4170 -248 4300 -226
rect 4170 -282 4218 -248
rect 4252 -282 4300 -248
rect 4170 -314 4300 -282
rect 4170 -330 4200 -314
rect 4270 -330 4300 -314
rect 4370 -226 4400 -210
rect 4470 -226 4500 -210
rect 4370 -248 4500 -226
rect 4370 -282 4418 -248
rect 4452 -282 4500 -248
rect 4370 -314 4500 -282
rect 4370 -330 4400 -314
rect 4470 -330 4500 -314
rect 4570 -226 4600 -210
rect 4670 -226 4700 -210
rect 4570 -248 4700 -226
rect 4570 -282 4618 -248
rect 4652 -282 4700 -248
rect 4570 -314 4700 -282
rect 4570 -330 4600 -314
rect 4670 -330 4700 -314
rect 4770 -226 4800 -210
rect 4870 -226 4900 -210
rect 4770 -248 4900 -226
rect 4770 -282 4818 -248
rect 4852 -282 4900 -248
rect 4770 -314 4900 -282
rect 4770 -330 4800 -314
rect 4870 -330 4900 -314
rect 4970 -226 5000 -210
rect 5070 -226 5100 -210
rect 4970 -248 5100 -226
rect 4970 -282 5018 -248
rect 5052 -282 5100 -248
rect 4970 -314 5100 -282
rect 4970 -330 5000 -314
rect 5070 -330 5100 -314
rect 5170 -226 5200 -210
rect 5270 -226 5300 -210
rect 5170 -248 5300 -226
rect 5170 -282 5218 -248
rect 5252 -282 5300 -248
rect 5170 -314 5300 -282
rect 5170 -330 5200 -314
rect 5270 -330 5300 -314
rect 5370 -226 5400 -210
rect 5470 -226 5500 -210
rect 5370 -248 5500 -226
rect 5370 -282 5418 -248
rect 5452 -282 5500 -248
rect 5370 -314 5500 -282
rect 5370 -330 5400 -314
rect 5470 -330 5500 -314
rect 5570 -226 5600 -210
rect 5670 -226 5700 -210
rect 5570 -248 5700 -226
rect 5570 -282 5618 -248
rect 5652 -282 5700 -248
rect 5570 -314 5700 -282
rect 5570 -330 5600 -314
rect 5670 -330 5700 -314
rect 5770 -226 5800 -210
rect 5870 -226 5900 -210
rect 5770 -248 5900 -226
rect 5770 -282 5818 -248
rect 5852 -282 5900 -248
rect 5770 -314 5900 -282
rect 5770 -330 5800 -314
rect 5870 -330 5900 -314
rect 5970 -226 6000 -210
rect 6070 -226 6100 -210
rect 5970 -248 6100 -226
rect 5970 -282 6018 -248
rect 6052 -282 6100 -248
rect 5970 -314 6100 -282
rect 5970 -330 6000 -314
rect 6070 -330 6100 -314
rect 6170 -226 6200 -210
rect 6270 -226 6300 -210
rect 6170 -248 6300 -226
rect 6170 -282 6218 -248
rect 6252 -282 6300 -248
rect 6170 -314 6300 -282
rect 8114 -290 8140 -260
rect 8290 -290 8416 -260
rect 8716 -290 8742 -260
rect 8800 -290 8826 -260
rect 9126 -290 9252 -260
rect 9402 -290 9428 -260
rect 6170 -330 6200 -314
rect 6270 -330 6300 -314
rect 8306 -309 8400 -290
rect 8306 -343 8334 -309
rect 8368 -343 8400 -309
rect 8306 -360 8400 -343
rect 9142 -309 9236 -290
rect 9142 -343 9174 -309
rect 9208 -343 9236 -309
rect 9142 -360 9236 -343
rect 8114 -390 8140 -360
rect 8290 -390 8416 -360
rect 8716 -390 8742 -360
rect 8800 -390 8826 -360
rect 9126 -390 9252 -360
rect 9402 -390 9428 -360
rect 8114 -490 8140 -460
rect 8290 -490 8416 -460
rect 8716 -490 8742 -460
rect 8800 -490 8826 -460
rect 9126 -490 9252 -460
rect 9402 -490 9428 -460
rect -30 -524 0 -498
rect 70 -524 100 -498
rect 170 -524 200 -498
rect 270 -524 300 -498
rect 370 -524 400 -498
rect 470 -524 500 -498
rect 570 -524 600 -498
rect 670 -524 700 -498
rect 770 -524 800 -498
rect 870 -524 900 -498
rect 970 -524 1000 -498
rect 1070 -524 1100 -498
rect 1170 -524 1200 -498
rect 1270 -524 1300 -498
rect 1370 -524 1400 -498
rect 1470 -524 1500 -498
rect 1570 -524 1600 -498
rect 1670 -524 1700 -498
rect 1770 -524 1800 -498
rect 1870 -524 1900 -498
rect 1970 -524 2000 -498
rect 2070 -524 2100 -498
rect 2170 -524 2200 -498
rect 2270 -524 2300 -498
rect 2370 -524 2400 -498
rect 2470 -524 2500 -498
rect 2570 -524 2600 -498
rect 2670 -524 2700 -498
rect 2770 -524 2800 -498
rect 2870 -524 2900 -498
rect 2970 -524 3000 -498
rect 3070 -524 3100 -498
rect 3170 -524 3200 -498
rect 3270 -524 3300 -498
rect 3370 -524 3400 -498
rect 3470 -524 3500 -498
rect 3570 -524 3600 -498
rect 3670 -524 3700 -498
rect 3770 -524 3800 -498
rect 3870 -524 3900 -498
rect 3970 -524 4000 -498
rect 4070 -524 4100 -498
rect 4170 -524 4200 -498
rect 4270 -524 4300 -498
rect 4370 -524 4400 -498
rect 4470 -524 4500 -498
rect 4570 -524 4600 -498
rect 4670 -524 4700 -498
rect 4770 -524 4800 -498
rect 4870 -524 4900 -498
rect 4970 -524 5000 -498
rect 5070 -524 5100 -498
rect 5170 -524 5200 -498
rect 5270 -524 5300 -498
rect 5370 -524 5400 -498
rect 5470 -524 5500 -498
rect 5570 -524 5600 -498
rect 5670 -524 5700 -498
rect 5770 -524 5800 -498
rect 5870 -524 5900 -498
rect 5970 -524 6000 -498
rect 6070 -524 6100 -498
rect 6170 -524 6200 -498
rect 6270 -524 6300 -498
rect 8306 -509 8400 -490
rect 8306 -543 8334 -509
rect 8368 -543 8400 -509
rect 8306 -560 8400 -543
rect 9142 -509 9236 -490
rect 9142 -543 9174 -509
rect 9208 -543 9236 -509
rect 9142 -560 9236 -543
rect 15 -577 107 -567
rect 15 -611 44 -577
rect 78 -611 107 -577
rect 15 -658 107 -611
rect 163 -577 255 -567
rect 163 -611 192 -577
rect 226 -611 255 -577
rect 415 -577 507 -567
rect 163 -658 255 -611
rect 415 -611 444 -577
rect 478 -611 507 -577
rect 415 -658 507 -611
rect 563 -577 655 -567
rect 563 -611 592 -577
rect 626 -611 655 -577
rect 815 -577 907 -567
rect 563 -658 655 -611
rect 815 -611 844 -577
rect 878 -611 907 -577
rect 815 -658 907 -611
rect 963 -577 1055 -567
rect 963 -611 992 -577
rect 1026 -611 1055 -577
rect 1215 -577 1307 -567
rect 963 -658 1055 -611
rect 1215 -611 1244 -577
rect 1278 -611 1307 -577
rect 1215 -658 1307 -611
rect 1363 -577 1455 -567
rect 1363 -611 1392 -577
rect 1426 -611 1455 -577
rect 1615 -577 1707 -567
rect 1363 -658 1455 -611
rect 1615 -611 1644 -577
rect 1678 -611 1707 -577
rect 1615 -658 1707 -611
rect 1763 -577 1855 -567
rect 1763 -611 1792 -577
rect 1826 -611 1855 -577
rect 2015 -577 2107 -567
rect 1763 -658 1855 -611
rect 2015 -611 2044 -577
rect 2078 -611 2107 -577
rect 2015 -658 2107 -611
rect 2163 -577 2255 -567
rect 2163 -611 2192 -577
rect 2226 -611 2255 -577
rect 2415 -577 2507 -567
rect 2163 -658 2255 -611
rect 2415 -611 2444 -577
rect 2478 -611 2507 -577
rect 2415 -658 2507 -611
rect 2563 -577 2655 -567
rect 2563 -611 2592 -577
rect 2626 -611 2655 -577
rect 2815 -577 2907 -567
rect 2563 -658 2655 -611
rect 2815 -611 2844 -577
rect 2878 -611 2907 -577
rect 2815 -658 2907 -611
rect 2963 -577 3055 -567
rect 2963 -611 2992 -577
rect 3026 -611 3055 -577
rect 3215 -577 3307 -567
rect 2963 -658 3055 -611
rect 3215 -611 3244 -577
rect 3278 -611 3307 -577
rect 3215 -658 3307 -611
rect 3363 -577 3455 -567
rect 3363 -611 3392 -577
rect 3426 -611 3455 -577
rect 3615 -577 3707 -567
rect 3363 -658 3455 -611
rect 3615 -611 3644 -577
rect 3678 -611 3707 -577
rect 3615 -658 3707 -611
rect 3763 -577 3855 -567
rect 3763 -611 3792 -577
rect 3826 -611 3855 -577
rect 4015 -577 4107 -567
rect 3763 -658 3855 -611
rect 4015 -611 4044 -577
rect 4078 -611 4107 -577
rect 4015 -658 4107 -611
rect 4163 -577 4255 -567
rect 4163 -611 4192 -577
rect 4226 -611 4255 -577
rect 4415 -577 4507 -567
rect 4163 -658 4255 -611
rect 4415 -611 4444 -577
rect 4478 -611 4507 -577
rect 4415 -658 4507 -611
rect 4563 -577 4655 -567
rect 4563 -611 4592 -577
rect 4626 -611 4655 -577
rect 4815 -577 4907 -567
rect 4563 -658 4655 -611
rect 4815 -611 4844 -577
rect 4878 -611 4907 -577
rect 4815 -658 4907 -611
rect 4963 -577 5055 -567
rect 4963 -611 4992 -577
rect 5026 -611 5055 -577
rect 5215 -577 5307 -567
rect 4963 -658 5055 -611
rect 5215 -611 5244 -577
rect 5278 -611 5307 -577
rect 5215 -658 5307 -611
rect 5363 -577 5455 -567
rect 5363 -611 5392 -577
rect 5426 -611 5455 -577
rect 5615 -577 5707 -567
rect 5363 -658 5455 -611
rect 5615 -611 5644 -577
rect 5678 -611 5707 -577
rect 5615 -658 5707 -611
rect 5763 -577 5855 -567
rect 5763 -611 5792 -577
rect 5826 -611 5855 -577
rect 6015 -577 6107 -567
rect 5763 -658 5855 -611
rect 6015 -611 6044 -577
rect 6078 -611 6107 -577
rect 6015 -658 6107 -611
rect 6163 -577 6255 -567
rect 6163 -611 6192 -577
rect 6226 -611 6255 -577
rect 8114 -590 8140 -560
rect 8290 -590 8416 -560
rect 8716 -590 8742 -560
rect 8800 -590 8826 -560
rect 9126 -590 9252 -560
rect 9402 -590 9428 -560
rect 6163 -658 6255 -611
rect 8114 -690 8140 -660
rect 8290 -690 8416 -660
rect 8716 -690 8742 -660
rect 8800 -690 8826 -660
rect 9126 -690 9252 -660
rect 9402 -690 9428 -660
rect 15 -768 107 -742
rect 163 -768 255 -742
rect 415 -768 507 -742
rect 563 -768 655 -742
rect 815 -768 907 -742
rect 963 -768 1055 -742
rect 1215 -768 1307 -742
rect 1363 -768 1455 -742
rect 1615 -768 1707 -742
rect 1763 -768 1855 -742
rect 2015 -768 2107 -742
rect 2163 -768 2255 -742
rect 2415 -768 2507 -742
rect 2563 -768 2655 -742
rect 2815 -768 2907 -742
rect 2963 -768 3055 -742
rect 3215 -768 3307 -742
rect 3363 -768 3455 -742
rect 3615 -768 3707 -742
rect 3763 -768 3855 -742
rect 4015 -768 4107 -742
rect 4163 -768 4255 -742
rect 4415 -768 4507 -742
rect 4563 -768 4655 -742
rect 4815 -768 4907 -742
rect 4963 -768 5055 -742
rect 5215 -768 5307 -742
rect 5363 -768 5455 -742
rect 5615 -768 5707 -742
rect 5763 -768 5855 -742
rect 6015 -768 6107 -742
rect 6163 -768 6255 -742
rect 8306 -709 8400 -690
rect 8306 -743 8334 -709
rect 8368 -743 8400 -709
rect 8306 -760 8400 -743
rect 9142 -709 9236 -690
rect 9142 -743 9174 -709
rect 9208 -743 9236 -709
rect 9142 -760 9236 -743
rect 8114 -790 8140 -760
rect 8290 -790 8416 -760
rect 8716 -790 8742 -760
rect 8800 -790 8826 -760
rect 9126 -790 9252 -760
rect 9402 -790 9428 -760
rect -98 -908 -32 -898
rect -98 -910 -82 -908
rect -106 -940 -82 -910
rect -98 -942 -82 -940
rect -48 -910 -32 -908
rect 702 -908 768 -898
rect 702 -910 718 -908
rect -48 -940 -10 -910
rect 108 -940 162 -910
rect 280 -940 390 -910
rect 508 -940 562 -910
rect 680 -940 718 -910
rect -48 -942 -32 -940
rect -98 -952 -32 -942
rect -98 -1008 -32 -998
rect -98 -1010 -82 -1008
rect -106 -1040 -82 -1010
rect -98 -1042 -82 -1040
rect -48 -1010 -32 -1008
rect 702 -942 718 -940
rect 752 -910 768 -908
rect 1502 -908 1568 -898
rect 1502 -910 1518 -908
rect 752 -940 790 -910
rect 908 -940 962 -910
rect 1080 -940 1190 -910
rect 1308 -940 1362 -910
rect 1480 -940 1518 -910
rect 752 -942 768 -940
rect 702 -952 768 -942
rect 702 -1008 768 -998
rect 702 -1010 718 -1008
rect -48 -1040 -10 -1010
rect 108 -1040 162 -1010
rect 280 -1040 390 -1010
rect 508 -1040 562 -1010
rect 680 -1040 718 -1010
rect -48 -1042 -32 -1040
rect -98 -1052 -32 -1042
rect -98 -1108 -32 -1098
rect -98 -1110 -82 -1108
rect -106 -1140 -82 -1110
rect -98 -1142 -82 -1140
rect -48 -1110 -32 -1108
rect 702 -1042 718 -1040
rect 752 -1010 768 -1008
rect 1502 -942 1518 -940
rect 1552 -910 1568 -908
rect 2302 -908 2368 -898
rect 2302 -910 2318 -908
rect 1552 -940 1590 -910
rect 1708 -940 1762 -910
rect 1880 -940 1990 -910
rect 2108 -940 2162 -910
rect 2280 -940 2318 -910
rect 1552 -942 1568 -940
rect 1502 -952 1568 -942
rect 1502 -1008 1568 -998
rect 1502 -1010 1518 -1008
rect 752 -1040 790 -1010
rect 908 -1040 962 -1010
rect 1080 -1040 1190 -1010
rect 1308 -1040 1362 -1010
rect 1480 -1040 1518 -1010
rect 752 -1042 768 -1040
rect 702 -1052 768 -1042
rect 702 -1108 768 -1098
rect 702 -1110 718 -1108
rect -48 -1140 -10 -1110
rect 108 -1140 162 -1110
rect 280 -1140 390 -1110
rect 508 -1140 562 -1110
rect 680 -1140 718 -1110
rect -48 -1142 -32 -1140
rect -98 -1152 -32 -1142
rect -98 -1208 -32 -1198
rect -98 -1210 -82 -1208
rect -106 -1240 -82 -1210
rect -98 -1242 -82 -1240
rect -48 -1210 -32 -1208
rect 702 -1142 718 -1140
rect 752 -1110 768 -1108
rect 1502 -1042 1518 -1040
rect 1552 -1010 1568 -1008
rect 2302 -942 2318 -940
rect 2352 -910 2368 -908
rect 3102 -908 3168 -898
rect 3102 -910 3118 -908
rect 2352 -940 2390 -910
rect 2508 -940 2562 -910
rect 2680 -940 2790 -910
rect 2908 -940 2962 -910
rect 3080 -940 3118 -910
rect 2352 -942 2368 -940
rect 2302 -952 2368 -942
rect 2302 -1008 2368 -998
rect 2302 -1010 2318 -1008
rect 1552 -1040 1590 -1010
rect 1708 -1040 1762 -1010
rect 1880 -1040 1990 -1010
rect 2108 -1040 2162 -1010
rect 2280 -1040 2318 -1010
rect 1552 -1042 1568 -1040
rect 1502 -1052 1568 -1042
rect 1502 -1108 1568 -1098
rect 1502 -1110 1518 -1108
rect 752 -1140 790 -1110
rect 908 -1140 962 -1110
rect 1080 -1140 1190 -1110
rect 1308 -1140 1362 -1110
rect 1480 -1140 1518 -1110
rect 752 -1142 768 -1140
rect 702 -1152 768 -1142
rect 702 -1208 768 -1198
rect 702 -1210 718 -1208
rect -48 -1240 -10 -1210
rect 108 -1240 162 -1210
rect 280 -1240 390 -1210
rect 508 -1240 562 -1210
rect 680 -1240 718 -1210
rect -48 -1242 -32 -1240
rect -98 -1252 -32 -1242
rect -98 -1308 -32 -1298
rect -98 -1310 -82 -1308
rect -106 -1340 -82 -1310
rect -98 -1342 -82 -1340
rect -48 -1310 -32 -1308
rect 702 -1242 718 -1240
rect 752 -1210 768 -1208
rect 1502 -1142 1518 -1140
rect 1552 -1110 1568 -1108
rect 2302 -1042 2318 -1040
rect 2352 -1010 2368 -1008
rect 3102 -942 3118 -940
rect 3152 -910 3168 -908
rect 3902 -908 3968 -898
rect 3902 -910 3918 -908
rect 3152 -940 3190 -910
rect 3308 -940 3362 -910
rect 3480 -940 3590 -910
rect 3708 -940 3762 -910
rect 3880 -940 3918 -910
rect 3152 -942 3168 -940
rect 3102 -952 3168 -942
rect 3102 -1008 3168 -998
rect 3102 -1010 3118 -1008
rect 2352 -1040 2390 -1010
rect 2508 -1040 2562 -1010
rect 2680 -1040 2790 -1010
rect 2908 -1040 2962 -1010
rect 3080 -1040 3118 -1010
rect 2352 -1042 2368 -1040
rect 2302 -1052 2368 -1042
rect 2302 -1108 2368 -1098
rect 2302 -1110 2318 -1108
rect 1552 -1140 1590 -1110
rect 1708 -1140 1762 -1110
rect 1880 -1140 1990 -1110
rect 2108 -1140 2162 -1110
rect 2280 -1140 2318 -1110
rect 1552 -1142 1568 -1140
rect 1502 -1152 1568 -1142
rect 1502 -1208 1568 -1198
rect 1502 -1210 1518 -1208
rect 752 -1240 790 -1210
rect 908 -1240 962 -1210
rect 1080 -1240 1190 -1210
rect 1308 -1240 1362 -1210
rect 1480 -1240 1518 -1210
rect 752 -1242 768 -1240
rect 702 -1252 768 -1242
rect 702 -1308 768 -1298
rect 702 -1310 718 -1308
rect -48 -1340 -10 -1310
rect 108 -1340 162 -1310
rect 280 -1340 390 -1310
rect 508 -1340 562 -1310
rect 680 -1340 718 -1310
rect -48 -1342 -32 -1340
rect -98 -1352 -32 -1342
rect -98 -1408 -32 -1398
rect -98 -1410 -82 -1408
rect -106 -1440 -82 -1410
rect -98 -1442 -82 -1440
rect -48 -1410 -32 -1408
rect 702 -1342 718 -1340
rect 752 -1310 768 -1308
rect 1502 -1242 1518 -1240
rect 1552 -1210 1568 -1208
rect 2302 -1142 2318 -1140
rect 2352 -1110 2368 -1108
rect 3102 -1042 3118 -1040
rect 3152 -1010 3168 -1008
rect 3902 -942 3918 -940
rect 3952 -910 3968 -908
rect 4702 -908 4768 -898
rect 4702 -910 4718 -908
rect 3952 -940 3990 -910
rect 4108 -940 4162 -910
rect 4280 -940 4390 -910
rect 4508 -940 4562 -910
rect 4680 -940 4718 -910
rect 3952 -942 3968 -940
rect 3902 -952 3968 -942
rect 3902 -1008 3968 -998
rect 3902 -1010 3918 -1008
rect 3152 -1040 3190 -1010
rect 3308 -1040 3362 -1010
rect 3480 -1040 3590 -1010
rect 3708 -1040 3762 -1010
rect 3880 -1040 3918 -1010
rect 3152 -1042 3168 -1040
rect 3102 -1052 3168 -1042
rect 3102 -1108 3168 -1098
rect 3102 -1110 3118 -1108
rect 2352 -1140 2390 -1110
rect 2508 -1140 2562 -1110
rect 2680 -1140 2790 -1110
rect 2908 -1140 2962 -1110
rect 3080 -1140 3118 -1110
rect 2352 -1142 2368 -1140
rect 2302 -1152 2368 -1142
rect 2302 -1208 2368 -1198
rect 2302 -1210 2318 -1208
rect 1552 -1240 1590 -1210
rect 1708 -1240 1762 -1210
rect 1880 -1240 1990 -1210
rect 2108 -1240 2162 -1210
rect 2280 -1240 2318 -1210
rect 1552 -1242 1568 -1240
rect 1502 -1252 1568 -1242
rect 1502 -1308 1568 -1298
rect 1502 -1310 1518 -1308
rect 752 -1340 790 -1310
rect 908 -1340 962 -1310
rect 1080 -1340 1190 -1310
rect 1308 -1340 1362 -1310
rect 1480 -1340 1518 -1310
rect 752 -1342 768 -1340
rect 702 -1352 768 -1342
rect 702 -1408 768 -1398
rect 702 -1410 718 -1408
rect -48 -1440 -10 -1410
rect 108 -1440 162 -1410
rect 280 -1440 390 -1410
rect 508 -1440 562 -1410
rect 680 -1440 718 -1410
rect -48 -1442 -32 -1440
rect -98 -1452 -32 -1442
rect -98 -1508 -32 -1498
rect -98 -1510 -82 -1508
rect -106 -1540 -82 -1510
rect -98 -1542 -82 -1540
rect -48 -1510 -32 -1508
rect 702 -1442 718 -1440
rect 752 -1410 768 -1408
rect 1502 -1342 1518 -1340
rect 1552 -1310 1568 -1308
rect 2302 -1242 2318 -1240
rect 2352 -1210 2368 -1208
rect 3102 -1142 3118 -1140
rect 3152 -1110 3168 -1108
rect 3902 -1042 3918 -1040
rect 3952 -1010 3968 -1008
rect 4702 -942 4718 -940
rect 4752 -910 4768 -908
rect 5502 -908 5568 -898
rect 5502 -910 5518 -908
rect 4752 -940 4790 -910
rect 4908 -940 4962 -910
rect 5080 -940 5190 -910
rect 5308 -940 5362 -910
rect 5480 -940 5518 -910
rect 4752 -942 4768 -940
rect 4702 -952 4768 -942
rect 4702 -1008 4768 -998
rect 4702 -1010 4718 -1008
rect 3952 -1040 3990 -1010
rect 4108 -1040 4162 -1010
rect 4280 -1040 4390 -1010
rect 4508 -1040 4562 -1010
rect 4680 -1040 4718 -1010
rect 3952 -1042 3968 -1040
rect 3902 -1052 3968 -1042
rect 3902 -1108 3968 -1098
rect 3902 -1110 3918 -1108
rect 3152 -1140 3190 -1110
rect 3308 -1140 3362 -1110
rect 3480 -1140 3590 -1110
rect 3708 -1140 3762 -1110
rect 3880 -1140 3918 -1110
rect 3152 -1142 3168 -1140
rect 3102 -1152 3168 -1142
rect 3102 -1208 3168 -1198
rect 3102 -1210 3118 -1208
rect 2352 -1240 2390 -1210
rect 2508 -1240 2562 -1210
rect 2680 -1240 2790 -1210
rect 2908 -1240 2962 -1210
rect 3080 -1240 3118 -1210
rect 2352 -1242 2368 -1240
rect 2302 -1252 2368 -1242
rect 2302 -1308 2368 -1298
rect 2302 -1310 2318 -1308
rect 1552 -1340 1590 -1310
rect 1708 -1340 1762 -1310
rect 1880 -1340 1990 -1310
rect 2108 -1340 2162 -1310
rect 2280 -1340 2318 -1310
rect 1552 -1342 1568 -1340
rect 1502 -1352 1568 -1342
rect 1502 -1408 1568 -1398
rect 1502 -1410 1518 -1408
rect 752 -1440 790 -1410
rect 908 -1440 962 -1410
rect 1080 -1440 1190 -1410
rect 1308 -1440 1362 -1410
rect 1480 -1440 1518 -1410
rect 752 -1442 768 -1440
rect 702 -1452 768 -1442
rect 702 -1508 768 -1498
rect 702 -1510 718 -1508
rect -48 -1540 -10 -1510
rect 108 -1540 162 -1510
rect 280 -1540 390 -1510
rect 508 -1540 562 -1510
rect 680 -1540 718 -1510
rect -48 -1542 -32 -1540
rect -98 -1552 -32 -1542
rect -98 -1608 -32 -1598
rect -98 -1610 -82 -1608
rect -106 -1640 -82 -1610
rect -98 -1642 -82 -1640
rect -48 -1610 -32 -1608
rect 702 -1542 718 -1540
rect 752 -1510 768 -1508
rect 1502 -1442 1518 -1440
rect 1552 -1410 1568 -1408
rect 2302 -1342 2318 -1340
rect 2352 -1310 2368 -1308
rect 3102 -1242 3118 -1240
rect 3152 -1210 3168 -1208
rect 3902 -1142 3918 -1140
rect 3952 -1110 3968 -1108
rect 4702 -1042 4718 -1040
rect 4752 -1010 4768 -1008
rect 5502 -942 5518 -940
rect 5552 -910 5568 -908
rect 8114 -890 8140 -860
rect 8290 -890 8416 -860
rect 8716 -890 8742 -860
rect 8800 -890 8826 -860
rect 9126 -890 9252 -860
rect 9402 -890 9428 -860
rect 6302 -908 6368 -898
rect 6302 -910 6318 -908
rect 5552 -940 5590 -910
rect 5708 -940 5762 -910
rect 5880 -940 5990 -910
rect 6108 -940 6162 -910
rect 6280 -940 6318 -910
rect 5552 -942 5568 -940
rect 5502 -952 5568 -942
rect 5502 -1008 5568 -998
rect 5502 -1010 5518 -1008
rect 4752 -1040 4790 -1010
rect 4908 -1040 4962 -1010
rect 5080 -1040 5190 -1010
rect 5308 -1040 5362 -1010
rect 5480 -1040 5518 -1010
rect 4752 -1042 4768 -1040
rect 4702 -1052 4768 -1042
rect 4702 -1108 4768 -1098
rect 4702 -1110 4718 -1108
rect 3952 -1140 3990 -1110
rect 4108 -1140 4162 -1110
rect 4280 -1140 4390 -1110
rect 4508 -1140 4562 -1110
rect 4680 -1140 4718 -1110
rect 3952 -1142 3968 -1140
rect 3902 -1152 3968 -1142
rect 3902 -1208 3968 -1198
rect 3902 -1210 3918 -1208
rect 3152 -1240 3190 -1210
rect 3308 -1240 3362 -1210
rect 3480 -1240 3590 -1210
rect 3708 -1240 3762 -1210
rect 3880 -1240 3918 -1210
rect 3152 -1242 3168 -1240
rect 3102 -1252 3168 -1242
rect 3102 -1308 3168 -1298
rect 3102 -1310 3118 -1308
rect 2352 -1340 2390 -1310
rect 2508 -1340 2562 -1310
rect 2680 -1340 2790 -1310
rect 2908 -1340 2962 -1310
rect 3080 -1340 3118 -1310
rect 2352 -1342 2368 -1340
rect 2302 -1352 2368 -1342
rect 2302 -1408 2368 -1398
rect 2302 -1410 2318 -1408
rect 1552 -1440 1590 -1410
rect 1708 -1440 1762 -1410
rect 1880 -1440 1990 -1410
rect 2108 -1440 2162 -1410
rect 2280 -1440 2318 -1410
rect 1552 -1442 1568 -1440
rect 1502 -1452 1568 -1442
rect 1502 -1508 1568 -1498
rect 1502 -1510 1518 -1508
rect 752 -1540 790 -1510
rect 908 -1540 962 -1510
rect 1080 -1540 1190 -1510
rect 1308 -1540 1362 -1510
rect 1480 -1540 1518 -1510
rect 752 -1542 768 -1540
rect 702 -1552 768 -1542
rect 702 -1608 768 -1598
rect 702 -1610 718 -1608
rect -48 -1640 -10 -1610
rect 108 -1640 162 -1610
rect 280 -1640 390 -1610
rect 508 -1640 562 -1610
rect 680 -1640 718 -1610
rect -48 -1642 -32 -1640
rect -98 -1652 -32 -1642
rect -98 -1708 -32 -1698
rect -98 -1710 -82 -1708
rect -106 -1740 -82 -1710
rect -98 -1742 -82 -1740
rect -48 -1710 -32 -1708
rect 702 -1642 718 -1640
rect 752 -1610 768 -1608
rect 1502 -1542 1518 -1540
rect 1552 -1510 1568 -1508
rect 2302 -1442 2318 -1440
rect 2352 -1410 2368 -1408
rect 3102 -1342 3118 -1340
rect 3152 -1310 3168 -1308
rect 3902 -1242 3918 -1240
rect 3952 -1210 3968 -1208
rect 4702 -1142 4718 -1140
rect 4752 -1110 4768 -1108
rect 5502 -1042 5518 -1040
rect 5552 -1010 5568 -1008
rect 6302 -942 6318 -940
rect 6352 -910 6368 -908
rect 6352 -940 6376 -910
rect 6352 -942 6368 -940
rect 6302 -952 6368 -942
rect 8306 -909 8400 -890
rect 8306 -943 8334 -909
rect 8368 -943 8400 -909
rect 8306 -960 8400 -943
rect 9142 -909 9236 -890
rect 9142 -943 9174 -909
rect 9208 -943 9236 -909
rect 9142 -960 9236 -943
rect 8114 -990 8140 -960
rect 8290 -990 8416 -960
rect 8716 -990 8742 -960
rect 8800 -990 8826 -960
rect 9126 -990 9252 -960
rect 9402 -990 9428 -960
rect 6302 -1008 6368 -998
rect 6302 -1010 6318 -1008
rect 5552 -1040 5590 -1010
rect 5708 -1040 5762 -1010
rect 5880 -1040 5990 -1010
rect 6108 -1040 6162 -1010
rect 6280 -1040 6318 -1010
rect 5552 -1042 5568 -1040
rect 5502 -1052 5568 -1042
rect 5502 -1108 5568 -1098
rect 5502 -1110 5518 -1108
rect 4752 -1140 4790 -1110
rect 4908 -1140 4962 -1110
rect 5080 -1140 5190 -1110
rect 5308 -1140 5362 -1110
rect 5480 -1140 5518 -1110
rect 4752 -1142 4768 -1140
rect 4702 -1152 4768 -1142
rect 4702 -1208 4768 -1198
rect 4702 -1210 4718 -1208
rect 3952 -1240 3990 -1210
rect 4108 -1240 4162 -1210
rect 4280 -1240 4390 -1210
rect 4508 -1240 4562 -1210
rect 4680 -1240 4718 -1210
rect 3952 -1242 3968 -1240
rect 3902 -1252 3968 -1242
rect 3902 -1308 3968 -1298
rect 3902 -1310 3918 -1308
rect 3152 -1340 3190 -1310
rect 3308 -1340 3362 -1310
rect 3480 -1340 3590 -1310
rect 3708 -1340 3762 -1310
rect 3880 -1340 3918 -1310
rect 3152 -1342 3168 -1340
rect 3102 -1352 3168 -1342
rect 3102 -1408 3168 -1398
rect 3102 -1410 3118 -1408
rect 2352 -1440 2390 -1410
rect 2508 -1440 2562 -1410
rect 2680 -1440 2790 -1410
rect 2908 -1440 2962 -1410
rect 3080 -1440 3118 -1410
rect 2352 -1442 2368 -1440
rect 2302 -1452 2368 -1442
rect 2302 -1508 2368 -1498
rect 2302 -1510 2318 -1508
rect 1552 -1540 1590 -1510
rect 1708 -1540 1762 -1510
rect 1880 -1540 1990 -1510
rect 2108 -1540 2162 -1510
rect 2280 -1540 2318 -1510
rect 1552 -1542 1568 -1540
rect 1502 -1552 1568 -1542
rect 1502 -1608 1568 -1598
rect 1502 -1610 1518 -1608
rect 752 -1640 790 -1610
rect 908 -1640 962 -1610
rect 1080 -1640 1190 -1610
rect 1308 -1640 1362 -1610
rect 1480 -1640 1518 -1610
rect 752 -1642 768 -1640
rect 702 -1652 768 -1642
rect 702 -1708 768 -1698
rect 702 -1710 718 -1708
rect -48 -1740 -10 -1710
rect 108 -1740 162 -1710
rect 280 -1740 390 -1710
rect 508 -1740 562 -1710
rect 680 -1740 718 -1710
rect -48 -1742 -32 -1740
rect -98 -1752 -32 -1742
rect -98 -1808 -32 -1798
rect -98 -1810 -82 -1808
rect -106 -1840 -82 -1810
rect -98 -1842 -82 -1840
rect -48 -1810 -32 -1808
rect 702 -1742 718 -1740
rect 752 -1710 768 -1708
rect 1502 -1642 1518 -1640
rect 1552 -1610 1568 -1608
rect 2302 -1542 2318 -1540
rect 2352 -1510 2368 -1508
rect 3102 -1442 3118 -1440
rect 3152 -1410 3168 -1408
rect 3902 -1342 3918 -1340
rect 3952 -1310 3968 -1308
rect 4702 -1242 4718 -1240
rect 4752 -1210 4768 -1208
rect 5502 -1142 5518 -1140
rect 5552 -1110 5568 -1108
rect 6302 -1042 6318 -1040
rect 6352 -1010 6368 -1008
rect 6352 -1040 6376 -1010
rect 6352 -1042 6368 -1040
rect 6302 -1052 6368 -1042
rect 8114 -1090 8140 -1060
rect 8290 -1090 8416 -1060
rect 8716 -1090 8742 -1060
rect 8800 -1090 8826 -1060
rect 9126 -1090 9252 -1060
rect 9402 -1090 9428 -1060
rect 6302 -1108 6368 -1098
rect 6302 -1110 6318 -1108
rect 5552 -1140 5590 -1110
rect 5708 -1140 5762 -1110
rect 5880 -1140 5990 -1110
rect 6108 -1140 6162 -1110
rect 6280 -1140 6318 -1110
rect 5552 -1142 5568 -1140
rect 5502 -1152 5568 -1142
rect 5502 -1208 5568 -1198
rect 5502 -1210 5518 -1208
rect 4752 -1240 4790 -1210
rect 4908 -1240 4962 -1210
rect 5080 -1240 5190 -1210
rect 5308 -1240 5362 -1210
rect 5480 -1240 5518 -1210
rect 4752 -1242 4768 -1240
rect 4702 -1252 4768 -1242
rect 4702 -1308 4768 -1298
rect 4702 -1310 4718 -1308
rect 3952 -1340 3990 -1310
rect 4108 -1340 4162 -1310
rect 4280 -1340 4390 -1310
rect 4508 -1340 4562 -1310
rect 4680 -1340 4718 -1310
rect 3952 -1342 3968 -1340
rect 3902 -1352 3968 -1342
rect 3902 -1408 3968 -1398
rect 3902 -1410 3918 -1408
rect 3152 -1440 3190 -1410
rect 3308 -1440 3362 -1410
rect 3480 -1440 3590 -1410
rect 3708 -1440 3762 -1410
rect 3880 -1440 3918 -1410
rect 3152 -1442 3168 -1440
rect 3102 -1452 3168 -1442
rect 3102 -1508 3168 -1498
rect 3102 -1510 3118 -1508
rect 2352 -1540 2390 -1510
rect 2508 -1540 2562 -1510
rect 2680 -1540 2790 -1510
rect 2908 -1540 2962 -1510
rect 3080 -1540 3118 -1510
rect 2352 -1542 2368 -1540
rect 2302 -1552 2368 -1542
rect 2302 -1608 2368 -1598
rect 2302 -1610 2318 -1608
rect 1552 -1640 1590 -1610
rect 1708 -1640 1762 -1610
rect 1880 -1640 1990 -1610
rect 2108 -1640 2162 -1610
rect 2280 -1640 2318 -1610
rect 1552 -1642 1568 -1640
rect 1502 -1652 1568 -1642
rect 1502 -1708 1568 -1698
rect 1502 -1710 1518 -1708
rect 752 -1740 790 -1710
rect 908 -1740 962 -1710
rect 1080 -1740 1190 -1710
rect 1308 -1740 1362 -1710
rect 1480 -1740 1518 -1710
rect 752 -1742 768 -1740
rect 702 -1752 768 -1742
rect 702 -1808 768 -1798
rect 702 -1810 718 -1808
rect -48 -1840 -10 -1810
rect 108 -1840 162 -1810
rect 280 -1840 390 -1810
rect 508 -1840 562 -1810
rect 680 -1840 718 -1810
rect -48 -1842 -32 -1840
rect -98 -1852 -32 -1842
rect 702 -1842 718 -1840
rect 752 -1810 768 -1808
rect 1502 -1742 1518 -1740
rect 1552 -1710 1568 -1708
rect 2302 -1642 2318 -1640
rect 2352 -1610 2368 -1608
rect 3102 -1542 3118 -1540
rect 3152 -1510 3168 -1508
rect 3902 -1442 3918 -1440
rect 3952 -1410 3968 -1408
rect 4702 -1342 4718 -1340
rect 4752 -1310 4768 -1308
rect 5502 -1242 5518 -1240
rect 5552 -1210 5568 -1208
rect 6302 -1142 6318 -1140
rect 6352 -1110 6368 -1108
rect 6352 -1140 6376 -1110
rect 6352 -1142 6368 -1140
rect 6302 -1152 6368 -1142
rect 8306 -1109 8400 -1090
rect 8306 -1143 8334 -1109
rect 8368 -1143 8400 -1109
rect 8306 -1160 8400 -1143
rect 9142 -1109 9236 -1090
rect 9142 -1143 9174 -1109
rect 9208 -1143 9236 -1109
rect 9142 -1160 9236 -1143
rect 8114 -1190 8140 -1160
rect 8290 -1190 8416 -1160
rect 8716 -1190 8742 -1160
rect 8800 -1190 8826 -1160
rect 9126 -1190 9252 -1160
rect 9402 -1190 9428 -1160
rect 6302 -1208 6368 -1198
rect 6302 -1210 6318 -1208
rect 5552 -1240 5590 -1210
rect 5708 -1240 5762 -1210
rect 5880 -1240 5990 -1210
rect 6108 -1240 6162 -1210
rect 6280 -1240 6318 -1210
rect 5552 -1242 5568 -1240
rect 5502 -1252 5568 -1242
rect 5502 -1308 5568 -1298
rect 5502 -1310 5518 -1308
rect 4752 -1340 4790 -1310
rect 4908 -1340 4962 -1310
rect 5080 -1340 5190 -1310
rect 5308 -1340 5362 -1310
rect 5480 -1340 5518 -1310
rect 4752 -1342 4768 -1340
rect 4702 -1352 4768 -1342
rect 4702 -1408 4768 -1398
rect 4702 -1410 4718 -1408
rect 3952 -1440 3990 -1410
rect 4108 -1440 4162 -1410
rect 4280 -1440 4390 -1410
rect 4508 -1440 4562 -1410
rect 4680 -1440 4718 -1410
rect 3952 -1442 3968 -1440
rect 3902 -1452 3968 -1442
rect 3902 -1508 3968 -1498
rect 3902 -1510 3918 -1508
rect 3152 -1540 3190 -1510
rect 3308 -1540 3362 -1510
rect 3480 -1540 3590 -1510
rect 3708 -1540 3762 -1510
rect 3880 -1540 3918 -1510
rect 3152 -1542 3168 -1540
rect 3102 -1552 3168 -1542
rect 3102 -1608 3168 -1598
rect 3102 -1610 3118 -1608
rect 2352 -1640 2390 -1610
rect 2508 -1640 2562 -1610
rect 2680 -1640 2790 -1610
rect 2908 -1640 2962 -1610
rect 3080 -1640 3118 -1610
rect 2352 -1642 2368 -1640
rect 2302 -1652 2368 -1642
rect 2302 -1708 2368 -1698
rect 2302 -1710 2318 -1708
rect 1552 -1740 1590 -1710
rect 1708 -1740 1762 -1710
rect 1880 -1740 1990 -1710
rect 2108 -1740 2162 -1710
rect 2280 -1740 2318 -1710
rect 1552 -1742 1568 -1740
rect 1502 -1752 1568 -1742
rect 1502 -1808 1568 -1798
rect 1502 -1810 1518 -1808
rect 752 -1840 790 -1810
rect 908 -1840 962 -1810
rect 1080 -1840 1190 -1810
rect 1308 -1840 1362 -1810
rect 1480 -1840 1518 -1810
rect 752 -1842 768 -1840
rect 702 -1852 768 -1842
rect 1502 -1842 1518 -1840
rect 1552 -1810 1568 -1808
rect 2302 -1742 2318 -1740
rect 2352 -1710 2368 -1708
rect 3102 -1642 3118 -1640
rect 3152 -1610 3168 -1608
rect 3902 -1542 3918 -1540
rect 3952 -1510 3968 -1508
rect 4702 -1442 4718 -1440
rect 4752 -1410 4768 -1408
rect 5502 -1342 5518 -1340
rect 5552 -1310 5568 -1308
rect 6302 -1242 6318 -1240
rect 6352 -1210 6368 -1208
rect 6352 -1240 6376 -1210
rect 6352 -1242 6368 -1240
rect 6302 -1252 6368 -1242
rect 8114 -1290 8140 -1260
rect 8290 -1290 8416 -1260
rect 8716 -1290 8742 -1260
rect 8800 -1290 8826 -1260
rect 9126 -1290 9252 -1260
rect 9402 -1290 9428 -1260
rect 6302 -1308 6368 -1298
rect 6302 -1310 6318 -1308
rect 5552 -1340 5590 -1310
rect 5708 -1340 5762 -1310
rect 5880 -1340 5990 -1310
rect 6108 -1340 6162 -1310
rect 6280 -1340 6318 -1310
rect 5552 -1342 5568 -1340
rect 5502 -1352 5568 -1342
rect 5502 -1408 5568 -1398
rect 5502 -1410 5518 -1408
rect 4752 -1440 4790 -1410
rect 4908 -1440 4962 -1410
rect 5080 -1440 5190 -1410
rect 5308 -1440 5362 -1410
rect 5480 -1440 5518 -1410
rect 4752 -1442 4768 -1440
rect 4702 -1452 4768 -1442
rect 4702 -1508 4768 -1498
rect 4702 -1510 4718 -1508
rect 3952 -1540 3990 -1510
rect 4108 -1540 4162 -1510
rect 4280 -1540 4390 -1510
rect 4508 -1540 4562 -1510
rect 4680 -1540 4718 -1510
rect 3952 -1542 3968 -1540
rect 3902 -1552 3968 -1542
rect 3902 -1608 3968 -1598
rect 3902 -1610 3918 -1608
rect 3152 -1640 3190 -1610
rect 3308 -1640 3362 -1610
rect 3480 -1640 3590 -1610
rect 3708 -1640 3762 -1610
rect 3880 -1640 3918 -1610
rect 3152 -1642 3168 -1640
rect 3102 -1652 3168 -1642
rect 3102 -1708 3168 -1698
rect 3102 -1710 3118 -1708
rect 2352 -1740 2390 -1710
rect 2508 -1740 2562 -1710
rect 2680 -1740 2790 -1710
rect 2908 -1740 2962 -1710
rect 3080 -1740 3118 -1710
rect 2352 -1742 2368 -1740
rect 2302 -1752 2368 -1742
rect 2302 -1808 2368 -1798
rect 2302 -1810 2318 -1808
rect 1552 -1840 1590 -1810
rect 1708 -1840 1762 -1810
rect 1880 -1840 1990 -1810
rect 2108 -1840 2162 -1810
rect 2280 -1840 2318 -1810
rect 1552 -1842 1568 -1840
rect 1502 -1852 1568 -1842
rect 2302 -1842 2318 -1840
rect 2352 -1810 2368 -1808
rect 3102 -1742 3118 -1740
rect 3152 -1710 3168 -1708
rect 3902 -1642 3918 -1640
rect 3952 -1610 3968 -1608
rect 4702 -1542 4718 -1540
rect 4752 -1510 4768 -1508
rect 5502 -1442 5518 -1440
rect 5552 -1410 5568 -1408
rect 6302 -1342 6318 -1340
rect 6352 -1310 6368 -1308
rect 6352 -1340 6376 -1310
rect 6352 -1342 6368 -1340
rect 6302 -1352 6368 -1342
rect 8306 -1309 8400 -1290
rect 8306 -1343 8334 -1309
rect 8368 -1343 8400 -1309
rect 8306 -1360 8400 -1343
rect 9142 -1309 9236 -1290
rect 9142 -1343 9174 -1309
rect 9208 -1343 9236 -1309
rect 9142 -1360 9236 -1343
rect 8114 -1390 8140 -1360
rect 8290 -1390 8416 -1360
rect 8716 -1390 8742 -1360
rect 8800 -1390 8826 -1360
rect 9126 -1390 9252 -1360
rect 9402 -1390 9428 -1360
rect 6302 -1408 6368 -1398
rect 6302 -1410 6318 -1408
rect 5552 -1440 5590 -1410
rect 5708 -1440 5762 -1410
rect 5880 -1440 5990 -1410
rect 6108 -1440 6162 -1410
rect 6280 -1440 6318 -1410
rect 5552 -1442 5568 -1440
rect 5502 -1452 5568 -1442
rect 5502 -1508 5568 -1498
rect 5502 -1510 5518 -1508
rect 4752 -1540 4790 -1510
rect 4908 -1540 4962 -1510
rect 5080 -1540 5190 -1510
rect 5308 -1540 5362 -1510
rect 5480 -1540 5518 -1510
rect 4752 -1542 4768 -1540
rect 4702 -1552 4768 -1542
rect 4702 -1608 4768 -1598
rect 4702 -1610 4718 -1608
rect 3952 -1640 3990 -1610
rect 4108 -1640 4162 -1610
rect 4280 -1640 4390 -1610
rect 4508 -1640 4562 -1610
rect 4680 -1640 4718 -1610
rect 3952 -1642 3968 -1640
rect 3902 -1652 3968 -1642
rect 3902 -1708 3968 -1698
rect 3902 -1710 3918 -1708
rect 3152 -1740 3190 -1710
rect 3308 -1740 3362 -1710
rect 3480 -1740 3590 -1710
rect 3708 -1740 3762 -1710
rect 3880 -1740 3918 -1710
rect 3152 -1742 3168 -1740
rect 3102 -1752 3168 -1742
rect 3102 -1808 3168 -1798
rect 3102 -1810 3118 -1808
rect 2352 -1840 2390 -1810
rect 2508 -1840 2562 -1810
rect 2680 -1840 2790 -1810
rect 2908 -1840 2962 -1810
rect 3080 -1840 3118 -1810
rect 2352 -1842 2368 -1840
rect 2302 -1852 2368 -1842
rect 3102 -1842 3118 -1840
rect 3152 -1810 3168 -1808
rect 3902 -1742 3918 -1740
rect 3952 -1710 3968 -1708
rect 4702 -1642 4718 -1640
rect 4752 -1610 4768 -1608
rect 5502 -1542 5518 -1540
rect 5552 -1510 5568 -1508
rect 6302 -1442 6318 -1440
rect 6352 -1410 6368 -1408
rect 6352 -1440 6376 -1410
rect 6352 -1442 6368 -1440
rect 6302 -1452 6368 -1442
rect 8114 -1490 8140 -1460
rect 8290 -1490 8416 -1460
rect 8716 -1490 8742 -1460
rect 8800 -1490 8826 -1460
rect 9126 -1490 9252 -1460
rect 9402 -1490 9428 -1460
rect 6302 -1508 6368 -1498
rect 6302 -1510 6318 -1508
rect 5552 -1540 5590 -1510
rect 5708 -1540 5762 -1510
rect 5880 -1540 5990 -1510
rect 6108 -1540 6162 -1510
rect 6280 -1540 6318 -1510
rect 5552 -1542 5568 -1540
rect 5502 -1552 5568 -1542
rect 5502 -1608 5568 -1598
rect 5502 -1610 5518 -1608
rect 4752 -1640 4790 -1610
rect 4908 -1640 4962 -1610
rect 5080 -1640 5190 -1610
rect 5308 -1640 5362 -1610
rect 5480 -1640 5518 -1610
rect 4752 -1642 4768 -1640
rect 4702 -1652 4768 -1642
rect 4702 -1708 4768 -1698
rect 4702 -1710 4718 -1708
rect 3952 -1740 3990 -1710
rect 4108 -1740 4162 -1710
rect 4280 -1740 4390 -1710
rect 4508 -1740 4562 -1710
rect 4680 -1740 4718 -1710
rect 3952 -1742 3968 -1740
rect 3902 -1752 3968 -1742
rect 3902 -1808 3968 -1798
rect 3902 -1810 3918 -1808
rect 3152 -1840 3190 -1810
rect 3308 -1840 3362 -1810
rect 3480 -1840 3590 -1810
rect 3708 -1840 3762 -1810
rect 3880 -1840 3918 -1810
rect 3152 -1842 3168 -1840
rect 3102 -1852 3168 -1842
rect 3902 -1842 3918 -1840
rect 3952 -1810 3968 -1808
rect 4702 -1742 4718 -1740
rect 4752 -1710 4768 -1708
rect 5502 -1642 5518 -1640
rect 5552 -1610 5568 -1608
rect 6302 -1542 6318 -1540
rect 6352 -1510 6368 -1508
rect 6352 -1540 6376 -1510
rect 6352 -1542 6368 -1540
rect 6302 -1552 6368 -1542
rect 8306 -1509 8400 -1490
rect 8306 -1543 8334 -1509
rect 8368 -1543 8400 -1509
rect 8306 -1560 8400 -1543
rect 9142 -1509 9236 -1490
rect 9142 -1543 9174 -1509
rect 9208 -1543 9236 -1509
rect 9142 -1560 9236 -1543
rect 8114 -1590 8140 -1560
rect 8290 -1590 8416 -1560
rect 8716 -1590 8742 -1560
rect 8800 -1590 8826 -1560
rect 9126 -1590 9252 -1560
rect 9402 -1590 9428 -1560
rect 6302 -1608 6368 -1598
rect 6302 -1610 6318 -1608
rect 5552 -1640 5590 -1610
rect 5708 -1640 5762 -1610
rect 5880 -1640 5990 -1610
rect 6108 -1640 6162 -1610
rect 6280 -1640 6318 -1610
rect 5552 -1642 5568 -1640
rect 5502 -1652 5568 -1642
rect 5502 -1708 5568 -1698
rect 5502 -1710 5518 -1708
rect 4752 -1740 4790 -1710
rect 4908 -1740 4962 -1710
rect 5080 -1740 5190 -1710
rect 5308 -1740 5362 -1710
rect 5480 -1740 5518 -1710
rect 4752 -1742 4768 -1740
rect 4702 -1752 4768 -1742
rect 4702 -1808 4768 -1798
rect 4702 -1810 4718 -1808
rect 3952 -1840 3990 -1810
rect 4108 -1840 4162 -1810
rect 4280 -1840 4390 -1810
rect 4508 -1840 4562 -1810
rect 4680 -1840 4718 -1810
rect 3952 -1842 3968 -1840
rect 3902 -1852 3968 -1842
rect 4702 -1842 4718 -1840
rect 4752 -1810 4768 -1808
rect 5502 -1742 5518 -1740
rect 5552 -1710 5568 -1708
rect 6302 -1642 6318 -1640
rect 6352 -1610 6368 -1608
rect 6352 -1640 6376 -1610
rect 6352 -1642 6368 -1640
rect 6302 -1652 6368 -1642
rect 8114 -1690 8140 -1660
rect 8290 -1690 8416 -1660
rect 8716 -1690 8742 -1660
rect 8800 -1690 8826 -1660
rect 9126 -1690 9252 -1660
rect 9402 -1690 9428 -1660
rect 6302 -1708 6368 -1698
rect 6302 -1710 6318 -1708
rect 5552 -1740 5590 -1710
rect 5708 -1740 5762 -1710
rect 5880 -1740 5990 -1710
rect 6108 -1740 6162 -1710
rect 6280 -1740 6318 -1710
rect 5552 -1742 5568 -1740
rect 5502 -1752 5568 -1742
rect 5502 -1808 5568 -1798
rect 5502 -1810 5518 -1808
rect 4752 -1840 4790 -1810
rect 4908 -1840 4962 -1810
rect 5080 -1840 5190 -1810
rect 5308 -1840 5362 -1810
rect 5480 -1840 5518 -1810
rect 4752 -1842 4768 -1840
rect 4702 -1852 4768 -1842
rect 5502 -1842 5518 -1840
rect 5552 -1810 5568 -1808
rect 6302 -1742 6318 -1740
rect 6352 -1710 6368 -1708
rect 6352 -1740 6376 -1710
rect 6352 -1742 6368 -1740
rect 6302 -1752 6368 -1742
rect 8306 -1709 8400 -1690
rect 8306 -1743 8334 -1709
rect 8368 -1743 8400 -1709
rect 8306 -1760 8400 -1743
rect 9142 -1709 9236 -1690
rect 9142 -1743 9174 -1709
rect 9208 -1743 9236 -1709
rect 9142 -1760 9236 -1743
rect 8114 -1790 8140 -1760
rect 8290 -1790 8416 -1760
rect 8716 -1790 8742 -1760
rect 8800 -1790 8826 -1760
rect 9126 -1790 9252 -1760
rect 9402 -1790 9428 -1760
rect 6302 -1808 6368 -1798
rect 6302 -1810 6318 -1808
rect 5552 -1840 5590 -1810
rect 5708 -1840 5762 -1810
rect 5880 -1840 5990 -1810
rect 6108 -1840 6162 -1810
rect 6280 -1840 6318 -1810
rect 5552 -1842 5568 -1840
rect 5502 -1852 5568 -1842
rect 6302 -1842 6318 -1840
rect 6352 -1810 6368 -1808
rect 6352 -1840 6376 -1810
rect 6352 -1842 6368 -1840
rect 6302 -1852 6368 -1842
<< polycont >>
rect 118 9840 152 9874
rect 318 9856 352 9890
rect 518 9840 552 9874
rect 718 9856 752 9890
rect 918 9840 952 9874
rect 1118 9856 1152 9890
rect 1318 9840 1352 9874
rect 1518 9856 1552 9890
rect 1718 9840 1752 9874
rect 1918 9856 1952 9890
rect 2118 9840 2152 9874
rect 2318 9856 2352 9890
rect 2518 9840 2552 9874
rect 2718 9856 2752 9890
rect 2918 9840 2952 9874
rect 3118 9856 3152 9890
rect 3318 9840 3352 9874
rect 3518 9856 3552 9890
rect 3718 9840 3752 9874
rect 3918 9856 3952 9890
rect 4118 9840 4152 9874
rect 4318 9856 4352 9890
rect 4518 9840 4552 9874
rect 4718 9856 4752 9890
rect 4918 9840 4952 9874
rect 5118 9856 5152 9890
rect 5318 9840 5352 9874
rect 5518 9856 5552 9890
rect 5718 9840 5752 9874
rect 5918 9856 5952 9890
rect 118 8630 152 8664
rect 318 8646 352 8680
rect 518 8630 552 8664
rect 718 8646 752 8680
rect 918 8630 952 8664
rect 1118 8646 1152 8680
rect 1318 8630 1352 8664
rect 1518 8646 1552 8680
rect 1718 8630 1752 8664
rect 1918 8646 1952 8680
rect 2118 8630 2152 8664
rect 2318 8646 2352 8680
rect 2518 8630 2552 8664
rect 6118 9840 6152 9874
rect 6318 9856 6352 9890
rect 6568 9854 6602 9888
rect 6668 9854 6702 9888
rect 6878 9854 6912 9888
rect 6978 9854 7012 9888
rect 7078 9854 7112 9888
rect 7178 9854 7212 9888
rect 7278 9854 7312 9888
rect 7378 9854 7412 9888
rect 2718 8646 2752 8680
rect 2918 8630 2952 8664
rect 3118 8646 3152 8680
rect 3318 8630 3352 8664
rect 3518 8646 3552 8680
rect 3718 8630 3752 8664
rect 3918 8646 3952 8680
rect 4118 8630 4152 8664
rect 118 7420 152 7454
rect 318 7436 352 7470
rect 518 7420 552 7454
rect 718 7436 752 7470
rect 918 7420 952 7454
rect 1118 7436 1152 7470
rect 4318 8646 4352 8680
rect 4518 8630 4552 8664
rect 4718 8646 4752 8680
rect 4918 8630 4952 8664
rect 5118 8646 5152 8680
rect 5318 8630 5352 8664
rect 5518 8646 5552 8680
rect 5718 8630 5752 8664
rect 5918 8646 5952 8680
rect 6118 8630 6152 8664
rect 6318 8646 6352 8680
rect 6568 8644 6602 8678
rect 6668 8644 6702 8678
rect 6878 8644 6912 8678
rect 6978 8644 7012 8678
rect 7078 8644 7112 8678
rect 7178 8644 7212 8678
rect 7278 8644 7312 8678
rect 7378 8644 7412 8678
rect 1318 7420 1352 7454
rect 1518 7436 1552 7470
rect 1718 7420 1752 7454
rect 1918 7436 1952 7470
rect 2118 7420 2152 7454
rect 2318 7436 2352 7470
rect 2518 7420 2552 7454
rect 2718 7436 2752 7470
rect 2918 7420 2952 7454
rect 3118 7436 3152 7470
rect 3318 7420 3352 7454
rect 3518 7436 3552 7470
rect 3718 7420 3752 7454
rect 3918 7436 3952 7470
rect 4118 7420 4152 7454
rect 4318 7436 4352 7470
rect 4518 7420 4552 7454
rect 4718 7436 4752 7470
rect 4918 7420 4952 7454
rect 5118 7436 5152 7470
rect 5318 7420 5352 7454
rect 5518 7436 5552 7470
rect 5718 7420 5752 7454
rect 5918 7436 5952 7470
rect 6118 7420 6152 7454
rect 6318 7436 6352 7470
rect 6568 7434 6602 7468
rect 6668 7434 6702 7468
rect 6878 7434 6912 7468
rect 6978 7434 7012 7468
rect 7078 7434 7112 7468
rect 7178 7434 7212 7468
rect 7278 7434 7312 7468
rect 7378 7434 7412 7468
rect 118 6210 152 6244
rect 318 6226 352 6260
rect 518 6210 552 6244
rect 718 6226 752 6260
rect 918 6210 952 6244
rect 1118 6226 1152 6260
rect 1318 6210 1352 6244
rect 1518 6226 1552 6260
rect 1718 6210 1752 6244
rect 1918 6226 1952 6260
rect 2118 6210 2152 6244
rect 2318 6226 2352 6260
rect 2518 6210 2552 6244
rect 2718 6226 2752 6260
rect 2918 6210 2952 6244
rect 3118 6226 3152 6260
rect 3318 6210 3352 6244
rect 3518 6226 3552 6260
rect 3718 6210 3752 6244
rect 3918 6226 3952 6260
rect 4118 6210 4152 6244
rect 4318 6226 4352 6260
rect 4518 6210 4552 6244
rect 4718 6226 4752 6260
rect 4918 6210 4952 6244
rect 5118 6226 5152 6260
rect 5318 6210 5352 6244
rect 5518 6226 5552 6260
rect 5718 6210 5752 6244
rect 5918 6226 5952 6260
rect 6118 6210 6152 6244
rect 118 4860 152 4894
rect 318 4876 352 4910
rect 518 4860 552 4894
rect 718 4876 752 4910
rect 918 4860 952 4894
rect 1118 4876 1152 4910
rect 1318 4860 1352 4894
rect 1518 4876 1552 4910
rect 1718 4860 1752 4894
rect 1918 4876 1952 4910
rect 6318 6226 6352 6260
rect 6568 6224 6602 6258
rect 6668 6224 6702 6258
rect 6878 6224 6912 6258
rect 6978 6224 7012 6258
rect 7078 6224 7112 6258
rect 7178 6224 7212 6258
rect 7278 6224 7312 6258
rect 7378 6224 7412 6258
rect 2118 4860 2152 4894
rect 2318 4876 2352 4910
rect 2518 4860 2552 4894
rect 2718 4876 2752 4910
rect 2918 4860 2952 4894
rect 3118 4876 3152 4910
rect 3318 4860 3352 4894
rect 3518 4876 3552 4910
rect 3718 4860 3752 4894
rect 3918 4876 3952 4910
rect 4118 4860 4152 4894
rect 4318 4876 4352 4910
rect 4518 4860 4552 4894
rect 4718 4876 4752 4910
rect 4918 4860 4952 4894
rect 5118 4876 5152 4910
rect 5318 4860 5352 4894
rect 5518 4876 5552 4910
rect 5718 4860 5752 4894
rect 5918 4876 5952 4910
rect 6118 4860 6152 4894
rect 118 3650 152 3684
rect 318 3666 352 3700
rect 518 3650 552 3684
rect 718 3666 752 3700
rect 918 3650 952 3684
rect 1118 3666 1152 3700
rect 1318 3650 1352 3684
rect 1518 3666 1552 3700
rect 1718 3650 1752 3684
rect 1918 3666 1952 3700
rect 2118 3650 2152 3684
rect 2318 3666 2352 3700
rect 2518 3650 2552 3684
rect 2718 3666 2752 3700
rect 2918 3650 2952 3684
rect 3118 3666 3152 3700
rect 3318 3650 3352 3684
rect 6318 4876 6352 4910
rect 6568 4874 6602 4908
rect 6668 4874 6702 4908
rect 6878 4874 6912 4908
rect 6978 4874 7012 4908
rect 7078 4874 7112 4908
rect 7178 4874 7212 4908
rect 7278 4874 7312 4908
rect 7378 4874 7412 4908
rect 3518 3666 3552 3700
rect 3718 3650 3752 3684
rect 3918 3666 3952 3700
rect 4118 3650 4152 3684
rect 4318 3666 4352 3700
rect 4518 3650 4552 3684
rect 4718 3666 4752 3700
rect 4918 3650 4952 3684
rect 5118 3666 5152 3700
rect 5318 3650 5352 3684
rect 5518 3666 5552 3700
rect 5718 3650 5752 3684
rect 5918 3666 5952 3700
rect 6118 3650 6152 3684
rect 6318 3666 6352 3700
rect 6568 3664 6602 3698
rect 6668 3664 6702 3698
rect 6878 3664 6912 3698
rect 6978 3664 7012 3698
rect 7078 3664 7112 3698
rect 7178 3664 7212 3698
rect 7278 3664 7312 3698
rect 7378 3664 7412 3698
rect 118 2440 152 2474
rect 318 2456 352 2490
rect 518 2440 552 2474
rect 718 2456 752 2490
rect 918 2440 952 2474
rect 1118 2456 1152 2490
rect 1318 2440 1352 2474
rect 1518 2456 1552 2490
rect 1718 2440 1752 2474
rect 1918 2456 1952 2490
rect 2118 2440 2152 2474
rect 2318 2456 2352 2490
rect 2518 2440 2552 2474
rect 2718 2456 2752 2490
rect 2918 2440 2952 2474
rect 3118 2456 3152 2490
rect 3318 2440 3352 2474
rect 3518 2456 3552 2490
rect 3718 2440 3752 2474
rect 3918 2456 3952 2490
rect 4118 2440 4152 2474
rect 4318 2456 4352 2490
rect 4518 2440 4552 2474
rect 4718 2456 4752 2490
rect 4918 2440 4952 2474
rect 5118 2456 5152 2490
rect 5318 2440 5352 2474
rect 5518 2456 5552 2490
rect 118 1230 152 1264
rect 318 1246 352 1280
rect 518 1230 552 1264
rect 718 1246 752 1280
rect 918 1230 952 1264
rect 1118 1246 1152 1280
rect 1318 1230 1352 1264
rect 5718 2440 5752 2474
rect 5918 2456 5952 2490
rect 6118 2440 6152 2474
rect 6318 2456 6352 2490
rect 6568 2454 6602 2488
rect 6668 2454 6702 2488
rect 6878 2454 6912 2488
rect 6978 2454 7012 2488
rect 7078 2454 7112 2488
rect 7178 2454 7212 2488
rect 7278 2454 7312 2488
rect 7378 2454 7412 2488
rect 1518 1246 1552 1280
rect 1718 1230 1752 1264
rect 1918 1246 1952 1280
rect 2118 1230 2152 1264
rect 2318 1246 2352 1280
rect 2518 1230 2552 1264
rect 2718 1246 2752 1280
rect 2918 1230 2952 1264
rect 3118 1246 3152 1280
rect 3318 1230 3352 1264
rect 3518 1246 3552 1280
rect 3718 1230 3752 1264
rect 3918 1246 3952 1280
rect 4118 1230 4152 1264
rect 4318 1246 4352 1280
rect 4518 1230 4552 1264
rect 4718 1246 4752 1280
rect 4918 1230 4952 1264
rect 5118 1246 5152 1280
rect 5318 1230 5352 1264
rect 5518 1246 5552 1280
rect 118 20 152 54
rect 318 36 352 70
rect 518 20 552 54
rect 718 36 752 70
rect 918 20 952 54
rect 1118 36 1152 70
rect 1318 20 1352 54
rect 1518 36 1552 70
rect 1718 20 1752 54
rect 1918 36 1952 70
rect 2118 20 2152 54
rect 2318 36 2352 70
rect 2518 20 2552 54
rect 2718 36 2752 70
rect 2918 20 2952 54
rect 3118 36 3152 70
rect 3318 20 3352 54
rect 5718 1230 5752 1264
rect 5918 1246 5952 1280
rect 6118 1230 6152 1264
rect 6318 1246 6352 1280
rect 6568 1244 6602 1278
rect 6668 1244 6702 1278
rect 6878 1244 6912 1278
rect 6978 1244 7012 1278
rect 7078 1244 7112 1278
rect 7178 1244 7212 1278
rect 7278 1244 7312 1278
rect 7378 1244 7412 1278
rect 3518 36 3552 70
rect 3718 20 3752 54
rect 3918 36 3952 70
rect 4118 20 4152 54
rect 4318 36 4352 70
rect 4518 20 4552 54
rect 4718 36 4752 70
rect 4918 20 4952 54
rect 5118 36 5152 70
rect 5318 20 5352 54
rect 5518 36 5552 70
rect 5718 20 5752 54
rect 5918 36 5952 70
rect 6118 20 6152 54
rect 6318 36 6352 70
rect 6568 34 6602 68
rect 6668 34 6702 68
rect 6878 34 6912 68
rect 6978 34 7012 68
rect 7078 34 7112 68
rect 7178 34 7212 68
rect 7278 34 7312 68
rect 7378 34 7412 68
rect 8334 -143 8368 -109
rect 9174 -143 9208 -109
rect 18 -282 52 -248
rect 218 -282 252 -248
rect 418 -282 452 -248
rect 618 -282 652 -248
rect 818 -282 852 -248
rect 1018 -282 1052 -248
rect 1218 -282 1252 -248
rect 1418 -282 1452 -248
rect 1618 -282 1652 -248
rect 1818 -282 1852 -248
rect 2018 -282 2052 -248
rect 2218 -282 2252 -248
rect 2418 -282 2452 -248
rect 2618 -282 2652 -248
rect 2818 -282 2852 -248
rect 3018 -282 3052 -248
rect 3218 -282 3252 -248
rect 3418 -282 3452 -248
rect 3618 -282 3652 -248
rect 3818 -282 3852 -248
rect 4018 -282 4052 -248
rect 4218 -282 4252 -248
rect 4418 -282 4452 -248
rect 4618 -282 4652 -248
rect 4818 -282 4852 -248
rect 5018 -282 5052 -248
rect 5218 -282 5252 -248
rect 5418 -282 5452 -248
rect 5618 -282 5652 -248
rect 5818 -282 5852 -248
rect 6018 -282 6052 -248
rect 6218 -282 6252 -248
rect 8334 -343 8368 -309
rect 9174 -343 9208 -309
rect 8334 -543 8368 -509
rect 9174 -543 9208 -509
rect 44 -611 78 -577
rect 192 -611 226 -577
rect 444 -611 478 -577
rect 592 -611 626 -577
rect 844 -611 878 -577
rect 992 -611 1026 -577
rect 1244 -611 1278 -577
rect 1392 -611 1426 -577
rect 1644 -611 1678 -577
rect 1792 -611 1826 -577
rect 2044 -611 2078 -577
rect 2192 -611 2226 -577
rect 2444 -611 2478 -577
rect 2592 -611 2626 -577
rect 2844 -611 2878 -577
rect 2992 -611 3026 -577
rect 3244 -611 3278 -577
rect 3392 -611 3426 -577
rect 3644 -611 3678 -577
rect 3792 -611 3826 -577
rect 4044 -611 4078 -577
rect 4192 -611 4226 -577
rect 4444 -611 4478 -577
rect 4592 -611 4626 -577
rect 4844 -611 4878 -577
rect 4992 -611 5026 -577
rect 5244 -611 5278 -577
rect 5392 -611 5426 -577
rect 5644 -611 5678 -577
rect 5792 -611 5826 -577
rect 6044 -611 6078 -577
rect 6192 -611 6226 -577
rect 8334 -743 8368 -709
rect 9174 -743 9208 -709
rect -82 -942 -48 -908
rect -82 -1042 -48 -1008
rect 718 -942 752 -908
rect -82 -1142 -48 -1108
rect 718 -1042 752 -1008
rect 1518 -942 1552 -908
rect -82 -1242 -48 -1208
rect 718 -1142 752 -1108
rect 1518 -1042 1552 -1008
rect 2318 -942 2352 -908
rect -82 -1342 -48 -1308
rect 718 -1242 752 -1208
rect 1518 -1142 1552 -1108
rect 2318 -1042 2352 -1008
rect 3118 -942 3152 -908
rect -82 -1442 -48 -1408
rect 718 -1342 752 -1308
rect 1518 -1242 1552 -1208
rect 2318 -1142 2352 -1108
rect 3118 -1042 3152 -1008
rect 3918 -942 3952 -908
rect -82 -1542 -48 -1508
rect 718 -1442 752 -1408
rect 1518 -1342 1552 -1308
rect 2318 -1242 2352 -1208
rect 3118 -1142 3152 -1108
rect 3918 -1042 3952 -1008
rect 4718 -942 4752 -908
rect -82 -1642 -48 -1608
rect 718 -1542 752 -1508
rect 1518 -1442 1552 -1408
rect 2318 -1342 2352 -1308
rect 3118 -1242 3152 -1208
rect 3918 -1142 3952 -1108
rect 4718 -1042 4752 -1008
rect 5518 -942 5552 -908
rect -82 -1742 -48 -1708
rect 718 -1642 752 -1608
rect 1518 -1542 1552 -1508
rect 2318 -1442 2352 -1408
rect 3118 -1342 3152 -1308
rect 3918 -1242 3952 -1208
rect 4718 -1142 4752 -1108
rect 5518 -1042 5552 -1008
rect 6318 -942 6352 -908
rect 8334 -943 8368 -909
rect 9174 -943 9208 -909
rect -82 -1842 -48 -1808
rect 718 -1742 752 -1708
rect 1518 -1642 1552 -1608
rect 2318 -1542 2352 -1508
rect 3118 -1442 3152 -1408
rect 3918 -1342 3952 -1308
rect 4718 -1242 4752 -1208
rect 5518 -1142 5552 -1108
rect 6318 -1042 6352 -1008
rect 718 -1842 752 -1808
rect 1518 -1742 1552 -1708
rect 2318 -1642 2352 -1608
rect 3118 -1542 3152 -1508
rect 3918 -1442 3952 -1408
rect 4718 -1342 4752 -1308
rect 5518 -1242 5552 -1208
rect 6318 -1142 6352 -1108
rect 8334 -1143 8368 -1109
rect 9174 -1143 9208 -1109
rect 1518 -1842 1552 -1808
rect 2318 -1742 2352 -1708
rect 3118 -1642 3152 -1608
rect 3918 -1542 3952 -1508
rect 4718 -1442 4752 -1408
rect 5518 -1342 5552 -1308
rect 6318 -1242 6352 -1208
rect 2318 -1842 2352 -1808
rect 3118 -1742 3152 -1708
rect 3918 -1642 3952 -1608
rect 4718 -1542 4752 -1508
rect 5518 -1442 5552 -1408
rect 6318 -1342 6352 -1308
rect 8334 -1343 8368 -1309
rect 9174 -1343 9208 -1309
rect 3118 -1842 3152 -1808
rect 3918 -1742 3952 -1708
rect 4718 -1642 4752 -1608
rect 5518 -1542 5552 -1508
rect 6318 -1442 6352 -1408
rect 3918 -1842 3952 -1808
rect 4718 -1742 4752 -1708
rect 5518 -1642 5552 -1608
rect 6318 -1542 6352 -1508
rect 8334 -1543 8368 -1509
rect 9174 -1543 9208 -1509
rect 4718 -1842 4752 -1808
rect 5518 -1742 5552 -1708
rect 6318 -1642 6352 -1608
rect 5518 -1842 5552 -1808
rect 6318 -1742 6352 -1708
rect 8334 -1743 8368 -1709
rect 9174 -1743 9208 -1709
rect 6318 -1842 6352 -1808
<< locali >>
rect 106 9997 164 10023
rect 106 9963 118 9997
rect 152 9963 164 9997
rect 106 9937 164 9963
rect 306 9997 364 10023
rect 306 9963 318 9997
rect 352 9963 364 9997
rect 306 9937 364 9963
rect 506 9997 564 10023
rect 506 9963 518 9997
rect 552 9963 564 9997
rect 506 9937 564 9963
rect 706 9997 764 10023
rect 706 9963 718 9997
rect 752 9963 764 9997
rect 706 9937 764 9963
rect 906 9997 964 10023
rect 906 9963 918 9997
rect 952 9963 964 9997
rect 906 9937 964 9963
rect 1106 9997 1164 10023
rect 1106 9963 1118 9997
rect 1152 9963 1164 9997
rect 1106 9937 1164 9963
rect 1306 9997 1364 10023
rect 1306 9963 1318 9997
rect 1352 9963 1364 9997
rect 1306 9937 1364 9963
rect 1506 9997 1564 10023
rect 1506 9963 1518 9997
rect 1552 9963 1564 9997
rect 1506 9937 1564 9963
rect 1706 9997 1764 10023
rect 1706 9963 1718 9997
rect 1752 9963 1764 9997
rect 1706 9937 1764 9963
rect 1906 9997 1964 10023
rect 1906 9963 1918 9997
rect 1952 9963 1964 9997
rect 1906 9937 1964 9963
rect 2106 9997 2164 10023
rect 2106 9963 2118 9997
rect 2152 9963 2164 9997
rect 2106 9937 2164 9963
rect 2306 9997 2364 10023
rect 2306 9963 2318 9997
rect 2352 9963 2364 9997
rect 2306 9937 2364 9963
rect 2506 9997 2564 10023
rect 2506 9963 2518 9997
rect 2552 9963 2564 9997
rect 2506 9937 2564 9963
rect 2706 9997 2764 10023
rect 2706 9963 2718 9997
rect 2752 9963 2764 9997
rect 2706 9937 2764 9963
rect 2906 9997 2964 10023
rect 2906 9963 2918 9997
rect 2952 9963 2964 9997
rect 2906 9937 2964 9963
rect 3106 9997 3164 10023
rect 3106 9963 3118 9997
rect 3152 9963 3164 9997
rect 3106 9937 3164 9963
rect 3306 9997 3364 10023
rect 3306 9963 3318 9997
rect 3352 9963 3364 9997
rect 3306 9937 3364 9963
rect 3506 9997 3564 10023
rect 3506 9963 3518 9997
rect 3552 9963 3564 9997
rect 3506 9937 3564 9963
rect 3706 9997 3764 10023
rect 3706 9963 3718 9997
rect 3752 9963 3764 9997
rect 3706 9937 3764 9963
rect 3906 9997 3964 10023
rect 3906 9963 3918 9997
rect 3952 9963 3964 9997
rect 3906 9937 3964 9963
rect 4106 9997 4164 10023
rect 4106 9963 4118 9997
rect 4152 9963 4164 9997
rect 4106 9937 4164 9963
rect 4306 9997 4364 10023
rect 4306 9963 4318 9997
rect 4352 9963 4364 9997
rect 4306 9937 4364 9963
rect 4506 9997 4564 10023
rect 4506 9963 4518 9997
rect 4552 9963 4564 9997
rect 4506 9937 4564 9963
rect 4706 9997 4764 10023
rect 4706 9963 4718 9997
rect 4752 9963 4764 9997
rect 4706 9937 4764 9963
rect 4906 9997 4964 10023
rect 4906 9963 4918 9997
rect 4952 9963 4964 9997
rect 4906 9937 4964 9963
rect 5106 9997 5164 10023
rect 5106 9963 5118 9997
rect 5152 9963 5164 9997
rect 5106 9937 5164 9963
rect 5306 9997 5364 10023
rect 5306 9963 5318 9997
rect 5352 9963 5364 9997
rect 5306 9937 5364 9963
rect 5506 9997 5564 10023
rect 5506 9963 5518 9997
rect 5552 9963 5564 9997
rect 5506 9937 5564 9963
rect 5706 9997 5764 10023
rect 5706 9963 5718 9997
rect 5752 9963 5764 9997
rect 5706 9937 5764 9963
rect 5906 9997 5964 10023
rect 5906 9963 5918 9997
rect 5952 9963 5964 9997
rect 5906 9937 5964 9963
rect 6106 9997 6164 10023
rect 6106 9963 6118 9997
rect 6152 9963 6164 9997
rect 6106 9937 6164 9963
rect 6306 9997 6364 10023
rect 6306 9963 6318 9997
rect 6352 9963 6364 9997
rect 6306 9937 6364 9963
rect 8 9840 18 9874
rect 52 9840 118 9874
rect 152 9840 168 9874
rect 208 9856 218 9890
rect 252 9856 318 9890
rect 352 9856 368 9890
rect 408 9840 418 9874
rect 452 9840 518 9874
rect 552 9840 568 9874
rect 608 9856 618 9890
rect 652 9856 718 9890
rect 752 9856 768 9890
rect 808 9840 818 9874
rect 852 9840 918 9874
rect 952 9840 968 9874
rect 1008 9856 1018 9890
rect 1052 9856 1118 9890
rect 1152 9856 1168 9890
rect 1208 9840 1218 9874
rect 1252 9840 1318 9874
rect 1352 9840 1368 9874
rect 1408 9856 1418 9890
rect 1452 9856 1518 9890
rect 1552 9856 1568 9890
rect 1608 9840 1618 9874
rect 1652 9840 1718 9874
rect 1752 9840 1768 9874
rect 1808 9856 1818 9890
rect 1852 9856 1918 9890
rect 1952 9856 1968 9890
rect 2008 9840 2018 9874
rect 2052 9840 2118 9874
rect 2152 9840 2168 9874
rect 2208 9856 2218 9890
rect 2252 9856 2318 9890
rect 2352 9856 2368 9890
rect 2408 9840 2418 9874
rect 2452 9840 2518 9874
rect 2552 9840 2568 9874
rect 2608 9856 2618 9890
rect 2652 9856 2718 9890
rect 2752 9856 2768 9890
rect 2808 9840 2818 9874
rect 2852 9840 2918 9874
rect 2952 9840 2968 9874
rect 3008 9856 3018 9890
rect 3052 9856 3118 9890
rect 3152 9856 3168 9890
rect 3208 9840 3218 9874
rect 3252 9840 3318 9874
rect 3352 9840 3368 9874
rect 3408 9856 3418 9890
rect 3452 9856 3518 9890
rect 3552 9856 3568 9890
rect 3608 9840 3618 9874
rect 3652 9840 3718 9874
rect 3752 9840 3768 9874
rect 3808 9856 3818 9890
rect 3852 9856 3918 9890
rect 3952 9856 3968 9890
rect 4008 9840 4018 9874
rect 4052 9840 4118 9874
rect 4152 9840 4168 9874
rect 4208 9856 4218 9890
rect 4252 9856 4318 9890
rect 4352 9856 4368 9890
rect 4408 9840 4418 9874
rect 4452 9840 4518 9874
rect 4552 9840 4568 9874
rect 4608 9856 4618 9890
rect 4652 9856 4718 9890
rect 4752 9856 4768 9890
rect 4808 9840 4818 9874
rect 4852 9840 4918 9874
rect 4952 9840 4968 9874
rect 5008 9856 5018 9890
rect 5052 9856 5118 9890
rect 5152 9856 5168 9890
rect 5208 9840 5218 9874
rect 5252 9840 5318 9874
rect 5352 9840 5368 9874
rect 5408 9856 5418 9890
rect 5452 9856 5518 9890
rect 5552 9856 5568 9890
rect 5608 9840 5618 9874
rect 5652 9840 5718 9874
rect 5752 9840 5768 9874
rect 5808 9856 5818 9890
rect 5852 9856 5918 9890
rect 5952 9856 5968 9890
rect 6008 9840 6018 9874
rect 6052 9840 6118 9874
rect 6152 9840 6168 9874
rect 6208 9856 6218 9890
rect 6252 9856 6318 9890
rect 6352 9856 6368 9890
rect 6516 9871 6568 9888
rect 6550 9854 6568 9871
rect 6602 9854 6618 9888
rect 6652 9854 6668 9888
rect 6702 9859 6720 9888
rect 6702 9854 6754 9859
rect 6862 9854 6878 9888
rect 6912 9854 6928 9888
rect 6962 9854 6978 9888
rect 7012 9854 7028 9888
rect 7062 9854 7078 9888
rect 7112 9854 7128 9888
rect 7162 9854 7178 9888
rect 7212 9854 7228 9888
rect 7262 9854 7278 9888
rect 7312 9854 7328 9888
rect 7362 9854 7378 9888
rect 7412 9854 7428 9888
rect 6 9767 64 9793
rect 6 9733 18 9767
rect 52 9733 64 9767
rect 6 9707 64 9733
rect 106 9767 164 9793
rect 106 9733 118 9767
rect 152 9733 164 9767
rect 106 9707 164 9733
rect 206 9767 264 9793
rect 206 9733 218 9767
rect 252 9733 264 9767
rect 206 9707 264 9733
rect 306 9767 364 9793
rect 306 9733 318 9767
rect 352 9733 364 9767
rect 306 9707 364 9733
rect 406 9767 464 9793
rect 406 9733 418 9767
rect 452 9733 464 9767
rect 406 9707 464 9733
rect 506 9767 564 9793
rect 506 9733 518 9767
rect 552 9733 564 9767
rect 506 9707 564 9733
rect 606 9767 664 9793
rect 606 9733 618 9767
rect 652 9733 664 9767
rect 606 9707 664 9733
rect 706 9767 764 9793
rect 706 9733 718 9767
rect 752 9733 764 9767
rect 706 9707 764 9733
rect 806 9767 864 9793
rect 806 9733 818 9767
rect 852 9733 864 9767
rect 806 9707 864 9733
rect 906 9767 964 9793
rect 906 9733 918 9767
rect 952 9733 964 9767
rect 906 9707 964 9733
rect 1006 9767 1064 9793
rect 1006 9733 1018 9767
rect 1052 9733 1064 9767
rect 1006 9707 1064 9733
rect 1106 9767 1164 9793
rect 1106 9733 1118 9767
rect 1152 9733 1164 9767
rect 1106 9707 1164 9733
rect 1206 9767 1264 9793
rect 1206 9733 1218 9767
rect 1252 9733 1264 9767
rect 1206 9707 1264 9733
rect 1306 9767 1364 9793
rect 1306 9733 1318 9767
rect 1352 9733 1364 9767
rect 1306 9707 1364 9733
rect 1406 9767 1464 9793
rect 1406 9733 1418 9767
rect 1452 9733 1464 9767
rect 1406 9707 1464 9733
rect 1506 9767 1564 9793
rect 1506 9733 1512 9767
rect 1552 9733 1564 9767
rect 1506 9707 1564 9733
rect 1606 9767 1664 9793
rect 1606 9733 1618 9767
rect 1658 9733 1664 9767
rect 1606 9707 1664 9733
rect 1706 9767 1764 9793
rect 1706 9733 1718 9767
rect 1752 9733 1764 9767
rect 1706 9707 1764 9733
rect 1806 9767 1864 9793
rect 1806 9733 1818 9767
rect 1852 9733 1864 9767
rect 1806 9707 1864 9733
rect 1906 9767 1964 9793
rect 1906 9733 1918 9767
rect 1952 9733 1964 9767
rect 1906 9707 1964 9733
rect 2006 9767 2064 9793
rect 2006 9733 2018 9767
rect 2052 9733 2064 9767
rect 2006 9707 2064 9733
rect 2106 9767 2164 9793
rect 2106 9733 2112 9767
rect 2152 9733 2164 9767
rect 2106 9707 2164 9733
rect 2206 9767 2264 9793
rect 2206 9733 2218 9767
rect 2258 9733 2264 9767
rect 2206 9707 2264 9733
rect 2306 9767 2364 9793
rect 2306 9733 2318 9767
rect 2352 9733 2364 9767
rect 2306 9707 2364 9733
rect 2406 9767 2464 9793
rect 2406 9733 2418 9767
rect 2452 9733 2464 9767
rect 2406 9707 2464 9733
rect 2506 9767 2564 9793
rect 2506 9733 2518 9767
rect 2552 9733 2564 9767
rect 2506 9707 2564 9733
rect 2606 9767 2664 9793
rect 2606 9733 2618 9767
rect 2652 9733 2664 9767
rect 2606 9707 2664 9733
rect 2706 9767 2764 9793
rect 2706 9733 2712 9767
rect 2752 9733 2764 9767
rect 2706 9707 2764 9733
rect 2806 9767 2864 9793
rect 2806 9733 2818 9767
rect 2858 9733 2864 9767
rect 2806 9707 2864 9733
rect 2906 9767 2964 9793
rect 2906 9733 2918 9767
rect 2952 9733 2964 9767
rect 2906 9707 2964 9733
rect 3006 9767 3064 9793
rect 3006 9733 3018 9767
rect 3052 9733 3064 9767
rect 3006 9707 3064 9733
rect 3106 9767 3164 9793
rect 3106 9733 3118 9767
rect 3152 9733 3164 9767
rect 3106 9707 3164 9733
rect 3206 9767 3264 9793
rect 3206 9733 3212 9767
rect 3252 9733 3264 9767
rect 3206 9707 3264 9733
rect 3306 9767 3364 9793
rect 3306 9733 3318 9767
rect 3358 9733 3364 9767
rect 3306 9707 3364 9733
rect 3406 9767 3464 9793
rect 3406 9733 3418 9767
rect 3452 9733 3464 9767
rect 3406 9707 3464 9733
rect 3506 9767 3564 9793
rect 3506 9733 3512 9767
rect 3552 9733 3564 9767
rect 3506 9707 3564 9733
rect 3606 9767 3664 9793
rect 3606 9733 3618 9767
rect 3658 9733 3664 9767
rect 3606 9707 3664 9733
rect 3706 9767 3764 9793
rect 3706 9733 3718 9767
rect 3752 9733 3764 9767
rect 3706 9707 3764 9733
rect 3806 9767 3864 9793
rect 3806 9733 3818 9767
rect 3852 9733 3864 9767
rect 3806 9707 3864 9733
rect 3906 9767 3964 9793
rect 3906 9733 3918 9767
rect 3952 9733 3964 9767
rect 3906 9707 3964 9733
rect 4006 9767 4064 9793
rect 4006 9733 4018 9767
rect 4052 9733 4064 9767
rect 4006 9707 4064 9733
rect 4106 9767 4164 9793
rect 4106 9733 4118 9767
rect 4152 9733 4164 9767
rect 4106 9707 4164 9733
rect 4206 9767 4264 9793
rect 4206 9733 4218 9767
rect 4252 9733 4264 9767
rect 4206 9707 4264 9733
rect 4306 9767 4364 9793
rect 4306 9733 4318 9767
rect 4352 9733 4364 9767
rect 4306 9707 4364 9733
rect 4406 9767 4464 9793
rect 4406 9733 4418 9767
rect 4452 9733 4464 9767
rect 4406 9707 4464 9733
rect 4506 9767 4564 9793
rect 4506 9733 4518 9767
rect 4552 9733 4564 9767
rect 4506 9707 4564 9733
rect 4606 9767 4664 9793
rect 4606 9733 4618 9767
rect 4652 9733 4664 9767
rect 4606 9707 4664 9733
rect 4706 9767 4764 9793
rect 4706 9733 4718 9767
rect 4752 9733 4764 9767
rect 4706 9707 4764 9733
rect 4806 9767 4864 9793
rect 4806 9733 4818 9767
rect 4852 9733 4864 9767
rect 4806 9707 4864 9733
rect 4906 9767 4964 9793
rect 4906 9733 4918 9767
rect 4952 9733 4964 9767
rect 4906 9707 4964 9733
rect 5006 9767 5064 9793
rect 5006 9733 5018 9767
rect 5052 9733 5064 9767
rect 5006 9707 5064 9733
rect 5106 9767 5164 9793
rect 5106 9733 5118 9767
rect 5152 9733 5164 9767
rect 5106 9707 5164 9733
rect 5206 9767 5264 9793
rect 5206 9733 5218 9767
rect 5252 9733 5264 9767
rect 5206 9707 5264 9733
rect 5306 9767 5364 9793
rect 5306 9733 5318 9767
rect 5352 9733 5364 9767
rect 5306 9707 5364 9733
rect 5406 9767 5464 9793
rect 5406 9733 5412 9767
rect 5452 9733 5464 9767
rect 5406 9707 5464 9733
rect 5506 9767 5564 9793
rect 5506 9733 5518 9767
rect 5558 9733 5564 9767
rect 5506 9707 5564 9733
rect 5606 9767 5664 9793
rect 5606 9733 5618 9767
rect 5652 9733 5664 9767
rect 5606 9707 5664 9733
rect 5706 9767 5764 9793
rect 5706 9733 5712 9767
rect 5752 9733 5764 9767
rect 5706 9707 5764 9733
rect 5806 9767 5864 9793
rect 5806 9733 5818 9767
rect 5858 9733 5864 9767
rect 5806 9707 5864 9733
rect 5906 9767 5964 9793
rect 5906 9733 5912 9767
rect 5952 9733 5964 9767
rect 5906 9707 5964 9733
rect 6006 9767 6064 9793
rect 6006 9733 6018 9767
rect 6058 9733 6064 9767
rect 6006 9707 6064 9733
rect 6106 9767 6164 9793
rect 6106 9733 6118 9767
rect 6152 9733 6164 9767
rect 6106 9707 6164 9733
rect 6206 9767 6264 9793
rect 6206 9733 6218 9767
rect 6252 9733 6264 9767
rect 6206 9707 6264 9733
rect 6306 9767 6364 9793
rect 6306 9733 6318 9767
rect 6352 9733 6364 9767
rect 6306 9707 6364 9733
rect 6406 9767 6464 9793
rect 6618 9786 6862 9820
rect 6406 9733 6412 9767
rect 6452 9733 6464 9767
rect 6508 9748 6516 9782
rect 6558 9748 6574 9782
rect 6618 9767 6652 9786
rect 6406 9707 6464 9733
rect 6828 9783 6862 9786
rect 6828 9767 6962 9783
rect 6618 9717 6652 9733
rect 6696 9718 6712 9752
rect 6754 9718 6762 9752
rect 6862 9733 6928 9767
rect 6828 9717 6962 9733
rect 7028 9767 7162 9783
rect 7062 9733 7128 9767
rect 7028 9717 7162 9733
rect 7228 9767 7362 9783
rect 7262 9733 7328 9767
rect 7228 9717 7362 9733
rect 7428 9767 7462 9783
rect 7428 9717 7462 9733
rect 6 9627 64 9653
rect 6 9593 18 9627
rect 52 9593 64 9627
rect 6 9567 64 9593
rect 106 9627 164 9653
rect 106 9593 118 9627
rect 152 9593 164 9627
rect 106 9567 164 9593
rect 206 9627 264 9653
rect 206 9593 218 9627
rect 252 9593 264 9627
rect 206 9567 264 9593
rect 306 9627 364 9653
rect 306 9593 318 9627
rect 352 9593 364 9627
rect 306 9567 364 9593
rect 406 9627 464 9653
rect 406 9593 418 9627
rect 452 9593 464 9627
rect 406 9567 464 9593
rect 506 9627 564 9653
rect 506 9593 518 9627
rect 552 9593 564 9627
rect 506 9567 564 9593
rect 606 9627 664 9653
rect 606 9593 612 9627
rect 652 9593 664 9627
rect 606 9567 664 9593
rect 706 9627 764 9653
rect 706 9593 718 9627
rect 758 9593 764 9627
rect 706 9567 764 9593
rect 806 9627 864 9653
rect 806 9593 818 9627
rect 852 9593 864 9627
rect 806 9567 864 9593
rect 906 9627 964 9653
rect 906 9593 918 9627
rect 952 9593 964 9627
rect 906 9567 964 9593
rect 1006 9627 1064 9653
rect 1006 9593 1018 9627
rect 1052 9593 1064 9627
rect 1006 9567 1064 9593
rect 1106 9627 1164 9653
rect 1106 9593 1118 9627
rect 1152 9593 1164 9627
rect 1106 9567 1164 9593
rect 1206 9627 1264 9653
rect 1206 9593 1218 9627
rect 1252 9593 1264 9627
rect 1206 9567 1264 9593
rect 1306 9627 1364 9653
rect 1306 9593 1318 9627
rect 1352 9593 1364 9627
rect 1306 9567 1364 9593
rect 1406 9627 1464 9653
rect 1406 9593 1418 9627
rect 1452 9593 1464 9627
rect 1406 9567 1464 9593
rect 1506 9627 1564 9653
rect 1506 9593 1518 9627
rect 1552 9593 1564 9627
rect 1506 9567 1564 9593
rect 1606 9627 1664 9653
rect 1606 9593 1618 9627
rect 1652 9593 1664 9627
rect 1606 9567 1664 9593
rect 1706 9627 1764 9653
rect 1706 9593 1718 9627
rect 1752 9593 1764 9627
rect 1706 9567 1764 9593
rect 1806 9627 1864 9653
rect 1806 9593 1818 9627
rect 1852 9593 1864 9627
rect 1806 9567 1864 9593
rect 1906 9627 1964 9653
rect 1906 9593 1918 9627
rect 1952 9593 1964 9627
rect 1906 9567 1964 9593
rect 2006 9627 2064 9653
rect 2006 9593 2018 9627
rect 2052 9593 2064 9627
rect 2006 9567 2064 9593
rect 2106 9627 2164 9653
rect 2106 9593 2112 9627
rect 2152 9593 2164 9627
rect 2106 9567 2164 9593
rect 2206 9627 2264 9653
rect 2206 9593 2218 9627
rect 2258 9593 2264 9627
rect 2206 9567 2264 9593
rect 2306 9627 2364 9653
rect 2306 9593 2312 9627
rect 2352 9593 2364 9627
rect 2306 9567 2364 9593
rect 2406 9627 2464 9653
rect 2406 9593 2418 9627
rect 2458 9593 2464 9627
rect 2406 9567 2464 9593
rect 2506 9627 2564 9653
rect 2506 9593 2518 9627
rect 2552 9593 2564 9627
rect 2506 9567 2564 9593
rect 2606 9627 2664 9653
rect 2606 9593 2618 9627
rect 2652 9593 2664 9627
rect 2606 9567 2664 9593
rect 2706 9627 2764 9653
rect 2706 9593 2718 9627
rect 2752 9593 2764 9627
rect 2706 9567 2764 9593
rect 2806 9627 2864 9653
rect 2806 9593 2818 9627
rect 2852 9593 2864 9627
rect 2806 9567 2864 9593
rect 2906 9627 2964 9653
rect 2906 9593 2912 9627
rect 2952 9593 2964 9627
rect 2906 9567 2964 9593
rect 3006 9627 3064 9653
rect 3006 9593 3018 9627
rect 3058 9593 3064 9627
rect 3006 9567 3064 9593
rect 3106 9627 3164 9653
rect 3106 9593 3118 9627
rect 3152 9593 3164 9627
rect 3106 9567 3164 9593
rect 3206 9627 3264 9653
rect 3206 9593 3218 9627
rect 3252 9593 3264 9627
rect 3206 9567 3264 9593
rect 3306 9627 3364 9653
rect 3306 9593 3318 9627
rect 3352 9593 3364 9627
rect 3306 9567 3364 9593
rect 3406 9627 3464 9653
rect 3406 9593 3418 9627
rect 3452 9593 3464 9627
rect 3406 9567 3464 9593
rect 3506 9627 3564 9653
rect 3506 9593 3518 9627
rect 3552 9593 3564 9627
rect 3506 9567 3564 9593
rect 3606 9627 3664 9653
rect 3606 9593 3618 9627
rect 3652 9593 3664 9627
rect 3606 9567 3664 9593
rect 3706 9627 3764 9653
rect 3706 9593 3718 9627
rect 3752 9593 3764 9627
rect 3706 9567 3764 9593
rect 3806 9627 3864 9653
rect 3806 9593 3818 9627
rect 3852 9593 3864 9627
rect 3806 9567 3864 9593
rect 3906 9627 3964 9653
rect 3906 9593 3918 9627
rect 3952 9593 3964 9627
rect 3906 9567 3964 9593
rect 4006 9627 4064 9653
rect 4006 9593 4012 9627
rect 4052 9593 4064 9627
rect 4006 9567 4064 9593
rect 4106 9627 4164 9653
rect 4106 9593 4118 9627
rect 4158 9593 4164 9627
rect 4106 9567 4164 9593
rect 4206 9627 4264 9653
rect 4206 9593 4218 9627
rect 4252 9593 4264 9627
rect 4206 9567 4264 9593
rect 4306 9627 4364 9653
rect 4306 9593 4318 9627
rect 4352 9593 4364 9627
rect 4306 9567 4364 9593
rect 4406 9627 4464 9653
rect 4406 9593 4418 9627
rect 4452 9593 4464 9627
rect 4406 9567 4464 9593
rect 4506 9627 4564 9653
rect 4506 9593 4518 9627
rect 4552 9593 4564 9627
rect 4506 9567 4564 9593
rect 4606 9627 4664 9653
rect 4606 9593 4618 9627
rect 4652 9593 4664 9627
rect 4606 9567 4664 9593
rect 4706 9627 4764 9653
rect 4706 9593 4718 9627
rect 4752 9593 4764 9627
rect 4706 9567 4764 9593
rect 4806 9627 4864 9653
rect 4806 9593 4818 9627
rect 4852 9593 4864 9627
rect 4806 9567 4864 9593
rect 4906 9627 4964 9653
rect 4906 9593 4918 9627
rect 4952 9593 4964 9627
rect 4906 9567 4964 9593
rect 5006 9627 5064 9653
rect 5006 9593 5018 9627
rect 5052 9593 5064 9627
rect 5006 9567 5064 9593
rect 5106 9627 5164 9653
rect 5106 9593 5118 9627
rect 5152 9593 5164 9627
rect 5106 9567 5164 9593
rect 5206 9627 5264 9653
rect 5206 9593 5218 9627
rect 5252 9593 5264 9627
rect 5206 9567 5264 9593
rect 5306 9627 5364 9653
rect 5306 9593 5318 9627
rect 5352 9593 5364 9627
rect 5306 9567 5364 9593
rect 5406 9627 5464 9653
rect 5406 9593 5418 9627
rect 5452 9593 5464 9627
rect 5406 9567 5464 9593
rect 5506 9627 5564 9653
rect 5506 9593 5518 9627
rect 5552 9593 5564 9627
rect 5506 9567 5564 9593
rect 5606 9627 5664 9653
rect 5606 9593 5618 9627
rect 5652 9593 5664 9627
rect 5606 9567 5664 9593
rect 5706 9627 5764 9653
rect 5706 9593 5718 9627
rect 5752 9593 5764 9627
rect 5706 9567 5764 9593
rect 5806 9627 5864 9653
rect 5806 9593 5818 9627
rect 5852 9593 5864 9627
rect 5806 9567 5864 9593
rect 5906 9627 5964 9653
rect 5906 9593 5912 9627
rect 5952 9593 5964 9627
rect 5906 9567 5964 9593
rect 6006 9627 6064 9653
rect 6006 9593 6018 9627
rect 6058 9593 6064 9627
rect 6006 9567 6064 9593
rect 6106 9627 6164 9653
rect 6106 9593 6118 9627
rect 6152 9593 6164 9627
rect 6106 9567 6164 9593
rect 6206 9627 6264 9653
rect 6206 9593 6218 9627
rect 6252 9593 6264 9627
rect 6206 9567 6264 9593
rect 6306 9627 6364 9653
rect 6306 9593 6318 9627
rect 6352 9593 6364 9627
rect 6306 9567 6364 9593
rect 6406 9627 6464 9653
rect 6618 9646 6862 9680
rect 6406 9593 6412 9627
rect 6452 9593 6464 9627
rect 6508 9608 6516 9642
rect 6558 9608 6574 9642
rect 6618 9627 6652 9646
rect 6406 9567 6464 9593
rect 6828 9627 6862 9646
rect 6618 9577 6652 9593
rect 6696 9578 6712 9612
rect 6754 9578 6762 9612
rect 6828 9577 6862 9593
rect 6928 9627 7162 9643
rect 6962 9593 7028 9627
rect 7062 9593 7128 9627
rect 6928 9577 7162 9593
rect 7228 9627 7362 9643
rect 7262 9593 7328 9627
rect 7228 9577 7362 9593
rect 7428 9627 7462 9643
rect 7428 9577 7462 9593
rect 6 9487 64 9513
rect 6 9453 18 9487
rect 52 9453 64 9487
rect 6 9427 64 9453
rect 106 9487 164 9513
rect 106 9453 118 9487
rect 152 9453 164 9487
rect 106 9427 164 9453
rect 206 9487 264 9513
rect 206 9453 218 9487
rect 252 9453 264 9487
rect 206 9427 264 9453
rect 306 9487 364 9513
rect 306 9453 318 9487
rect 352 9453 364 9487
rect 306 9427 364 9453
rect 406 9487 464 9513
rect 406 9453 412 9487
rect 452 9453 464 9487
rect 406 9427 464 9453
rect 506 9487 564 9513
rect 506 9453 518 9487
rect 558 9453 564 9487
rect 506 9427 564 9453
rect 606 9487 664 9513
rect 606 9453 618 9487
rect 652 9453 664 9487
rect 606 9427 664 9453
rect 706 9487 764 9513
rect 706 9453 718 9487
rect 752 9453 764 9487
rect 706 9427 764 9453
rect 806 9487 864 9513
rect 806 9453 818 9487
rect 852 9453 864 9487
rect 806 9427 864 9453
rect 906 9487 964 9513
rect 906 9453 912 9487
rect 952 9453 964 9487
rect 906 9427 964 9453
rect 1006 9487 1064 9513
rect 1006 9453 1018 9487
rect 1058 9453 1064 9487
rect 1006 9427 1064 9453
rect 1106 9487 1164 9513
rect 1106 9453 1112 9487
rect 1152 9453 1164 9487
rect 1106 9427 1164 9453
rect 1206 9487 1264 9513
rect 1206 9453 1218 9487
rect 1258 9453 1264 9487
rect 1206 9427 1264 9453
rect 1306 9487 1364 9513
rect 1306 9453 1318 9487
rect 1352 9453 1364 9487
rect 1306 9427 1364 9453
rect 1406 9487 1464 9513
rect 1406 9453 1418 9487
rect 1452 9453 1464 9487
rect 1406 9427 1464 9453
rect 1506 9487 1564 9513
rect 1506 9453 1518 9487
rect 1552 9453 1564 9487
rect 1506 9427 1564 9453
rect 1606 9487 1664 9513
rect 1606 9453 1618 9487
rect 1652 9453 1664 9487
rect 1606 9427 1664 9453
rect 1706 9487 1764 9513
rect 1706 9453 1712 9487
rect 1752 9453 1764 9487
rect 1706 9427 1764 9453
rect 1806 9487 1864 9513
rect 1806 9453 1818 9487
rect 1858 9453 1864 9487
rect 1806 9427 1864 9453
rect 1906 9487 1964 9513
rect 1906 9453 1918 9487
rect 1952 9453 1964 9487
rect 1906 9427 1964 9453
rect 2006 9487 2064 9513
rect 2006 9453 2012 9487
rect 2052 9453 2064 9487
rect 2006 9427 2064 9453
rect 2106 9487 2164 9513
rect 2106 9453 2118 9487
rect 2158 9453 2164 9487
rect 2106 9427 2164 9453
rect 2206 9487 2264 9513
rect 2206 9453 2218 9487
rect 2252 9453 2264 9487
rect 2206 9427 2264 9453
rect 2306 9487 2364 9513
rect 2306 9453 2312 9487
rect 2352 9453 2364 9487
rect 2306 9427 2364 9453
rect 2406 9487 2464 9513
rect 2406 9453 2418 9487
rect 2458 9453 2464 9487
rect 2406 9427 2464 9453
rect 2506 9487 2564 9513
rect 2506 9453 2512 9487
rect 2552 9453 2564 9487
rect 2506 9427 2564 9453
rect 2606 9487 2664 9513
rect 2606 9453 2618 9487
rect 2658 9453 2664 9487
rect 2606 9427 2664 9453
rect 2706 9487 2764 9513
rect 2706 9453 2712 9487
rect 2752 9453 2764 9487
rect 2706 9427 2764 9453
rect 2806 9487 2864 9513
rect 2806 9453 2818 9487
rect 2858 9453 2864 9487
rect 2806 9427 2864 9453
rect 2906 9487 2964 9513
rect 2906 9453 2918 9487
rect 2952 9453 2964 9487
rect 2906 9427 2964 9453
rect 3006 9487 3064 9513
rect 3006 9453 3018 9487
rect 3052 9453 3064 9487
rect 3006 9427 3064 9453
rect 3106 9487 3164 9513
rect 3106 9453 3118 9487
rect 3152 9453 3164 9487
rect 3106 9427 3164 9453
rect 3206 9487 3264 9513
rect 3206 9453 3218 9487
rect 3252 9453 3264 9487
rect 3206 9427 3264 9453
rect 3306 9487 3364 9513
rect 3306 9453 3318 9487
rect 3352 9453 3364 9487
rect 3306 9427 3364 9453
rect 3406 9487 3464 9513
rect 3406 9453 3418 9487
rect 3452 9453 3464 9487
rect 3406 9427 3464 9453
rect 3506 9487 3564 9513
rect 3506 9453 3518 9487
rect 3552 9453 3564 9487
rect 3506 9427 3564 9453
rect 3606 9487 3664 9513
rect 3606 9453 3618 9487
rect 3652 9453 3664 9487
rect 3606 9427 3664 9453
rect 3706 9487 3764 9513
rect 3706 9453 3718 9487
rect 3752 9453 3764 9487
rect 3706 9427 3764 9453
rect 3806 9487 3864 9513
rect 3806 9453 3818 9487
rect 3852 9453 3864 9487
rect 3806 9427 3864 9453
rect 3906 9487 3964 9513
rect 3906 9453 3918 9487
rect 3952 9453 3964 9487
rect 3906 9427 3964 9453
rect 4006 9487 4064 9513
rect 4006 9453 4012 9487
rect 4052 9453 4064 9487
rect 4006 9427 4064 9453
rect 4106 9487 4164 9513
rect 4106 9453 4118 9487
rect 4158 9453 4164 9487
rect 4106 9427 4164 9453
rect 4206 9487 4264 9513
rect 4206 9453 4218 9487
rect 4252 9453 4264 9487
rect 4206 9427 4264 9453
rect 4306 9487 4364 9513
rect 4306 9453 4318 9487
rect 4352 9453 4364 9487
rect 4306 9427 4364 9453
rect 4406 9487 4464 9513
rect 4406 9453 4418 9487
rect 4452 9453 4464 9487
rect 4406 9427 4464 9453
rect 4506 9487 4564 9513
rect 4506 9453 4512 9487
rect 4552 9453 4564 9487
rect 4506 9427 4564 9453
rect 4606 9487 4664 9513
rect 4606 9453 4618 9487
rect 4658 9453 4664 9487
rect 4606 9427 4664 9453
rect 4706 9487 4764 9513
rect 4706 9453 4718 9487
rect 4752 9453 4764 9487
rect 4706 9427 4764 9453
rect 4806 9487 4864 9513
rect 4806 9453 4812 9487
rect 4852 9453 4864 9487
rect 4806 9427 4864 9453
rect 4906 9487 4964 9513
rect 4906 9453 4918 9487
rect 4958 9453 4964 9487
rect 4906 9427 4964 9453
rect 5006 9487 5064 9513
rect 5006 9453 5012 9487
rect 5052 9453 5064 9487
rect 5006 9427 5064 9453
rect 5106 9487 5164 9513
rect 5106 9453 5118 9487
rect 5158 9453 5164 9487
rect 5106 9427 5164 9453
rect 5206 9487 5264 9513
rect 5206 9453 5212 9487
rect 5252 9453 5264 9487
rect 5206 9427 5264 9453
rect 5306 9487 5364 9513
rect 5306 9453 5318 9487
rect 5358 9453 5364 9487
rect 5306 9427 5364 9453
rect 5406 9487 5464 9513
rect 5406 9453 5418 9487
rect 5452 9453 5464 9487
rect 5406 9427 5464 9453
rect 5506 9487 5564 9513
rect 5506 9453 5518 9487
rect 5552 9453 5564 9487
rect 5506 9427 5564 9453
rect 5606 9487 5664 9513
rect 5606 9453 5612 9487
rect 5652 9453 5664 9487
rect 5606 9427 5664 9453
rect 5706 9487 5764 9513
rect 5706 9453 5718 9487
rect 5758 9453 5764 9487
rect 5706 9427 5764 9453
rect 5806 9487 5864 9513
rect 5806 9453 5812 9487
rect 5852 9453 5864 9487
rect 5806 9427 5864 9453
rect 5906 9487 5964 9513
rect 5906 9453 5918 9487
rect 5958 9453 5964 9487
rect 5906 9427 5964 9453
rect 6006 9487 6064 9513
rect 6006 9453 6018 9487
rect 6052 9453 6064 9487
rect 6006 9427 6064 9453
rect 6106 9487 6164 9513
rect 6106 9453 6112 9487
rect 6152 9453 6164 9487
rect 6106 9427 6164 9453
rect 6206 9487 6264 9513
rect 6206 9453 6218 9487
rect 6258 9453 6264 9487
rect 6206 9427 6264 9453
rect 6306 9487 6364 9513
rect 6306 9453 6318 9487
rect 6352 9453 6364 9487
rect 6306 9427 6364 9453
rect 6406 9487 6464 9513
rect 6618 9506 6862 9540
rect 6406 9453 6412 9487
rect 6452 9453 6464 9487
rect 6508 9468 6516 9502
rect 6558 9468 6574 9502
rect 6618 9487 6652 9506
rect 6406 9427 6464 9453
rect 6828 9503 6862 9506
rect 6828 9487 6962 9503
rect 6618 9437 6652 9453
rect 6696 9438 6712 9472
rect 6754 9438 6762 9472
rect 6862 9453 6928 9487
rect 6828 9437 6962 9453
rect 7028 9487 7062 9503
rect 7028 9437 7062 9453
rect 7128 9487 7362 9503
rect 7162 9453 7228 9487
rect 7262 9453 7328 9487
rect 7128 9437 7362 9453
rect 7428 9487 7462 9503
rect 7428 9437 7462 9453
rect 6 9347 64 9373
rect 6 9313 18 9347
rect 52 9313 64 9347
rect 6 9287 64 9313
rect 106 9347 164 9373
rect 106 9313 118 9347
rect 152 9313 164 9347
rect 106 9287 164 9313
rect 206 9347 264 9373
rect 206 9313 218 9347
rect 252 9313 264 9347
rect 206 9287 264 9313
rect 306 9347 364 9373
rect 306 9313 318 9347
rect 352 9313 364 9347
rect 306 9287 364 9313
rect 406 9347 464 9373
rect 406 9313 418 9347
rect 452 9313 464 9347
rect 406 9287 464 9313
rect 506 9347 564 9373
rect 506 9313 518 9347
rect 552 9313 564 9347
rect 506 9287 564 9313
rect 606 9347 664 9373
rect 606 9313 618 9347
rect 652 9313 664 9347
rect 606 9287 664 9313
rect 706 9347 764 9373
rect 706 9313 718 9347
rect 752 9313 764 9347
rect 706 9287 764 9313
rect 806 9347 864 9373
rect 806 9313 818 9347
rect 852 9313 864 9347
rect 806 9287 864 9313
rect 906 9347 964 9373
rect 906 9313 918 9347
rect 952 9313 964 9347
rect 906 9287 964 9313
rect 1006 9347 1064 9373
rect 1006 9313 1018 9347
rect 1052 9313 1064 9347
rect 1006 9287 1064 9313
rect 1106 9347 1164 9373
rect 1106 9313 1118 9347
rect 1152 9313 1164 9347
rect 1106 9287 1164 9313
rect 1206 9347 1264 9373
rect 1206 9313 1218 9347
rect 1252 9313 1264 9347
rect 1206 9287 1264 9313
rect 1306 9347 1364 9373
rect 1306 9313 1318 9347
rect 1352 9313 1364 9347
rect 1306 9287 1364 9313
rect 1406 9347 1464 9373
rect 1406 9313 1418 9347
rect 1452 9313 1464 9347
rect 1406 9287 1464 9313
rect 1506 9347 1564 9373
rect 1506 9313 1518 9347
rect 1552 9313 1564 9347
rect 1506 9287 1564 9313
rect 1606 9347 1664 9373
rect 1606 9313 1618 9347
rect 1652 9313 1664 9347
rect 1606 9287 1664 9313
rect 1706 9347 1764 9373
rect 1706 9313 1712 9347
rect 1752 9313 1764 9347
rect 1706 9287 1764 9313
rect 1806 9347 1864 9373
rect 1806 9313 1818 9347
rect 1858 9313 1864 9347
rect 1806 9287 1864 9313
rect 1906 9347 1964 9373
rect 1906 9313 1918 9347
rect 1952 9313 1964 9347
rect 1906 9287 1964 9313
rect 2006 9347 2064 9373
rect 2006 9313 2018 9347
rect 2052 9313 2064 9347
rect 2006 9287 2064 9313
rect 2106 9347 2164 9373
rect 2106 9313 2118 9347
rect 2152 9313 2164 9347
rect 2106 9287 2164 9313
rect 2206 9347 2264 9373
rect 2206 9313 2218 9347
rect 2252 9313 2264 9347
rect 2206 9287 2264 9313
rect 2306 9347 2364 9373
rect 2306 9313 2318 9347
rect 2352 9313 2364 9347
rect 2306 9287 2364 9313
rect 2406 9347 2464 9373
rect 2406 9313 2418 9347
rect 2452 9313 2464 9347
rect 2406 9287 2464 9313
rect 2506 9347 2564 9373
rect 2506 9313 2518 9347
rect 2552 9313 2564 9347
rect 2506 9287 2564 9313
rect 2606 9347 2664 9373
rect 2606 9313 2618 9347
rect 2652 9313 2664 9347
rect 2606 9287 2664 9313
rect 2706 9347 2764 9373
rect 2706 9313 2718 9347
rect 2752 9313 2764 9347
rect 2706 9287 2764 9313
rect 2806 9347 2864 9373
rect 2806 9313 2818 9347
rect 2852 9313 2864 9347
rect 2806 9287 2864 9313
rect 2906 9347 2964 9373
rect 2906 9313 2918 9347
rect 2952 9313 2964 9347
rect 2906 9287 2964 9313
rect 3006 9347 3064 9373
rect 3006 9313 3018 9347
rect 3052 9313 3064 9347
rect 3006 9287 3064 9313
rect 3106 9347 3164 9373
rect 3106 9313 3118 9347
rect 3152 9313 3164 9347
rect 3106 9287 3164 9313
rect 3206 9347 3264 9373
rect 3206 9313 3218 9347
rect 3252 9313 3264 9347
rect 3206 9287 3264 9313
rect 3306 9347 3364 9373
rect 3306 9313 3318 9347
rect 3352 9313 3364 9347
rect 3306 9287 3364 9313
rect 3406 9347 3464 9373
rect 3406 9313 3418 9347
rect 3452 9313 3464 9347
rect 3406 9287 3464 9313
rect 3506 9347 3564 9373
rect 3506 9313 3518 9347
rect 3552 9313 3564 9347
rect 3506 9287 3564 9313
rect 3606 9347 3664 9373
rect 3606 9313 3618 9347
rect 3652 9313 3664 9347
rect 3606 9287 3664 9313
rect 3706 9347 3764 9373
rect 3706 9313 3718 9347
rect 3752 9313 3764 9347
rect 3706 9287 3764 9313
rect 3806 9347 3864 9373
rect 3806 9313 3818 9347
rect 3852 9313 3864 9347
rect 3806 9287 3864 9313
rect 3906 9347 3964 9373
rect 3906 9313 3918 9347
rect 3952 9313 3964 9347
rect 3906 9287 3964 9313
rect 4006 9347 4064 9373
rect 4006 9313 4018 9347
rect 4052 9313 4064 9347
rect 4006 9287 4064 9313
rect 4106 9347 4164 9373
rect 4106 9313 4112 9347
rect 4152 9313 4164 9347
rect 4106 9287 4164 9313
rect 4206 9347 4264 9373
rect 4206 9313 4218 9347
rect 4258 9313 4264 9347
rect 4206 9287 4264 9313
rect 4306 9347 4364 9373
rect 4306 9313 4318 9347
rect 4352 9313 4364 9347
rect 4306 9287 4364 9313
rect 4406 9347 4464 9373
rect 4406 9313 4418 9347
rect 4452 9313 4464 9347
rect 4406 9287 4464 9313
rect 4506 9347 4564 9373
rect 4506 9313 4518 9347
rect 4552 9313 4564 9347
rect 4506 9287 4564 9313
rect 4606 9347 4664 9373
rect 4606 9313 4618 9347
rect 4652 9313 4664 9347
rect 4606 9287 4664 9313
rect 4706 9347 4764 9373
rect 4706 9313 4718 9347
rect 4752 9313 4764 9347
rect 4706 9287 4764 9313
rect 4806 9347 4864 9373
rect 4806 9313 4818 9347
rect 4852 9313 4864 9347
rect 4806 9287 4864 9313
rect 4906 9347 4964 9373
rect 4906 9313 4918 9347
rect 4952 9313 4964 9347
rect 4906 9287 4964 9313
rect 5006 9347 5064 9373
rect 5006 9313 5018 9347
rect 5052 9313 5064 9347
rect 5006 9287 5064 9313
rect 5106 9347 5164 9373
rect 5106 9313 5118 9347
rect 5152 9313 5164 9347
rect 5106 9287 5164 9313
rect 5206 9347 5264 9373
rect 5206 9313 5218 9347
rect 5252 9313 5264 9347
rect 5206 9287 5264 9313
rect 5306 9347 5364 9373
rect 5306 9313 5318 9347
rect 5352 9313 5364 9347
rect 5306 9287 5364 9313
rect 5406 9347 5464 9373
rect 5406 9313 5418 9347
rect 5452 9313 5464 9347
rect 5406 9287 5464 9313
rect 5506 9347 5564 9373
rect 5506 9313 5518 9347
rect 5552 9313 5564 9347
rect 5506 9287 5564 9313
rect 5606 9347 5664 9373
rect 5606 9313 5618 9347
rect 5652 9313 5664 9347
rect 5606 9287 5664 9313
rect 5706 9347 5764 9373
rect 5706 9313 5718 9347
rect 5752 9313 5764 9347
rect 5706 9287 5764 9313
rect 5806 9347 5864 9373
rect 5806 9313 5818 9347
rect 5852 9313 5864 9347
rect 5806 9287 5864 9313
rect 5906 9347 5964 9373
rect 5906 9313 5918 9347
rect 5952 9313 5964 9347
rect 5906 9287 5964 9313
rect 6006 9347 6064 9373
rect 6006 9313 6018 9347
rect 6052 9313 6064 9347
rect 6006 9287 6064 9313
rect 6106 9347 6164 9373
rect 6106 9313 6118 9347
rect 6152 9313 6164 9347
rect 6106 9287 6164 9313
rect 6206 9347 6264 9373
rect 6206 9313 6218 9347
rect 6252 9313 6264 9347
rect 6206 9287 6264 9313
rect 6306 9347 6364 9373
rect 6306 9313 6318 9347
rect 6352 9313 6364 9347
rect 6306 9287 6364 9313
rect 6406 9347 6464 9373
rect 6618 9366 6862 9400
rect 6406 9313 6412 9347
rect 6452 9313 6464 9347
rect 6508 9328 6516 9362
rect 6558 9328 6574 9362
rect 6618 9347 6652 9366
rect 6406 9287 6464 9313
rect 6828 9347 6862 9366
rect 6618 9297 6652 9313
rect 6696 9298 6712 9332
rect 6754 9298 6762 9332
rect 6828 9297 6862 9313
rect 6928 9347 7062 9363
rect 6962 9313 7028 9347
rect 6928 9297 7062 9313
rect 7128 9347 7362 9363
rect 7162 9313 7228 9347
rect 7262 9313 7328 9347
rect 7128 9297 7362 9313
rect 7428 9347 7462 9363
rect 7428 9297 7462 9313
rect 6 9207 64 9233
rect 6 9173 18 9207
rect 58 9173 64 9207
rect 6 9147 64 9173
rect 106 9207 164 9233
rect 106 9173 118 9207
rect 152 9173 164 9207
rect 106 9147 164 9173
rect 206 9207 264 9233
rect 206 9173 218 9207
rect 252 9173 264 9207
rect 206 9147 264 9173
rect 306 9207 364 9233
rect 306 9173 318 9207
rect 352 9173 364 9207
rect 306 9147 364 9173
rect 406 9207 464 9233
rect 406 9173 418 9207
rect 452 9173 464 9207
rect 406 9147 464 9173
rect 506 9207 564 9233
rect 506 9173 518 9207
rect 552 9173 564 9207
rect 506 9147 564 9173
rect 606 9207 664 9233
rect 606 9173 618 9207
rect 652 9173 664 9207
rect 606 9147 664 9173
rect 706 9207 764 9233
rect 706 9173 718 9207
rect 752 9173 764 9207
rect 706 9147 764 9173
rect 806 9207 864 9233
rect 806 9173 818 9207
rect 852 9173 864 9207
rect 806 9147 864 9173
rect 906 9207 964 9233
rect 906 9173 918 9207
rect 952 9173 964 9207
rect 906 9147 964 9173
rect 1006 9207 1064 9233
rect 1006 9173 1018 9207
rect 1052 9173 1064 9207
rect 1006 9147 1064 9173
rect 1106 9207 1164 9233
rect 1106 9173 1118 9207
rect 1152 9173 1164 9207
rect 1106 9147 1164 9173
rect 1206 9207 1264 9233
rect 1206 9173 1218 9207
rect 1252 9173 1264 9207
rect 1206 9147 1264 9173
rect 1306 9207 1364 9233
rect 1306 9173 1318 9207
rect 1352 9173 1364 9207
rect 1306 9147 1364 9173
rect 1406 9207 1464 9233
rect 1406 9173 1418 9207
rect 1452 9173 1464 9207
rect 1406 9147 1464 9173
rect 1506 9207 1564 9233
rect 1506 9173 1512 9207
rect 1552 9173 1564 9207
rect 1506 9147 1564 9173
rect 1606 9207 1664 9233
rect 1606 9173 1618 9207
rect 1658 9173 1664 9207
rect 1606 9147 1664 9173
rect 1706 9207 1764 9233
rect 1706 9173 1718 9207
rect 1752 9173 1764 9207
rect 1706 9147 1764 9173
rect 1806 9207 1864 9233
rect 1806 9173 1818 9207
rect 1852 9173 1864 9207
rect 1806 9147 1864 9173
rect 1906 9207 1964 9233
rect 1906 9173 1918 9207
rect 1952 9173 1964 9207
rect 1906 9147 1964 9173
rect 2006 9207 2064 9233
rect 2006 9173 2018 9207
rect 2052 9173 2064 9207
rect 2006 9147 2064 9173
rect 2106 9207 2164 9233
rect 2106 9173 2118 9207
rect 2152 9173 2164 9207
rect 2106 9147 2164 9173
rect 2206 9207 2264 9233
rect 2206 9173 2218 9207
rect 2252 9173 2264 9207
rect 2206 9147 2264 9173
rect 2306 9207 2364 9233
rect 2306 9173 2318 9207
rect 2352 9173 2364 9207
rect 2306 9147 2364 9173
rect 2406 9207 2464 9233
rect 2406 9173 2412 9207
rect 2452 9173 2464 9207
rect 2406 9147 2464 9173
rect 2506 9207 2564 9233
rect 2506 9173 2518 9207
rect 2558 9173 2564 9207
rect 2506 9147 2564 9173
rect 2606 9207 2664 9233
rect 2606 9173 2618 9207
rect 2652 9173 2664 9207
rect 2606 9147 2664 9173
rect 2706 9207 2764 9233
rect 2706 9173 2718 9207
rect 2752 9173 2764 9207
rect 2706 9147 2764 9173
rect 2806 9207 2864 9233
rect 2806 9173 2818 9207
rect 2852 9173 2864 9207
rect 2806 9147 2864 9173
rect 2906 9207 2964 9233
rect 2906 9173 2918 9207
rect 2952 9173 2964 9207
rect 2906 9147 2964 9173
rect 3006 9207 3064 9233
rect 3006 9173 3018 9207
rect 3052 9173 3064 9207
rect 3006 9147 3064 9173
rect 3106 9207 3164 9233
rect 3106 9173 3118 9207
rect 3152 9173 3164 9207
rect 3106 9147 3164 9173
rect 3206 9207 3264 9233
rect 3206 9173 3218 9207
rect 3252 9173 3264 9207
rect 3206 9147 3264 9173
rect 3306 9207 3364 9233
rect 3306 9173 3318 9207
rect 3352 9173 3364 9207
rect 3306 9147 3364 9173
rect 3406 9207 3464 9233
rect 3406 9173 3418 9207
rect 3452 9173 3464 9207
rect 3406 9147 3464 9173
rect 3506 9207 3564 9233
rect 3506 9173 3518 9207
rect 3552 9173 3564 9207
rect 3506 9147 3564 9173
rect 3606 9207 3664 9233
rect 3606 9173 3618 9207
rect 3652 9173 3664 9207
rect 3606 9147 3664 9173
rect 3706 9207 3764 9233
rect 3706 9173 3718 9207
rect 3752 9173 3764 9207
rect 3706 9147 3764 9173
rect 3806 9207 3864 9233
rect 3806 9173 3818 9207
rect 3852 9173 3864 9207
rect 3806 9147 3864 9173
rect 3906 9207 3964 9233
rect 3906 9173 3918 9207
rect 3952 9173 3964 9207
rect 3906 9147 3964 9173
rect 4006 9207 4064 9233
rect 4006 9173 4012 9207
rect 4052 9173 4064 9207
rect 4006 9147 4064 9173
rect 4106 9207 4164 9233
rect 4106 9173 4118 9207
rect 4158 9173 4164 9207
rect 4106 9147 4164 9173
rect 4206 9207 4264 9233
rect 4206 9173 4218 9207
rect 4252 9173 4264 9207
rect 4206 9147 4264 9173
rect 4306 9207 4364 9233
rect 4306 9173 4318 9207
rect 4352 9173 4364 9207
rect 4306 9147 4364 9173
rect 4406 9207 4464 9233
rect 4406 9173 4418 9207
rect 4452 9173 4464 9207
rect 4406 9147 4464 9173
rect 4506 9207 4564 9233
rect 4506 9173 4518 9207
rect 4552 9173 4564 9207
rect 4506 9147 4564 9173
rect 4606 9207 4664 9233
rect 4606 9173 4618 9207
rect 4652 9173 4664 9207
rect 4606 9147 4664 9173
rect 4706 9207 4764 9233
rect 4706 9173 4718 9207
rect 4752 9173 4764 9207
rect 4706 9147 4764 9173
rect 4806 9207 4864 9233
rect 4806 9173 4818 9207
rect 4852 9173 4864 9207
rect 4806 9147 4864 9173
rect 4906 9207 4964 9233
rect 4906 9173 4918 9207
rect 4952 9173 4964 9207
rect 4906 9147 4964 9173
rect 5006 9207 5064 9233
rect 5006 9173 5012 9207
rect 5052 9173 5064 9207
rect 5006 9147 5064 9173
rect 5106 9207 5164 9233
rect 5106 9173 5118 9207
rect 5158 9173 5164 9207
rect 5106 9147 5164 9173
rect 5206 9207 5264 9233
rect 5206 9173 5218 9207
rect 5252 9173 5264 9207
rect 5206 9147 5264 9173
rect 5306 9207 5364 9233
rect 5306 9173 5318 9207
rect 5352 9173 5364 9207
rect 5306 9147 5364 9173
rect 5406 9207 5464 9233
rect 5406 9173 5412 9207
rect 5452 9173 5464 9207
rect 5406 9147 5464 9173
rect 5506 9207 5564 9233
rect 5506 9173 5518 9207
rect 5558 9173 5564 9207
rect 5506 9147 5564 9173
rect 5606 9207 5664 9233
rect 5606 9173 5618 9207
rect 5652 9173 5664 9207
rect 5606 9147 5664 9173
rect 5706 9207 5764 9233
rect 5706 9173 5712 9207
rect 5752 9173 5764 9207
rect 5706 9147 5764 9173
rect 5806 9207 5864 9233
rect 5806 9173 5818 9207
rect 5858 9173 5864 9207
rect 5806 9147 5864 9173
rect 5906 9207 5964 9233
rect 5906 9173 5918 9207
rect 5952 9173 5964 9207
rect 5906 9147 5964 9173
rect 6006 9207 6064 9233
rect 6006 9173 6018 9207
rect 6052 9173 6064 9207
rect 6006 9147 6064 9173
rect 6106 9207 6164 9233
rect 6106 9173 6118 9207
rect 6152 9173 6164 9207
rect 6106 9147 6164 9173
rect 6206 9207 6264 9233
rect 6206 9173 6218 9207
rect 6252 9173 6264 9207
rect 6206 9147 6264 9173
rect 6306 9207 6364 9233
rect 6306 9173 6318 9207
rect 6352 9173 6364 9207
rect 6306 9147 6364 9173
rect 6406 9207 6464 9233
rect 6618 9226 6862 9260
rect 6406 9173 6418 9207
rect 6452 9173 6464 9207
rect 6508 9188 6516 9222
rect 6558 9188 6574 9222
rect 6618 9207 6652 9226
rect 6406 9147 6464 9173
rect 6828 9223 6862 9226
rect 6828 9207 6962 9223
rect 6618 9157 6652 9173
rect 6696 9158 6712 9192
rect 6754 9158 6762 9192
rect 6862 9173 6928 9207
rect 6828 9157 6962 9173
rect 7028 9207 7162 9223
rect 7062 9173 7128 9207
rect 7028 9157 7162 9173
rect 7228 9207 7262 9223
rect 7228 9157 7262 9173
rect 7328 9207 7462 9223
rect 7362 9173 7428 9207
rect 7328 9157 7462 9173
rect 6 9067 64 9093
rect 6 9033 18 9067
rect 52 9033 64 9067
rect 6 9007 64 9033
rect 106 9067 164 9093
rect 106 9033 118 9067
rect 152 9033 164 9067
rect 106 9007 164 9033
rect 206 9067 264 9093
rect 206 9033 218 9067
rect 252 9033 264 9067
rect 206 9007 264 9033
rect 306 9067 364 9093
rect 306 9033 318 9067
rect 352 9033 364 9067
rect 306 9007 364 9033
rect 406 9067 464 9093
rect 406 9033 418 9067
rect 452 9033 464 9067
rect 406 9007 464 9033
rect 506 9067 564 9093
rect 506 9033 518 9067
rect 552 9033 564 9067
rect 506 9007 564 9033
rect 606 9067 664 9093
rect 606 9033 612 9067
rect 652 9033 664 9067
rect 606 9007 664 9033
rect 706 9067 764 9093
rect 706 9033 718 9067
rect 758 9033 764 9067
rect 706 9007 764 9033
rect 806 9067 864 9093
rect 806 9033 818 9067
rect 852 9033 864 9067
rect 806 9007 864 9033
rect 906 9067 964 9093
rect 906 9033 918 9067
rect 952 9033 964 9067
rect 906 9007 964 9033
rect 1006 9067 1064 9093
rect 1006 9033 1018 9067
rect 1052 9033 1064 9067
rect 1006 9007 1064 9033
rect 1106 9067 1164 9093
rect 1106 9033 1118 9067
rect 1152 9033 1164 9067
rect 1106 9007 1164 9033
rect 1206 9067 1264 9093
rect 1206 9033 1218 9067
rect 1252 9033 1264 9067
rect 1206 9007 1264 9033
rect 1306 9067 1364 9093
rect 1306 9033 1318 9067
rect 1352 9033 1364 9067
rect 1306 9007 1364 9033
rect 1406 9067 1464 9093
rect 1406 9033 1418 9067
rect 1452 9033 1464 9067
rect 1406 9007 1464 9033
rect 1506 9067 1564 9093
rect 1506 9033 1518 9067
rect 1552 9033 1564 9067
rect 1506 9007 1564 9033
rect 1606 9067 1664 9093
rect 1606 9033 1618 9067
rect 1652 9033 1664 9067
rect 1606 9007 1664 9033
rect 1706 9067 1764 9093
rect 1706 9033 1712 9067
rect 1752 9033 1764 9067
rect 1706 9007 1764 9033
rect 1806 9067 1864 9093
rect 1806 9033 1818 9067
rect 1858 9033 1864 9067
rect 1806 9007 1864 9033
rect 1906 9067 1964 9093
rect 1906 9033 1912 9067
rect 1952 9033 1964 9067
rect 1906 9007 1964 9033
rect 2006 9067 2064 9093
rect 2006 9033 2018 9067
rect 2058 9033 2064 9067
rect 2006 9007 2064 9033
rect 2106 9067 2164 9093
rect 2106 9033 2118 9067
rect 2152 9033 2164 9067
rect 2106 9007 2164 9033
rect 2206 9067 2264 9093
rect 2206 9033 2218 9067
rect 2252 9033 2264 9067
rect 2206 9007 2264 9033
rect 2306 9067 2364 9093
rect 2306 9033 2318 9067
rect 2352 9033 2364 9067
rect 2306 9007 2364 9033
rect 2406 9067 2464 9093
rect 2406 9033 2418 9067
rect 2452 9033 2464 9067
rect 2406 9007 2464 9033
rect 2506 9067 2564 9093
rect 2506 9033 2518 9067
rect 2552 9033 2564 9067
rect 2506 9007 2564 9033
rect 2606 9067 2664 9093
rect 2606 9033 2612 9067
rect 2652 9033 2664 9067
rect 2606 9007 2664 9033
rect 2706 9067 2764 9093
rect 2706 9033 2718 9067
rect 2758 9033 2764 9067
rect 2706 9007 2764 9033
rect 2806 9067 2864 9093
rect 2806 9033 2812 9067
rect 2852 9033 2864 9067
rect 2806 9007 2864 9033
rect 2906 9067 2964 9093
rect 2906 9033 2918 9067
rect 2958 9033 2964 9067
rect 2906 9007 2964 9033
rect 3006 9067 3064 9093
rect 3006 9033 3018 9067
rect 3052 9033 3064 9067
rect 3006 9007 3064 9033
rect 3106 9067 3164 9093
rect 3106 9033 3118 9067
rect 3152 9033 3164 9067
rect 3106 9007 3164 9033
rect 3206 9067 3264 9093
rect 3206 9033 3212 9067
rect 3252 9033 3264 9067
rect 3206 9007 3264 9033
rect 3306 9067 3364 9093
rect 3306 9033 3318 9067
rect 3358 9033 3364 9067
rect 3306 9007 3364 9033
rect 3406 9067 3464 9093
rect 3406 9033 3418 9067
rect 3452 9033 3464 9067
rect 3406 9007 3464 9033
rect 3506 9067 3564 9093
rect 3506 9033 3518 9067
rect 3552 9033 3564 9067
rect 3506 9007 3564 9033
rect 3606 9067 3664 9093
rect 3606 9033 3618 9067
rect 3652 9033 3664 9067
rect 3606 9007 3664 9033
rect 3706 9067 3764 9093
rect 3706 9033 3718 9067
rect 3752 9033 3764 9067
rect 3706 9007 3764 9033
rect 3806 9067 3864 9093
rect 3806 9033 3818 9067
rect 3852 9033 3864 9067
rect 3806 9007 3864 9033
rect 3906 9067 3964 9093
rect 3906 9033 3918 9067
rect 3952 9033 3964 9067
rect 3906 9007 3964 9033
rect 4006 9067 4064 9093
rect 4006 9033 4018 9067
rect 4052 9033 4064 9067
rect 4006 9007 4064 9033
rect 4106 9067 4164 9093
rect 4106 9033 4118 9067
rect 4152 9033 4164 9067
rect 4106 9007 4164 9033
rect 4206 9067 4264 9093
rect 4206 9033 4218 9067
rect 4252 9033 4264 9067
rect 4206 9007 4264 9033
rect 4306 9067 4364 9093
rect 4306 9033 4318 9067
rect 4352 9033 4364 9067
rect 4306 9007 4364 9033
rect 4406 9067 4464 9093
rect 4406 9033 4418 9067
rect 4452 9033 4464 9067
rect 4406 9007 4464 9033
rect 4506 9067 4564 9093
rect 4506 9033 4512 9067
rect 4552 9033 4564 9067
rect 4506 9007 4564 9033
rect 4606 9067 4664 9093
rect 4606 9033 4618 9067
rect 4658 9033 4664 9067
rect 4606 9007 4664 9033
rect 4706 9067 4764 9093
rect 4706 9033 4712 9067
rect 4752 9033 4764 9067
rect 4706 9007 4764 9033
rect 4806 9067 4864 9093
rect 4806 9033 4818 9067
rect 4858 9033 4864 9067
rect 4806 9007 4864 9033
rect 4906 9067 4964 9093
rect 4906 9033 4918 9067
rect 4952 9033 4964 9067
rect 4906 9007 4964 9033
rect 5006 9067 5064 9093
rect 5006 9033 5018 9067
rect 5052 9033 5064 9067
rect 5006 9007 5064 9033
rect 5106 9067 5164 9093
rect 5106 9033 5118 9067
rect 5152 9033 5164 9067
rect 5106 9007 5164 9033
rect 5206 9067 5264 9093
rect 5206 9033 5212 9067
rect 5252 9033 5264 9067
rect 5206 9007 5264 9033
rect 5306 9067 5364 9093
rect 5306 9033 5318 9067
rect 5358 9033 5364 9067
rect 5306 9007 5364 9033
rect 5406 9067 5464 9093
rect 5406 9033 5418 9067
rect 5452 9033 5464 9067
rect 5406 9007 5464 9033
rect 5506 9067 5564 9093
rect 5506 9033 5518 9067
rect 5552 9033 5564 9067
rect 5506 9007 5564 9033
rect 5606 9067 5664 9093
rect 5606 9033 5618 9067
rect 5652 9033 5664 9067
rect 5606 9007 5664 9033
rect 5706 9067 5764 9093
rect 5706 9033 5718 9067
rect 5752 9033 5764 9067
rect 5706 9007 5764 9033
rect 5806 9067 5864 9093
rect 5806 9033 5818 9067
rect 5852 9033 5864 9067
rect 5806 9007 5864 9033
rect 5906 9067 5964 9093
rect 5906 9033 5918 9067
rect 5952 9033 5964 9067
rect 5906 9007 5964 9033
rect 6006 9067 6064 9093
rect 6006 9033 6018 9067
rect 6052 9033 6064 9067
rect 6006 9007 6064 9033
rect 6106 9067 6164 9093
rect 6106 9033 6118 9067
rect 6152 9033 6164 9067
rect 6106 9007 6164 9033
rect 6206 9067 6264 9093
rect 6206 9033 6218 9067
rect 6252 9033 6264 9067
rect 6206 9007 6264 9033
rect 6306 9067 6364 9093
rect 6306 9033 6318 9067
rect 6352 9033 6364 9067
rect 6306 9007 6364 9033
rect 6406 9067 6464 9093
rect 6618 9086 6862 9120
rect 6406 9033 6412 9067
rect 6452 9033 6464 9067
rect 6508 9048 6516 9082
rect 6558 9048 6574 9082
rect 6618 9067 6652 9086
rect 6406 9007 6464 9033
rect 6828 9067 6862 9086
rect 6618 9017 6652 9033
rect 6696 9018 6712 9052
rect 6754 9018 6762 9052
rect 6828 9017 6862 9033
rect 6928 9067 7162 9083
rect 6962 9033 7028 9067
rect 7062 9033 7128 9067
rect 6928 9017 7162 9033
rect 7228 9067 7262 9083
rect 7228 9017 7262 9033
rect 7328 9067 7462 9083
rect 7362 9033 7428 9067
rect 7328 9017 7462 9033
rect 6 8927 64 8953
rect 6 8893 18 8927
rect 52 8893 64 8927
rect 6 8867 64 8893
rect 106 8927 164 8953
rect 106 8893 118 8927
rect 152 8893 164 8927
rect 106 8867 164 8893
rect 206 8927 264 8953
rect 206 8893 218 8927
rect 252 8893 264 8927
rect 206 8867 264 8893
rect 306 8927 364 8953
rect 306 8893 318 8927
rect 352 8893 364 8927
rect 306 8867 364 8893
rect 406 8927 464 8953
rect 406 8893 418 8927
rect 452 8893 464 8927
rect 406 8867 464 8893
rect 506 8927 564 8953
rect 506 8893 518 8927
rect 552 8893 564 8927
rect 506 8867 564 8893
rect 606 8927 664 8953
rect 606 8893 618 8927
rect 652 8893 664 8927
rect 606 8867 664 8893
rect 706 8927 764 8953
rect 706 8893 718 8927
rect 752 8893 764 8927
rect 706 8867 764 8893
rect 806 8927 864 8953
rect 806 8893 818 8927
rect 852 8893 864 8927
rect 806 8867 864 8893
rect 906 8927 964 8953
rect 906 8893 918 8927
rect 952 8893 964 8927
rect 906 8867 964 8893
rect 1006 8927 1064 8953
rect 1006 8893 1018 8927
rect 1052 8893 1064 8927
rect 1006 8867 1064 8893
rect 1106 8927 1164 8953
rect 1106 8893 1118 8927
rect 1152 8893 1164 8927
rect 1106 8867 1164 8893
rect 1206 8927 1264 8953
rect 1206 8893 1218 8927
rect 1252 8893 1264 8927
rect 1206 8867 1264 8893
rect 1306 8927 1364 8953
rect 1306 8893 1318 8927
rect 1352 8893 1364 8927
rect 1306 8867 1364 8893
rect 1406 8927 1464 8953
rect 1406 8893 1418 8927
rect 1452 8893 1464 8927
rect 1406 8867 1464 8893
rect 1506 8927 1564 8953
rect 1506 8893 1518 8927
rect 1552 8893 1564 8927
rect 1506 8867 1564 8893
rect 1606 8927 1664 8953
rect 1606 8893 1618 8927
rect 1652 8893 1664 8927
rect 1606 8867 1664 8893
rect 1706 8927 1764 8953
rect 1706 8893 1718 8927
rect 1752 8893 1764 8927
rect 1706 8867 1764 8893
rect 1806 8927 1864 8953
rect 1806 8893 1818 8927
rect 1852 8893 1864 8927
rect 1806 8867 1864 8893
rect 1906 8927 1964 8953
rect 1906 8893 1918 8927
rect 1952 8893 1964 8927
rect 1906 8867 1964 8893
rect 2006 8927 2064 8953
rect 2006 8893 2018 8927
rect 2052 8893 2064 8927
rect 2006 8867 2064 8893
rect 2106 8927 2164 8953
rect 2106 8893 2118 8927
rect 2152 8893 2164 8927
rect 2106 8867 2164 8893
rect 2206 8927 2264 8953
rect 2206 8893 2218 8927
rect 2252 8893 2264 8927
rect 2206 8867 2264 8893
rect 2306 8927 2364 8953
rect 2306 8893 2318 8927
rect 2352 8893 2364 8927
rect 2306 8867 2364 8893
rect 2406 8927 2464 8953
rect 2406 8893 2418 8927
rect 2452 8893 2464 8927
rect 2406 8867 2464 8893
rect 2506 8927 2564 8953
rect 2506 8893 2518 8927
rect 2552 8893 2564 8927
rect 2506 8867 2564 8893
rect 2606 8927 2664 8953
rect 2606 8893 2612 8927
rect 2652 8893 2664 8927
rect 2606 8867 2664 8893
rect 2706 8927 2764 8953
rect 2706 8893 2718 8927
rect 2758 8893 2764 8927
rect 2706 8867 2764 8893
rect 2806 8927 2864 8953
rect 2806 8893 2818 8927
rect 2852 8893 2864 8927
rect 2806 8867 2864 8893
rect 2906 8927 2964 8953
rect 2906 8893 2918 8927
rect 2952 8893 2964 8927
rect 2906 8867 2964 8893
rect 3006 8927 3064 8953
rect 3006 8893 3018 8927
rect 3052 8893 3064 8927
rect 3006 8867 3064 8893
rect 3106 8927 3164 8953
rect 3106 8893 3118 8927
rect 3152 8893 3164 8927
rect 3106 8867 3164 8893
rect 3206 8927 3264 8953
rect 3206 8893 3218 8927
rect 3252 8893 3264 8927
rect 3206 8867 3264 8893
rect 3306 8927 3364 8953
rect 3306 8893 3318 8927
rect 3352 8893 3364 8927
rect 3306 8867 3364 8893
rect 3406 8927 3464 8953
rect 3406 8893 3418 8927
rect 3452 8893 3464 8927
rect 3406 8867 3464 8893
rect 3506 8927 3564 8953
rect 3506 8893 3518 8927
rect 3552 8893 3564 8927
rect 3506 8867 3564 8893
rect 3606 8927 3664 8953
rect 3606 8893 3618 8927
rect 3652 8893 3664 8927
rect 3606 8867 3664 8893
rect 3706 8927 3764 8953
rect 3706 8893 3718 8927
rect 3752 8893 3764 8927
rect 3706 8867 3764 8893
rect 3806 8927 3864 8953
rect 3806 8893 3818 8927
rect 3852 8893 3864 8927
rect 3806 8867 3864 8893
rect 3906 8927 3964 8953
rect 3906 8893 3918 8927
rect 3952 8893 3964 8927
rect 3906 8867 3964 8893
rect 4006 8927 4064 8953
rect 4006 8893 4018 8927
rect 4052 8893 4064 8927
rect 4006 8867 4064 8893
rect 4106 8927 4164 8953
rect 4106 8893 4118 8927
rect 4152 8893 4164 8927
rect 4106 8867 4164 8893
rect 4206 8927 4264 8953
rect 4206 8893 4218 8927
rect 4252 8893 4264 8927
rect 4206 8867 4264 8893
rect 4306 8927 4364 8953
rect 4306 8893 4318 8927
rect 4352 8893 4364 8927
rect 4306 8867 4364 8893
rect 4406 8927 4464 8953
rect 4406 8893 4412 8927
rect 4452 8893 4464 8927
rect 4406 8867 4464 8893
rect 4506 8927 4564 8953
rect 4506 8893 4518 8927
rect 4558 8893 4564 8927
rect 4506 8867 4564 8893
rect 4606 8927 4664 8953
rect 4606 8893 4612 8927
rect 4652 8893 4664 8927
rect 4606 8867 4664 8893
rect 4706 8927 4764 8953
rect 4706 8893 4718 8927
rect 4758 8893 4764 8927
rect 4706 8867 4764 8893
rect 4806 8927 4864 8953
rect 4806 8893 4812 8927
rect 4852 8893 4864 8927
rect 4806 8867 4864 8893
rect 4906 8927 4964 8953
rect 4906 8893 4918 8927
rect 4958 8893 4964 8927
rect 4906 8867 4964 8893
rect 5006 8927 5064 8953
rect 5006 8893 5018 8927
rect 5052 8893 5064 8927
rect 5006 8867 5064 8893
rect 5106 8927 5164 8953
rect 5106 8893 5118 8927
rect 5152 8893 5164 8927
rect 5106 8867 5164 8893
rect 5206 8927 5264 8953
rect 5206 8893 5218 8927
rect 5252 8893 5264 8927
rect 5206 8867 5264 8893
rect 5306 8927 5364 8953
rect 5306 8893 5318 8927
rect 5352 8893 5364 8927
rect 5306 8867 5364 8893
rect 5406 8927 5464 8953
rect 5406 8893 5418 8927
rect 5452 8893 5464 8927
rect 5406 8867 5464 8893
rect 5506 8927 5564 8953
rect 5506 8893 5518 8927
rect 5552 8893 5564 8927
rect 5506 8867 5564 8893
rect 5606 8927 5664 8953
rect 5606 8893 5612 8927
rect 5652 8893 5664 8927
rect 5606 8867 5664 8893
rect 5706 8927 5764 8953
rect 5706 8893 5718 8927
rect 5758 8893 5764 8927
rect 5706 8867 5764 8893
rect 5806 8927 5864 8953
rect 5806 8893 5818 8927
rect 5852 8893 5864 8927
rect 5806 8867 5864 8893
rect 5906 8927 5964 8953
rect 5906 8893 5918 8927
rect 5952 8893 5964 8927
rect 5906 8867 5964 8893
rect 6006 8927 6064 8953
rect 6006 8893 6018 8927
rect 6052 8893 6064 8927
rect 6006 8867 6064 8893
rect 6106 8927 6164 8953
rect 6106 8893 6112 8927
rect 6152 8893 6164 8927
rect 6106 8867 6164 8893
rect 6206 8927 6264 8953
rect 6206 8893 6218 8927
rect 6258 8893 6264 8927
rect 6206 8867 6264 8893
rect 6306 8927 6364 8953
rect 6306 8893 6318 8927
rect 6352 8893 6364 8927
rect 6306 8867 6364 8893
rect 6406 8927 6464 8953
rect 6618 8946 6862 8980
rect 6406 8893 6418 8927
rect 6452 8893 6464 8927
rect 6508 8908 6516 8942
rect 6558 8908 6574 8942
rect 6618 8927 6652 8946
rect 6406 8867 6464 8893
rect 6828 8943 6862 8946
rect 6828 8927 6962 8943
rect 6618 8877 6652 8893
rect 6696 8878 6712 8912
rect 6754 8878 6762 8912
rect 6862 8893 6928 8927
rect 6828 8877 6962 8893
rect 7028 8927 7062 8943
rect 7028 8877 7062 8893
rect 7128 8927 7262 8943
rect 7162 8893 7228 8927
rect 7128 8877 7262 8893
rect 7328 8927 7462 8943
rect 7362 8893 7428 8927
rect 7328 8877 7462 8893
rect 6 8787 64 8813
rect 6 8753 18 8787
rect 58 8753 64 8787
rect 6 8727 64 8753
rect 106 8787 164 8813
rect 106 8753 118 8787
rect 152 8753 164 8787
rect 106 8727 164 8753
rect 206 8787 264 8813
rect 206 8753 212 8787
rect 252 8753 264 8787
rect 206 8727 264 8753
rect 306 8787 364 8813
rect 306 8753 318 8787
rect 358 8753 364 8787
rect 306 8727 364 8753
rect 406 8787 464 8813
rect 406 8753 418 8787
rect 452 8753 464 8787
rect 406 8727 464 8753
rect 506 8787 564 8813
rect 506 8753 518 8787
rect 552 8753 564 8787
rect 506 8727 564 8753
rect 606 8787 664 8813
rect 606 8753 618 8787
rect 652 8753 664 8787
rect 606 8727 664 8753
rect 706 8787 764 8813
rect 706 8753 718 8787
rect 752 8753 764 8787
rect 706 8727 764 8753
rect 806 8787 864 8813
rect 806 8753 818 8787
rect 852 8753 864 8787
rect 806 8727 864 8753
rect 906 8787 964 8813
rect 906 8753 918 8787
rect 952 8753 964 8787
rect 906 8727 964 8753
rect 1006 8787 1064 8813
rect 1006 8753 1018 8787
rect 1052 8753 1064 8787
rect 1006 8727 1064 8753
rect 1106 8787 1164 8813
rect 1106 8753 1118 8787
rect 1152 8753 1164 8787
rect 1106 8727 1164 8753
rect 1206 8787 1264 8813
rect 1206 8753 1218 8787
rect 1252 8753 1264 8787
rect 1206 8727 1264 8753
rect 1306 8787 1364 8813
rect 1306 8753 1318 8787
rect 1352 8753 1364 8787
rect 1306 8727 1364 8753
rect 1406 8787 1464 8813
rect 1406 8753 1418 8787
rect 1452 8753 1464 8787
rect 1406 8727 1464 8753
rect 1506 8787 1564 8813
rect 1506 8753 1518 8787
rect 1552 8753 1564 8787
rect 1506 8727 1564 8753
rect 1606 8787 1664 8813
rect 1606 8753 1618 8787
rect 1652 8753 1664 8787
rect 1606 8727 1664 8753
rect 1706 8787 1764 8813
rect 1706 8753 1718 8787
rect 1752 8753 1764 8787
rect 1706 8727 1764 8753
rect 1806 8787 1864 8813
rect 1806 8753 1818 8787
rect 1852 8753 1864 8787
rect 1806 8727 1864 8753
rect 1906 8787 1964 8813
rect 1906 8753 1918 8787
rect 1952 8753 1964 8787
rect 1906 8727 1964 8753
rect 2006 8787 2064 8813
rect 2006 8753 2018 8787
rect 2052 8753 2064 8787
rect 2006 8727 2064 8753
rect 2106 8787 2164 8813
rect 2106 8753 2118 8787
rect 2152 8753 2164 8787
rect 2106 8727 2164 8753
rect 2206 8787 2264 8813
rect 2206 8753 2218 8787
rect 2252 8753 2264 8787
rect 2206 8727 2264 8753
rect 2306 8787 2364 8813
rect 2306 8753 2318 8787
rect 2352 8753 2364 8787
rect 2306 8727 2364 8753
rect 2406 8787 2464 8813
rect 2406 8753 2418 8787
rect 2452 8753 2464 8787
rect 2406 8727 2464 8753
rect 2506 8787 2564 8813
rect 2506 8753 2518 8787
rect 2552 8753 2564 8787
rect 2506 8727 2564 8753
rect 2606 8787 2664 8813
rect 2606 8753 2612 8787
rect 2652 8753 2664 8787
rect 2606 8727 2664 8753
rect 2706 8787 2764 8813
rect 2706 8753 2718 8787
rect 2758 8753 2764 8787
rect 2706 8727 2764 8753
rect 2806 8787 2864 8813
rect 2806 8753 2818 8787
rect 2852 8753 2864 8787
rect 2806 8727 2864 8753
rect 2906 8787 2964 8813
rect 2906 8753 2918 8787
rect 2952 8753 2964 8787
rect 2906 8727 2964 8753
rect 3006 8787 3064 8813
rect 3006 8753 3018 8787
rect 3052 8753 3064 8787
rect 3006 8727 3064 8753
rect 3106 8787 3164 8813
rect 3106 8753 3112 8787
rect 3152 8753 3164 8787
rect 3106 8727 3164 8753
rect 3206 8787 3264 8813
rect 3206 8753 3218 8787
rect 3258 8753 3264 8787
rect 3206 8727 3264 8753
rect 3306 8787 3364 8813
rect 3306 8753 3318 8787
rect 3352 8753 3364 8787
rect 3306 8727 3364 8753
rect 3406 8787 3464 8813
rect 3406 8753 3418 8787
rect 3452 8753 3464 8787
rect 3406 8727 3464 8753
rect 3506 8787 3564 8813
rect 3506 8753 3518 8787
rect 3552 8753 3564 8787
rect 3506 8727 3564 8753
rect 3606 8787 3664 8813
rect 3606 8753 3618 8787
rect 3652 8753 3664 8787
rect 3606 8727 3664 8753
rect 3706 8787 3764 8813
rect 3706 8753 3718 8787
rect 3752 8753 3764 8787
rect 3706 8727 3764 8753
rect 3806 8787 3864 8813
rect 3806 8753 3818 8787
rect 3852 8753 3864 8787
rect 3806 8727 3864 8753
rect 3906 8787 3964 8813
rect 3906 8753 3918 8787
rect 3952 8753 3964 8787
rect 3906 8727 3964 8753
rect 4006 8787 4064 8813
rect 4006 8753 4018 8787
rect 4052 8753 4064 8787
rect 4006 8727 4064 8753
rect 4106 8787 4164 8813
rect 4106 8753 4118 8787
rect 4152 8753 4164 8787
rect 4106 8727 4164 8753
rect 4206 8787 4264 8813
rect 4206 8753 4218 8787
rect 4252 8753 4264 8787
rect 4206 8727 4264 8753
rect 4306 8787 4364 8813
rect 4306 8753 4318 8787
rect 4352 8753 4364 8787
rect 4306 8727 4364 8753
rect 4406 8787 4464 8813
rect 4406 8753 4418 8787
rect 4452 8753 4464 8787
rect 4406 8727 4464 8753
rect 4506 8787 4564 8813
rect 4506 8753 4518 8787
rect 4552 8753 4564 8787
rect 4506 8727 4564 8753
rect 4606 8787 4664 8813
rect 4606 8753 4618 8787
rect 4652 8753 4664 8787
rect 4606 8727 4664 8753
rect 4706 8787 4764 8813
rect 4706 8753 4718 8787
rect 4752 8753 4764 8787
rect 4706 8727 4764 8753
rect 4806 8787 4864 8813
rect 4806 8753 4818 8787
rect 4852 8753 4864 8787
rect 4806 8727 4864 8753
rect 4906 8787 4964 8813
rect 4906 8753 4918 8787
rect 4952 8753 4964 8787
rect 4906 8727 4964 8753
rect 5006 8787 5064 8813
rect 5006 8753 5018 8787
rect 5052 8753 5064 8787
rect 5006 8727 5064 8753
rect 5106 8787 5164 8813
rect 5106 8753 5118 8787
rect 5152 8753 5164 8787
rect 5106 8727 5164 8753
rect 5206 8787 5264 8813
rect 5206 8753 5218 8787
rect 5252 8753 5264 8787
rect 5206 8727 5264 8753
rect 5306 8787 5364 8813
rect 5306 8753 5318 8787
rect 5352 8753 5364 8787
rect 5306 8727 5364 8753
rect 5406 8787 5464 8813
rect 5406 8753 5418 8787
rect 5452 8753 5464 8787
rect 5406 8727 5464 8753
rect 5506 8787 5564 8813
rect 5506 8753 5512 8787
rect 5552 8753 5564 8787
rect 5506 8727 5564 8753
rect 5606 8787 5664 8813
rect 5606 8753 5618 8787
rect 5658 8753 5664 8787
rect 5606 8727 5664 8753
rect 5706 8787 5764 8813
rect 5706 8753 5718 8787
rect 5752 8753 5764 8787
rect 5706 8727 5764 8753
rect 5806 8787 5864 8813
rect 5806 8753 5818 8787
rect 5852 8753 5864 8787
rect 5806 8727 5864 8753
rect 5906 8787 5964 8813
rect 5906 8753 5912 8787
rect 5952 8753 5964 8787
rect 5906 8727 5964 8753
rect 6006 8787 6064 8813
rect 6006 8753 6018 8787
rect 6058 8753 6064 8787
rect 6006 8727 6064 8753
rect 6106 8787 6164 8813
rect 6106 8753 6118 8787
rect 6152 8753 6164 8787
rect 6106 8727 6164 8753
rect 6206 8787 6264 8813
rect 6206 8753 6218 8787
rect 6252 8753 6264 8787
rect 6206 8727 6264 8753
rect 6306 8787 6364 8813
rect 6306 8753 6318 8787
rect 6352 8753 6364 8787
rect 6306 8727 6364 8753
rect 6406 8787 6464 8813
rect 6618 8806 6862 8840
rect 6406 8753 6418 8787
rect 6452 8753 6464 8787
rect 6508 8768 6516 8802
rect 6558 8768 6574 8802
rect 6618 8787 6652 8806
rect 6406 8727 6464 8753
rect 6828 8787 6862 8806
rect 6618 8737 6652 8753
rect 6696 8738 6712 8772
rect 6754 8738 6762 8772
rect 6828 8737 6862 8753
rect 6928 8787 7062 8803
rect 6962 8753 7028 8787
rect 6928 8737 7062 8753
rect 7128 8787 7262 8803
rect 7162 8753 7228 8787
rect 7128 8737 7262 8753
rect 7328 8787 7462 8803
rect 7362 8753 7428 8787
rect 7328 8737 7462 8753
rect 8 8630 18 8664
rect 52 8630 118 8664
rect 152 8630 168 8664
rect 208 8646 218 8680
rect 252 8646 318 8680
rect 352 8646 368 8680
rect 408 8630 418 8664
rect 452 8630 518 8664
rect 552 8630 568 8664
rect 608 8646 618 8680
rect 652 8646 718 8680
rect 752 8646 768 8680
rect 808 8630 818 8664
rect 852 8630 918 8664
rect 952 8630 968 8664
rect 1008 8646 1018 8680
rect 1052 8646 1118 8680
rect 1152 8646 1168 8680
rect 1208 8630 1218 8664
rect 1252 8630 1318 8664
rect 1352 8630 1368 8664
rect 1408 8646 1418 8680
rect 1452 8646 1518 8680
rect 1552 8646 1568 8680
rect 1608 8630 1618 8664
rect 1652 8630 1718 8664
rect 1752 8630 1768 8664
rect 1808 8646 1818 8680
rect 1852 8646 1918 8680
rect 1952 8646 1968 8680
rect 2008 8630 2018 8664
rect 2052 8630 2118 8664
rect 2152 8630 2168 8664
rect 2208 8646 2218 8680
rect 2252 8646 2318 8680
rect 2352 8646 2368 8680
rect 2408 8630 2418 8664
rect 2452 8630 2518 8664
rect 2552 8630 2568 8664
rect 2608 8646 2618 8680
rect 2652 8646 2718 8680
rect 2752 8646 2768 8680
rect 2808 8630 2818 8664
rect 2852 8630 2918 8664
rect 2952 8630 2968 8664
rect 3008 8646 3018 8680
rect 3052 8646 3118 8680
rect 3152 8646 3168 8680
rect 3208 8630 3218 8664
rect 3252 8630 3318 8664
rect 3352 8630 3368 8664
rect 3408 8646 3418 8680
rect 3452 8646 3518 8680
rect 3552 8646 3568 8680
rect 3608 8630 3618 8664
rect 3652 8630 3718 8664
rect 3752 8630 3768 8664
rect 3808 8646 3818 8680
rect 3852 8646 3918 8680
rect 3952 8646 3968 8680
rect 4008 8630 4018 8664
rect 4052 8630 4118 8664
rect 4152 8630 4168 8664
rect 4208 8646 4218 8680
rect 4252 8646 4318 8680
rect 4352 8646 4368 8680
rect 4408 8630 4418 8664
rect 4452 8630 4518 8664
rect 4552 8630 4568 8664
rect 4608 8646 4618 8680
rect 4652 8646 4718 8680
rect 4752 8646 4768 8680
rect 4808 8630 4818 8664
rect 4852 8630 4918 8664
rect 4952 8630 4968 8664
rect 5008 8646 5018 8680
rect 5052 8646 5118 8680
rect 5152 8646 5168 8680
rect 5208 8630 5218 8664
rect 5252 8630 5318 8664
rect 5352 8630 5368 8664
rect 5408 8646 5418 8680
rect 5452 8646 5518 8680
rect 5552 8646 5568 8680
rect 5608 8630 5618 8664
rect 5652 8630 5718 8664
rect 5752 8630 5768 8664
rect 5808 8646 5818 8680
rect 5852 8646 5918 8680
rect 5952 8646 5968 8680
rect 6008 8630 6018 8664
rect 6052 8630 6118 8664
rect 6152 8630 6168 8664
rect 6208 8646 6218 8680
rect 6252 8646 6318 8680
rect 6352 8646 6368 8680
rect 6516 8661 6568 8678
rect 6550 8644 6568 8661
rect 6602 8644 6618 8678
rect 6652 8644 6668 8678
rect 6702 8649 6720 8678
rect 6702 8644 6754 8649
rect 6862 8644 6878 8678
rect 6912 8644 6928 8678
rect 6962 8644 6978 8678
rect 7012 8644 7028 8678
rect 7062 8644 7078 8678
rect 7112 8644 7128 8678
rect 7162 8644 7178 8678
rect 7212 8644 7228 8678
rect 7262 8644 7278 8678
rect 7312 8644 7328 8678
rect 7362 8644 7378 8678
rect 7412 8644 7428 8678
rect 6 8557 64 8583
rect 6 8523 18 8557
rect 52 8523 64 8557
rect 6 8497 64 8523
rect 106 8557 164 8583
rect 106 8523 118 8557
rect 152 8523 164 8557
rect 106 8497 164 8523
rect 206 8557 264 8583
rect 206 8523 218 8557
rect 252 8523 264 8557
rect 206 8497 264 8523
rect 306 8557 364 8583
rect 306 8523 318 8557
rect 352 8523 364 8557
rect 306 8497 364 8523
rect 406 8557 464 8583
rect 406 8523 418 8557
rect 452 8523 464 8557
rect 406 8497 464 8523
rect 506 8557 564 8583
rect 506 8523 518 8557
rect 552 8523 564 8557
rect 506 8497 564 8523
rect 606 8557 664 8583
rect 606 8523 618 8557
rect 652 8523 664 8557
rect 606 8497 664 8523
rect 706 8557 764 8583
rect 706 8523 718 8557
rect 752 8523 764 8557
rect 706 8497 764 8523
rect 806 8557 864 8583
rect 806 8523 812 8557
rect 852 8523 864 8557
rect 806 8497 864 8523
rect 906 8557 964 8583
rect 906 8523 918 8557
rect 958 8523 964 8557
rect 906 8497 964 8523
rect 1006 8557 1064 8583
rect 1006 8523 1012 8557
rect 1052 8523 1064 8557
rect 1006 8497 1064 8523
rect 1106 8557 1164 8583
rect 1106 8523 1118 8557
rect 1158 8523 1164 8557
rect 1106 8497 1164 8523
rect 1206 8557 1264 8583
rect 1206 8523 1218 8557
rect 1252 8523 1264 8557
rect 1206 8497 1264 8523
rect 1306 8557 1364 8583
rect 1306 8523 1318 8557
rect 1352 8523 1364 8557
rect 1306 8497 1364 8523
rect 1406 8557 1464 8583
rect 1406 8523 1418 8557
rect 1452 8523 1464 8557
rect 1406 8497 1464 8523
rect 1506 8557 1564 8583
rect 1506 8523 1518 8557
rect 1552 8523 1564 8557
rect 1506 8497 1564 8523
rect 1606 8557 1664 8583
rect 1606 8523 1618 8557
rect 1652 8523 1664 8557
rect 1606 8497 1664 8523
rect 1706 8557 1764 8583
rect 1706 8523 1718 8557
rect 1752 8523 1764 8557
rect 1706 8497 1764 8523
rect 1806 8557 1864 8583
rect 1806 8523 1818 8557
rect 1852 8523 1864 8557
rect 1806 8497 1864 8523
rect 1906 8557 1964 8583
rect 1906 8523 1918 8557
rect 1952 8523 1964 8557
rect 1906 8497 1964 8523
rect 2006 8557 2064 8583
rect 2006 8523 2018 8557
rect 2052 8523 2064 8557
rect 2006 8497 2064 8523
rect 2106 8557 2164 8583
rect 2106 8523 2118 8557
rect 2152 8523 2164 8557
rect 2106 8497 2164 8523
rect 2206 8557 2264 8583
rect 2206 8523 2218 8557
rect 2252 8523 2264 8557
rect 2206 8497 2264 8523
rect 2306 8557 2364 8583
rect 2306 8523 2318 8557
rect 2352 8523 2364 8557
rect 2306 8497 2364 8523
rect 2406 8557 2464 8583
rect 2406 8523 2418 8557
rect 2452 8523 2464 8557
rect 2406 8497 2464 8523
rect 2506 8557 2564 8583
rect 2506 8523 2518 8557
rect 2552 8523 2564 8557
rect 2506 8497 2564 8523
rect 2606 8557 2664 8583
rect 2606 8523 2618 8557
rect 2652 8523 2664 8557
rect 2606 8497 2664 8523
rect 2706 8557 2764 8583
rect 2706 8523 2712 8557
rect 2752 8523 2764 8557
rect 2706 8497 2764 8523
rect 2806 8557 2864 8583
rect 2806 8523 2818 8557
rect 2858 8523 2864 8557
rect 2806 8497 2864 8523
rect 2906 8557 2964 8583
rect 2906 8523 2918 8557
rect 2952 8523 2964 8557
rect 2906 8497 2964 8523
rect 3006 8557 3064 8583
rect 3006 8523 3018 8557
rect 3052 8523 3064 8557
rect 3006 8497 3064 8523
rect 3106 8557 3164 8583
rect 3106 8523 3118 8557
rect 3152 8523 3164 8557
rect 3106 8497 3164 8523
rect 3206 8557 3264 8583
rect 3206 8523 3218 8557
rect 3252 8523 3264 8557
rect 3206 8497 3264 8523
rect 3306 8557 3364 8583
rect 3306 8523 3312 8557
rect 3352 8523 3364 8557
rect 3306 8497 3364 8523
rect 3406 8557 3464 8583
rect 3406 8523 3418 8557
rect 3458 8523 3464 8557
rect 3406 8497 3464 8523
rect 3506 8557 3564 8583
rect 3506 8523 3512 8557
rect 3552 8523 3564 8557
rect 3506 8497 3564 8523
rect 3606 8557 3664 8583
rect 3606 8523 3618 8557
rect 3658 8523 3664 8557
rect 3606 8497 3664 8523
rect 3706 8557 3764 8583
rect 3706 8523 3718 8557
rect 3752 8523 3764 8557
rect 3706 8497 3764 8523
rect 3806 8557 3864 8583
rect 3806 8523 3818 8557
rect 3852 8523 3864 8557
rect 3806 8497 3864 8523
rect 3906 8557 3964 8583
rect 3906 8523 3918 8557
rect 3952 8523 3964 8557
rect 3906 8497 3964 8523
rect 4006 8557 4064 8583
rect 4006 8523 4012 8557
rect 4052 8523 4064 8557
rect 4006 8497 4064 8523
rect 4106 8557 4164 8583
rect 4106 8523 4118 8557
rect 4158 8523 4164 8557
rect 4106 8497 4164 8523
rect 4206 8557 4264 8583
rect 4206 8523 4218 8557
rect 4252 8523 4264 8557
rect 4206 8497 4264 8523
rect 4306 8557 4364 8583
rect 4306 8523 4312 8557
rect 4352 8523 4364 8557
rect 4306 8497 4364 8523
rect 4406 8557 4464 8583
rect 4406 8523 4418 8557
rect 4458 8523 4464 8557
rect 4406 8497 4464 8523
rect 4506 8557 4564 8583
rect 4506 8523 4518 8557
rect 4552 8523 4564 8557
rect 4506 8497 4564 8523
rect 4606 8557 4664 8583
rect 4606 8523 4618 8557
rect 4652 8523 4664 8557
rect 4606 8497 4664 8523
rect 4706 8557 4764 8583
rect 4706 8523 4712 8557
rect 4752 8523 4764 8557
rect 4706 8497 4764 8523
rect 4806 8557 4864 8583
rect 4806 8523 4818 8557
rect 4858 8523 4864 8557
rect 4806 8497 4864 8523
rect 4906 8557 4964 8583
rect 4906 8523 4918 8557
rect 4952 8523 4964 8557
rect 4906 8497 4964 8523
rect 5006 8557 5064 8583
rect 5006 8523 5018 8557
rect 5052 8523 5064 8557
rect 5006 8497 5064 8523
rect 5106 8557 5164 8583
rect 5106 8523 5118 8557
rect 5152 8523 5164 8557
rect 5106 8497 5164 8523
rect 5206 8557 5264 8583
rect 5206 8523 5218 8557
rect 5252 8523 5264 8557
rect 5206 8497 5264 8523
rect 5306 8557 5364 8583
rect 5306 8523 5318 8557
rect 5352 8523 5364 8557
rect 5306 8497 5364 8523
rect 5406 8557 5464 8583
rect 5406 8523 5418 8557
rect 5452 8523 5464 8557
rect 5406 8497 5464 8523
rect 5506 8557 5564 8583
rect 5506 8523 5518 8557
rect 5552 8523 5564 8557
rect 5506 8497 5564 8523
rect 5606 8557 5664 8583
rect 5606 8523 5612 8557
rect 5652 8523 5664 8557
rect 5606 8497 5664 8523
rect 5706 8557 5764 8583
rect 5706 8523 5718 8557
rect 5758 8523 5764 8557
rect 5706 8497 5764 8523
rect 5806 8557 5864 8583
rect 5806 8523 5818 8557
rect 5852 8523 5864 8557
rect 5806 8497 5864 8523
rect 5906 8557 5964 8583
rect 5906 8523 5918 8557
rect 5952 8523 5964 8557
rect 5906 8497 5964 8523
rect 6006 8557 6064 8583
rect 6006 8523 6018 8557
rect 6052 8523 6064 8557
rect 6006 8497 6064 8523
rect 6106 8557 6164 8583
rect 6106 8523 6118 8557
rect 6152 8523 6164 8557
rect 6106 8497 6164 8523
rect 6206 8557 6264 8583
rect 6206 8523 6218 8557
rect 6252 8523 6264 8557
rect 6206 8497 6264 8523
rect 6306 8557 6364 8583
rect 6306 8523 6318 8557
rect 6352 8523 6364 8557
rect 6306 8497 6364 8523
rect 6406 8557 6464 8583
rect 6618 8576 6862 8610
rect 6406 8523 6418 8557
rect 6452 8523 6464 8557
rect 6508 8538 6516 8572
rect 6558 8538 6574 8572
rect 6618 8557 6652 8576
rect 6406 8497 6464 8523
rect 6828 8573 6862 8576
rect 6828 8557 6962 8573
rect 6618 8507 6652 8523
rect 6696 8508 6712 8542
rect 6754 8508 6762 8542
rect 6862 8523 6928 8557
rect 6828 8507 6962 8523
rect 7028 8557 7162 8573
rect 7062 8523 7128 8557
rect 7028 8507 7162 8523
rect 7228 8557 7362 8573
rect 7262 8523 7328 8557
rect 7228 8507 7362 8523
rect 7428 8557 7462 8573
rect 7428 8507 7462 8523
rect 6 8417 64 8443
rect 6 8383 18 8417
rect 58 8383 64 8417
rect 6 8357 64 8383
rect 106 8417 164 8443
rect 106 8383 118 8417
rect 152 8383 164 8417
rect 106 8357 164 8383
rect 206 8417 264 8443
rect 206 8383 218 8417
rect 252 8383 264 8417
rect 206 8357 264 8383
rect 306 8417 364 8443
rect 306 8383 318 8417
rect 352 8383 364 8417
rect 306 8357 364 8383
rect 406 8417 464 8443
rect 406 8383 418 8417
rect 452 8383 464 8417
rect 406 8357 464 8383
rect 506 8417 564 8443
rect 506 8383 518 8417
rect 552 8383 564 8417
rect 506 8357 564 8383
rect 606 8417 664 8443
rect 606 8383 618 8417
rect 652 8383 664 8417
rect 606 8357 664 8383
rect 706 8417 764 8443
rect 706 8383 718 8417
rect 752 8383 764 8417
rect 706 8357 764 8383
rect 806 8417 864 8443
rect 806 8383 818 8417
rect 852 8383 864 8417
rect 806 8357 864 8383
rect 906 8417 964 8443
rect 906 8383 918 8417
rect 952 8383 964 8417
rect 906 8357 964 8383
rect 1006 8417 1064 8443
rect 1006 8383 1018 8417
rect 1052 8383 1064 8417
rect 1006 8357 1064 8383
rect 1106 8417 1164 8443
rect 1106 8383 1118 8417
rect 1152 8383 1164 8417
rect 1106 8357 1164 8383
rect 1206 8417 1264 8443
rect 1206 8383 1218 8417
rect 1252 8383 1264 8417
rect 1206 8357 1264 8383
rect 1306 8417 1364 8443
rect 1306 8383 1312 8417
rect 1352 8383 1364 8417
rect 1306 8357 1364 8383
rect 1406 8417 1464 8443
rect 1406 8383 1418 8417
rect 1458 8383 1464 8417
rect 1406 8357 1464 8383
rect 1506 8417 1564 8443
rect 1506 8383 1518 8417
rect 1552 8383 1564 8417
rect 1506 8357 1564 8383
rect 1606 8417 1664 8443
rect 1606 8383 1618 8417
rect 1652 8383 1664 8417
rect 1606 8357 1664 8383
rect 1706 8417 1764 8443
rect 1706 8383 1718 8417
rect 1752 8383 1764 8417
rect 1706 8357 1764 8383
rect 1806 8417 1864 8443
rect 1806 8383 1812 8417
rect 1852 8383 1864 8417
rect 1806 8357 1864 8383
rect 1906 8417 1964 8443
rect 1906 8383 1918 8417
rect 1958 8383 1964 8417
rect 1906 8357 1964 8383
rect 2006 8417 2064 8443
rect 2006 8383 2012 8417
rect 2052 8383 2064 8417
rect 2006 8357 2064 8383
rect 2106 8417 2164 8443
rect 2106 8383 2118 8417
rect 2158 8383 2164 8417
rect 2106 8357 2164 8383
rect 2206 8417 2264 8443
rect 2206 8383 2218 8417
rect 2252 8383 2264 8417
rect 2206 8357 2264 8383
rect 2306 8417 2364 8443
rect 2306 8383 2312 8417
rect 2352 8383 2364 8417
rect 2306 8357 2364 8383
rect 2406 8417 2464 8443
rect 2406 8383 2418 8417
rect 2458 8383 2464 8417
rect 2406 8357 2464 8383
rect 2506 8417 2564 8443
rect 2506 8383 2518 8417
rect 2552 8383 2564 8417
rect 2506 8357 2564 8383
rect 2606 8417 2664 8443
rect 2606 8383 2618 8417
rect 2652 8383 2664 8417
rect 2606 8357 2664 8383
rect 2706 8417 2764 8443
rect 2706 8383 2718 8417
rect 2752 8383 2764 8417
rect 2706 8357 2764 8383
rect 2806 8417 2864 8443
rect 2806 8383 2818 8417
rect 2852 8383 2864 8417
rect 2806 8357 2864 8383
rect 2906 8417 2964 8443
rect 2906 8383 2918 8417
rect 2952 8383 2964 8417
rect 2906 8357 2964 8383
rect 3006 8417 3064 8443
rect 3006 8383 3018 8417
rect 3052 8383 3064 8417
rect 3006 8357 3064 8383
rect 3106 8417 3164 8443
rect 3106 8383 3118 8417
rect 3152 8383 3164 8417
rect 3106 8357 3164 8383
rect 3206 8417 3264 8443
rect 3206 8383 3218 8417
rect 3252 8383 3264 8417
rect 3206 8357 3264 8383
rect 3306 8417 3364 8443
rect 3306 8383 3318 8417
rect 3352 8383 3364 8417
rect 3306 8357 3364 8383
rect 3406 8417 3464 8443
rect 3406 8383 3418 8417
rect 3452 8383 3464 8417
rect 3406 8357 3464 8383
rect 3506 8417 3564 8443
rect 3506 8383 3518 8417
rect 3552 8383 3564 8417
rect 3506 8357 3564 8383
rect 3606 8417 3664 8443
rect 3606 8383 3618 8417
rect 3652 8383 3664 8417
rect 3606 8357 3664 8383
rect 3706 8417 3764 8443
rect 3706 8383 3718 8417
rect 3752 8383 3764 8417
rect 3706 8357 3764 8383
rect 3806 8417 3864 8443
rect 3806 8383 3812 8417
rect 3852 8383 3864 8417
rect 3806 8357 3864 8383
rect 3906 8417 3964 8443
rect 3906 8383 3918 8417
rect 3958 8383 3964 8417
rect 3906 8357 3964 8383
rect 4006 8417 4064 8443
rect 4006 8383 4018 8417
rect 4052 8383 4064 8417
rect 4006 8357 4064 8383
rect 4106 8417 4164 8443
rect 4106 8383 4118 8417
rect 4152 8383 4164 8417
rect 4106 8357 4164 8383
rect 4206 8417 4264 8443
rect 4206 8383 4218 8417
rect 4252 8383 4264 8417
rect 4206 8357 4264 8383
rect 4306 8417 4364 8443
rect 4306 8383 4318 8417
rect 4352 8383 4364 8417
rect 4306 8357 4364 8383
rect 4406 8417 4464 8443
rect 4406 8383 4418 8417
rect 4452 8383 4464 8417
rect 4406 8357 4464 8383
rect 4506 8417 4564 8443
rect 4506 8383 4518 8417
rect 4552 8383 4564 8417
rect 4506 8357 4564 8383
rect 4606 8417 4664 8443
rect 4606 8383 4618 8417
rect 4652 8383 4664 8417
rect 4606 8357 4664 8383
rect 4706 8417 4764 8443
rect 4706 8383 4712 8417
rect 4752 8383 4764 8417
rect 4706 8357 4764 8383
rect 4806 8417 4864 8443
rect 4806 8383 4818 8417
rect 4858 8383 4864 8417
rect 4806 8357 4864 8383
rect 4906 8417 4964 8443
rect 4906 8383 4912 8417
rect 4952 8383 4964 8417
rect 4906 8357 4964 8383
rect 5006 8417 5064 8443
rect 5006 8383 5018 8417
rect 5058 8383 5064 8417
rect 5006 8357 5064 8383
rect 5106 8417 5164 8443
rect 5106 8383 5118 8417
rect 5152 8383 5164 8417
rect 5106 8357 5164 8383
rect 5206 8417 5264 8443
rect 5206 8383 5218 8417
rect 5252 8383 5264 8417
rect 5206 8357 5264 8383
rect 5306 8417 5364 8443
rect 5306 8383 5318 8417
rect 5352 8383 5364 8417
rect 5306 8357 5364 8383
rect 5406 8417 5464 8443
rect 5406 8383 5418 8417
rect 5452 8383 5464 8417
rect 5406 8357 5464 8383
rect 5506 8417 5564 8443
rect 5506 8383 5518 8417
rect 5552 8383 5564 8417
rect 5506 8357 5564 8383
rect 5606 8417 5664 8443
rect 5606 8383 5618 8417
rect 5652 8383 5664 8417
rect 5606 8357 5664 8383
rect 5706 8417 5764 8443
rect 5706 8383 5718 8417
rect 5752 8383 5764 8417
rect 5706 8357 5764 8383
rect 5806 8417 5864 8443
rect 5806 8383 5812 8417
rect 5852 8383 5864 8417
rect 5806 8357 5864 8383
rect 5906 8417 5964 8443
rect 5906 8383 5918 8417
rect 5958 8383 5964 8417
rect 5906 8357 5964 8383
rect 6006 8417 6064 8443
rect 6006 8383 6018 8417
rect 6052 8383 6064 8417
rect 6006 8357 6064 8383
rect 6106 8417 6164 8443
rect 6106 8383 6118 8417
rect 6152 8383 6164 8417
rect 6106 8357 6164 8383
rect 6206 8417 6264 8443
rect 6206 8383 6218 8417
rect 6252 8383 6264 8417
rect 6206 8357 6264 8383
rect 6306 8417 6364 8443
rect 6306 8383 6318 8417
rect 6352 8383 6364 8417
rect 6306 8357 6364 8383
rect 6406 8417 6464 8443
rect 6618 8436 6862 8470
rect 6406 8383 6412 8417
rect 6452 8383 6464 8417
rect 6508 8398 6516 8432
rect 6558 8398 6574 8432
rect 6618 8417 6652 8436
rect 6406 8357 6464 8383
rect 6828 8417 6862 8436
rect 6618 8367 6652 8383
rect 6696 8368 6712 8402
rect 6754 8368 6762 8402
rect 6828 8367 6862 8383
rect 6928 8417 7162 8433
rect 6962 8383 7028 8417
rect 7062 8383 7128 8417
rect 6928 8367 7162 8383
rect 7228 8417 7362 8433
rect 7262 8383 7328 8417
rect 7228 8367 7362 8383
rect 7428 8417 7462 8433
rect 7428 8367 7462 8383
rect 6 8277 64 8303
rect 6 8243 18 8277
rect 52 8243 64 8277
rect 6 8217 64 8243
rect 106 8277 164 8303
rect 106 8243 118 8277
rect 152 8243 164 8277
rect 106 8217 164 8243
rect 206 8277 264 8303
rect 206 8243 218 8277
rect 252 8243 264 8277
rect 206 8217 264 8243
rect 306 8277 364 8303
rect 306 8243 318 8277
rect 352 8243 364 8277
rect 306 8217 364 8243
rect 406 8277 464 8303
rect 406 8243 418 8277
rect 452 8243 464 8277
rect 406 8217 464 8243
rect 506 8277 564 8303
rect 506 8243 518 8277
rect 552 8243 564 8277
rect 506 8217 564 8243
rect 606 8277 664 8303
rect 606 8243 612 8277
rect 652 8243 664 8277
rect 606 8217 664 8243
rect 706 8277 764 8303
rect 706 8243 718 8277
rect 758 8243 764 8277
rect 706 8217 764 8243
rect 806 8277 864 8303
rect 806 8243 812 8277
rect 852 8243 864 8277
rect 806 8217 864 8243
rect 906 8277 964 8303
rect 906 8243 918 8277
rect 958 8243 964 8277
rect 906 8217 964 8243
rect 1006 8277 1064 8303
rect 1006 8243 1018 8277
rect 1052 8243 1064 8277
rect 1006 8217 1064 8243
rect 1106 8277 1164 8303
rect 1106 8243 1118 8277
rect 1152 8243 1164 8277
rect 1106 8217 1164 8243
rect 1206 8277 1264 8303
rect 1206 8243 1218 8277
rect 1252 8243 1264 8277
rect 1206 8217 1264 8243
rect 1306 8277 1364 8303
rect 1306 8243 1318 8277
rect 1352 8243 1364 8277
rect 1306 8217 1364 8243
rect 1406 8277 1464 8303
rect 1406 8243 1418 8277
rect 1452 8243 1464 8277
rect 1406 8217 1464 8243
rect 1506 8277 1564 8303
rect 1506 8243 1518 8277
rect 1552 8243 1564 8277
rect 1506 8217 1564 8243
rect 1606 8277 1664 8303
rect 1606 8243 1618 8277
rect 1652 8243 1664 8277
rect 1606 8217 1664 8243
rect 1706 8277 1764 8303
rect 1706 8243 1718 8277
rect 1752 8243 1764 8277
rect 1706 8217 1764 8243
rect 1806 8277 1864 8303
rect 1806 8243 1818 8277
rect 1852 8243 1864 8277
rect 1806 8217 1864 8243
rect 1906 8277 1964 8303
rect 1906 8243 1912 8277
rect 1952 8243 1964 8277
rect 1906 8217 1964 8243
rect 2006 8277 2064 8303
rect 2006 8243 2018 8277
rect 2058 8243 2064 8277
rect 2006 8217 2064 8243
rect 2106 8277 2164 8303
rect 2106 8243 2118 8277
rect 2152 8243 2164 8277
rect 2106 8217 2164 8243
rect 2206 8277 2264 8303
rect 2206 8243 2218 8277
rect 2252 8243 2264 8277
rect 2206 8217 2264 8243
rect 2306 8277 2364 8303
rect 2306 8243 2312 8277
rect 2352 8243 2364 8277
rect 2306 8217 2364 8243
rect 2406 8277 2464 8303
rect 2406 8243 2418 8277
rect 2458 8243 2464 8277
rect 2406 8217 2464 8243
rect 2506 8277 2564 8303
rect 2506 8243 2512 8277
rect 2552 8243 2564 8277
rect 2506 8217 2564 8243
rect 2606 8277 2664 8303
rect 2606 8243 2618 8277
rect 2658 8243 2664 8277
rect 2606 8217 2664 8243
rect 2706 8277 2764 8303
rect 2706 8243 2718 8277
rect 2752 8243 2764 8277
rect 2706 8217 2764 8243
rect 2806 8277 2864 8303
rect 2806 8243 2818 8277
rect 2852 8243 2864 8277
rect 2806 8217 2864 8243
rect 2906 8277 2964 8303
rect 2906 8243 2918 8277
rect 2952 8243 2964 8277
rect 2906 8217 2964 8243
rect 3006 8277 3064 8303
rect 3006 8243 3018 8277
rect 3052 8243 3064 8277
rect 3006 8217 3064 8243
rect 3106 8277 3164 8303
rect 3106 8243 3112 8277
rect 3152 8243 3164 8277
rect 3106 8217 3164 8243
rect 3206 8277 3264 8303
rect 3206 8243 3218 8277
rect 3258 8243 3264 8277
rect 3206 8217 3264 8243
rect 3306 8277 3364 8303
rect 3306 8243 3318 8277
rect 3352 8243 3364 8277
rect 3306 8217 3364 8243
rect 3406 8277 3464 8303
rect 3406 8243 3418 8277
rect 3452 8243 3464 8277
rect 3406 8217 3464 8243
rect 3506 8277 3564 8303
rect 3506 8243 3512 8277
rect 3552 8243 3564 8277
rect 3506 8217 3564 8243
rect 3606 8277 3664 8303
rect 3606 8243 3618 8277
rect 3658 8243 3664 8277
rect 3606 8217 3664 8243
rect 3706 8277 3764 8303
rect 3706 8243 3718 8277
rect 3752 8243 3764 8277
rect 3706 8217 3764 8243
rect 3806 8277 3864 8303
rect 3806 8243 3818 8277
rect 3852 8243 3864 8277
rect 3806 8217 3864 8243
rect 3906 8277 3964 8303
rect 3906 8243 3918 8277
rect 3952 8243 3964 8277
rect 3906 8217 3964 8243
rect 4006 8277 4064 8303
rect 4006 8243 4018 8277
rect 4052 8243 4064 8277
rect 4006 8217 4064 8243
rect 4106 8277 4164 8303
rect 4106 8243 4118 8277
rect 4152 8243 4164 8277
rect 4106 8217 4164 8243
rect 4206 8277 4264 8303
rect 4206 8243 4218 8277
rect 4252 8243 4264 8277
rect 4206 8217 4264 8243
rect 4306 8277 4364 8303
rect 4306 8243 4318 8277
rect 4352 8243 4364 8277
rect 4306 8217 4364 8243
rect 4406 8277 4464 8303
rect 4406 8243 4418 8277
rect 4452 8243 4464 8277
rect 4406 8217 4464 8243
rect 4506 8277 4564 8303
rect 4506 8243 4518 8277
rect 4552 8243 4564 8277
rect 4506 8217 4564 8243
rect 4606 8277 4664 8303
rect 4606 8243 4618 8277
rect 4652 8243 4664 8277
rect 4606 8217 4664 8243
rect 4706 8277 4764 8303
rect 4706 8243 4718 8277
rect 4752 8243 4764 8277
rect 4706 8217 4764 8243
rect 4806 8277 4864 8303
rect 4806 8243 4818 8277
rect 4852 8243 4864 8277
rect 4806 8217 4864 8243
rect 4906 8277 4964 8303
rect 4906 8243 4918 8277
rect 4952 8243 4964 8277
rect 4906 8217 4964 8243
rect 5006 8277 5064 8303
rect 5006 8243 5018 8277
rect 5052 8243 5064 8277
rect 5006 8217 5064 8243
rect 5106 8277 5164 8303
rect 5106 8243 5118 8277
rect 5152 8243 5164 8277
rect 5106 8217 5164 8243
rect 5206 8277 5264 8303
rect 5206 8243 5218 8277
rect 5252 8243 5264 8277
rect 5206 8217 5264 8243
rect 5306 8277 5364 8303
rect 5306 8243 5318 8277
rect 5352 8243 5364 8277
rect 5306 8217 5364 8243
rect 5406 8277 5464 8303
rect 5406 8243 5418 8277
rect 5452 8243 5464 8277
rect 5406 8217 5464 8243
rect 5506 8277 5564 8303
rect 5506 8243 5518 8277
rect 5552 8243 5564 8277
rect 5506 8217 5564 8243
rect 5606 8277 5664 8303
rect 5606 8243 5618 8277
rect 5652 8243 5664 8277
rect 5606 8217 5664 8243
rect 5706 8277 5764 8303
rect 5706 8243 5718 8277
rect 5752 8243 5764 8277
rect 5706 8217 5764 8243
rect 5806 8277 5864 8303
rect 5806 8243 5818 8277
rect 5852 8243 5864 8277
rect 5806 8217 5864 8243
rect 5906 8277 5964 8303
rect 5906 8243 5918 8277
rect 5952 8243 5964 8277
rect 5906 8217 5964 8243
rect 6006 8277 6064 8303
rect 6006 8243 6018 8277
rect 6052 8243 6064 8277
rect 6006 8217 6064 8243
rect 6106 8277 6164 8303
rect 6106 8243 6118 8277
rect 6152 8243 6164 8277
rect 6106 8217 6164 8243
rect 6206 8277 6264 8303
rect 6206 8243 6218 8277
rect 6252 8243 6264 8277
rect 6206 8217 6264 8243
rect 6306 8277 6364 8303
rect 6306 8243 6318 8277
rect 6352 8243 6364 8277
rect 6306 8217 6364 8243
rect 6406 8277 6464 8303
rect 6618 8296 6862 8330
rect 6406 8243 6412 8277
rect 6452 8243 6464 8277
rect 6508 8258 6516 8292
rect 6558 8258 6574 8292
rect 6618 8277 6652 8296
rect 6406 8217 6464 8243
rect 6828 8293 6862 8296
rect 6828 8277 6962 8293
rect 6618 8227 6652 8243
rect 6696 8228 6712 8262
rect 6754 8228 6762 8262
rect 6862 8243 6928 8277
rect 6828 8227 6962 8243
rect 7028 8277 7062 8293
rect 7028 8227 7062 8243
rect 7128 8277 7362 8293
rect 7162 8243 7228 8277
rect 7262 8243 7328 8277
rect 7128 8227 7362 8243
rect 7428 8277 7462 8293
rect 7428 8227 7462 8243
rect 6 8137 64 8163
rect 6 8103 18 8137
rect 52 8103 64 8137
rect 6 8077 64 8103
rect 106 8137 164 8163
rect 106 8103 118 8137
rect 152 8103 164 8137
rect 106 8077 164 8103
rect 206 8137 264 8163
rect 206 8103 218 8137
rect 252 8103 264 8137
rect 206 8077 264 8103
rect 306 8137 364 8163
rect 306 8103 318 8137
rect 352 8103 364 8137
rect 306 8077 364 8103
rect 406 8137 464 8163
rect 406 8103 418 8137
rect 452 8103 464 8137
rect 406 8077 464 8103
rect 506 8137 564 8163
rect 506 8103 518 8137
rect 552 8103 564 8137
rect 506 8077 564 8103
rect 606 8137 664 8163
rect 606 8103 618 8137
rect 652 8103 664 8137
rect 606 8077 664 8103
rect 706 8137 764 8163
rect 706 8103 718 8137
rect 752 8103 764 8137
rect 706 8077 764 8103
rect 806 8137 864 8163
rect 806 8103 818 8137
rect 852 8103 864 8137
rect 806 8077 864 8103
rect 906 8137 964 8163
rect 906 8103 918 8137
rect 952 8103 964 8137
rect 906 8077 964 8103
rect 1006 8137 1064 8163
rect 1006 8103 1018 8137
rect 1052 8103 1064 8137
rect 1006 8077 1064 8103
rect 1106 8137 1164 8163
rect 1106 8103 1118 8137
rect 1152 8103 1164 8137
rect 1106 8077 1164 8103
rect 1206 8137 1264 8163
rect 1206 8103 1212 8137
rect 1252 8103 1264 8137
rect 1206 8077 1264 8103
rect 1306 8137 1364 8163
rect 1306 8103 1318 8137
rect 1358 8103 1364 8137
rect 1306 8077 1364 8103
rect 1406 8137 1464 8163
rect 1406 8103 1418 8137
rect 1452 8103 1464 8137
rect 1406 8077 1464 8103
rect 1506 8137 1564 8163
rect 1506 8103 1518 8137
rect 1552 8103 1564 8137
rect 1506 8077 1564 8103
rect 1606 8137 1664 8163
rect 1606 8103 1618 8137
rect 1652 8103 1664 8137
rect 1606 8077 1664 8103
rect 1706 8137 1764 8163
rect 1706 8103 1718 8137
rect 1752 8103 1764 8137
rect 1706 8077 1764 8103
rect 1806 8137 1864 8163
rect 1806 8103 1818 8137
rect 1852 8103 1864 8137
rect 1806 8077 1864 8103
rect 1906 8137 1964 8163
rect 1906 8103 1918 8137
rect 1952 8103 1964 8137
rect 1906 8077 1964 8103
rect 2006 8137 2064 8163
rect 2006 8103 2018 8137
rect 2052 8103 2064 8137
rect 2006 8077 2064 8103
rect 2106 8137 2164 8163
rect 2106 8103 2118 8137
rect 2152 8103 2164 8137
rect 2106 8077 2164 8103
rect 2206 8137 2264 8163
rect 2206 8103 2218 8137
rect 2252 8103 2264 8137
rect 2206 8077 2264 8103
rect 2306 8137 2364 8163
rect 2306 8103 2318 8137
rect 2352 8103 2364 8137
rect 2306 8077 2364 8103
rect 2406 8137 2464 8163
rect 2406 8103 2418 8137
rect 2452 8103 2464 8137
rect 2406 8077 2464 8103
rect 2506 8137 2564 8163
rect 2506 8103 2518 8137
rect 2552 8103 2564 8137
rect 2506 8077 2564 8103
rect 2606 8137 2664 8163
rect 2606 8103 2612 8137
rect 2652 8103 2664 8137
rect 2606 8077 2664 8103
rect 2706 8137 2764 8163
rect 2706 8103 2718 8137
rect 2758 8103 2764 8137
rect 2706 8077 2764 8103
rect 2806 8137 2864 8163
rect 2806 8103 2812 8137
rect 2852 8103 2864 8137
rect 2806 8077 2864 8103
rect 2906 8137 2964 8163
rect 2906 8103 2918 8137
rect 2958 8103 2964 8137
rect 2906 8077 2964 8103
rect 3006 8137 3064 8163
rect 3006 8103 3018 8137
rect 3052 8103 3064 8137
rect 3006 8077 3064 8103
rect 3106 8137 3164 8163
rect 3106 8103 3118 8137
rect 3152 8103 3164 8137
rect 3106 8077 3164 8103
rect 3206 8137 3264 8163
rect 3206 8103 3218 8137
rect 3252 8103 3264 8137
rect 3206 8077 3264 8103
rect 3306 8137 3364 8163
rect 3306 8103 3318 8137
rect 3352 8103 3364 8137
rect 3306 8077 3364 8103
rect 3406 8137 3464 8163
rect 3406 8103 3418 8137
rect 3452 8103 3464 8137
rect 3406 8077 3464 8103
rect 3506 8137 3564 8163
rect 3506 8103 3518 8137
rect 3552 8103 3564 8137
rect 3506 8077 3564 8103
rect 3606 8137 3664 8163
rect 3606 8103 3618 8137
rect 3652 8103 3664 8137
rect 3606 8077 3664 8103
rect 3706 8137 3764 8163
rect 3706 8103 3712 8137
rect 3752 8103 3764 8137
rect 3706 8077 3764 8103
rect 3806 8137 3864 8163
rect 3806 8103 3818 8137
rect 3858 8103 3864 8137
rect 3806 8077 3864 8103
rect 3906 8137 3964 8163
rect 3906 8103 3918 8137
rect 3952 8103 3964 8137
rect 3906 8077 3964 8103
rect 4006 8137 4064 8163
rect 4006 8103 4018 8137
rect 4052 8103 4064 8137
rect 4006 8077 4064 8103
rect 4106 8137 4164 8163
rect 4106 8103 4118 8137
rect 4152 8103 4164 8137
rect 4106 8077 4164 8103
rect 4206 8137 4264 8163
rect 4206 8103 4218 8137
rect 4252 8103 4264 8137
rect 4206 8077 4264 8103
rect 4306 8137 4364 8163
rect 4306 8103 4318 8137
rect 4352 8103 4364 8137
rect 4306 8077 4364 8103
rect 4406 8137 4464 8163
rect 4406 8103 4418 8137
rect 4452 8103 4464 8137
rect 4406 8077 4464 8103
rect 4506 8137 4564 8163
rect 4506 8103 4518 8137
rect 4552 8103 4564 8137
rect 4506 8077 4564 8103
rect 4606 8137 4664 8163
rect 4606 8103 4618 8137
rect 4652 8103 4664 8137
rect 4606 8077 4664 8103
rect 4706 8137 4764 8163
rect 4706 8103 4718 8137
rect 4752 8103 4764 8137
rect 4706 8077 4764 8103
rect 4806 8137 4864 8163
rect 4806 8103 4818 8137
rect 4852 8103 4864 8137
rect 4806 8077 4864 8103
rect 4906 8137 4964 8163
rect 4906 8103 4918 8137
rect 4952 8103 4964 8137
rect 4906 8077 4964 8103
rect 5006 8137 5064 8163
rect 5006 8103 5018 8137
rect 5052 8103 5064 8137
rect 5006 8077 5064 8103
rect 5106 8137 5164 8163
rect 5106 8103 5118 8137
rect 5152 8103 5164 8137
rect 5106 8077 5164 8103
rect 5206 8137 5264 8163
rect 5206 8103 5218 8137
rect 5252 8103 5264 8137
rect 5206 8077 5264 8103
rect 5306 8137 5364 8163
rect 5306 8103 5318 8137
rect 5352 8103 5364 8137
rect 5306 8077 5364 8103
rect 5406 8137 5464 8163
rect 5406 8103 5418 8137
rect 5452 8103 5464 8137
rect 5406 8077 5464 8103
rect 5506 8137 5564 8163
rect 5506 8103 5518 8137
rect 5552 8103 5564 8137
rect 5506 8077 5564 8103
rect 5606 8137 5664 8163
rect 5606 8103 5618 8137
rect 5652 8103 5664 8137
rect 5606 8077 5664 8103
rect 5706 8137 5764 8163
rect 5706 8103 5718 8137
rect 5752 8103 5764 8137
rect 5706 8077 5764 8103
rect 5806 8137 5864 8163
rect 5806 8103 5818 8137
rect 5852 8103 5864 8137
rect 5806 8077 5864 8103
rect 5906 8137 5964 8163
rect 5906 8103 5918 8137
rect 5952 8103 5964 8137
rect 5906 8077 5964 8103
rect 6006 8137 6064 8163
rect 6006 8103 6018 8137
rect 6052 8103 6064 8137
rect 6006 8077 6064 8103
rect 6106 8137 6164 8163
rect 6106 8103 6118 8137
rect 6152 8103 6164 8137
rect 6106 8077 6164 8103
rect 6206 8137 6264 8163
rect 6206 8103 6218 8137
rect 6252 8103 6264 8137
rect 6206 8077 6264 8103
rect 6306 8137 6364 8163
rect 6306 8103 6318 8137
rect 6352 8103 6364 8137
rect 6306 8077 6364 8103
rect 6406 8137 6464 8163
rect 6618 8156 6862 8190
rect 6406 8103 6418 8137
rect 6452 8103 6464 8137
rect 6508 8118 6516 8152
rect 6558 8118 6574 8152
rect 6618 8137 6652 8156
rect 6406 8077 6464 8103
rect 6828 8137 6862 8156
rect 6618 8087 6652 8103
rect 6696 8088 6712 8122
rect 6754 8088 6762 8122
rect 6828 8087 6862 8103
rect 6928 8137 7062 8153
rect 6962 8103 7028 8137
rect 6928 8087 7062 8103
rect 7128 8137 7362 8153
rect 7162 8103 7228 8137
rect 7262 8103 7328 8137
rect 7128 8087 7362 8103
rect 7428 8137 7462 8153
rect 7428 8087 7462 8103
rect 6 7997 64 8023
rect 6 7963 18 7997
rect 52 7963 64 7997
rect 6 7937 64 7963
rect 106 7997 164 8023
rect 106 7963 118 7997
rect 152 7963 164 7997
rect 106 7937 164 7963
rect 206 7997 264 8023
rect 206 7963 212 7997
rect 252 7963 264 7997
rect 206 7937 264 7963
rect 306 7997 364 8023
rect 306 7963 318 7997
rect 358 7963 364 7997
rect 306 7937 364 7963
rect 406 7997 464 8023
rect 406 7963 418 7997
rect 452 7963 464 7997
rect 406 7937 464 7963
rect 506 7997 564 8023
rect 506 7963 518 7997
rect 552 7963 564 7997
rect 506 7937 564 7963
rect 606 7997 664 8023
rect 606 7963 618 7997
rect 652 7963 664 7997
rect 606 7937 664 7963
rect 706 7997 764 8023
rect 706 7963 718 7997
rect 752 7963 764 7997
rect 706 7937 764 7963
rect 806 7997 864 8023
rect 806 7963 818 7997
rect 852 7963 864 7997
rect 806 7937 864 7963
rect 906 7997 964 8023
rect 906 7963 918 7997
rect 952 7963 964 7997
rect 906 7937 964 7963
rect 1006 7997 1064 8023
rect 1006 7963 1012 7997
rect 1052 7963 1064 7997
rect 1006 7937 1064 7963
rect 1106 7997 1164 8023
rect 1106 7963 1118 7997
rect 1158 7963 1164 7997
rect 1106 7937 1164 7963
rect 1206 7997 1264 8023
rect 1206 7963 1218 7997
rect 1252 7963 1264 7997
rect 1206 7937 1264 7963
rect 1306 7997 1364 8023
rect 1306 7963 1312 7997
rect 1352 7963 1364 7997
rect 1306 7937 1364 7963
rect 1406 7997 1464 8023
rect 1406 7963 1418 7997
rect 1458 7963 1464 7997
rect 1406 7937 1464 7963
rect 1506 7997 1564 8023
rect 1506 7963 1518 7997
rect 1552 7963 1564 7997
rect 1506 7937 1564 7963
rect 1606 7997 1664 8023
rect 1606 7963 1618 7997
rect 1652 7963 1664 7997
rect 1606 7937 1664 7963
rect 1706 7997 1764 8023
rect 1706 7963 1712 7997
rect 1752 7963 1764 7997
rect 1706 7937 1764 7963
rect 1806 7997 1864 8023
rect 1806 7963 1818 7997
rect 1858 7963 1864 7997
rect 1806 7937 1864 7963
rect 1906 7997 1964 8023
rect 1906 7963 1918 7997
rect 1952 7963 1964 7997
rect 1906 7937 1964 7963
rect 2006 7997 2064 8023
rect 2006 7963 2012 7997
rect 2052 7963 2064 7997
rect 2006 7937 2064 7963
rect 2106 7997 2164 8023
rect 2106 7963 2118 7997
rect 2158 7963 2164 7997
rect 2106 7937 2164 7963
rect 2206 7997 2264 8023
rect 2206 7963 2218 7997
rect 2252 7963 2264 7997
rect 2206 7937 2264 7963
rect 2306 7997 2364 8023
rect 2306 7963 2318 7997
rect 2352 7963 2364 7997
rect 2306 7937 2364 7963
rect 2406 7997 2464 8023
rect 2406 7963 2418 7997
rect 2452 7963 2464 7997
rect 2406 7937 2464 7963
rect 2506 7997 2564 8023
rect 2506 7963 2518 7997
rect 2552 7963 2564 7997
rect 2506 7937 2564 7963
rect 2606 7997 2664 8023
rect 2606 7963 2618 7997
rect 2652 7963 2664 7997
rect 2606 7937 2664 7963
rect 2706 7997 2764 8023
rect 2706 7963 2712 7997
rect 2752 7963 2764 7997
rect 2706 7937 2764 7963
rect 2806 7997 2864 8023
rect 2806 7963 2818 7997
rect 2858 7963 2864 7997
rect 2806 7937 2864 7963
rect 2906 7997 2964 8023
rect 2906 7963 2912 7997
rect 2952 7963 2964 7997
rect 2906 7937 2964 7963
rect 3006 7997 3064 8023
rect 3006 7963 3018 7997
rect 3058 7963 3064 7997
rect 3006 7937 3064 7963
rect 3106 7997 3164 8023
rect 3106 7963 3118 7997
rect 3152 7963 3164 7997
rect 3106 7937 3164 7963
rect 3206 7997 3264 8023
rect 3206 7963 3218 7997
rect 3252 7963 3264 7997
rect 3206 7937 3264 7963
rect 3306 7997 3364 8023
rect 3306 7963 3318 7997
rect 3352 7963 3364 7997
rect 3306 7937 3364 7963
rect 3406 7997 3464 8023
rect 3406 7963 3418 7997
rect 3452 7963 3464 7997
rect 3406 7937 3464 7963
rect 3506 7997 3564 8023
rect 3506 7963 3518 7997
rect 3552 7963 3564 7997
rect 3506 7937 3564 7963
rect 3606 7997 3664 8023
rect 3606 7963 3618 7997
rect 3652 7963 3664 7997
rect 3606 7937 3664 7963
rect 3706 7997 3764 8023
rect 3706 7963 3718 7997
rect 3752 7963 3764 7997
rect 3706 7937 3764 7963
rect 3806 7997 3864 8023
rect 3806 7963 3818 7997
rect 3852 7963 3864 7997
rect 3806 7937 3864 7963
rect 3906 7997 3964 8023
rect 3906 7963 3918 7997
rect 3952 7963 3964 7997
rect 3906 7937 3964 7963
rect 4006 7997 4064 8023
rect 4006 7963 4018 7997
rect 4052 7963 4064 7997
rect 4006 7937 4064 7963
rect 4106 7997 4164 8023
rect 4106 7963 4118 7997
rect 4152 7963 4164 7997
rect 4106 7937 4164 7963
rect 4206 7997 4264 8023
rect 4206 7963 4218 7997
rect 4252 7963 4264 7997
rect 4206 7937 4264 7963
rect 4306 7997 4364 8023
rect 4306 7963 4318 7997
rect 4352 7963 4364 7997
rect 4306 7937 4364 7963
rect 4406 7997 4464 8023
rect 4406 7963 4418 7997
rect 4452 7963 4464 7997
rect 4406 7937 4464 7963
rect 4506 7997 4564 8023
rect 4506 7963 4518 7997
rect 4552 7963 4564 7997
rect 4506 7937 4564 7963
rect 4606 7997 4664 8023
rect 4606 7963 4618 7997
rect 4652 7963 4664 7997
rect 4606 7937 4664 7963
rect 4706 7997 4764 8023
rect 4706 7963 4718 7997
rect 4752 7963 4764 7997
rect 4706 7937 4764 7963
rect 4806 7997 4864 8023
rect 4806 7963 4818 7997
rect 4852 7963 4864 7997
rect 4806 7937 4864 7963
rect 4906 7997 4964 8023
rect 4906 7963 4912 7997
rect 4952 7963 4964 7997
rect 4906 7937 4964 7963
rect 5006 7997 5064 8023
rect 5006 7963 5018 7997
rect 5058 7963 5064 7997
rect 5006 7937 5064 7963
rect 5106 7997 5164 8023
rect 5106 7963 5118 7997
rect 5152 7963 5164 7997
rect 5106 7937 5164 7963
rect 5206 7997 5264 8023
rect 5206 7963 5218 7997
rect 5252 7963 5264 7997
rect 5206 7937 5264 7963
rect 5306 7997 5364 8023
rect 5306 7963 5318 7997
rect 5352 7963 5364 7997
rect 5306 7937 5364 7963
rect 5406 7997 5464 8023
rect 5406 7963 5418 7997
rect 5452 7963 5464 7997
rect 5406 7937 5464 7963
rect 5506 7997 5564 8023
rect 5506 7963 5518 7997
rect 5552 7963 5564 7997
rect 5506 7937 5564 7963
rect 5606 7997 5664 8023
rect 5606 7963 5618 7997
rect 5652 7963 5664 7997
rect 5606 7937 5664 7963
rect 5706 7997 5764 8023
rect 5706 7963 5718 7997
rect 5752 7963 5764 7997
rect 5706 7937 5764 7963
rect 5806 7997 5864 8023
rect 5806 7963 5818 7997
rect 5852 7963 5864 7997
rect 5806 7937 5864 7963
rect 5906 7997 5964 8023
rect 5906 7963 5918 7997
rect 5952 7963 5964 7997
rect 5906 7937 5964 7963
rect 6006 7997 6064 8023
rect 6006 7963 6018 7997
rect 6052 7963 6064 7997
rect 6006 7937 6064 7963
rect 6106 7997 6164 8023
rect 6106 7963 6118 7997
rect 6152 7963 6164 7997
rect 6106 7937 6164 7963
rect 6206 7997 6264 8023
rect 6206 7963 6218 7997
rect 6252 7963 6264 7997
rect 6206 7937 6264 7963
rect 6306 7997 6364 8023
rect 6306 7963 6318 7997
rect 6352 7963 6364 7997
rect 6306 7937 6364 7963
rect 6406 7997 6464 8023
rect 6618 8016 6862 8050
rect 6406 7963 6418 7997
rect 6452 7963 6464 7997
rect 6508 7978 6516 8012
rect 6558 7978 6574 8012
rect 6618 7997 6652 8016
rect 6406 7937 6464 7963
rect 6828 8013 6862 8016
rect 6828 7997 6962 8013
rect 6618 7947 6652 7963
rect 6696 7948 6712 7982
rect 6754 7948 6762 7982
rect 6862 7963 6928 7997
rect 6828 7947 6962 7963
rect 7028 7997 7162 8013
rect 7062 7963 7128 7997
rect 7028 7947 7162 7963
rect 7228 7997 7262 8013
rect 7228 7947 7262 7963
rect 7328 7997 7462 8013
rect 7362 7963 7428 7997
rect 7328 7947 7462 7963
rect 6 7857 64 7883
rect 6 7823 18 7857
rect 58 7823 64 7857
rect 6 7797 64 7823
rect 106 7857 164 7883
rect 106 7823 118 7857
rect 152 7823 164 7857
rect 106 7797 164 7823
rect 206 7857 264 7883
rect 206 7823 218 7857
rect 252 7823 264 7857
rect 206 7797 264 7823
rect 306 7857 364 7883
rect 306 7823 318 7857
rect 352 7823 364 7857
rect 306 7797 364 7823
rect 406 7857 464 7883
rect 406 7823 418 7857
rect 452 7823 464 7857
rect 406 7797 464 7823
rect 506 7857 564 7883
rect 506 7823 518 7857
rect 552 7823 564 7857
rect 506 7797 564 7823
rect 606 7857 664 7883
rect 606 7823 612 7857
rect 652 7823 664 7857
rect 606 7797 664 7823
rect 706 7857 764 7883
rect 706 7823 718 7857
rect 758 7823 764 7857
rect 706 7797 764 7823
rect 806 7857 864 7883
rect 806 7823 812 7857
rect 852 7823 864 7857
rect 806 7797 864 7823
rect 906 7857 964 7883
rect 906 7823 918 7857
rect 958 7823 964 7857
rect 906 7797 964 7823
rect 1006 7857 1064 7883
rect 1006 7823 1018 7857
rect 1052 7823 1064 7857
rect 1006 7797 1064 7823
rect 1106 7857 1164 7883
rect 1106 7823 1118 7857
rect 1152 7823 1164 7857
rect 1106 7797 1164 7823
rect 1206 7857 1264 7883
rect 1206 7823 1218 7857
rect 1252 7823 1264 7857
rect 1206 7797 1264 7823
rect 1306 7857 1364 7883
rect 1306 7823 1318 7857
rect 1352 7823 1364 7857
rect 1306 7797 1364 7823
rect 1406 7857 1464 7883
rect 1406 7823 1412 7857
rect 1452 7823 1464 7857
rect 1406 7797 1464 7823
rect 1506 7857 1564 7883
rect 1506 7823 1518 7857
rect 1558 7823 1564 7857
rect 1506 7797 1564 7823
rect 1606 7857 1664 7883
rect 1606 7823 1612 7857
rect 1652 7823 1664 7857
rect 1606 7797 1664 7823
rect 1706 7857 1764 7883
rect 1706 7823 1718 7857
rect 1758 7823 1764 7857
rect 1706 7797 1764 7823
rect 1806 7857 1864 7883
rect 1806 7823 1818 7857
rect 1852 7823 1864 7857
rect 1806 7797 1864 7823
rect 1906 7857 1964 7883
rect 1906 7823 1918 7857
rect 1952 7823 1964 7857
rect 1906 7797 1964 7823
rect 2006 7857 2064 7883
rect 2006 7823 2018 7857
rect 2052 7823 2064 7857
rect 2006 7797 2064 7823
rect 2106 7857 2164 7883
rect 2106 7823 2118 7857
rect 2152 7823 2164 7857
rect 2106 7797 2164 7823
rect 2206 7857 2264 7883
rect 2206 7823 2218 7857
rect 2252 7823 2264 7857
rect 2206 7797 2264 7823
rect 2306 7857 2364 7883
rect 2306 7823 2318 7857
rect 2352 7823 2364 7857
rect 2306 7797 2364 7823
rect 2406 7857 2464 7883
rect 2406 7823 2418 7857
rect 2452 7823 2464 7857
rect 2406 7797 2464 7823
rect 2506 7857 2564 7883
rect 2506 7823 2512 7857
rect 2552 7823 2564 7857
rect 2506 7797 2564 7823
rect 2606 7857 2664 7883
rect 2606 7823 2618 7857
rect 2658 7823 2664 7857
rect 2606 7797 2664 7823
rect 2706 7857 2764 7883
rect 2706 7823 2718 7857
rect 2752 7823 2764 7857
rect 2706 7797 2764 7823
rect 2806 7857 2864 7883
rect 2806 7823 2818 7857
rect 2852 7823 2864 7857
rect 2806 7797 2864 7823
rect 2906 7857 2964 7883
rect 2906 7823 2918 7857
rect 2952 7823 2964 7857
rect 2906 7797 2964 7823
rect 3006 7857 3064 7883
rect 3006 7823 3018 7857
rect 3052 7823 3064 7857
rect 3006 7797 3064 7823
rect 3106 7857 3164 7883
rect 3106 7823 3118 7857
rect 3152 7823 3164 7857
rect 3106 7797 3164 7823
rect 3206 7857 3264 7883
rect 3206 7823 3218 7857
rect 3252 7823 3264 7857
rect 3206 7797 3264 7823
rect 3306 7857 3364 7883
rect 3306 7823 3312 7857
rect 3352 7823 3364 7857
rect 3306 7797 3364 7823
rect 3406 7857 3464 7883
rect 3406 7823 3418 7857
rect 3458 7823 3464 7857
rect 3406 7797 3464 7823
rect 3506 7857 3564 7883
rect 3506 7823 3518 7857
rect 3552 7823 3564 7857
rect 3506 7797 3564 7823
rect 3606 7857 3664 7883
rect 3606 7823 3618 7857
rect 3652 7823 3664 7857
rect 3606 7797 3664 7823
rect 3706 7857 3764 7883
rect 3706 7823 3712 7857
rect 3752 7823 3764 7857
rect 3706 7797 3764 7823
rect 3806 7857 3864 7883
rect 3806 7823 3818 7857
rect 3858 7823 3864 7857
rect 3806 7797 3864 7823
rect 3906 7857 3964 7883
rect 3906 7823 3912 7857
rect 3952 7823 3964 7857
rect 3906 7797 3964 7823
rect 4006 7857 4064 7883
rect 4006 7823 4018 7857
rect 4058 7823 4064 7857
rect 4006 7797 4064 7823
rect 4106 7857 4164 7883
rect 4106 7823 4112 7857
rect 4152 7823 4164 7857
rect 4106 7797 4164 7823
rect 4206 7857 4264 7883
rect 4206 7823 4218 7857
rect 4258 7823 4264 7857
rect 4206 7797 4264 7823
rect 4306 7857 4364 7883
rect 4306 7823 4318 7857
rect 4352 7823 4364 7857
rect 4306 7797 4364 7823
rect 4406 7857 4464 7883
rect 4406 7823 4418 7857
rect 4452 7823 4464 7857
rect 4406 7797 4464 7823
rect 4506 7857 4564 7883
rect 4506 7823 4512 7857
rect 4552 7823 4564 7857
rect 4506 7797 4564 7823
rect 4606 7857 4664 7883
rect 4606 7823 4618 7857
rect 4658 7823 4664 7857
rect 4606 7797 4664 7823
rect 4706 7857 4764 7883
rect 4706 7823 4712 7857
rect 4752 7823 4764 7857
rect 4706 7797 4764 7823
rect 4806 7857 4864 7883
rect 4806 7823 4818 7857
rect 4858 7823 4864 7857
rect 4806 7797 4864 7823
rect 4906 7857 4964 7883
rect 4906 7823 4912 7857
rect 4952 7823 4964 7857
rect 4906 7797 4964 7823
rect 5006 7857 5064 7883
rect 5006 7823 5018 7857
rect 5058 7823 5064 7857
rect 5006 7797 5064 7823
rect 5106 7857 5164 7883
rect 5106 7823 5118 7857
rect 5152 7823 5164 7857
rect 5106 7797 5164 7823
rect 5206 7857 5264 7883
rect 5206 7823 5218 7857
rect 5252 7823 5264 7857
rect 5206 7797 5264 7823
rect 5306 7857 5364 7883
rect 5306 7823 5318 7857
rect 5352 7823 5364 7857
rect 5306 7797 5364 7823
rect 5406 7857 5464 7883
rect 5406 7823 5418 7857
rect 5452 7823 5464 7857
rect 5406 7797 5464 7823
rect 5506 7857 5564 7883
rect 5506 7823 5512 7857
rect 5552 7823 5564 7857
rect 5506 7797 5564 7823
rect 5606 7857 5664 7883
rect 5606 7823 5618 7857
rect 5658 7823 5664 7857
rect 5606 7797 5664 7823
rect 5706 7857 5764 7883
rect 5706 7823 5712 7857
rect 5752 7823 5764 7857
rect 5706 7797 5764 7823
rect 5806 7857 5864 7883
rect 5806 7823 5818 7857
rect 5858 7823 5864 7857
rect 5806 7797 5864 7823
rect 5906 7857 5964 7883
rect 5906 7823 5918 7857
rect 5952 7823 5964 7857
rect 5906 7797 5964 7823
rect 6006 7857 6064 7883
rect 6006 7823 6018 7857
rect 6052 7823 6064 7857
rect 6006 7797 6064 7823
rect 6106 7857 6164 7883
rect 6106 7823 6118 7857
rect 6152 7823 6164 7857
rect 6106 7797 6164 7823
rect 6206 7857 6264 7883
rect 6206 7823 6218 7857
rect 6252 7823 6264 7857
rect 6206 7797 6264 7823
rect 6306 7857 6364 7883
rect 6306 7823 6318 7857
rect 6352 7823 6364 7857
rect 6306 7797 6364 7823
rect 6406 7857 6464 7883
rect 6618 7876 6862 7910
rect 6406 7823 6412 7857
rect 6452 7823 6464 7857
rect 6508 7838 6516 7872
rect 6558 7838 6574 7872
rect 6618 7857 6652 7876
rect 6406 7797 6464 7823
rect 6828 7857 6862 7876
rect 6618 7807 6652 7823
rect 6696 7808 6712 7842
rect 6754 7808 6762 7842
rect 6828 7807 6862 7823
rect 6928 7857 7162 7873
rect 6962 7823 7028 7857
rect 7062 7823 7128 7857
rect 6928 7807 7162 7823
rect 7228 7857 7262 7873
rect 7228 7807 7262 7823
rect 7328 7857 7462 7873
rect 7362 7823 7428 7857
rect 7328 7807 7462 7823
rect 6 7717 64 7743
rect 6 7683 18 7717
rect 58 7683 64 7717
rect 6 7657 64 7683
rect 106 7717 164 7743
rect 106 7683 118 7717
rect 152 7683 164 7717
rect 106 7657 164 7683
rect 206 7717 264 7743
rect 206 7683 218 7717
rect 252 7683 264 7717
rect 206 7657 264 7683
rect 306 7717 364 7743
rect 306 7683 318 7717
rect 352 7683 364 7717
rect 306 7657 364 7683
rect 406 7717 464 7743
rect 406 7683 418 7717
rect 452 7683 464 7717
rect 406 7657 464 7683
rect 506 7717 564 7743
rect 506 7683 518 7717
rect 552 7683 564 7717
rect 506 7657 564 7683
rect 606 7717 664 7743
rect 606 7683 618 7717
rect 652 7683 664 7717
rect 606 7657 664 7683
rect 706 7717 764 7743
rect 706 7683 718 7717
rect 752 7683 764 7717
rect 706 7657 764 7683
rect 806 7717 864 7743
rect 806 7683 818 7717
rect 852 7683 864 7717
rect 806 7657 864 7683
rect 906 7717 964 7743
rect 906 7683 918 7717
rect 952 7683 964 7717
rect 906 7657 964 7683
rect 1006 7717 1064 7743
rect 1006 7683 1018 7717
rect 1052 7683 1064 7717
rect 1006 7657 1064 7683
rect 1106 7717 1164 7743
rect 1106 7683 1118 7717
rect 1152 7683 1164 7717
rect 1106 7657 1164 7683
rect 1206 7717 1264 7743
rect 1206 7683 1218 7717
rect 1252 7683 1264 7717
rect 1206 7657 1264 7683
rect 1306 7717 1364 7743
rect 1306 7683 1318 7717
rect 1352 7683 1364 7717
rect 1306 7657 1364 7683
rect 1406 7717 1464 7743
rect 1406 7683 1418 7717
rect 1452 7683 1464 7717
rect 1406 7657 1464 7683
rect 1506 7717 1564 7743
rect 1506 7683 1512 7717
rect 1552 7683 1564 7717
rect 1506 7657 1564 7683
rect 1606 7717 1664 7743
rect 1606 7683 1618 7717
rect 1658 7683 1664 7717
rect 1606 7657 1664 7683
rect 1706 7717 1764 7743
rect 1706 7683 1712 7717
rect 1752 7683 1764 7717
rect 1706 7657 1764 7683
rect 1806 7717 1864 7743
rect 1806 7683 1818 7717
rect 1858 7683 1864 7717
rect 1806 7657 1864 7683
rect 1906 7717 1964 7743
rect 1906 7683 1918 7717
rect 1952 7683 1964 7717
rect 1906 7657 1964 7683
rect 2006 7717 2064 7743
rect 2006 7683 2018 7717
rect 2052 7683 2064 7717
rect 2006 7657 2064 7683
rect 2106 7717 2164 7743
rect 2106 7683 2118 7717
rect 2152 7683 2164 7717
rect 2106 7657 2164 7683
rect 2206 7717 2264 7743
rect 2206 7683 2218 7717
rect 2252 7683 2264 7717
rect 2206 7657 2264 7683
rect 2306 7717 2364 7743
rect 2306 7683 2318 7717
rect 2352 7683 2364 7717
rect 2306 7657 2364 7683
rect 2406 7717 2464 7743
rect 2406 7683 2418 7717
rect 2452 7683 2464 7717
rect 2406 7657 2464 7683
rect 2506 7717 2564 7743
rect 2506 7683 2518 7717
rect 2552 7683 2564 7717
rect 2506 7657 2564 7683
rect 2606 7717 2664 7743
rect 2606 7683 2618 7717
rect 2652 7683 2664 7717
rect 2606 7657 2664 7683
rect 2706 7717 2764 7743
rect 2706 7683 2712 7717
rect 2752 7683 2764 7717
rect 2706 7657 2764 7683
rect 2806 7717 2864 7743
rect 2806 7683 2818 7717
rect 2858 7683 2864 7717
rect 2806 7657 2864 7683
rect 2906 7717 2964 7743
rect 2906 7683 2918 7717
rect 2952 7683 2964 7717
rect 2906 7657 2964 7683
rect 3006 7717 3064 7743
rect 3006 7683 3018 7717
rect 3052 7683 3064 7717
rect 3006 7657 3064 7683
rect 3106 7717 3164 7743
rect 3106 7683 3118 7717
rect 3152 7683 3164 7717
rect 3106 7657 3164 7683
rect 3206 7717 3264 7743
rect 3206 7683 3218 7717
rect 3252 7683 3264 7717
rect 3206 7657 3264 7683
rect 3306 7717 3364 7743
rect 3306 7683 3318 7717
rect 3352 7683 3364 7717
rect 3306 7657 3364 7683
rect 3406 7717 3464 7743
rect 3406 7683 3418 7717
rect 3452 7683 3464 7717
rect 3406 7657 3464 7683
rect 3506 7717 3564 7743
rect 3506 7683 3518 7717
rect 3552 7683 3564 7717
rect 3506 7657 3564 7683
rect 3606 7717 3664 7743
rect 3606 7683 3618 7717
rect 3652 7683 3664 7717
rect 3606 7657 3664 7683
rect 3706 7717 3764 7743
rect 3706 7683 3718 7717
rect 3752 7683 3764 7717
rect 3706 7657 3764 7683
rect 3806 7717 3864 7743
rect 3806 7683 3818 7717
rect 3852 7683 3864 7717
rect 3806 7657 3864 7683
rect 3906 7717 3964 7743
rect 3906 7683 3918 7717
rect 3952 7683 3964 7717
rect 3906 7657 3964 7683
rect 4006 7717 4064 7743
rect 4006 7683 4018 7717
rect 4052 7683 4064 7717
rect 4006 7657 4064 7683
rect 4106 7717 4164 7743
rect 4106 7683 4112 7717
rect 4152 7683 4164 7717
rect 4106 7657 4164 7683
rect 4206 7717 4264 7743
rect 4206 7683 4218 7717
rect 4258 7683 4264 7717
rect 4206 7657 4264 7683
rect 4306 7717 4364 7743
rect 4306 7683 4312 7717
rect 4352 7683 4364 7717
rect 4306 7657 4364 7683
rect 4406 7717 4464 7743
rect 4406 7683 4418 7717
rect 4458 7683 4464 7717
rect 4406 7657 4464 7683
rect 4506 7717 4564 7743
rect 4506 7683 4518 7717
rect 4552 7683 4564 7717
rect 4506 7657 4564 7683
rect 4606 7717 4664 7743
rect 4606 7683 4618 7717
rect 4652 7683 4664 7717
rect 4606 7657 4664 7683
rect 4706 7717 4764 7743
rect 4706 7683 4718 7717
rect 4752 7683 4764 7717
rect 4706 7657 4764 7683
rect 4806 7717 4864 7743
rect 4806 7683 4818 7717
rect 4852 7683 4864 7717
rect 4806 7657 4864 7683
rect 4906 7717 4964 7743
rect 4906 7683 4918 7717
rect 4952 7683 4964 7717
rect 4906 7657 4964 7683
rect 5006 7717 5064 7743
rect 5006 7683 5018 7717
rect 5052 7683 5064 7717
rect 5006 7657 5064 7683
rect 5106 7717 5164 7743
rect 5106 7683 5118 7717
rect 5152 7683 5164 7717
rect 5106 7657 5164 7683
rect 5206 7717 5264 7743
rect 5206 7683 5218 7717
rect 5252 7683 5264 7717
rect 5206 7657 5264 7683
rect 5306 7717 5364 7743
rect 5306 7683 5318 7717
rect 5352 7683 5364 7717
rect 5306 7657 5364 7683
rect 5406 7717 5464 7743
rect 5406 7683 5418 7717
rect 5452 7683 5464 7717
rect 5406 7657 5464 7683
rect 5506 7717 5564 7743
rect 5506 7683 5512 7717
rect 5552 7683 5564 7717
rect 5506 7657 5564 7683
rect 5606 7717 5664 7743
rect 5606 7683 5618 7717
rect 5658 7683 5664 7717
rect 5606 7657 5664 7683
rect 5706 7717 5764 7743
rect 5706 7683 5712 7717
rect 5752 7683 5764 7717
rect 5706 7657 5764 7683
rect 5806 7717 5864 7743
rect 5806 7683 5818 7717
rect 5858 7683 5864 7717
rect 5806 7657 5864 7683
rect 5906 7717 5964 7743
rect 5906 7683 5918 7717
rect 5952 7683 5964 7717
rect 5906 7657 5964 7683
rect 6006 7717 6064 7743
rect 6006 7683 6018 7717
rect 6052 7683 6064 7717
rect 6006 7657 6064 7683
rect 6106 7717 6164 7743
rect 6106 7683 6118 7717
rect 6152 7683 6164 7717
rect 6106 7657 6164 7683
rect 6206 7717 6264 7743
rect 6206 7683 6218 7717
rect 6252 7683 6264 7717
rect 6206 7657 6264 7683
rect 6306 7717 6364 7743
rect 6306 7683 6318 7717
rect 6352 7683 6364 7717
rect 6306 7657 6364 7683
rect 6406 7717 6464 7743
rect 6618 7736 6862 7770
rect 6406 7683 6418 7717
rect 6452 7683 6464 7717
rect 6508 7698 6516 7732
rect 6558 7698 6574 7732
rect 6618 7717 6652 7736
rect 6406 7657 6464 7683
rect 6828 7733 6862 7736
rect 6828 7717 6962 7733
rect 6618 7667 6652 7683
rect 6696 7668 6712 7702
rect 6754 7668 6762 7702
rect 6862 7683 6928 7717
rect 6828 7667 6962 7683
rect 7028 7717 7062 7733
rect 7028 7667 7062 7683
rect 7128 7717 7262 7733
rect 7162 7683 7228 7717
rect 7128 7667 7262 7683
rect 7328 7717 7462 7733
rect 7362 7683 7428 7717
rect 7328 7667 7462 7683
rect 6 7577 64 7603
rect 6 7543 18 7577
rect 58 7543 64 7577
rect 6 7517 64 7543
rect 106 7577 164 7603
rect 106 7543 118 7577
rect 152 7543 164 7577
rect 106 7517 164 7543
rect 206 7577 264 7603
rect 206 7543 218 7577
rect 252 7543 264 7577
rect 206 7517 264 7543
rect 306 7577 364 7603
rect 306 7543 318 7577
rect 352 7543 364 7577
rect 306 7517 364 7543
rect 406 7577 464 7603
rect 406 7543 418 7577
rect 452 7543 464 7577
rect 406 7517 464 7543
rect 506 7577 564 7603
rect 506 7543 518 7577
rect 552 7543 564 7577
rect 506 7517 564 7543
rect 606 7577 664 7603
rect 606 7543 618 7577
rect 652 7543 664 7577
rect 606 7517 664 7543
rect 706 7577 764 7603
rect 706 7543 718 7577
rect 752 7543 764 7577
rect 706 7517 764 7543
rect 806 7577 864 7603
rect 806 7543 818 7577
rect 852 7543 864 7577
rect 806 7517 864 7543
rect 906 7577 964 7603
rect 906 7543 918 7577
rect 952 7543 964 7577
rect 906 7517 964 7543
rect 1006 7577 1064 7603
rect 1006 7543 1012 7577
rect 1052 7543 1064 7577
rect 1006 7517 1064 7543
rect 1106 7577 1164 7603
rect 1106 7543 1118 7577
rect 1158 7543 1164 7577
rect 1106 7517 1164 7543
rect 1206 7577 1264 7603
rect 1206 7543 1218 7577
rect 1252 7543 1264 7577
rect 1206 7517 1264 7543
rect 1306 7577 1364 7603
rect 1306 7543 1312 7577
rect 1352 7543 1364 7577
rect 1306 7517 1364 7543
rect 1406 7577 1464 7603
rect 1406 7543 1418 7577
rect 1458 7543 1464 7577
rect 1406 7517 1464 7543
rect 1506 7577 1564 7603
rect 1506 7543 1518 7577
rect 1552 7543 1564 7577
rect 1506 7517 1564 7543
rect 1606 7577 1664 7603
rect 1606 7543 1618 7577
rect 1652 7543 1664 7577
rect 1606 7517 1664 7543
rect 1706 7577 1764 7603
rect 1706 7543 1718 7577
rect 1752 7543 1764 7577
rect 1706 7517 1764 7543
rect 1806 7577 1864 7603
rect 1806 7543 1818 7577
rect 1852 7543 1864 7577
rect 1806 7517 1864 7543
rect 1906 7577 1964 7603
rect 1906 7543 1918 7577
rect 1952 7543 1964 7577
rect 1906 7517 1964 7543
rect 2006 7577 2064 7603
rect 2006 7543 2018 7577
rect 2052 7543 2064 7577
rect 2006 7517 2064 7543
rect 2106 7577 2164 7603
rect 2106 7543 2118 7577
rect 2152 7543 2164 7577
rect 2106 7517 2164 7543
rect 2206 7577 2264 7603
rect 2206 7543 2218 7577
rect 2252 7543 2264 7577
rect 2206 7517 2264 7543
rect 2306 7577 2364 7603
rect 2306 7543 2318 7577
rect 2352 7543 2364 7577
rect 2306 7517 2364 7543
rect 2406 7577 2464 7603
rect 2406 7543 2418 7577
rect 2452 7543 2464 7577
rect 2406 7517 2464 7543
rect 2506 7577 2564 7603
rect 2506 7543 2518 7577
rect 2552 7543 2564 7577
rect 2506 7517 2564 7543
rect 2606 7577 2664 7603
rect 2606 7543 2618 7577
rect 2652 7543 2664 7577
rect 2606 7517 2664 7543
rect 2706 7577 2764 7603
rect 2706 7543 2712 7577
rect 2752 7543 2764 7577
rect 2706 7517 2764 7543
rect 2806 7577 2864 7603
rect 2806 7543 2818 7577
rect 2858 7543 2864 7577
rect 2806 7517 2864 7543
rect 2906 7577 2964 7603
rect 2906 7543 2918 7577
rect 2952 7543 2964 7577
rect 2906 7517 2964 7543
rect 3006 7577 3064 7603
rect 3006 7543 3012 7577
rect 3052 7543 3064 7577
rect 3006 7517 3064 7543
rect 3106 7577 3164 7603
rect 3106 7543 3118 7577
rect 3158 7543 3164 7577
rect 3106 7517 3164 7543
rect 3206 7577 3264 7603
rect 3206 7543 3212 7577
rect 3252 7543 3264 7577
rect 3206 7517 3264 7543
rect 3306 7577 3364 7603
rect 3306 7543 3318 7577
rect 3358 7543 3364 7577
rect 3306 7517 3364 7543
rect 3406 7577 3464 7603
rect 3406 7543 3418 7577
rect 3452 7543 3464 7577
rect 3406 7517 3464 7543
rect 3506 7577 3564 7603
rect 3506 7543 3518 7577
rect 3552 7543 3564 7577
rect 3506 7517 3564 7543
rect 3606 7577 3664 7603
rect 3606 7543 3618 7577
rect 3652 7543 3664 7577
rect 3606 7517 3664 7543
rect 3706 7577 3764 7603
rect 3706 7543 3718 7577
rect 3752 7543 3764 7577
rect 3706 7517 3764 7543
rect 3806 7577 3864 7603
rect 3806 7543 3818 7577
rect 3852 7543 3864 7577
rect 3806 7517 3864 7543
rect 3906 7577 3964 7603
rect 3906 7543 3912 7577
rect 3952 7543 3964 7577
rect 3906 7517 3964 7543
rect 4006 7577 4064 7603
rect 4006 7543 4018 7577
rect 4058 7543 4064 7577
rect 4006 7517 4064 7543
rect 4106 7577 4164 7603
rect 4106 7543 4118 7577
rect 4152 7543 4164 7577
rect 4106 7517 4164 7543
rect 4206 7577 4264 7603
rect 4206 7543 4218 7577
rect 4252 7543 4264 7577
rect 4206 7517 4264 7543
rect 4306 7577 4364 7603
rect 4306 7543 4318 7577
rect 4352 7543 4364 7577
rect 4306 7517 4364 7543
rect 4406 7577 4464 7603
rect 4406 7543 4418 7577
rect 4452 7543 4464 7577
rect 4406 7517 4464 7543
rect 4506 7577 4564 7603
rect 4506 7543 4518 7577
rect 4552 7543 4564 7577
rect 4506 7517 4564 7543
rect 4606 7577 4664 7603
rect 4606 7543 4618 7577
rect 4652 7543 4664 7577
rect 4606 7517 4664 7543
rect 4706 7577 4764 7603
rect 4706 7543 4718 7577
rect 4752 7543 4764 7577
rect 4706 7517 4764 7543
rect 4806 7577 4864 7603
rect 4806 7543 4818 7577
rect 4852 7543 4864 7577
rect 4806 7517 4864 7543
rect 4906 7577 4964 7603
rect 4906 7543 4912 7577
rect 4952 7543 4964 7577
rect 4906 7517 4964 7543
rect 5006 7577 5064 7603
rect 5006 7543 5018 7577
rect 5058 7543 5064 7577
rect 5006 7517 5064 7543
rect 5106 7577 5164 7603
rect 5106 7543 5112 7577
rect 5152 7543 5164 7577
rect 5106 7517 5164 7543
rect 5206 7577 5264 7603
rect 5206 7543 5218 7577
rect 5258 7543 5264 7577
rect 5206 7517 5264 7543
rect 5306 7577 5364 7603
rect 5306 7543 5318 7577
rect 5352 7543 5364 7577
rect 5306 7517 5364 7543
rect 5406 7577 5464 7603
rect 5406 7543 5418 7577
rect 5452 7543 5464 7577
rect 5406 7517 5464 7543
rect 5506 7577 5564 7603
rect 5506 7543 5518 7577
rect 5552 7543 5564 7577
rect 5506 7517 5564 7543
rect 5606 7577 5664 7603
rect 5606 7543 5618 7577
rect 5652 7543 5664 7577
rect 5606 7517 5664 7543
rect 5706 7577 5764 7603
rect 5706 7543 5718 7577
rect 5752 7543 5764 7577
rect 5706 7517 5764 7543
rect 5806 7577 5864 7603
rect 5806 7543 5818 7577
rect 5852 7543 5864 7577
rect 5806 7517 5864 7543
rect 5906 7577 5964 7603
rect 5906 7543 5918 7577
rect 5952 7543 5964 7577
rect 5906 7517 5964 7543
rect 6006 7577 6064 7603
rect 6006 7543 6018 7577
rect 6052 7543 6064 7577
rect 6006 7517 6064 7543
rect 6106 7577 6164 7603
rect 6106 7543 6118 7577
rect 6152 7543 6164 7577
rect 6106 7517 6164 7543
rect 6206 7577 6264 7603
rect 6206 7543 6218 7577
rect 6252 7543 6264 7577
rect 6206 7517 6264 7543
rect 6306 7577 6364 7603
rect 6306 7543 6318 7577
rect 6352 7543 6364 7577
rect 6306 7517 6364 7543
rect 6406 7577 6464 7603
rect 6618 7596 6862 7630
rect 6406 7543 6412 7577
rect 6452 7543 6464 7577
rect 6508 7558 6516 7592
rect 6558 7558 6574 7592
rect 6618 7577 6652 7596
rect 6406 7517 6464 7543
rect 6828 7577 6862 7596
rect 6618 7527 6652 7543
rect 6696 7528 6712 7562
rect 6754 7528 6762 7562
rect 6828 7527 6862 7543
rect 6928 7577 7062 7593
rect 6962 7543 7028 7577
rect 6928 7527 7062 7543
rect 7128 7577 7262 7593
rect 7162 7543 7228 7577
rect 7128 7527 7262 7543
rect 7328 7577 7462 7593
rect 7362 7543 7428 7577
rect 7328 7527 7462 7543
rect 8 7420 18 7454
rect 52 7420 118 7454
rect 152 7420 168 7454
rect 208 7436 218 7470
rect 252 7436 318 7470
rect 352 7436 368 7470
rect 408 7420 418 7454
rect 452 7420 518 7454
rect 552 7420 568 7454
rect 608 7436 618 7470
rect 652 7436 718 7470
rect 752 7436 768 7470
rect 808 7420 818 7454
rect 852 7420 918 7454
rect 952 7420 968 7454
rect 1008 7436 1018 7470
rect 1052 7436 1118 7470
rect 1152 7436 1168 7470
rect 1208 7420 1218 7454
rect 1252 7420 1318 7454
rect 1352 7420 1368 7454
rect 1408 7436 1418 7470
rect 1452 7436 1518 7470
rect 1552 7436 1568 7470
rect 1608 7420 1618 7454
rect 1652 7420 1718 7454
rect 1752 7420 1768 7454
rect 1808 7436 1818 7470
rect 1852 7436 1918 7470
rect 1952 7436 1968 7470
rect 2008 7420 2018 7454
rect 2052 7420 2118 7454
rect 2152 7420 2168 7454
rect 2208 7436 2218 7470
rect 2252 7436 2318 7470
rect 2352 7436 2368 7470
rect 2408 7420 2418 7454
rect 2452 7420 2518 7454
rect 2552 7420 2568 7454
rect 2608 7436 2618 7470
rect 2652 7436 2718 7470
rect 2752 7436 2768 7470
rect 2808 7420 2818 7454
rect 2852 7420 2918 7454
rect 2952 7420 2968 7454
rect 3008 7436 3018 7470
rect 3052 7436 3118 7470
rect 3152 7436 3168 7470
rect 3208 7420 3218 7454
rect 3252 7420 3318 7454
rect 3352 7420 3368 7454
rect 3408 7436 3418 7470
rect 3452 7436 3518 7470
rect 3552 7436 3568 7470
rect 3608 7420 3618 7454
rect 3652 7420 3718 7454
rect 3752 7420 3768 7454
rect 3808 7436 3818 7470
rect 3852 7436 3918 7470
rect 3952 7436 3968 7470
rect 4008 7420 4018 7454
rect 4052 7420 4118 7454
rect 4152 7420 4168 7454
rect 4208 7436 4218 7470
rect 4252 7436 4318 7470
rect 4352 7436 4368 7470
rect 4408 7420 4418 7454
rect 4452 7420 4518 7454
rect 4552 7420 4568 7454
rect 4608 7436 4618 7470
rect 4652 7436 4718 7470
rect 4752 7436 4768 7470
rect 4808 7420 4818 7454
rect 4852 7420 4918 7454
rect 4952 7420 4968 7454
rect 5008 7436 5018 7470
rect 5052 7436 5118 7470
rect 5152 7436 5168 7470
rect 5208 7420 5218 7454
rect 5252 7420 5318 7454
rect 5352 7420 5368 7454
rect 5408 7436 5418 7470
rect 5452 7436 5518 7470
rect 5552 7436 5568 7470
rect 5608 7420 5618 7454
rect 5652 7420 5718 7454
rect 5752 7420 5768 7454
rect 5808 7436 5818 7470
rect 5852 7436 5918 7470
rect 5952 7436 5968 7470
rect 6008 7420 6018 7454
rect 6052 7420 6118 7454
rect 6152 7420 6168 7454
rect 6208 7436 6218 7470
rect 6252 7436 6318 7470
rect 6352 7436 6368 7470
rect 6516 7451 6568 7468
rect 6550 7434 6568 7451
rect 6602 7434 6618 7468
rect 6652 7434 6668 7468
rect 6702 7439 6720 7468
rect 6702 7434 6754 7439
rect 6862 7434 6878 7468
rect 6912 7434 6928 7468
rect 6962 7434 6978 7468
rect 7012 7434 7028 7468
rect 7062 7434 7078 7468
rect 7112 7434 7128 7468
rect 7162 7434 7178 7468
rect 7212 7434 7228 7468
rect 7262 7434 7278 7468
rect 7312 7434 7328 7468
rect 7362 7434 7378 7468
rect 7412 7434 7428 7468
rect 6 7347 64 7373
rect 6 7313 18 7347
rect 52 7313 64 7347
rect 6 7287 64 7313
rect 106 7347 164 7373
rect 106 7313 118 7347
rect 152 7313 164 7347
rect 106 7287 164 7313
rect 206 7347 264 7373
rect 206 7313 218 7347
rect 252 7313 264 7347
rect 206 7287 264 7313
rect 306 7347 364 7373
rect 306 7313 318 7347
rect 352 7313 364 7347
rect 306 7287 364 7313
rect 406 7347 464 7373
rect 406 7313 418 7347
rect 452 7313 464 7347
rect 406 7287 464 7313
rect 506 7347 564 7373
rect 506 7313 518 7347
rect 552 7313 564 7347
rect 506 7287 564 7313
rect 606 7347 664 7373
rect 606 7313 618 7347
rect 652 7313 664 7347
rect 606 7287 664 7313
rect 706 7347 764 7373
rect 706 7313 718 7347
rect 752 7313 764 7347
rect 706 7287 764 7313
rect 806 7347 864 7373
rect 806 7313 818 7347
rect 852 7313 864 7347
rect 806 7287 864 7313
rect 906 7347 964 7373
rect 906 7313 918 7347
rect 952 7313 964 7347
rect 906 7287 964 7313
rect 1006 7347 1064 7373
rect 1006 7313 1018 7347
rect 1052 7313 1064 7347
rect 1006 7287 1064 7313
rect 1106 7347 1164 7373
rect 1106 7313 1118 7347
rect 1152 7313 1164 7347
rect 1106 7287 1164 7313
rect 1206 7347 1264 7373
rect 1206 7313 1212 7347
rect 1252 7313 1264 7347
rect 1206 7287 1264 7313
rect 1306 7347 1364 7373
rect 1306 7313 1318 7347
rect 1358 7313 1364 7347
rect 1306 7287 1364 7313
rect 1406 7347 1464 7373
rect 1406 7313 1418 7347
rect 1452 7313 1464 7347
rect 1406 7287 1464 7313
rect 1506 7347 1564 7373
rect 1506 7313 1512 7347
rect 1552 7313 1564 7347
rect 1506 7287 1564 7313
rect 1606 7347 1664 7373
rect 1606 7313 1618 7347
rect 1658 7313 1664 7347
rect 1606 7287 1664 7313
rect 1706 7347 1764 7373
rect 1706 7313 1718 7347
rect 1752 7313 1764 7347
rect 1706 7287 1764 7313
rect 1806 7347 1864 7373
rect 1806 7313 1818 7347
rect 1852 7313 1864 7347
rect 1806 7287 1864 7313
rect 1906 7347 1964 7373
rect 1906 7313 1918 7347
rect 1952 7313 1964 7347
rect 1906 7287 1964 7313
rect 2006 7347 2064 7373
rect 2006 7313 2018 7347
rect 2052 7313 2064 7347
rect 2006 7287 2064 7313
rect 2106 7347 2164 7373
rect 2106 7313 2112 7347
rect 2152 7313 2164 7347
rect 2106 7287 2164 7313
rect 2206 7347 2264 7373
rect 2206 7313 2218 7347
rect 2258 7313 2264 7347
rect 2206 7287 2264 7313
rect 2306 7347 2364 7373
rect 2306 7313 2312 7347
rect 2352 7313 2364 7347
rect 2306 7287 2364 7313
rect 2406 7347 2464 7373
rect 2406 7313 2418 7347
rect 2458 7313 2464 7347
rect 2406 7287 2464 7313
rect 2506 7347 2564 7373
rect 2506 7313 2512 7347
rect 2552 7313 2564 7347
rect 2506 7287 2564 7313
rect 2606 7347 2664 7373
rect 2606 7313 2618 7347
rect 2658 7313 2664 7347
rect 2606 7287 2664 7313
rect 2706 7347 2764 7373
rect 2706 7313 2718 7347
rect 2752 7313 2764 7347
rect 2706 7287 2764 7313
rect 2806 7347 2864 7373
rect 2806 7313 2818 7347
rect 2852 7313 2864 7347
rect 2806 7287 2864 7313
rect 2906 7347 2964 7373
rect 2906 7313 2918 7347
rect 2952 7313 2964 7347
rect 2906 7287 2964 7313
rect 3006 7347 3064 7373
rect 3006 7313 3018 7347
rect 3052 7313 3064 7347
rect 3006 7287 3064 7313
rect 3106 7347 3164 7373
rect 3106 7313 3118 7347
rect 3152 7313 3164 7347
rect 3106 7287 3164 7313
rect 3206 7347 3264 7373
rect 3206 7313 3218 7347
rect 3252 7313 3264 7347
rect 3206 7287 3264 7313
rect 3306 7347 3364 7373
rect 3306 7313 3318 7347
rect 3352 7313 3364 7347
rect 3306 7287 3364 7313
rect 3406 7347 3464 7373
rect 3406 7313 3418 7347
rect 3452 7313 3464 7347
rect 3406 7287 3464 7313
rect 3506 7347 3564 7373
rect 3506 7313 3518 7347
rect 3552 7313 3564 7347
rect 3506 7287 3564 7313
rect 3606 7347 3664 7373
rect 3606 7313 3618 7347
rect 3652 7313 3664 7347
rect 3606 7287 3664 7313
rect 3706 7347 3764 7373
rect 3706 7313 3718 7347
rect 3752 7313 3764 7347
rect 3706 7287 3764 7313
rect 3806 7347 3864 7373
rect 3806 7313 3818 7347
rect 3852 7313 3864 7347
rect 3806 7287 3864 7313
rect 3906 7347 3964 7373
rect 3906 7313 3918 7347
rect 3952 7313 3964 7347
rect 3906 7287 3964 7313
rect 4006 7347 4064 7373
rect 4006 7313 4018 7347
rect 4052 7313 4064 7347
rect 4006 7287 4064 7313
rect 4106 7347 4164 7373
rect 4106 7313 4118 7347
rect 4152 7313 4164 7347
rect 4106 7287 4164 7313
rect 4206 7347 4264 7373
rect 4206 7313 4218 7347
rect 4252 7313 4264 7347
rect 4206 7287 4264 7313
rect 4306 7347 4364 7373
rect 4306 7313 4318 7347
rect 4352 7313 4364 7347
rect 4306 7287 4364 7313
rect 4406 7347 4464 7373
rect 4406 7313 4418 7347
rect 4452 7313 4464 7347
rect 4406 7287 4464 7313
rect 4506 7347 4564 7373
rect 4506 7313 4518 7347
rect 4552 7313 4564 7347
rect 4506 7287 4564 7313
rect 4606 7347 4664 7373
rect 4606 7313 4618 7347
rect 4652 7313 4664 7347
rect 4606 7287 4664 7313
rect 4706 7347 4764 7373
rect 4706 7313 4718 7347
rect 4752 7313 4764 7347
rect 4706 7287 4764 7313
rect 4806 7347 4864 7373
rect 4806 7313 4818 7347
rect 4852 7313 4864 7347
rect 4806 7287 4864 7313
rect 4906 7347 4964 7373
rect 4906 7313 4918 7347
rect 4952 7313 4964 7347
rect 4906 7287 4964 7313
rect 5006 7347 5064 7373
rect 5006 7313 5018 7347
rect 5052 7313 5064 7347
rect 5006 7287 5064 7313
rect 5106 7347 5164 7373
rect 5106 7313 5118 7347
rect 5152 7313 5164 7347
rect 5106 7287 5164 7313
rect 5206 7347 5264 7373
rect 5206 7313 5218 7347
rect 5252 7313 5264 7347
rect 5206 7287 5264 7313
rect 5306 7347 5364 7373
rect 5306 7313 5318 7347
rect 5352 7313 5364 7347
rect 5306 7287 5364 7313
rect 5406 7347 5464 7373
rect 5406 7313 5418 7347
rect 5452 7313 5464 7347
rect 5406 7287 5464 7313
rect 5506 7347 5564 7373
rect 5506 7313 5518 7347
rect 5552 7313 5564 7347
rect 5506 7287 5564 7313
rect 5606 7347 5664 7373
rect 5606 7313 5618 7347
rect 5652 7313 5664 7347
rect 5606 7287 5664 7313
rect 5706 7347 5764 7373
rect 5706 7313 5718 7347
rect 5752 7313 5764 7347
rect 5706 7287 5764 7313
rect 5806 7347 5864 7373
rect 5806 7313 5818 7347
rect 5852 7313 5864 7347
rect 5806 7287 5864 7313
rect 5906 7347 5964 7373
rect 5906 7313 5918 7347
rect 5952 7313 5964 7347
rect 5906 7287 5964 7313
rect 6006 7347 6064 7373
rect 6006 7313 6018 7347
rect 6052 7313 6064 7347
rect 6006 7287 6064 7313
rect 6106 7347 6164 7373
rect 6106 7313 6118 7347
rect 6152 7313 6164 7347
rect 6106 7287 6164 7313
rect 6206 7347 6264 7373
rect 6206 7313 6218 7347
rect 6252 7313 6264 7347
rect 6206 7287 6264 7313
rect 6306 7347 6364 7373
rect 6306 7313 6318 7347
rect 6352 7313 6364 7347
rect 6306 7287 6364 7313
rect 6406 7347 6464 7373
rect 6618 7366 6862 7400
rect 6406 7313 6418 7347
rect 6452 7313 6464 7347
rect 6508 7328 6516 7362
rect 6558 7328 6574 7362
rect 6618 7347 6652 7366
rect 6406 7287 6464 7313
rect 6828 7363 6862 7366
rect 6828 7347 6962 7363
rect 6618 7297 6652 7313
rect 6696 7298 6712 7332
rect 6754 7298 6762 7332
rect 6862 7313 6928 7347
rect 6828 7297 6962 7313
rect 7028 7347 7162 7363
rect 7062 7313 7128 7347
rect 7028 7297 7162 7313
rect 7228 7347 7362 7363
rect 7262 7313 7328 7347
rect 7228 7297 7362 7313
rect 7428 7347 7462 7363
rect 7428 7297 7462 7313
rect 6 7207 64 7233
rect 6 7173 18 7207
rect 52 7173 64 7207
rect 6 7147 64 7173
rect 106 7207 164 7233
rect 106 7173 118 7207
rect 152 7173 164 7207
rect 106 7147 164 7173
rect 206 7207 264 7233
rect 206 7173 218 7207
rect 252 7173 264 7207
rect 206 7147 264 7173
rect 306 7207 364 7233
rect 306 7173 312 7207
rect 352 7173 364 7207
rect 306 7147 364 7173
rect 406 7207 464 7233
rect 406 7173 418 7207
rect 458 7173 464 7207
rect 406 7147 464 7173
rect 506 7207 564 7233
rect 506 7173 518 7207
rect 552 7173 564 7207
rect 506 7147 564 7173
rect 606 7207 664 7233
rect 606 7173 618 7207
rect 652 7173 664 7207
rect 606 7147 664 7173
rect 706 7207 764 7233
rect 706 7173 718 7207
rect 752 7173 764 7207
rect 706 7147 764 7173
rect 806 7207 864 7233
rect 806 7173 818 7207
rect 852 7173 864 7207
rect 806 7147 864 7173
rect 906 7207 964 7233
rect 906 7173 918 7207
rect 952 7173 964 7207
rect 906 7147 964 7173
rect 1006 7207 1064 7233
rect 1006 7173 1018 7207
rect 1052 7173 1064 7207
rect 1006 7147 1064 7173
rect 1106 7207 1164 7233
rect 1106 7173 1118 7207
rect 1152 7173 1164 7207
rect 1106 7147 1164 7173
rect 1206 7207 1264 7233
rect 1206 7173 1218 7207
rect 1252 7173 1264 7207
rect 1206 7147 1264 7173
rect 1306 7207 1364 7233
rect 1306 7173 1318 7207
rect 1352 7173 1364 7207
rect 1306 7147 1364 7173
rect 1406 7207 1464 7233
rect 1406 7173 1418 7207
rect 1452 7173 1464 7207
rect 1406 7147 1464 7173
rect 1506 7207 1564 7233
rect 1506 7173 1518 7207
rect 1552 7173 1564 7207
rect 1506 7147 1564 7173
rect 1606 7207 1664 7233
rect 1606 7173 1618 7207
rect 1652 7173 1664 7207
rect 1606 7147 1664 7173
rect 1706 7207 1764 7233
rect 1706 7173 1718 7207
rect 1752 7173 1764 7207
rect 1706 7147 1764 7173
rect 1806 7207 1864 7233
rect 1806 7173 1818 7207
rect 1852 7173 1864 7207
rect 1806 7147 1864 7173
rect 1906 7207 1964 7233
rect 1906 7173 1918 7207
rect 1952 7173 1964 7207
rect 1906 7147 1964 7173
rect 2006 7207 2064 7233
rect 2006 7173 2018 7207
rect 2052 7173 2064 7207
rect 2006 7147 2064 7173
rect 2106 7207 2164 7233
rect 2106 7173 2118 7207
rect 2152 7173 2164 7207
rect 2106 7147 2164 7173
rect 2206 7207 2264 7233
rect 2206 7173 2218 7207
rect 2252 7173 2264 7207
rect 2206 7147 2264 7173
rect 2306 7207 2364 7233
rect 2306 7173 2318 7207
rect 2352 7173 2364 7207
rect 2306 7147 2364 7173
rect 2406 7207 2464 7233
rect 2406 7173 2418 7207
rect 2452 7173 2464 7207
rect 2406 7147 2464 7173
rect 2506 7207 2564 7233
rect 2506 7173 2512 7207
rect 2552 7173 2564 7207
rect 2506 7147 2564 7173
rect 2606 7207 2664 7233
rect 2606 7173 2618 7207
rect 2658 7173 2664 7207
rect 2606 7147 2664 7173
rect 2706 7207 2764 7233
rect 2706 7173 2718 7207
rect 2752 7173 2764 7207
rect 2706 7147 2764 7173
rect 2806 7207 2864 7233
rect 2806 7173 2818 7207
rect 2852 7173 2864 7207
rect 2806 7147 2864 7173
rect 2906 7207 2964 7233
rect 2906 7173 2912 7207
rect 2952 7173 2964 7207
rect 2906 7147 2964 7173
rect 3006 7207 3064 7233
rect 3006 7173 3018 7207
rect 3058 7173 3064 7207
rect 3006 7147 3064 7173
rect 3106 7207 3164 7233
rect 3106 7173 3118 7207
rect 3152 7173 3164 7207
rect 3106 7147 3164 7173
rect 3206 7207 3264 7233
rect 3206 7173 3212 7207
rect 3252 7173 3264 7207
rect 3206 7147 3264 7173
rect 3306 7207 3364 7233
rect 3306 7173 3318 7207
rect 3358 7173 3364 7207
rect 3306 7147 3364 7173
rect 3406 7207 3464 7233
rect 3406 7173 3418 7207
rect 3452 7173 3464 7207
rect 3406 7147 3464 7173
rect 3506 7207 3564 7233
rect 3506 7173 3518 7207
rect 3552 7173 3564 7207
rect 3506 7147 3564 7173
rect 3606 7207 3664 7233
rect 3606 7173 3618 7207
rect 3652 7173 3664 7207
rect 3606 7147 3664 7173
rect 3706 7207 3764 7233
rect 3706 7173 3718 7207
rect 3752 7173 3764 7207
rect 3706 7147 3764 7173
rect 3806 7207 3864 7233
rect 3806 7173 3818 7207
rect 3852 7173 3864 7207
rect 3806 7147 3864 7173
rect 3906 7207 3964 7233
rect 3906 7173 3918 7207
rect 3952 7173 3964 7207
rect 3906 7147 3964 7173
rect 4006 7207 4064 7233
rect 4006 7173 4018 7207
rect 4052 7173 4064 7207
rect 4006 7147 4064 7173
rect 4106 7207 4164 7233
rect 4106 7173 4118 7207
rect 4152 7173 4164 7207
rect 4106 7147 4164 7173
rect 4206 7207 4264 7233
rect 4206 7173 4218 7207
rect 4252 7173 4264 7207
rect 4206 7147 4264 7173
rect 4306 7207 4364 7233
rect 4306 7173 4312 7207
rect 4352 7173 4364 7207
rect 4306 7147 4364 7173
rect 4406 7207 4464 7233
rect 4406 7173 4418 7207
rect 4458 7173 4464 7207
rect 4406 7147 4464 7173
rect 4506 7207 4564 7233
rect 4506 7173 4518 7207
rect 4552 7173 4564 7207
rect 4506 7147 4564 7173
rect 4606 7207 4664 7233
rect 4606 7173 4612 7207
rect 4652 7173 4664 7207
rect 4606 7147 4664 7173
rect 4706 7207 4764 7233
rect 4706 7173 4718 7207
rect 4758 7173 4764 7207
rect 4706 7147 4764 7173
rect 4806 7207 4864 7233
rect 4806 7173 4818 7207
rect 4852 7173 4864 7207
rect 4806 7147 4864 7173
rect 4906 7207 4964 7233
rect 4906 7173 4918 7207
rect 4952 7173 4964 7207
rect 4906 7147 4964 7173
rect 5006 7207 5064 7233
rect 5006 7173 5012 7207
rect 5052 7173 5064 7207
rect 5006 7147 5064 7173
rect 5106 7207 5164 7233
rect 5106 7173 5118 7207
rect 5158 7173 5164 7207
rect 5106 7147 5164 7173
rect 5206 7207 5264 7233
rect 5206 7173 5218 7207
rect 5252 7173 5264 7207
rect 5206 7147 5264 7173
rect 5306 7207 5364 7233
rect 5306 7173 5318 7207
rect 5352 7173 5364 7207
rect 5306 7147 5364 7173
rect 5406 7207 5464 7233
rect 5406 7173 5418 7207
rect 5452 7173 5464 7207
rect 5406 7147 5464 7173
rect 5506 7207 5564 7233
rect 5506 7173 5518 7207
rect 5552 7173 5564 7207
rect 5506 7147 5564 7173
rect 5606 7207 5664 7233
rect 5606 7173 5618 7207
rect 5652 7173 5664 7207
rect 5606 7147 5664 7173
rect 5706 7207 5764 7233
rect 5706 7173 5718 7207
rect 5752 7173 5764 7207
rect 5706 7147 5764 7173
rect 5806 7207 5864 7233
rect 5806 7173 5818 7207
rect 5852 7173 5864 7207
rect 5806 7147 5864 7173
rect 5906 7207 5964 7233
rect 5906 7173 5918 7207
rect 5952 7173 5964 7207
rect 5906 7147 5964 7173
rect 6006 7207 6064 7233
rect 6006 7173 6012 7207
rect 6052 7173 6064 7207
rect 6006 7147 6064 7173
rect 6106 7207 6164 7233
rect 6106 7173 6118 7207
rect 6158 7173 6164 7207
rect 6106 7147 6164 7173
rect 6206 7207 6264 7233
rect 6206 7173 6218 7207
rect 6252 7173 6264 7207
rect 6206 7147 6264 7173
rect 6306 7207 6364 7233
rect 6306 7173 6318 7207
rect 6352 7173 6364 7207
rect 6306 7147 6364 7173
rect 6406 7207 6464 7233
rect 6618 7226 6862 7260
rect 6406 7173 6412 7207
rect 6452 7173 6464 7207
rect 6508 7188 6516 7222
rect 6558 7188 6574 7222
rect 6618 7207 6652 7226
rect 6406 7147 6464 7173
rect 6828 7207 6862 7226
rect 6618 7157 6652 7173
rect 6696 7158 6712 7192
rect 6754 7158 6762 7192
rect 6828 7157 6862 7173
rect 6928 7207 7162 7223
rect 6962 7173 7028 7207
rect 7062 7173 7128 7207
rect 6928 7157 7162 7173
rect 7228 7207 7362 7223
rect 7262 7173 7328 7207
rect 7228 7157 7362 7173
rect 7428 7207 7462 7223
rect 7428 7157 7462 7173
rect 6 7067 64 7093
rect 6 7033 18 7067
rect 58 7033 64 7067
rect 6 7007 64 7033
rect 106 7067 164 7093
rect 106 7033 118 7067
rect 152 7033 164 7067
rect 106 7007 164 7033
rect 206 7067 264 7093
rect 206 7033 218 7067
rect 252 7033 264 7067
rect 206 7007 264 7033
rect 306 7067 364 7093
rect 306 7033 312 7067
rect 352 7033 364 7067
rect 306 7007 364 7033
rect 406 7067 464 7093
rect 406 7033 418 7067
rect 458 7033 464 7067
rect 406 7007 464 7033
rect 506 7067 564 7093
rect 506 7033 518 7067
rect 552 7033 564 7067
rect 506 7007 564 7033
rect 606 7067 664 7093
rect 606 7033 618 7067
rect 652 7033 664 7067
rect 606 7007 664 7033
rect 706 7067 764 7093
rect 706 7033 718 7067
rect 752 7033 764 7067
rect 706 7007 764 7033
rect 806 7067 864 7093
rect 806 7033 818 7067
rect 852 7033 864 7067
rect 806 7007 864 7033
rect 906 7067 964 7093
rect 906 7033 918 7067
rect 952 7033 964 7067
rect 906 7007 964 7033
rect 1006 7067 1064 7093
rect 1006 7033 1018 7067
rect 1052 7033 1064 7067
rect 1006 7007 1064 7033
rect 1106 7067 1164 7093
rect 1106 7033 1118 7067
rect 1152 7033 1164 7067
rect 1106 7007 1164 7033
rect 1206 7067 1264 7093
rect 1206 7033 1212 7067
rect 1252 7033 1264 7067
rect 1206 7007 1264 7033
rect 1306 7067 1364 7093
rect 1306 7033 1318 7067
rect 1358 7033 1364 7067
rect 1306 7007 1364 7033
rect 1406 7067 1464 7093
rect 1406 7033 1418 7067
rect 1452 7033 1464 7067
rect 1406 7007 1464 7033
rect 1506 7067 1564 7093
rect 1506 7033 1518 7067
rect 1552 7033 1564 7067
rect 1506 7007 1564 7033
rect 1606 7067 1664 7093
rect 1606 7033 1618 7067
rect 1652 7033 1664 7067
rect 1606 7007 1664 7033
rect 1706 7067 1764 7093
rect 1706 7033 1718 7067
rect 1752 7033 1764 7067
rect 1706 7007 1764 7033
rect 1806 7067 1864 7093
rect 1806 7033 1818 7067
rect 1852 7033 1864 7067
rect 1806 7007 1864 7033
rect 1906 7067 1964 7093
rect 1906 7033 1918 7067
rect 1952 7033 1964 7067
rect 1906 7007 1964 7033
rect 2006 7067 2064 7093
rect 2006 7033 2018 7067
rect 2052 7033 2064 7067
rect 2006 7007 2064 7033
rect 2106 7067 2164 7093
rect 2106 7033 2118 7067
rect 2152 7033 2164 7067
rect 2106 7007 2164 7033
rect 2206 7067 2264 7093
rect 2206 7033 2212 7067
rect 2252 7033 2264 7067
rect 2206 7007 2264 7033
rect 2306 7067 2364 7093
rect 2306 7033 2318 7067
rect 2358 7033 2364 7067
rect 2306 7007 2364 7033
rect 2406 7067 2464 7093
rect 2406 7033 2418 7067
rect 2452 7033 2464 7067
rect 2406 7007 2464 7033
rect 2506 7067 2564 7093
rect 2506 7033 2518 7067
rect 2552 7033 2564 7067
rect 2506 7007 2564 7033
rect 2606 7067 2664 7093
rect 2606 7033 2618 7067
rect 2652 7033 2664 7067
rect 2606 7007 2664 7033
rect 2706 7067 2764 7093
rect 2706 7033 2718 7067
rect 2752 7033 2764 7067
rect 2706 7007 2764 7033
rect 2806 7067 2864 7093
rect 2806 7033 2818 7067
rect 2852 7033 2864 7067
rect 2806 7007 2864 7033
rect 2906 7067 2964 7093
rect 2906 7033 2918 7067
rect 2952 7033 2964 7067
rect 2906 7007 2964 7033
rect 3006 7067 3064 7093
rect 3006 7033 3012 7067
rect 3052 7033 3064 7067
rect 3006 7007 3064 7033
rect 3106 7067 3164 7093
rect 3106 7033 3118 7067
rect 3158 7033 3164 7067
rect 3106 7007 3164 7033
rect 3206 7067 3264 7093
rect 3206 7033 3218 7067
rect 3252 7033 3264 7067
rect 3206 7007 3264 7033
rect 3306 7067 3364 7093
rect 3306 7033 3318 7067
rect 3352 7033 3364 7067
rect 3306 7007 3364 7033
rect 3406 7067 3464 7093
rect 3406 7033 3412 7067
rect 3452 7033 3464 7067
rect 3406 7007 3464 7033
rect 3506 7067 3564 7093
rect 3506 7033 3518 7067
rect 3558 7033 3564 7067
rect 3506 7007 3564 7033
rect 3606 7067 3664 7093
rect 3606 7033 3618 7067
rect 3652 7033 3664 7067
rect 3606 7007 3664 7033
rect 3706 7067 3764 7093
rect 3706 7033 3718 7067
rect 3752 7033 3764 7067
rect 3706 7007 3764 7033
rect 3806 7067 3864 7093
rect 3806 7033 3818 7067
rect 3852 7033 3864 7067
rect 3806 7007 3864 7033
rect 3906 7067 3964 7093
rect 3906 7033 3918 7067
rect 3952 7033 3964 7067
rect 3906 7007 3964 7033
rect 4006 7067 4064 7093
rect 4006 7033 4012 7067
rect 4052 7033 4064 7067
rect 4006 7007 4064 7033
rect 4106 7067 4164 7093
rect 4106 7033 4118 7067
rect 4158 7033 4164 7067
rect 4106 7007 4164 7033
rect 4206 7067 4264 7093
rect 4206 7033 4218 7067
rect 4252 7033 4264 7067
rect 4206 7007 4264 7033
rect 4306 7067 4364 7093
rect 4306 7033 4318 7067
rect 4352 7033 4364 7067
rect 4306 7007 4364 7033
rect 4406 7067 4464 7093
rect 4406 7033 4418 7067
rect 4452 7033 4464 7067
rect 4406 7007 4464 7033
rect 4506 7067 4564 7093
rect 4506 7033 4518 7067
rect 4552 7033 4564 7067
rect 4506 7007 4564 7033
rect 4606 7067 4664 7093
rect 4606 7033 4618 7067
rect 4652 7033 4664 7067
rect 4606 7007 4664 7033
rect 4706 7067 4764 7093
rect 4706 7033 4718 7067
rect 4752 7033 4764 7067
rect 4706 7007 4764 7033
rect 4806 7067 4864 7093
rect 4806 7033 4818 7067
rect 4852 7033 4864 7067
rect 4806 7007 4864 7033
rect 4906 7067 4964 7093
rect 4906 7033 4918 7067
rect 4952 7033 4964 7067
rect 4906 7007 4964 7033
rect 5006 7067 5064 7093
rect 5006 7033 5018 7067
rect 5052 7033 5064 7067
rect 5006 7007 5064 7033
rect 5106 7067 5164 7093
rect 5106 7033 5112 7067
rect 5152 7033 5164 7067
rect 5106 7007 5164 7033
rect 5206 7067 5264 7093
rect 5206 7033 5218 7067
rect 5258 7033 5264 7067
rect 5206 7007 5264 7033
rect 5306 7067 5364 7093
rect 5306 7033 5318 7067
rect 5352 7033 5364 7067
rect 5306 7007 5364 7033
rect 5406 7067 5464 7093
rect 5406 7033 5418 7067
rect 5452 7033 5464 7067
rect 5406 7007 5464 7033
rect 5506 7067 5564 7093
rect 5506 7033 5518 7067
rect 5552 7033 5564 7067
rect 5506 7007 5564 7033
rect 5606 7067 5664 7093
rect 5606 7033 5618 7067
rect 5652 7033 5664 7067
rect 5606 7007 5664 7033
rect 5706 7067 5764 7093
rect 5706 7033 5718 7067
rect 5752 7033 5764 7067
rect 5706 7007 5764 7033
rect 5806 7067 5864 7093
rect 5806 7033 5818 7067
rect 5852 7033 5864 7067
rect 5806 7007 5864 7033
rect 5906 7067 5964 7093
rect 5906 7033 5918 7067
rect 5952 7033 5964 7067
rect 5906 7007 5964 7033
rect 6006 7067 6064 7093
rect 6006 7033 6018 7067
rect 6052 7033 6064 7067
rect 6006 7007 6064 7033
rect 6106 7067 6164 7093
rect 6106 7033 6112 7067
rect 6152 7033 6164 7067
rect 6106 7007 6164 7033
rect 6206 7067 6264 7093
rect 6206 7033 6218 7067
rect 6258 7033 6264 7067
rect 6206 7007 6264 7033
rect 6306 7067 6364 7093
rect 6306 7033 6318 7067
rect 6352 7033 6364 7067
rect 6306 7007 6364 7033
rect 6406 7067 6464 7093
rect 6618 7086 6862 7120
rect 6406 7033 6418 7067
rect 6452 7033 6464 7067
rect 6508 7048 6516 7082
rect 6558 7048 6574 7082
rect 6618 7067 6652 7086
rect 6406 7007 6464 7033
rect 6828 7083 6862 7086
rect 6828 7067 6962 7083
rect 6618 7017 6652 7033
rect 6696 7018 6712 7052
rect 6754 7018 6762 7052
rect 6862 7033 6928 7067
rect 6828 7017 6962 7033
rect 7028 7067 7062 7083
rect 7028 7017 7062 7033
rect 7128 7067 7362 7083
rect 7162 7033 7228 7067
rect 7262 7033 7328 7067
rect 7128 7017 7362 7033
rect 7428 7067 7462 7083
rect 7428 7017 7462 7033
rect 6 6927 64 6953
rect 6 6893 18 6927
rect 58 6893 64 6927
rect 6 6867 64 6893
rect 106 6927 164 6953
rect 106 6893 118 6927
rect 152 6893 164 6927
rect 106 6867 164 6893
rect 206 6927 264 6953
rect 206 6893 218 6927
rect 252 6893 264 6927
rect 206 6867 264 6893
rect 306 6927 364 6953
rect 306 6893 318 6927
rect 352 6893 364 6927
rect 306 6867 364 6893
rect 406 6927 464 6953
rect 406 6893 418 6927
rect 452 6893 464 6927
rect 406 6867 464 6893
rect 506 6927 564 6953
rect 506 6893 518 6927
rect 552 6893 564 6927
rect 506 6867 564 6893
rect 606 6927 664 6953
rect 606 6893 618 6927
rect 652 6893 664 6927
rect 606 6867 664 6893
rect 706 6927 764 6953
rect 706 6893 718 6927
rect 752 6893 764 6927
rect 706 6867 764 6893
rect 806 6927 864 6953
rect 806 6893 818 6927
rect 852 6893 864 6927
rect 806 6867 864 6893
rect 906 6927 964 6953
rect 906 6893 918 6927
rect 952 6893 964 6927
rect 906 6867 964 6893
rect 1006 6927 1064 6953
rect 1006 6893 1018 6927
rect 1052 6893 1064 6927
rect 1006 6867 1064 6893
rect 1106 6927 1164 6953
rect 1106 6893 1118 6927
rect 1152 6893 1164 6927
rect 1106 6867 1164 6893
rect 1206 6927 1264 6953
rect 1206 6893 1218 6927
rect 1252 6893 1264 6927
rect 1206 6867 1264 6893
rect 1306 6927 1364 6953
rect 1306 6893 1318 6927
rect 1352 6893 1364 6927
rect 1306 6867 1364 6893
rect 1406 6927 1464 6953
rect 1406 6893 1412 6927
rect 1452 6893 1464 6927
rect 1406 6867 1464 6893
rect 1506 6927 1564 6953
rect 1506 6893 1518 6927
rect 1558 6893 1564 6927
rect 1506 6867 1564 6893
rect 1606 6927 1664 6953
rect 1606 6893 1618 6927
rect 1652 6893 1664 6927
rect 1606 6867 1664 6893
rect 1706 6927 1764 6953
rect 1706 6893 1718 6927
rect 1752 6893 1764 6927
rect 1706 6867 1764 6893
rect 1806 6927 1864 6953
rect 1806 6893 1818 6927
rect 1852 6893 1864 6927
rect 1806 6867 1864 6893
rect 1906 6927 1964 6953
rect 1906 6893 1918 6927
rect 1952 6893 1964 6927
rect 1906 6867 1964 6893
rect 2006 6927 2064 6953
rect 2006 6893 2012 6927
rect 2052 6893 2064 6927
rect 2006 6867 2064 6893
rect 2106 6927 2164 6953
rect 2106 6893 2118 6927
rect 2158 6893 2164 6927
rect 2106 6867 2164 6893
rect 2206 6927 2264 6953
rect 2206 6893 2218 6927
rect 2252 6893 2264 6927
rect 2206 6867 2264 6893
rect 2306 6927 2364 6953
rect 2306 6893 2318 6927
rect 2352 6893 2364 6927
rect 2306 6867 2364 6893
rect 2406 6927 2464 6953
rect 2406 6893 2418 6927
rect 2452 6893 2464 6927
rect 2406 6867 2464 6893
rect 2506 6927 2564 6953
rect 2506 6893 2518 6927
rect 2552 6893 2564 6927
rect 2506 6867 2564 6893
rect 2606 6927 2664 6953
rect 2606 6893 2618 6927
rect 2652 6893 2664 6927
rect 2606 6867 2664 6893
rect 2706 6927 2764 6953
rect 2706 6893 2718 6927
rect 2752 6893 2764 6927
rect 2706 6867 2764 6893
rect 2806 6927 2864 6953
rect 2806 6893 2818 6927
rect 2852 6893 2864 6927
rect 2806 6867 2864 6893
rect 2906 6927 2964 6953
rect 2906 6893 2912 6927
rect 2952 6893 2964 6927
rect 2906 6867 2964 6893
rect 3006 6927 3064 6953
rect 3006 6893 3018 6927
rect 3058 6893 3064 6927
rect 3006 6867 3064 6893
rect 3106 6927 3164 6953
rect 3106 6893 3112 6927
rect 3152 6893 3164 6927
rect 3106 6867 3164 6893
rect 3206 6927 3264 6953
rect 3206 6893 3218 6927
rect 3258 6893 3264 6927
rect 3206 6867 3264 6893
rect 3306 6927 3364 6953
rect 3306 6893 3318 6927
rect 3352 6893 3364 6927
rect 3306 6867 3364 6893
rect 3406 6927 3464 6953
rect 3406 6893 3412 6927
rect 3452 6893 3464 6927
rect 3406 6867 3464 6893
rect 3506 6927 3564 6953
rect 3506 6893 3518 6927
rect 3558 6893 3564 6927
rect 3506 6867 3564 6893
rect 3606 6927 3664 6953
rect 3606 6893 3618 6927
rect 3652 6893 3664 6927
rect 3606 6867 3664 6893
rect 3706 6927 3764 6953
rect 3706 6893 3718 6927
rect 3752 6893 3764 6927
rect 3706 6867 3764 6893
rect 3806 6927 3864 6953
rect 3806 6893 3818 6927
rect 3852 6893 3864 6927
rect 3806 6867 3864 6893
rect 3906 6927 3964 6953
rect 3906 6893 3918 6927
rect 3952 6893 3964 6927
rect 3906 6867 3964 6893
rect 4006 6927 4064 6953
rect 4006 6893 4018 6927
rect 4052 6893 4064 6927
rect 4006 6867 4064 6893
rect 4106 6927 4164 6953
rect 4106 6893 4118 6927
rect 4152 6893 4164 6927
rect 4106 6867 4164 6893
rect 4206 6927 4264 6953
rect 4206 6893 4212 6927
rect 4252 6893 4264 6927
rect 4206 6867 4264 6893
rect 4306 6927 4364 6953
rect 4306 6893 4318 6927
rect 4358 6893 4364 6927
rect 4306 6867 4364 6893
rect 4406 6927 4464 6953
rect 4406 6893 4418 6927
rect 4452 6893 4464 6927
rect 4406 6867 4464 6893
rect 4506 6927 4564 6953
rect 4506 6893 4518 6927
rect 4552 6893 4564 6927
rect 4506 6867 4564 6893
rect 4606 6927 4664 6953
rect 4606 6893 4618 6927
rect 4652 6893 4664 6927
rect 4606 6867 4664 6893
rect 4706 6927 4764 6953
rect 4706 6893 4718 6927
rect 4752 6893 4764 6927
rect 4706 6867 4764 6893
rect 4806 6927 4864 6953
rect 4806 6893 4812 6927
rect 4852 6893 4864 6927
rect 4806 6867 4864 6893
rect 4906 6927 4964 6953
rect 4906 6893 4918 6927
rect 4958 6893 4964 6927
rect 4906 6867 4964 6893
rect 5006 6927 5064 6953
rect 5006 6893 5018 6927
rect 5052 6893 5064 6927
rect 5006 6867 5064 6893
rect 5106 6927 5164 6953
rect 5106 6893 5112 6927
rect 5152 6893 5164 6927
rect 5106 6867 5164 6893
rect 5206 6927 5264 6953
rect 5206 6893 5218 6927
rect 5258 6893 5264 6927
rect 5206 6867 5264 6893
rect 5306 6927 5364 6953
rect 5306 6893 5312 6927
rect 5352 6893 5364 6927
rect 5306 6867 5364 6893
rect 5406 6927 5464 6953
rect 5406 6893 5418 6927
rect 5458 6893 5464 6927
rect 5406 6867 5464 6893
rect 5506 6927 5564 6953
rect 5506 6893 5518 6927
rect 5552 6893 5564 6927
rect 5506 6867 5564 6893
rect 5606 6927 5664 6953
rect 5606 6893 5618 6927
rect 5652 6893 5664 6927
rect 5606 6867 5664 6893
rect 5706 6927 5764 6953
rect 5706 6893 5718 6927
rect 5752 6893 5764 6927
rect 5706 6867 5764 6893
rect 5806 6927 5864 6953
rect 5806 6893 5818 6927
rect 5852 6893 5864 6927
rect 5806 6867 5864 6893
rect 5906 6927 5964 6953
rect 5906 6893 5918 6927
rect 5952 6893 5964 6927
rect 5906 6867 5964 6893
rect 6006 6927 6064 6953
rect 6006 6893 6018 6927
rect 6052 6893 6064 6927
rect 6006 6867 6064 6893
rect 6106 6927 6164 6953
rect 6106 6893 6112 6927
rect 6152 6893 6164 6927
rect 6106 6867 6164 6893
rect 6206 6927 6264 6953
rect 6206 6893 6218 6927
rect 6258 6893 6264 6927
rect 6206 6867 6264 6893
rect 6306 6927 6364 6953
rect 6306 6893 6318 6927
rect 6352 6893 6364 6927
rect 6306 6867 6364 6893
rect 6406 6927 6464 6953
rect 6618 6946 6862 6980
rect 6406 6893 6418 6927
rect 6452 6893 6464 6927
rect 6508 6908 6516 6942
rect 6558 6908 6574 6942
rect 6618 6927 6652 6946
rect 6406 6867 6464 6893
rect 6828 6927 6862 6946
rect 6618 6877 6652 6893
rect 6696 6878 6712 6912
rect 6754 6878 6762 6912
rect 6828 6877 6862 6893
rect 6928 6927 7062 6943
rect 6962 6893 7028 6927
rect 6928 6877 7062 6893
rect 7128 6927 7362 6943
rect 7162 6893 7228 6927
rect 7262 6893 7328 6927
rect 7128 6877 7362 6893
rect 7428 6927 7462 6943
rect 7428 6877 7462 6893
rect 6 6787 64 6813
rect 6 6753 18 6787
rect 52 6753 64 6787
rect 6 6727 64 6753
rect 106 6787 164 6813
rect 106 6753 118 6787
rect 152 6753 164 6787
rect 106 6727 164 6753
rect 206 6787 264 6813
rect 206 6753 218 6787
rect 252 6753 264 6787
rect 206 6727 264 6753
rect 306 6787 364 6813
rect 306 6753 318 6787
rect 352 6753 364 6787
rect 306 6727 364 6753
rect 406 6787 464 6813
rect 406 6753 418 6787
rect 452 6753 464 6787
rect 406 6727 464 6753
rect 506 6787 564 6813
rect 506 6753 518 6787
rect 552 6753 564 6787
rect 506 6727 564 6753
rect 606 6787 664 6813
rect 606 6753 618 6787
rect 652 6753 664 6787
rect 606 6727 664 6753
rect 706 6787 764 6813
rect 706 6753 718 6787
rect 752 6753 764 6787
rect 706 6727 764 6753
rect 806 6787 864 6813
rect 806 6753 818 6787
rect 852 6753 864 6787
rect 806 6727 864 6753
rect 906 6787 964 6813
rect 906 6753 918 6787
rect 952 6753 964 6787
rect 906 6727 964 6753
rect 1006 6787 1064 6813
rect 1006 6753 1018 6787
rect 1052 6753 1064 6787
rect 1006 6727 1064 6753
rect 1106 6787 1164 6813
rect 1106 6753 1118 6787
rect 1152 6753 1164 6787
rect 1106 6727 1164 6753
rect 1206 6787 1264 6813
rect 1206 6753 1218 6787
rect 1252 6753 1264 6787
rect 1206 6727 1264 6753
rect 1306 6787 1364 6813
rect 1306 6753 1312 6787
rect 1352 6753 1364 6787
rect 1306 6727 1364 6753
rect 1406 6787 1464 6813
rect 1406 6753 1418 6787
rect 1458 6753 1464 6787
rect 1406 6727 1464 6753
rect 1506 6787 1564 6813
rect 1506 6753 1512 6787
rect 1552 6753 1564 6787
rect 1506 6727 1564 6753
rect 1606 6787 1664 6813
rect 1606 6753 1618 6787
rect 1658 6753 1664 6787
rect 1606 6727 1664 6753
rect 1706 6787 1764 6813
rect 1706 6753 1718 6787
rect 1752 6753 1764 6787
rect 1706 6727 1764 6753
rect 1806 6787 1864 6813
rect 1806 6753 1818 6787
rect 1852 6753 1864 6787
rect 1806 6727 1864 6753
rect 1906 6787 1964 6813
rect 1906 6753 1918 6787
rect 1952 6753 1964 6787
rect 1906 6727 1964 6753
rect 2006 6787 2064 6813
rect 2006 6753 2018 6787
rect 2052 6753 2064 6787
rect 2006 6727 2064 6753
rect 2106 6787 2164 6813
rect 2106 6753 2112 6787
rect 2152 6753 2164 6787
rect 2106 6727 2164 6753
rect 2206 6787 2264 6813
rect 2206 6753 2218 6787
rect 2258 6753 2264 6787
rect 2206 6727 2264 6753
rect 2306 6787 2364 6813
rect 2306 6753 2318 6787
rect 2352 6753 2364 6787
rect 2306 6727 2364 6753
rect 2406 6787 2464 6813
rect 2406 6753 2418 6787
rect 2452 6753 2464 6787
rect 2406 6727 2464 6753
rect 2506 6787 2564 6813
rect 2506 6753 2518 6787
rect 2552 6753 2564 6787
rect 2506 6727 2564 6753
rect 2606 6787 2664 6813
rect 2606 6753 2618 6787
rect 2652 6753 2664 6787
rect 2606 6727 2664 6753
rect 2706 6787 2764 6813
rect 2706 6753 2718 6787
rect 2752 6753 2764 6787
rect 2706 6727 2764 6753
rect 2806 6787 2864 6813
rect 2806 6753 2818 6787
rect 2852 6753 2864 6787
rect 2806 6727 2864 6753
rect 2906 6787 2964 6813
rect 2906 6753 2918 6787
rect 2952 6753 2964 6787
rect 2906 6727 2964 6753
rect 3006 6787 3064 6813
rect 3006 6753 3018 6787
rect 3052 6753 3064 6787
rect 3006 6727 3064 6753
rect 3106 6787 3164 6813
rect 3106 6753 3118 6787
rect 3152 6753 3164 6787
rect 3106 6727 3164 6753
rect 3206 6787 3264 6813
rect 3206 6753 3218 6787
rect 3252 6753 3264 6787
rect 3206 6727 3264 6753
rect 3306 6787 3364 6813
rect 3306 6753 3318 6787
rect 3352 6753 3364 6787
rect 3306 6727 3364 6753
rect 3406 6787 3464 6813
rect 3406 6753 3418 6787
rect 3452 6753 3464 6787
rect 3406 6727 3464 6753
rect 3506 6787 3564 6813
rect 3506 6753 3518 6787
rect 3552 6753 3564 6787
rect 3506 6727 3564 6753
rect 3606 6787 3664 6813
rect 3606 6753 3618 6787
rect 3652 6753 3664 6787
rect 3606 6727 3664 6753
rect 3706 6787 3764 6813
rect 3706 6753 3718 6787
rect 3752 6753 3764 6787
rect 3706 6727 3764 6753
rect 3806 6787 3864 6813
rect 3806 6753 3818 6787
rect 3852 6753 3864 6787
rect 3806 6727 3864 6753
rect 3906 6787 3964 6813
rect 3906 6753 3918 6787
rect 3952 6753 3964 6787
rect 3906 6727 3964 6753
rect 4006 6787 4064 6813
rect 4006 6753 4018 6787
rect 4052 6753 4064 6787
rect 4006 6727 4064 6753
rect 4106 6787 4164 6813
rect 4106 6753 4118 6787
rect 4152 6753 4164 6787
rect 4106 6727 4164 6753
rect 4206 6787 4264 6813
rect 4206 6753 4218 6787
rect 4252 6753 4264 6787
rect 4206 6727 4264 6753
rect 4306 6787 4364 6813
rect 4306 6753 4318 6787
rect 4352 6753 4364 6787
rect 4306 6727 4364 6753
rect 4406 6787 4464 6813
rect 4406 6753 4418 6787
rect 4452 6753 4464 6787
rect 4406 6727 4464 6753
rect 4506 6787 4564 6813
rect 4506 6753 4518 6787
rect 4552 6753 4564 6787
rect 4506 6727 4564 6753
rect 4606 6787 4664 6813
rect 4606 6753 4618 6787
rect 4652 6753 4664 6787
rect 4606 6727 4664 6753
rect 4706 6787 4764 6813
rect 4706 6753 4718 6787
rect 4752 6753 4764 6787
rect 4706 6727 4764 6753
rect 4806 6787 4864 6813
rect 4806 6753 4818 6787
rect 4852 6753 4864 6787
rect 4806 6727 4864 6753
rect 4906 6787 4964 6813
rect 4906 6753 4918 6787
rect 4952 6753 4964 6787
rect 4906 6727 4964 6753
rect 5006 6787 5064 6813
rect 5006 6753 5018 6787
rect 5052 6753 5064 6787
rect 5006 6727 5064 6753
rect 5106 6787 5164 6813
rect 5106 6753 5118 6787
rect 5152 6753 5164 6787
rect 5106 6727 5164 6753
rect 5206 6787 5264 6813
rect 5206 6753 5218 6787
rect 5252 6753 5264 6787
rect 5206 6727 5264 6753
rect 5306 6787 5364 6813
rect 5306 6753 5318 6787
rect 5352 6753 5364 6787
rect 5306 6727 5364 6753
rect 5406 6787 5464 6813
rect 5406 6753 5412 6787
rect 5452 6753 5464 6787
rect 5406 6727 5464 6753
rect 5506 6787 5564 6813
rect 5506 6753 5518 6787
rect 5558 6753 5564 6787
rect 5506 6727 5564 6753
rect 5606 6787 5664 6813
rect 5606 6753 5612 6787
rect 5652 6753 5664 6787
rect 5606 6727 5664 6753
rect 5706 6787 5764 6813
rect 5706 6753 5718 6787
rect 5758 6753 5764 6787
rect 5706 6727 5764 6753
rect 5806 6787 5864 6813
rect 5806 6753 5812 6787
rect 5852 6753 5864 6787
rect 5806 6727 5864 6753
rect 5906 6787 5964 6813
rect 5906 6753 5918 6787
rect 5958 6753 5964 6787
rect 5906 6727 5964 6753
rect 6006 6787 6064 6813
rect 6006 6753 6018 6787
rect 6052 6753 6064 6787
rect 6006 6727 6064 6753
rect 6106 6787 6164 6813
rect 6106 6753 6118 6787
rect 6152 6753 6164 6787
rect 6106 6727 6164 6753
rect 6206 6787 6264 6813
rect 6206 6753 6218 6787
rect 6252 6753 6264 6787
rect 6206 6727 6264 6753
rect 6306 6787 6364 6813
rect 6306 6753 6318 6787
rect 6352 6753 6364 6787
rect 6306 6727 6364 6753
rect 6406 6787 6464 6813
rect 6618 6806 6862 6840
rect 6406 6753 6418 6787
rect 6452 6753 6464 6787
rect 6508 6768 6516 6802
rect 6558 6768 6574 6802
rect 6618 6787 6652 6806
rect 6406 6727 6464 6753
rect 6828 6803 6862 6806
rect 6828 6787 6962 6803
rect 6618 6737 6652 6753
rect 6696 6738 6712 6772
rect 6754 6738 6762 6772
rect 6862 6753 6928 6787
rect 6828 6737 6962 6753
rect 7028 6787 7162 6803
rect 7062 6753 7128 6787
rect 7028 6737 7162 6753
rect 7228 6787 7262 6803
rect 7228 6737 7262 6753
rect 7328 6787 7462 6803
rect 7362 6753 7428 6787
rect 7328 6737 7462 6753
rect 6 6647 64 6673
rect 6 6613 18 6647
rect 58 6613 64 6647
rect 6 6587 64 6613
rect 106 6647 164 6673
rect 106 6613 118 6647
rect 152 6613 164 6647
rect 106 6587 164 6613
rect 206 6647 264 6673
rect 206 6613 212 6647
rect 252 6613 264 6647
rect 206 6587 264 6613
rect 306 6647 364 6673
rect 306 6613 318 6647
rect 358 6613 364 6647
rect 306 6587 364 6613
rect 406 6647 464 6673
rect 406 6613 418 6647
rect 452 6613 464 6647
rect 406 6587 464 6613
rect 506 6647 564 6673
rect 506 6613 518 6647
rect 552 6613 564 6647
rect 506 6587 564 6613
rect 606 6647 664 6673
rect 606 6613 618 6647
rect 652 6613 664 6647
rect 606 6587 664 6613
rect 706 6647 764 6673
rect 706 6613 718 6647
rect 752 6613 764 6647
rect 706 6587 764 6613
rect 806 6647 864 6673
rect 806 6613 818 6647
rect 852 6613 864 6647
rect 806 6587 864 6613
rect 906 6647 964 6673
rect 906 6613 918 6647
rect 952 6613 964 6647
rect 906 6587 964 6613
rect 1006 6647 1064 6673
rect 1006 6613 1012 6647
rect 1052 6613 1064 6647
rect 1006 6587 1064 6613
rect 1106 6647 1164 6673
rect 1106 6613 1118 6647
rect 1158 6613 1164 6647
rect 1106 6587 1164 6613
rect 1206 6647 1264 6673
rect 1206 6613 1212 6647
rect 1252 6613 1264 6647
rect 1206 6587 1264 6613
rect 1306 6647 1364 6673
rect 1306 6613 1318 6647
rect 1358 6613 1364 6647
rect 1306 6587 1364 6613
rect 1406 6647 1464 6673
rect 1406 6613 1418 6647
rect 1452 6613 1464 6647
rect 1406 6587 1464 6613
rect 1506 6647 1564 6673
rect 1506 6613 1518 6647
rect 1552 6613 1564 6647
rect 1506 6587 1564 6613
rect 1606 6647 1664 6673
rect 1606 6613 1618 6647
rect 1652 6613 1664 6647
rect 1606 6587 1664 6613
rect 1706 6647 1764 6673
rect 1706 6613 1718 6647
rect 1752 6613 1764 6647
rect 1706 6587 1764 6613
rect 1806 6647 1864 6673
rect 1806 6613 1818 6647
rect 1852 6613 1864 6647
rect 1806 6587 1864 6613
rect 1906 6647 1964 6673
rect 1906 6613 1918 6647
rect 1952 6613 1964 6647
rect 1906 6587 1964 6613
rect 2006 6647 2064 6673
rect 2006 6613 2018 6647
rect 2052 6613 2064 6647
rect 2006 6587 2064 6613
rect 2106 6647 2164 6673
rect 2106 6613 2118 6647
rect 2152 6613 2164 6647
rect 2106 6587 2164 6613
rect 2206 6647 2264 6673
rect 2206 6613 2218 6647
rect 2252 6613 2264 6647
rect 2206 6587 2264 6613
rect 2306 6647 2364 6673
rect 2306 6613 2318 6647
rect 2352 6613 2364 6647
rect 2306 6587 2364 6613
rect 2406 6647 2464 6673
rect 2406 6613 2418 6647
rect 2452 6613 2464 6647
rect 2406 6587 2464 6613
rect 2506 6647 2564 6673
rect 2506 6613 2518 6647
rect 2552 6613 2564 6647
rect 2506 6587 2564 6613
rect 2606 6647 2664 6673
rect 2606 6613 2618 6647
rect 2652 6613 2664 6647
rect 2606 6587 2664 6613
rect 2706 6647 2764 6673
rect 2706 6613 2718 6647
rect 2752 6613 2764 6647
rect 2706 6587 2764 6613
rect 2806 6647 2864 6673
rect 2806 6613 2818 6647
rect 2852 6613 2864 6647
rect 2806 6587 2864 6613
rect 2906 6647 2964 6673
rect 2906 6613 2918 6647
rect 2952 6613 2964 6647
rect 2906 6587 2964 6613
rect 3006 6647 3064 6673
rect 3006 6613 3018 6647
rect 3052 6613 3064 6647
rect 3006 6587 3064 6613
rect 3106 6647 3164 6673
rect 3106 6613 3118 6647
rect 3152 6613 3164 6647
rect 3106 6587 3164 6613
rect 3206 6647 3264 6673
rect 3206 6613 3218 6647
rect 3252 6613 3264 6647
rect 3206 6587 3264 6613
rect 3306 6647 3364 6673
rect 3306 6613 3318 6647
rect 3352 6613 3364 6647
rect 3306 6587 3364 6613
rect 3406 6647 3464 6673
rect 3406 6613 3412 6647
rect 3452 6613 3464 6647
rect 3406 6587 3464 6613
rect 3506 6647 3564 6673
rect 3506 6613 3518 6647
rect 3558 6613 3564 6647
rect 3506 6587 3564 6613
rect 3606 6647 3664 6673
rect 3606 6613 3612 6647
rect 3652 6613 3664 6647
rect 3606 6587 3664 6613
rect 3706 6647 3764 6673
rect 3706 6613 3718 6647
rect 3758 6613 3764 6647
rect 3706 6587 3764 6613
rect 3806 6647 3864 6673
rect 3806 6613 3818 6647
rect 3852 6613 3864 6647
rect 3806 6587 3864 6613
rect 3906 6647 3964 6673
rect 3906 6613 3918 6647
rect 3952 6613 3964 6647
rect 3906 6587 3964 6613
rect 4006 6647 4064 6673
rect 4006 6613 4018 6647
rect 4052 6613 4064 6647
rect 4006 6587 4064 6613
rect 4106 6647 4164 6673
rect 4106 6613 4118 6647
rect 4152 6613 4164 6647
rect 4106 6587 4164 6613
rect 4206 6647 4264 6673
rect 4206 6613 4218 6647
rect 4252 6613 4264 6647
rect 4206 6587 4264 6613
rect 4306 6647 4364 6673
rect 4306 6613 4318 6647
rect 4352 6613 4364 6647
rect 4306 6587 4364 6613
rect 4406 6647 4464 6673
rect 4406 6613 4412 6647
rect 4452 6613 4464 6647
rect 4406 6587 4464 6613
rect 4506 6647 4564 6673
rect 4506 6613 4518 6647
rect 4558 6613 4564 6647
rect 4506 6587 4564 6613
rect 4606 6647 4664 6673
rect 4606 6613 4618 6647
rect 4652 6613 4664 6647
rect 4606 6587 4664 6613
rect 4706 6647 4764 6673
rect 4706 6613 4718 6647
rect 4752 6613 4764 6647
rect 4706 6587 4764 6613
rect 4806 6647 4864 6673
rect 4806 6613 4818 6647
rect 4852 6613 4864 6647
rect 4806 6587 4864 6613
rect 4906 6647 4964 6673
rect 4906 6613 4918 6647
rect 4952 6613 4964 6647
rect 4906 6587 4964 6613
rect 5006 6647 5064 6673
rect 5006 6613 5018 6647
rect 5052 6613 5064 6647
rect 5006 6587 5064 6613
rect 5106 6647 5164 6673
rect 5106 6613 5118 6647
rect 5152 6613 5164 6647
rect 5106 6587 5164 6613
rect 5206 6647 5264 6673
rect 5206 6613 5218 6647
rect 5252 6613 5264 6647
rect 5206 6587 5264 6613
rect 5306 6647 5364 6673
rect 5306 6613 5318 6647
rect 5352 6613 5364 6647
rect 5306 6587 5364 6613
rect 5406 6647 5464 6673
rect 5406 6613 5418 6647
rect 5452 6613 5464 6647
rect 5406 6587 5464 6613
rect 5506 6647 5564 6673
rect 5506 6613 5518 6647
rect 5552 6613 5564 6647
rect 5506 6587 5564 6613
rect 5606 6647 5664 6673
rect 5606 6613 5618 6647
rect 5652 6613 5664 6647
rect 5606 6587 5664 6613
rect 5706 6647 5764 6673
rect 5706 6613 5718 6647
rect 5752 6613 5764 6647
rect 5706 6587 5764 6613
rect 5806 6647 5864 6673
rect 5806 6613 5812 6647
rect 5852 6613 5864 6647
rect 5806 6587 5864 6613
rect 5906 6647 5964 6673
rect 5906 6613 5918 6647
rect 5958 6613 5964 6647
rect 5906 6587 5964 6613
rect 6006 6647 6064 6673
rect 6006 6613 6018 6647
rect 6052 6613 6064 6647
rect 6006 6587 6064 6613
rect 6106 6647 6164 6673
rect 6106 6613 6118 6647
rect 6152 6613 6164 6647
rect 6106 6587 6164 6613
rect 6206 6647 6264 6673
rect 6206 6613 6218 6647
rect 6252 6613 6264 6647
rect 6206 6587 6264 6613
rect 6306 6647 6364 6673
rect 6306 6613 6318 6647
rect 6352 6613 6364 6647
rect 6306 6587 6364 6613
rect 6406 6647 6464 6673
rect 6618 6666 6862 6700
rect 6406 6613 6418 6647
rect 6452 6613 6464 6647
rect 6508 6628 6516 6662
rect 6558 6628 6574 6662
rect 6618 6647 6652 6666
rect 6406 6587 6464 6613
rect 6828 6647 6862 6666
rect 6618 6597 6652 6613
rect 6696 6598 6712 6632
rect 6754 6598 6762 6632
rect 6828 6597 6862 6613
rect 6928 6647 7162 6663
rect 6962 6613 7028 6647
rect 7062 6613 7128 6647
rect 6928 6597 7162 6613
rect 7228 6647 7262 6663
rect 7228 6597 7262 6613
rect 7328 6647 7462 6663
rect 7362 6613 7428 6647
rect 7328 6597 7462 6613
rect 6 6507 64 6533
rect 6 6473 18 6507
rect 52 6473 64 6507
rect 6 6447 64 6473
rect 106 6507 164 6533
rect 106 6473 118 6507
rect 152 6473 164 6507
rect 106 6447 164 6473
rect 206 6507 264 6533
rect 206 6473 218 6507
rect 252 6473 264 6507
rect 206 6447 264 6473
rect 306 6507 364 6533
rect 306 6473 318 6507
rect 352 6473 364 6507
rect 306 6447 364 6473
rect 406 6507 464 6533
rect 406 6473 418 6507
rect 452 6473 464 6507
rect 406 6447 464 6473
rect 506 6507 564 6533
rect 506 6473 512 6507
rect 552 6473 564 6507
rect 506 6447 564 6473
rect 606 6507 664 6533
rect 606 6473 618 6507
rect 658 6473 664 6507
rect 606 6447 664 6473
rect 706 6507 764 6533
rect 706 6473 718 6507
rect 752 6473 764 6507
rect 706 6447 764 6473
rect 806 6507 864 6533
rect 806 6473 818 6507
rect 852 6473 864 6507
rect 806 6447 864 6473
rect 906 6507 964 6533
rect 906 6473 918 6507
rect 952 6473 964 6507
rect 906 6447 964 6473
rect 1006 6507 1064 6533
rect 1006 6473 1018 6507
rect 1052 6473 1064 6507
rect 1006 6447 1064 6473
rect 1106 6507 1164 6533
rect 1106 6473 1118 6507
rect 1152 6473 1164 6507
rect 1106 6447 1164 6473
rect 1206 6507 1264 6533
rect 1206 6473 1218 6507
rect 1252 6473 1264 6507
rect 1206 6447 1264 6473
rect 1306 6507 1364 6533
rect 1306 6473 1318 6507
rect 1352 6473 1364 6507
rect 1306 6447 1364 6473
rect 1406 6507 1464 6533
rect 1406 6473 1418 6507
rect 1452 6473 1464 6507
rect 1406 6447 1464 6473
rect 1506 6507 1564 6533
rect 1506 6473 1518 6507
rect 1552 6473 1564 6507
rect 1506 6447 1564 6473
rect 1606 6507 1664 6533
rect 1606 6473 1612 6507
rect 1652 6473 1664 6507
rect 1606 6447 1664 6473
rect 1706 6507 1764 6533
rect 1706 6473 1718 6507
rect 1758 6473 1764 6507
rect 1706 6447 1764 6473
rect 1806 6507 1864 6533
rect 1806 6473 1818 6507
rect 1852 6473 1864 6507
rect 1806 6447 1864 6473
rect 1906 6507 1964 6533
rect 1906 6473 1918 6507
rect 1952 6473 1964 6507
rect 1906 6447 1964 6473
rect 2006 6507 2064 6533
rect 2006 6473 2018 6507
rect 2052 6473 2064 6507
rect 2006 6447 2064 6473
rect 2106 6507 2164 6533
rect 2106 6473 2118 6507
rect 2152 6473 2164 6507
rect 2106 6447 2164 6473
rect 2206 6507 2264 6533
rect 2206 6473 2218 6507
rect 2252 6473 2264 6507
rect 2206 6447 2264 6473
rect 2306 6507 2364 6533
rect 2306 6473 2318 6507
rect 2352 6473 2364 6507
rect 2306 6447 2364 6473
rect 2406 6507 2464 6533
rect 2406 6473 2418 6507
rect 2452 6473 2464 6507
rect 2406 6447 2464 6473
rect 2506 6507 2564 6533
rect 2506 6473 2518 6507
rect 2552 6473 2564 6507
rect 2506 6447 2564 6473
rect 2606 6507 2664 6533
rect 2606 6473 2618 6507
rect 2652 6473 2664 6507
rect 2606 6447 2664 6473
rect 2706 6507 2764 6533
rect 2706 6473 2718 6507
rect 2752 6473 2764 6507
rect 2706 6447 2764 6473
rect 2806 6507 2864 6533
rect 2806 6473 2818 6507
rect 2852 6473 2864 6507
rect 2806 6447 2864 6473
rect 2906 6507 2964 6533
rect 2906 6473 2918 6507
rect 2952 6473 2964 6507
rect 2906 6447 2964 6473
rect 3006 6507 3064 6533
rect 3006 6473 3018 6507
rect 3052 6473 3064 6507
rect 3006 6447 3064 6473
rect 3106 6507 3164 6533
rect 3106 6473 3118 6507
rect 3152 6473 3164 6507
rect 3106 6447 3164 6473
rect 3206 6507 3264 6533
rect 3206 6473 3218 6507
rect 3252 6473 3264 6507
rect 3206 6447 3264 6473
rect 3306 6507 3364 6533
rect 3306 6473 3318 6507
rect 3352 6473 3364 6507
rect 3306 6447 3364 6473
rect 3406 6507 3464 6533
rect 3406 6473 3418 6507
rect 3452 6473 3464 6507
rect 3406 6447 3464 6473
rect 3506 6507 3564 6533
rect 3506 6473 3518 6507
rect 3552 6473 3564 6507
rect 3506 6447 3564 6473
rect 3606 6507 3664 6533
rect 3606 6473 3618 6507
rect 3652 6473 3664 6507
rect 3606 6447 3664 6473
rect 3706 6507 3764 6533
rect 3706 6473 3712 6507
rect 3752 6473 3764 6507
rect 3706 6447 3764 6473
rect 3806 6507 3864 6533
rect 3806 6473 3818 6507
rect 3858 6473 3864 6507
rect 3806 6447 3864 6473
rect 3906 6507 3964 6533
rect 3906 6473 3918 6507
rect 3952 6473 3964 6507
rect 3906 6447 3964 6473
rect 4006 6507 4064 6533
rect 4006 6473 4018 6507
rect 4052 6473 4064 6507
rect 4006 6447 4064 6473
rect 4106 6507 4164 6533
rect 4106 6473 4118 6507
rect 4152 6473 4164 6507
rect 4106 6447 4164 6473
rect 4206 6507 4264 6533
rect 4206 6473 4218 6507
rect 4252 6473 4264 6507
rect 4206 6447 4264 6473
rect 4306 6507 4364 6533
rect 4306 6473 4318 6507
rect 4352 6473 4364 6507
rect 4306 6447 4364 6473
rect 4406 6507 4464 6533
rect 4406 6473 4418 6507
rect 4452 6473 4464 6507
rect 4406 6447 4464 6473
rect 4506 6507 4564 6533
rect 4506 6473 4518 6507
rect 4552 6473 4564 6507
rect 4506 6447 4564 6473
rect 4606 6507 4664 6533
rect 4606 6473 4618 6507
rect 4652 6473 4664 6507
rect 4606 6447 4664 6473
rect 4706 6507 4764 6533
rect 4706 6473 4718 6507
rect 4752 6473 4764 6507
rect 4706 6447 4764 6473
rect 4806 6507 4864 6533
rect 4806 6473 4818 6507
rect 4852 6473 4864 6507
rect 4806 6447 4864 6473
rect 4906 6507 4964 6533
rect 4906 6473 4918 6507
rect 4952 6473 4964 6507
rect 4906 6447 4964 6473
rect 5006 6507 5064 6533
rect 5006 6473 5018 6507
rect 5052 6473 5064 6507
rect 5006 6447 5064 6473
rect 5106 6507 5164 6533
rect 5106 6473 5112 6507
rect 5152 6473 5164 6507
rect 5106 6447 5164 6473
rect 5206 6507 5264 6533
rect 5206 6473 5218 6507
rect 5258 6473 5264 6507
rect 5206 6447 5264 6473
rect 5306 6507 5364 6533
rect 5306 6473 5312 6507
rect 5352 6473 5364 6507
rect 5306 6447 5364 6473
rect 5406 6507 5464 6533
rect 5406 6473 5418 6507
rect 5458 6473 5464 6507
rect 5406 6447 5464 6473
rect 5506 6507 5564 6533
rect 5506 6473 5518 6507
rect 5552 6473 5564 6507
rect 5506 6447 5564 6473
rect 5606 6507 5664 6533
rect 5606 6473 5618 6507
rect 5652 6473 5664 6507
rect 5606 6447 5664 6473
rect 5706 6507 5764 6533
rect 5706 6473 5718 6507
rect 5752 6473 5764 6507
rect 5706 6447 5764 6473
rect 5806 6507 5864 6533
rect 5806 6473 5818 6507
rect 5852 6473 5864 6507
rect 5806 6447 5864 6473
rect 5906 6507 5964 6533
rect 5906 6473 5918 6507
rect 5952 6473 5964 6507
rect 5906 6447 5964 6473
rect 6006 6507 6064 6533
rect 6006 6473 6018 6507
rect 6052 6473 6064 6507
rect 6006 6447 6064 6473
rect 6106 6507 6164 6533
rect 6106 6473 6118 6507
rect 6152 6473 6164 6507
rect 6106 6447 6164 6473
rect 6206 6507 6264 6533
rect 6206 6473 6218 6507
rect 6252 6473 6264 6507
rect 6206 6447 6264 6473
rect 6306 6507 6364 6533
rect 6306 6473 6318 6507
rect 6352 6473 6364 6507
rect 6306 6447 6364 6473
rect 6406 6507 6464 6533
rect 6618 6526 6862 6560
rect 6406 6473 6418 6507
rect 6452 6473 6464 6507
rect 6508 6488 6516 6522
rect 6558 6488 6574 6522
rect 6618 6507 6652 6526
rect 6406 6447 6464 6473
rect 6828 6523 6862 6526
rect 6828 6507 6962 6523
rect 6618 6457 6652 6473
rect 6696 6458 6712 6492
rect 6754 6458 6762 6492
rect 6862 6473 6928 6507
rect 6828 6457 6962 6473
rect 7028 6507 7062 6523
rect 7028 6457 7062 6473
rect 7128 6507 7262 6523
rect 7162 6473 7228 6507
rect 7128 6457 7262 6473
rect 7328 6507 7462 6523
rect 7362 6473 7428 6507
rect 7328 6457 7462 6473
rect 6 6367 64 6393
rect 6 6333 18 6367
rect 58 6333 64 6367
rect 6 6307 64 6333
rect 106 6367 164 6393
rect 106 6333 112 6367
rect 152 6333 164 6367
rect 106 6307 164 6333
rect 206 6367 264 6393
rect 206 6333 218 6367
rect 258 6333 264 6367
rect 206 6307 264 6333
rect 306 6367 364 6393
rect 306 6333 318 6367
rect 352 6333 364 6367
rect 306 6307 364 6333
rect 406 6367 464 6393
rect 406 6333 418 6367
rect 452 6333 464 6367
rect 406 6307 464 6333
rect 506 6367 564 6393
rect 506 6333 518 6367
rect 552 6333 564 6367
rect 506 6307 564 6333
rect 606 6367 664 6393
rect 606 6333 618 6367
rect 652 6333 664 6367
rect 606 6307 664 6333
rect 706 6367 764 6393
rect 706 6333 718 6367
rect 752 6333 764 6367
rect 706 6307 764 6333
rect 806 6367 864 6393
rect 806 6333 812 6367
rect 852 6333 864 6367
rect 806 6307 864 6333
rect 906 6367 964 6393
rect 906 6333 918 6367
rect 958 6333 964 6367
rect 906 6307 964 6333
rect 1006 6367 1064 6393
rect 1006 6333 1012 6367
rect 1052 6333 1064 6367
rect 1006 6307 1064 6333
rect 1106 6367 1164 6393
rect 1106 6333 1118 6367
rect 1158 6333 1164 6367
rect 1106 6307 1164 6333
rect 1206 6367 1264 6393
rect 1206 6333 1218 6367
rect 1252 6333 1264 6367
rect 1206 6307 1264 6333
rect 1306 6367 1364 6393
rect 1306 6333 1318 6367
rect 1352 6333 1364 6367
rect 1306 6307 1364 6333
rect 1406 6367 1464 6393
rect 1406 6333 1418 6367
rect 1452 6333 1464 6367
rect 1406 6307 1464 6333
rect 1506 6367 1564 6393
rect 1506 6333 1518 6367
rect 1552 6333 1564 6367
rect 1506 6307 1564 6333
rect 1606 6367 1664 6393
rect 1606 6333 1612 6367
rect 1652 6333 1664 6367
rect 1606 6307 1664 6333
rect 1706 6367 1764 6393
rect 1706 6333 1718 6367
rect 1758 6333 1764 6367
rect 1706 6307 1764 6333
rect 1806 6367 1864 6393
rect 1806 6333 1818 6367
rect 1852 6333 1864 6367
rect 1806 6307 1864 6333
rect 1906 6367 1964 6393
rect 1906 6333 1912 6367
rect 1952 6333 1964 6367
rect 1906 6307 1964 6333
rect 2006 6367 2064 6393
rect 2006 6333 2018 6367
rect 2058 6333 2064 6367
rect 2006 6307 2064 6333
rect 2106 6367 2164 6393
rect 2106 6333 2118 6367
rect 2152 6333 2164 6367
rect 2106 6307 2164 6333
rect 2206 6367 2264 6393
rect 2206 6333 2218 6367
rect 2252 6333 2264 6367
rect 2206 6307 2264 6333
rect 2306 6367 2364 6393
rect 2306 6333 2318 6367
rect 2352 6333 2364 6367
rect 2306 6307 2364 6333
rect 2406 6367 2464 6393
rect 2406 6333 2418 6367
rect 2452 6333 2464 6367
rect 2406 6307 2464 6333
rect 2506 6367 2564 6393
rect 2506 6333 2518 6367
rect 2552 6333 2564 6367
rect 2506 6307 2564 6333
rect 2606 6367 2664 6393
rect 2606 6333 2618 6367
rect 2652 6333 2664 6367
rect 2606 6307 2664 6333
rect 2706 6367 2764 6393
rect 2706 6333 2718 6367
rect 2752 6333 2764 6367
rect 2706 6307 2764 6333
rect 2806 6367 2864 6393
rect 2806 6333 2812 6367
rect 2852 6333 2864 6367
rect 2806 6307 2864 6333
rect 2906 6367 2964 6393
rect 2906 6333 2918 6367
rect 2958 6333 2964 6367
rect 2906 6307 2964 6333
rect 3006 6367 3064 6393
rect 3006 6333 3018 6367
rect 3052 6333 3064 6367
rect 3006 6307 3064 6333
rect 3106 6367 3164 6393
rect 3106 6333 3118 6367
rect 3152 6333 3164 6367
rect 3106 6307 3164 6333
rect 3206 6367 3264 6393
rect 3206 6333 3218 6367
rect 3252 6333 3264 6367
rect 3206 6307 3264 6333
rect 3306 6367 3364 6393
rect 3306 6333 3312 6367
rect 3352 6333 3364 6367
rect 3306 6307 3364 6333
rect 3406 6367 3464 6393
rect 3406 6333 3418 6367
rect 3458 6333 3464 6367
rect 3406 6307 3464 6333
rect 3506 6367 3564 6393
rect 3506 6333 3518 6367
rect 3552 6333 3564 6367
rect 3506 6307 3564 6333
rect 3606 6367 3664 6393
rect 3606 6333 3618 6367
rect 3652 6333 3664 6367
rect 3606 6307 3664 6333
rect 3706 6367 3764 6393
rect 3706 6333 3718 6367
rect 3752 6333 3764 6367
rect 3706 6307 3764 6333
rect 3806 6367 3864 6393
rect 3806 6333 3818 6367
rect 3852 6333 3864 6367
rect 3806 6307 3864 6333
rect 3906 6367 3964 6393
rect 3906 6333 3918 6367
rect 3952 6333 3964 6367
rect 3906 6307 3964 6333
rect 4006 6367 4064 6393
rect 4006 6333 4018 6367
rect 4052 6333 4064 6367
rect 4006 6307 4064 6333
rect 4106 6367 4164 6393
rect 4106 6333 4118 6367
rect 4152 6333 4164 6367
rect 4106 6307 4164 6333
rect 4206 6367 4264 6393
rect 4206 6333 4218 6367
rect 4252 6333 4264 6367
rect 4206 6307 4264 6333
rect 4306 6367 4364 6393
rect 4306 6333 4318 6367
rect 4352 6333 4364 6367
rect 4306 6307 4364 6333
rect 4406 6367 4464 6393
rect 4406 6333 4418 6367
rect 4452 6333 4464 6367
rect 4406 6307 4464 6333
rect 4506 6367 4564 6393
rect 4506 6333 4518 6367
rect 4552 6333 4564 6367
rect 4506 6307 4564 6333
rect 4606 6367 4664 6393
rect 4606 6333 4618 6367
rect 4652 6333 4664 6367
rect 4606 6307 4664 6333
rect 4706 6367 4764 6393
rect 4706 6333 4718 6367
rect 4752 6333 4764 6367
rect 4706 6307 4764 6333
rect 4806 6367 4864 6393
rect 4806 6333 4818 6367
rect 4852 6333 4864 6367
rect 4806 6307 4864 6333
rect 4906 6367 4964 6393
rect 4906 6333 4918 6367
rect 4952 6333 4964 6367
rect 4906 6307 4964 6333
rect 5006 6367 5064 6393
rect 5006 6333 5012 6367
rect 5052 6333 5064 6367
rect 5006 6307 5064 6333
rect 5106 6367 5164 6393
rect 5106 6333 5118 6367
rect 5158 6333 5164 6367
rect 5106 6307 5164 6333
rect 5206 6367 5264 6393
rect 5206 6333 5218 6367
rect 5252 6333 5264 6367
rect 5206 6307 5264 6333
rect 5306 6367 5364 6393
rect 5306 6333 5312 6367
rect 5352 6333 5364 6367
rect 5306 6307 5364 6333
rect 5406 6367 5464 6393
rect 5406 6333 5418 6367
rect 5458 6333 5464 6367
rect 5406 6307 5464 6333
rect 5506 6367 5564 6393
rect 5506 6333 5518 6367
rect 5552 6333 5564 6367
rect 5506 6307 5564 6333
rect 5606 6367 5664 6393
rect 5606 6333 5618 6367
rect 5652 6333 5664 6367
rect 5606 6307 5664 6333
rect 5706 6367 5764 6393
rect 5706 6333 5718 6367
rect 5752 6333 5764 6367
rect 5706 6307 5764 6333
rect 5806 6367 5864 6393
rect 5806 6333 5818 6367
rect 5852 6333 5864 6367
rect 5806 6307 5864 6333
rect 5906 6367 5964 6393
rect 5906 6333 5918 6367
rect 5952 6333 5964 6367
rect 5906 6307 5964 6333
rect 6006 6367 6064 6393
rect 6006 6333 6018 6367
rect 6052 6333 6064 6367
rect 6006 6307 6064 6333
rect 6106 6367 6164 6393
rect 6106 6333 6112 6367
rect 6152 6333 6164 6367
rect 6106 6307 6164 6333
rect 6206 6367 6264 6393
rect 6206 6333 6218 6367
rect 6258 6333 6264 6367
rect 6206 6307 6264 6333
rect 6306 6367 6364 6393
rect 6306 6333 6318 6367
rect 6352 6333 6364 6367
rect 6306 6307 6364 6333
rect 6406 6367 6464 6393
rect 6618 6386 6862 6420
rect 6406 6333 6412 6367
rect 6452 6333 6464 6367
rect 6508 6348 6516 6382
rect 6558 6348 6574 6382
rect 6618 6367 6652 6386
rect 6406 6307 6464 6333
rect 6828 6367 6862 6386
rect 6618 6317 6652 6333
rect 6696 6318 6712 6352
rect 6754 6318 6762 6352
rect 6828 6317 6862 6333
rect 6928 6367 7062 6383
rect 6962 6333 7028 6367
rect 6928 6317 7062 6333
rect 7128 6367 7262 6383
rect 7162 6333 7228 6367
rect 7128 6317 7262 6333
rect 7328 6367 7462 6383
rect 7362 6333 7428 6367
rect 7328 6317 7462 6333
rect 8 6210 18 6244
rect 52 6210 118 6244
rect 152 6210 168 6244
rect 208 6226 218 6260
rect 252 6226 318 6260
rect 352 6226 368 6260
rect 408 6210 418 6244
rect 452 6210 518 6244
rect 552 6210 568 6244
rect 608 6226 618 6260
rect 652 6226 718 6260
rect 752 6226 768 6260
rect 808 6210 818 6244
rect 852 6210 918 6244
rect 952 6210 968 6244
rect 1008 6226 1018 6260
rect 1052 6226 1118 6260
rect 1152 6226 1168 6260
rect 1208 6210 1218 6244
rect 1252 6210 1318 6244
rect 1352 6210 1368 6244
rect 1408 6226 1418 6260
rect 1452 6226 1518 6260
rect 1552 6226 1568 6260
rect 1608 6210 1618 6244
rect 1652 6210 1718 6244
rect 1752 6210 1768 6244
rect 1808 6226 1818 6260
rect 1852 6226 1918 6260
rect 1952 6226 1968 6260
rect 2008 6210 2018 6244
rect 2052 6210 2118 6244
rect 2152 6210 2168 6244
rect 2208 6226 2218 6260
rect 2252 6226 2318 6260
rect 2352 6226 2368 6260
rect 2408 6210 2418 6244
rect 2452 6210 2518 6244
rect 2552 6210 2568 6244
rect 2608 6226 2618 6260
rect 2652 6226 2718 6260
rect 2752 6226 2768 6260
rect 2808 6210 2818 6244
rect 2852 6210 2918 6244
rect 2952 6210 2968 6244
rect 3008 6226 3018 6260
rect 3052 6226 3118 6260
rect 3152 6226 3168 6260
rect 3208 6210 3218 6244
rect 3252 6210 3318 6244
rect 3352 6210 3368 6244
rect 3408 6226 3418 6260
rect 3452 6226 3518 6260
rect 3552 6226 3568 6260
rect 3608 6210 3618 6244
rect 3652 6210 3718 6244
rect 3752 6210 3768 6244
rect 3808 6226 3818 6260
rect 3852 6226 3918 6260
rect 3952 6226 3968 6260
rect 4008 6210 4018 6244
rect 4052 6210 4118 6244
rect 4152 6210 4168 6244
rect 4208 6226 4218 6260
rect 4252 6226 4318 6260
rect 4352 6226 4368 6260
rect 4408 6210 4418 6244
rect 4452 6210 4518 6244
rect 4552 6210 4568 6244
rect 4608 6226 4618 6260
rect 4652 6226 4718 6260
rect 4752 6226 4768 6260
rect 4808 6210 4818 6244
rect 4852 6210 4918 6244
rect 4952 6210 4968 6244
rect 5008 6226 5018 6260
rect 5052 6226 5118 6260
rect 5152 6226 5168 6260
rect 5208 6210 5218 6244
rect 5252 6210 5318 6244
rect 5352 6210 5368 6244
rect 5408 6226 5418 6260
rect 5452 6226 5518 6260
rect 5552 6226 5568 6260
rect 5608 6210 5618 6244
rect 5652 6210 5718 6244
rect 5752 6210 5768 6244
rect 5808 6226 5818 6260
rect 5852 6226 5918 6260
rect 5952 6226 5968 6260
rect 6008 6210 6018 6244
rect 6052 6210 6118 6244
rect 6152 6210 6168 6244
rect 6208 6226 6218 6260
rect 6252 6226 6318 6260
rect 6352 6226 6368 6260
rect 6516 6241 6568 6258
rect 6550 6224 6568 6241
rect 6602 6224 6618 6258
rect 6652 6224 6668 6258
rect 6702 6229 6720 6258
rect 6702 6224 6754 6229
rect 6862 6224 6878 6258
rect 6912 6224 6928 6258
rect 6962 6224 6978 6258
rect 7012 6224 7028 6258
rect 7062 6224 7078 6258
rect 7112 6224 7128 6258
rect 7162 6224 7178 6258
rect 7212 6224 7228 6258
rect 7262 6224 7278 6258
rect 7312 6224 7328 6258
rect 7362 6224 7378 6258
rect 7412 6224 7428 6258
rect 6 6137 64 6163
rect 6 6103 18 6137
rect 52 6103 64 6137
rect 6 6077 64 6103
rect 106 6137 164 6163
rect 106 6103 118 6137
rect 152 6103 164 6137
rect 106 6077 164 6103
rect 206 6137 264 6163
rect 206 6103 218 6137
rect 252 6103 264 6137
rect 206 6077 264 6103
rect 306 6137 364 6163
rect 306 6103 318 6137
rect 352 6103 364 6137
rect 306 6077 364 6103
rect 406 6137 464 6163
rect 406 6103 418 6137
rect 452 6103 464 6137
rect 406 6077 464 6103
rect 506 6137 564 6163
rect 506 6103 518 6137
rect 552 6103 564 6137
rect 506 6077 564 6103
rect 606 6137 664 6163
rect 606 6103 618 6137
rect 652 6103 664 6137
rect 606 6077 664 6103
rect 706 6137 764 6163
rect 706 6103 718 6137
rect 752 6103 764 6137
rect 706 6077 764 6103
rect 806 6137 864 6163
rect 806 6103 818 6137
rect 852 6103 864 6137
rect 806 6077 864 6103
rect 906 6137 964 6163
rect 906 6103 918 6137
rect 952 6103 964 6137
rect 906 6077 964 6103
rect 1006 6137 1064 6163
rect 1006 6103 1018 6137
rect 1052 6103 1064 6137
rect 1006 6077 1064 6103
rect 1106 6137 1164 6163
rect 1106 6103 1118 6137
rect 1152 6103 1164 6137
rect 1106 6077 1164 6103
rect 1206 6137 1264 6163
rect 1206 6103 1218 6137
rect 1252 6103 1264 6137
rect 1206 6077 1264 6103
rect 1306 6137 1364 6163
rect 1306 6103 1318 6137
rect 1352 6103 1364 6137
rect 1306 6077 1364 6103
rect 1406 6137 1464 6163
rect 1406 6103 1418 6137
rect 1452 6103 1464 6137
rect 1406 6077 1464 6103
rect 1506 6137 1564 6163
rect 1506 6103 1518 6137
rect 1552 6103 1564 6137
rect 1506 6077 1564 6103
rect 1606 6137 1664 6163
rect 1606 6103 1618 6137
rect 1652 6103 1664 6137
rect 1606 6077 1664 6103
rect 1706 6137 1764 6163
rect 1706 6103 1718 6137
rect 1752 6103 1764 6137
rect 1706 6077 1764 6103
rect 1806 6137 1864 6163
rect 1806 6103 1818 6137
rect 1852 6103 1864 6137
rect 1806 6077 1864 6103
rect 1906 6137 1964 6163
rect 1906 6103 1918 6137
rect 1952 6103 1964 6137
rect 1906 6077 1964 6103
rect 2006 6137 2064 6163
rect 2006 6103 2018 6137
rect 2052 6103 2064 6137
rect 2006 6077 2064 6103
rect 2106 6137 2164 6163
rect 2106 6103 2118 6137
rect 2152 6103 2164 6137
rect 2106 6077 2164 6103
rect 2206 6137 2264 6163
rect 2206 6103 2218 6137
rect 2252 6103 2264 6137
rect 2206 6077 2264 6103
rect 2306 6137 2364 6163
rect 2306 6103 2318 6137
rect 2352 6103 2364 6137
rect 2306 6077 2364 6103
rect 2406 6137 2464 6163
rect 2406 6103 2412 6137
rect 2452 6103 2464 6137
rect 2406 6077 2464 6103
rect 2506 6137 2564 6163
rect 2506 6103 2518 6137
rect 2558 6103 2564 6137
rect 2506 6077 2564 6103
rect 2606 6137 2664 6163
rect 2606 6103 2618 6137
rect 2652 6103 2664 6137
rect 2606 6077 2664 6103
rect 2706 6137 2764 6163
rect 2706 6103 2718 6137
rect 2752 6103 2764 6137
rect 2706 6077 2764 6103
rect 2806 6137 2864 6163
rect 2806 6103 2818 6137
rect 2852 6103 2864 6137
rect 2806 6077 2864 6103
rect 2906 6137 2964 6163
rect 2906 6103 2918 6137
rect 2952 6103 2964 6137
rect 2906 6077 2964 6103
rect 3006 6137 3064 6163
rect 3006 6103 3018 6137
rect 3052 6103 3064 6137
rect 3006 6077 3064 6103
rect 3106 6137 3164 6163
rect 3106 6103 3118 6137
rect 3152 6103 3164 6137
rect 3106 6077 3164 6103
rect 3206 6137 3264 6163
rect 3206 6103 3218 6137
rect 3252 6103 3264 6137
rect 3206 6077 3264 6103
rect 3306 6137 3364 6163
rect 3306 6103 3318 6137
rect 3352 6103 3364 6137
rect 3306 6077 3364 6103
rect 3406 6137 3464 6163
rect 3406 6103 3418 6137
rect 3452 6103 3464 6137
rect 3406 6077 3464 6103
rect 3506 6137 3564 6163
rect 3506 6103 3518 6137
rect 3552 6103 3564 6137
rect 3506 6077 3564 6103
rect 3606 6137 3664 6163
rect 3606 6103 3618 6137
rect 3652 6103 3664 6137
rect 3606 6077 3664 6103
rect 3706 6137 3764 6163
rect 3706 6103 3712 6137
rect 3752 6103 3764 6137
rect 3706 6077 3764 6103
rect 3806 6137 3864 6163
rect 3806 6103 3818 6137
rect 3858 6103 3864 6137
rect 3806 6077 3864 6103
rect 3906 6137 3964 6163
rect 3906 6103 3918 6137
rect 3952 6103 3964 6137
rect 3906 6077 3964 6103
rect 4006 6137 4064 6163
rect 4006 6103 4012 6137
rect 4052 6103 4064 6137
rect 4006 6077 4064 6103
rect 4106 6137 4164 6163
rect 4106 6103 4118 6137
rect 4158 6103 4164 6137
rect 4106 6077 4164 6103
rect 4206 6137 4264 6163
rect 4206 6103 4218 6137
rect 4252 6103 4264 6137
rect 4206 6077 4264 6103
rect 4306 6137 4364 6163
rect 4306 6103 4318 6137
rect 4352 6103 4364 6137
rect 4306 6077 4364 6103
rect 4406 6137 4464 6163
rect 4406 6103 4412 6137
rect 4452 6103 4464 6137
rect 4406 6077 4464 6103
rect 4506 6137 4564 6163
rect 4506 6103 4518 6137
rect 4558 6103 4564 6137
rect 4506 6077 4564 6103
rect 4606 6137 4664 6163
rect 4606 6103 4612 6137
rect 4652 6103 4664 6137
rect 4606 6077 4664 6103
rect 4706 6137 4764 6163
rect 4706 6103 4718 6137
rect 4758 6103 4764 6137
rect 4706 6077 4764 6103
rect 4806 6137 4864 6163
rect 4806 6103 4818 6137
rect 4852 6103 4864 6137
rect 4806 6077 4864 6103
rect 4906 6137 4964 6163
rect 4906 6103 4918 6137
rect 4952 6103 4964 6137
rect 4906 6077 4964 6103
rect 5006 6137 5064 6163
rect 5006 6103 5018 6137
rect 5052 6103 5064 6137
rect 5006 6077 5064 6103
rect 5106 6137 5164 6163
rect 5106 6103 5118 6137
rect 5152 6103 5164 6137
rect 5106 6077 5164 6103
rect 5206 6137 5264 6163
rect 5206 6103 5218 6137
rect 5252 6103 5264 6137
rect 5206 6077 5264 6103
rect 5306 6137 5364 6163
rect 5306 6103 5318 6137
rect 5352 6103 5364 6137
rect 5306 6077 5364 6103
rect 5406 6137 5464 6163
rect 5406 6103 5418 6137
rect 5452 6103 5464 6137
rect 5406 6077 5464 6103
rect 5506 6137 5564 6163
rect 5506 6103 5518 6137
rect 5552 6103 5564 6137
rect 5506 6077 5564 6103
rect 5606 6137 5664 6163
rect 5606 6103 5618 6137
rect 5652 6103 5664 6137
rect 5606 6077 5664 6103
rect 5706 6137 5764 6163
rect 5706 6103 5718 6137
rect 5752 6103 5764 6137
rect 5706 6077 5764 6103
rect 5806 6137 5864 6163
rect 5806 6103 5818 6137
rect 5852 6103 5864 6137
rect 5806 6077 5864 6103
rect 5906 6137 5964 6163
rect 5906 6103 5918 6137
rect 5952 6103 5964 6137
rect 5906 6077 5964 6103
rect 6006 6137 6064 6163
rect 6006 6103 6012 6137
rect 6052 6103 6064 6137
rect 6006 6077 6064 6103
rect 6106 6137 6164 6163
rect 6106 6103 6118 6137
rect 6158 6103 6164 6137
rect 6106 6077 6164 6103
rect 6206 6137 6264 6163
rect 6206 6103 6212 6137
rect 6252 6103 6264 6137
rect 6206 6077 6264 6103
rect 6306 6137 6364 6163
rect 6306 6103 6318 6137
rect 6358 6103 6364 6137
rect 6306 6077 6364 6103
rect 6406 6137 6464 6163
rect 6618 6156 6862 6190
rect 6406 6103 6412 6137
rect 6452 6103 6464 6137
rect 6508 6118 6516 6152
rect 6558 6118 6574 6152
rect 6618 6137 6652 6156
rect 6406 6077 6464 6103
rect 6828 6153 6862 6156
rect 6828 6137 6962 6153
rect 6618 6087 6652 6103
rect 6696 6088 6712 6122
rect 6754 6088 6762 6122
rect 6862 6103 6928 6137
rect 6828 6087 6962 6103
rect 7028 6137 7162 6153
rect 7062 6103 7128 6137
rect 7028 6087 7162 6103
rect 7228 6137 7362 6153
rect 7262 6103 7328 6137
rect 7228 6087 7362 6103
rect 7428 6137 7462 6153
rect 7428 6087 7462 6103
rect 6 5997 64 6023
rect 6 5963 18 5997
rect 52 5963 64 5997
rect 6 5937 64 5963
rect 106 5997 164 6023
rect 106 5963 118 5997
rect 152 5963 164 5997
rect 106 5937 164 5963
rect 206 5997 264 6023
rect 206 5963 218 5997
rect 252 5963 264 5997
rect 206 5937 264 5963
rect 306 5997 364 6023
rect 306 5963 318 5997
rect 352 5963 364 5997
rect 306 5937 364 5963
rect 406 5997 464 6023
rect 406 5963 412 5997
rect 452 5963 464 5997
rect 406 5937 464 5963
rect 506 5997 564 6023
rect 506 5963 518 5997
rect 558 5963 564 5997
rect 506 5937 564 5963
rect 606 5997 664 6023
rect 606 5963 618 5997
rect 652 5963 664 5997
rect 606 5937 664 5963
rect 706 5997 764 6023
rect 706 5963 718 5997
rect 752 5963 764 5997
rect 706 5937 764 5963
rect 806 5997 864 6023
rect 806 5963 818 5997
rect 852 5963 864 5997
rect 806 5937 864 5963
rect 906 5997 964 6023
rect 906 5963 918 5997
rect 952 5963 964 5997
rect 906 5937 964 5963
rect 1006 5997 1064 6023
rect 1006 5963 1018 5997
rect 1052 5963 1064 5997
rect 1006 5937 1064 5963
rect 1106 5997 1164 6023
rect 1106 5963 1118 5997
rect 1152 5963 1164 5997
rect 1106 5937 1164 5963
rect 1206 5997 1264 6023
rect 1206 5963 1218 5997
rect 1252 5963 1264 5997
rect 1206 5937 1264 5963
rect 1306 5997 1364 6023
rect 1306 5963 1312 5997
rect 1352 5963 1364 5997
rect 1306 5937 1364 5963
rect 1406 5997 1464 6023
rect 1406 5963 1418 5997
rect 1458 5963 1464 5997
rect 1406 5937 1464 5963
rect 1506 5997 1564 6023
rect 1506 5963 1518 5997
rect 1552 5963 1564 5997
rect 1506 5937 1564 5963
rect 1606 5997 1664 6023
rect 1606 5963 1618 5997
rect 1652 5963 1664 5997
rect 1606 5937 1664 5963
rect 1706 5997 1764 6023
rect 1706 5963 1718 5997
rect 1752 5963 1764 5997
rect 1706 5937 1764 5963
rect 1806 5997 1864 6023
rect 1806 5963 1818 5997
rect 1852 5963 1864 5997
rect 1806 5937 1864 5963
rect 1906 5997 1964 6023
rect 1906 5963 1918 5997
rect 1952 5963 1964 5997
rect 1906 5937 1964 5963
rect 2006 5997 2064 6023
rect 2006 5963 2018 5997
rect 2052 5963 2064 5997
rect 2006 5937 2064 5963
rect 2106 5997 2164 6023
rect 2106 5963 2118 5997
rect 2152 5963 2164 5997
rect 2106 5937 2164 5963
rect 2206 5997 2264 6023
rect 2206 5963 2218 5997
rect 2252 5963 2264 5997
rect 2206 5937 2264 5963
rect 2306 5997 2364 6023
rect 2306 5963 2318 5997
rect 2352 5963 2364 5997
rect 2306 5937 2364 5963
rect 2406 5997 2464 6023
rect 2406 5963 2418 5997
rect 2452 5963 2464 5997
rect 2406 5937 2464 5963
rect 2506 5997 2564 6023
rect 2506 5963 2518 5997
rect 2552 5963 2564 5997
rect 2506 5937 2564 5963
rect 2606 5997 2664 6023
rect 2606 5963 2618 5997
rect 2652 5963 2664 5997
rect 2606 5937 2664 5963
rect 2706 5997 2764 6023
rect 2706 5963 2718 5997
rect 2752 5963 2764 5997
rect 2706 5937 2764 5963
rect 2806 5997 2864 6023
rect 2806 5963 2818 5997
rect 2852 5963 2864 5997
rect 2806 5937 2864 5963
rect 2906 5997 2964 6023
rect 2906 5963 2918 5997
rect 2952 5963 2964 5997
rect 2906 5937 2964 5963
rect 3006 5997 3064 6023
rect 3006 5963 3018 5997
rect 3052 5963 3064 5997
rect 3006 5937 3064 5963
rect 3106 5997 3164 6023
rect 3106 5963 3118 5997
rect 3152 5963 3164 5997
rect 3106 5937 3164 5963
rect 3206 5997 3264 6023
rect 3206 5963 3218 5997
rect 3252 5963 3264 5997
rect 3206 5937 3264 5963
rect 3306 5997 3364 6023
rect 3306 5963 3312 5997
rect 3352 5963 3364 5997
rect 3306 5937 3364 5963
rect 3406 5997 3464 6023
rect 3406 5963 3418 5997
rect 3458 5963 3464 5997
rect 3406 5937 3464 5963
rect 3506 5997 3564 6023
rect 3506 5963 3518 5997
rect 3552 5963 3564 5997
rect 3506 5937 3564 5963
rect 3606 5997 3664 6023
rect 3606 5963 3618 5997
rect 3652 5963 3664 5997
rect 3606 5937 3664 5963
rect 3706 5997 3764 6023
rect 3706 5963 3718 5997
rect 3752 5963 3764 5997
rect 3706 5937 3764 5963
rect 3806 5997 3864 6023
rect 3806 5963 3818 5997
rect 3852 5963 3864 5997
rect 3806 5937 3864 5963
rect 3906 5997 3964 6023
rect 3906 5963 3918 5997
rect 3952 5963 3964 5997
rect 3906 5937 3964 5963
rect 4006 5997 4064 6023
rect 4006 5963 4018 5997
rect 4052 5963 4064 5997
rect 4006 5937 4064 5963
rect 4106 5997 4164 6023
rect 4106 5963 4118 5997
rect 4152 5963 4164 5997
rect 4106 5937 4164 5963
rect 4206 5997 4264 6023
rect 4206 5963 4218 5997
rect 4252 5963 4264 5997
rect 4206 5937 4264 5963
rect 4306 5997 4364 6023
rect 4306 5963 4318 5997
rect 4352 5963 4364 5997
rect 4306 5937 4364 5963
rect 4406 5997 4464 6023
rect 4406 5963 4418 5997
rect 4452 5963 4464 5997
rect 4406 5937 4464 5963
rect 4506 5997 4564 6023
rect 4506 5963 4518 5997
rect 4552 5963 4564 5997
rect 4506 5937 4564 5963
rect 4606 5997 4664 6023
rect 4606 5963 4618 5997
rect 4652 5963 4664 5997
rect 4606 5937 4664 5963
rect 4706 5997 4764 6023
rect 4706 5963 4718 5997
rect 4752 5963 4764 5997
rect 4706 5937 4764 5963
rect 4806 5997 4864 6023
rect 4806 5963 4818 5997
rect 4852 5963 4864 5997
rect 4806 5937 4864 5963
rect 4906 5997 4964 6023
rect 4906 5963 4918 5997
rect 4952 5963 4964 5997
rect 4906 5937 4964 5963
rect 5006 5997 5064 6023
rect 5006 5963 5018 5997
rect 5052 5963 5064 5997
rect 5006 5937 5064 5963
rect 5106 5997 5164 6023
rect 5106 5963 5118 5997
rect 5152 5963 5164 5997
rect 5106 5937 5164 5963
rect 5206 5997 5264 6023
rect 5206 5963 5212 5997
rect 5252 5963 5264 5997
rect 5206 5937 5264 5963
rect 5306 5997 5364 6023
rect 5306 5963 5318 5997
rect 5358 5963 5364 5997
rect 5306 5937 5364 5963
rect 5406 5997 5464 6023
rect 5406 5963 5418 5997
rect 5452 5963 5464 5997
rect 5406 5937 5464 5963
rect 5506 5997 5564 6023
rect 5506 5963 5518 5997
rect 5552 5963 5564 5997
rect 5506 5937 5564 5963
rect 5606 5997 5664 6023
rect 5606 5963 5618 5997
rect 5652 5963 5664 5997
rect 5606 5937 5664 5963
rect 5706 5997 5764 6023
rect 5706 5963 5718 5997
rect 5752 5963 5764 5997
rect 5706 5937 5764 5963
rect 5806 5997 5864 6023
rect 5806 5963 5812 5997
rect 5852 5963 5864 5997
rect 5806 5937 5864 5963
rect 5906 5997 5964 6023
rect 5906 5963 5918 5997
rect 5958 5963 5964 5997
rect 5906 5937 5964 5963
rect 6006 5997 6064 6023
rect 6006 5963 6018 5997
rect 6052 5963 6064 5997
rect 6006 5937 6064 5963
rect 6106 5997 6164 6023
rect 6106 5963 6118 5997
rect 6152 5963 6164 5997
rect 6106 5937 6164 5963
rect 6206 5997 6264 6023
rect 6206 5963 6218 5997
rect 6252 5963 6264 5997
rect 6206 5937 6264 5963
rect 6306 5997 6364 6023
rect 6306 5963 6318 5997
rect 6352 5963 6364 5997
rect 6306 5937 6364 5963
rect 6406 5997 6464 6023
rect 6618 6016 6862 6050
rect 6406 5963 6412 5997
rect 6452 5963 6464 5997
rect 6508 5978 6516 6012
rect 6558 5978 6574 6012
rect 6618 5997 6652 6016
rect 6406 5937 6464 5963
rect 6828 5997 6862 6016
rect 6618 5947 6652 5963
rect 6696 5948 6712 5982
rect 6754 5948 6762 5982
rect 6828 5947 6862 5963
rect 6928 5997 7162 6013
rect 6962 5963 7028 5997
rect 7062 5963 7128 5997
rect 6928 5947 7162 5963
rect 7228 5997 7362 6013
rect 7262 5963 7328 5997
rect 7228 5947 7362 5963
rect 7428 5997 7462 6013
rect 7428 5947 7462 5963
rect 6 5857 64 5883
rect 6 5823 18 5857
rect 58 5823 64 5857
rect 6 5797 64 5823
rect 106 5857 164 5883
rect 106 5823 118 5857
rect 152 5823 164 5857
rect 106 5797 164 5823
rect 206 5857 264 5883
rect 206 5823 218 5857
rect 252 5823 264 5857
rect 206 5797 264 5823
rect 306 5857 364 5883
rect 306 5823 318 5857
rect 352 5823 364 5857
rect 306 5797 364 5823
rect 406 5857 464 5883
rect 406 5823 418 5857
rect 452 5823 464 5857
rect 406 5797 464 5823
rect 506 5857 564 5883
rect 506 5823 518 5857
rect 552 5823 564 5857
rect 506 5797 564 5823
rect 606 5857 664 5883
rect 606 5823 618 5857
rect 652 5823 664 5857
rect 606 5797 664 5823
rect 706 5857 764 5883
rect 706 5823 718 5857
rect 752 5823 764 5857
rect 706 5797 764 5823
rect 806 5857 864 5883
rect 806 5823 818 5857
rect 852 5823 864 5857
rect 806 5797 864 5823
rect 906 5857 964 5883
rect 906 5823 918 5857
rect 952 5823 964 5857
rect 906 5797 964 5823
rect 1006 5857 1064 5883
rect 1006 5823 1018 5857
rect 1052 5823 1064 5857
rect 1006 5797 1064 5823
rect 1106 5857 1164 5883
rect 1106 5823 1118 5857
rect 1152 5823 1164 5857
rect 1106 5797 1164 5823
rect 1206 5857 1264 5883
rect 1206 5823 1218 5857
rect 1252 5823 1264 5857
rect 1206 5797 1264 5823
rect 1306 5857 1364 5883
rect 1306 5823 1318 5857
rect 1352 5823 1364 5857
rect 1306 5797 1364 5823
rect 1406 5857 1464 5883
rect 1406 5823 1418 5857
rect 1452 5823 1464 5857
rect 1406 5797 1464 5823
rect 1506 5857 1564 5883
rect 1506 5823 1518 5857
rect 1552 5823 1564 5857
rect 1506 5797 1564 5823
rect 1606 5857 1664 5883
rect 1606 5823 1618 5857
rect 1652 5823 1664 5857
rect 1606 5797 1664 5823
rect 1706 5857 1764 5883
rect 1706 5823 1718 5857
rect 1752 5823 1764 5857
rect 1706 5797 1764 5823
rect 1806 5857 1864 5883
rect 1806 5823 1818 5857
rect 1852 5823 1864 5857
rect 1806 5797 1864 5823
rect 1906 5857 1964 5883
rect 1906 5823 1918 5857
rect 1952 5823 1964 5857
rect 1906 5797 1964 5823
rect 2006 5857 2064 5883
rect 2006 5823 2012 5857
rect 2052 5823 2064 5857
rect 2006 5797 2064 5823
rect 2106 5857 2164 5883
rect 2106 5823 2118 5857
rect 2158 5823 2164 5857
rect 2106 5797 2164 5823
rect 2206 5857 2264 5883
rect 2206 5823 2218 5857
rect 2252 5823 2264 5857
rect 2206 5797 2264 5823
rect 2306 5857 2364 5883
rect 2306 5823 2318 5857
rect 2352 5823 2364 5857
rect 2306 5797 2364 5823
rect 2406 5857 2464 5883
rect 2406 5823 2418 5857
rect 2452 5823 2464 5857
rect 2406 5797 2464 5823
rect 2506 5857 2564 5883
rect 2506 5823 2518 5857
rect 2552 5823 2564 5857
rect 2506 5797 2564 5823
rect 2606 5857 2664 5883
rect 2606 5823 2618 5857
rect 2652 5823 2664 5857
rect 2606 5797 2664 5823
rect 2706 5857 2764 5883
rect 2706 5823 2718 5857
rect 2752 5823 2764 5857
rect 2706 5797 2764 5823
rect 2806 5857 2864 5883
rect 2806 5823 2818 5857
rect 2852 5823 2864 5857
rect 2806 5797 2864 5823
rect 2906 5857 2964 5883
rect 2906 5823 2918 5857
rect 2952 5823 2964 5857
rect 2906 5797 2964 5823
rect 3006 5857 3064 5883
rect 3006 5823 3018 5857
rect 3052 5823 3064 5857
rect 3006 5797 3064 5823
rect 3106 5857 3164 5883
rect 3106 5823 3118 5857
rect 3152 5823 3164 5857
rect 3106 5797 3164 5823
rect 3206 5857 3264 5883
rect 3206 5823 3218 5857
rect 3252 5823 3264 5857
rect 3206 5797 3264 5823
rect 3306 5857 3364 5883
rect 3306 5823 3318 5857
rect 3352 5823 3364 5857
rect 3306 5797 3364 5823
rect 3406 5857 3464 5883
rect 3406 5823 3412 5857
rect 3452 5823 3464 5857
rect 3406 5797 3464 5823
rect 3506 5857 3564 5883
rect 3506 5823 3518 5857
rect 3558 5823 3564 5857
rect 3506 5797 3564 5823
rect 3606 5857 3664 5883
rect 3606 5823 3618 5857
rect 3652 5823 3664 5857
rect 3606 5797 3664 5823
rect 3706 5857 3764 5883
rect 3706 5823 3718 5857
rect 3752 5823 3764 5857
rect 3706 5797 3764 5823
rect 3806 5857 3864 5883
rect 3806 5823 3818 5857
rect 3852 5823 3864 5857
rect 3806 5797 3864 5823
rect 3906 5857 3964 5883
rect 3906 5823 3918 5857
rect 3952 5823 3964 5857
rect 3906 5797 3964 5823
rect 4006 5857 4064 5883
rect 4006 5823 4018 5857
rect 4052 5823 4064 5857
rect 4006 5797 4064 5823
rect 4106 5857 4164 5883
rect 4106 5823 4112 5857
rect 4152 5823 4164 5857
rect 4106 5797 4164 5823
rect 4206 5857 4264 5883
rect 4206 5823 4218 5857
rect 4258 5823 4264 5857
rect 4206 5797 4264 5823
rect 4306 5857 4364 5883
rect 4306 5823 4318 5857
rect 4352 5823 4364 5857
rect 4306 5797 4364 5823
rect 4406 5857 4464 5883
rect 4406 5823 4418 5857
rect 4452 5823 4464 5857
rect 4406 5797 4464 5823
rect 4506 5857 4564 5883
rect 4506 5823 4518 5857
rect 4552 5823 4564 5857
rect 4506 5797 4564 5823
rect 4606 5857 4664 5883
rect 4606 5823 4618 5857
rect 4652 5823 4664 5857
rect 4606 5797 4664 5823
rect 4706 5857 4764 5883
rect 4706 5823 4718 5857
rect 4752 5823 4764 5857
rect 4706 5797 4764 5823
rect 4806 5857 4864 5883
rect 4806 5823 4818 5857
rect 4852 5823 4864 5857
rect 4806 5797 4864 5823
rect 4906 5857 4964 5883
rect 4906 5823 4918 5857
rect 4952 5823 4964 5857
rect 4906 5797 4964 5823
rect 5006 5857 5064 5883
rect 5006 5823 5018 5857
rect 5052 5823 5064 5857
rect 5006 5797 5064 5823
rect 5106 5857 5164 5883
rect 5106 5823 5118 5857
rect 5152 5823 5164 5857
rect 5106 5797 5164 5823
rect 5206 5857 5264 5883
rect 5206 5823 5218 5857
rect 5252 5823 5264 5857
rect 5206 5797 5264 5823
rect 5306 5857 5364 5883
rect 5306 5823 5318 5857
rect 5352 5823 5364 5857
rect 5306 5797 5364 5823
rect 5406 5857 5464 5883
rect 5406 5823 5418 5857
rect 5452 5823 5464 5857
rect 5406 5797 5464 5823
rect 5506 5857 5564 5883
rect 5506 5823 5518 5857
rect 5552 5823 5564 5857
rect 5506 5797 5564 5823
rect 5606 5857 5664 5883
rect 5606 5823 5618 5857
rect 5652 5823 5664 5857
rect 5606 5797 5664 5823
rect 5706 5857 5764 5883
rect 5706 5823 5712 5857
rect 5752 5823 5764 5857
rect 5706 5797 5764 5823
rect 5806 5857 5864 5883
rect 5806 5823 5818 5857
rect 5858 5823 5864 5857
rect 5806 5797 5864 5823
rect 5906 5857 5964 5883
rect 5906 5823 5912 5857
rect 5952 5823 5964 5857
rect 5906 5797 5964 5823
rect 6006 5857 6064 5883
rect 6006 5823 6018 5857
rect 6058 5823 6064 5857
rect 6006 5797 6064 5823
rect 6106 5857 6164 5883
rect 6106 5823 6118 5857
rect 6152 5823 6164 5857
rect 6106 5797 6164 5823
rect 6206 5857 6264 5883
rect 6206 5823 6218 5857
rect 6252 5823 6264 5857
rect 6206 5797 6264 5823
rect 6306 5857 6364 5883
rect 6306 5823 6318 5857
rect 6352 5823 6364 5857
rect 6306 5797 6364 5823
rect 6406 5857 6464 5883
rect 6618 5876 6862 5910
rect 6406 5823 6418 5857
rect 6452 5823 6464 5857
rect 6508 5838 6516 5872
rect 6558 5838 6574 5872
rect 6618 5857 6652 5876
rect 6406 5797 6464 5823
rect 6828 5873 6862 5876
rect 6828 5857 6962 5873
rect 6618 5807 6652 5823
rect 6696 5808 6712 5842
rect 6754 5808 6762 5842
rect 6862 5823 6928 5857
rect 6828 5807 6962 5823
rect 7028 5857 7062 5873
rect 7028 5807 7062 5823
rect 7128 5857 7362 5873
rect 7162 5823 7228 5857
rect 7262 5823 7328 5857
rect 7128 5807 7362 5823
rect 7428 5857 7462 5873
rect 7428 5807 7462 5823
rect 6 5717 64 5743
rect 6 5683 18 5717
rect 52 5683 64 5717
rect 6 5657 64 5683
rect 106 5717 164 5743
rect 106 5683 118 5717
rect 152 5683 164 5717
rect 106 5657 164 5683
rect 206 5717 264 5743
rect 206 5683 218 5717
rect 252 5683 264 5717
rect 206 5657 264 5683
rect 306 5717 364 5743
rect 306 5683 312 5717
rect 352 5683 364 5717
rect 306 5657 364 5683
rect 406 5717 464 5743
rect 406 5683 418 5717
rect 458 5683 464 5717
rect 406 5657 464 5683
rect 506 5717 564 5743
rect 506 5683 518 5717
rect 552 5683 564 5717
rect 506 5657 564 5683
rect 606 5717 664 5743
rect 606 5683 618 5717
rect 652 5683 664 5717
rect 606 5657 664 5683
rect 706 5717 764 5743
rect 706 5683 718 5717
rect 752 5683 764 5717
rect 706 5657 764 5683
rect 806 5717 864 5743
rect 806 5683 818 5717
rect 852 5683 864 5717
rect 806 5657 864 5683
rect 906 5717 964 5743
rect 906 5683 918 5717
rect 952 5683 964 5717
rect 906 5657 964 5683
rect 1006 5717 1064 5743
rect 1006 5683 1012 5717
rect 1052 5683 1064 5717
rect 1006 5657 1064 5683
rect 1106 5717 1164 5743
rect 1106 5683 1118 5717
rect 1158 5683 1164 5717
rect 1106 5657 1164 5683
rect 1206 5717 1264 5743
rect 1206 5683 1218 5717
rect 1252 5683 1264 5717
rect 1206 5657 1264 5683
rect 1306 5717 1364 5743
rect 1306 5683 1318 5717
rect 1352 5683 1364 5717
rect 1306 5657 1364 5683
rect 1406 5717 1464 5743
rect 1406 5683 1418 5717
rect 1452 5683 1464 5717
rect 1406 5657 1464 5683
rect 1506 5717 1564 5743
rect 1506 5683 1518 5717
rect 1552 5683 1564 5717
rect 1506 5657 1564 5683
rect 1606 5717 1664 5743
rect 1606 5683 1618 5717
rect 1652 5683 1664 5717
rect 1606 5657 1664 5683
rect 1706 5717 1764 5743
rect 1706 5683 1718 5717
rect 1752 5683 1764 5717
rect 1706 5657 1764 5683
rect 1806 5717 1864 5743
rect 1806 5683 1818 5717
rect 1852 5683 1864 5717
rect 1806 5657 1864 5683
rect 1906 5717 1964 5743
rect 1906 5683 1918 5717
rect 1952 5683 1964 5717
rect 1906 5657 1964 5683
rect 2006 5717 2064 5743
rect 2006 5683 2018 5717
rect 2052 5683 2064 5717
rect 2006 5657 2064 5683
rect 2106 5717 2164 5743
rect 2106 5683 2118 5717
rect 2152 5683 2164 5717
rect 2106 5657 2164 5683
rect 2206 5717 2264 5743
rect 2206 5683 2218 5717
rect 2252 5683 2264 5717
rect 2206 5657 2264 5683
rect 2306 5717 2364 5743
rect 2306 5683 2318 5717
rect 2352 5683 2364 5717
rect 2306 5657 2364 5683
rect 2406 5717 2464 5743
rect 2406 5683 2418 5717
rect 2452 5683 2464 5717
rect 2406 5657 2464 5683
rect 2506 5717 2564 5743
rect 2506 5683 2518 5717
rect 2552 5683 2564 5717
rect 2506 5657 2564 5683
rect 2606 5717 2664 5743
rect 2606 5683 2618 5717
rect 2652 5683 2664 5717
rect 2606 5657 2664 5683
rect 2706 5717 2764 5743
rect 2706 5683 2718 5717
rect 2752 5683 2764 5717
rect 2706 5657 2764 5683
rect 2806 5717 2864 5743
rect 2806 5683 2812 5717
rect 2852 5683 2864 5717
rect 2806 5657 2864 5683
rect 2906 5717 2964 5743
rect 2906 5683 2918 5717
rect 2958 5683 2964 5717
rect 2906 5657 2964 5683
rect 3006 5717 3064 5743
rect 3006 5683 3012 5717
rect 3052 5683 3064 5717
rect 3006 5657 3064 5683
rect 3106 5717 3164 5743
rect 3106 5683 3118 5717
rect 3158 5683 3164 5717
rect 3106 5657 3164 5683
rect 3206 5717 3264 5743
rect 3206 5683 3212 5717
rect 3252 5683 3264 5717
rect 3206 5657 3264 5683
rect 3306 5717 3364 5743
rect 3306 5683 3318 5717
rect 3358 5683 3364 5717
rect 3306 5657 3364 5683
rect 3406 5717 3464 5743
rect 3406 5683 3412 5717
rect 3452 5683 3464 5717
rect 3406 5657 3464 5683
rect 3506 5717 3564 5743
rect 3506 5683 3518 5717
rect 3558 5683 3564 5717
rect 3506 5657 3564 5683
rect 3606 5717 3664 5743
rect 3606 5683 3612 5717
rect 3652 5683 3664 5717
rect 3606 5657 3664 5683
rect 3706 5717 3764 5743
rect 3706 5683 3718 5717
rect 3758 5683 3764 5717
rect 3706 5657 3764 5683
rect 3806 5717 3864 5743
rect 3806 5683 3818 5717
rect 3852 5683 3864 5717
rect 3806 5657 3864 5683
rect 3906 5717 3964 5743
rect 3906 5683 3918 5717
rect 3952 5683 3964 5717
rect 3906 5657 3964 5683
rect 4006 5717 4064 5743
rect 4006 5683 4018 5717
rect 4052 5683 4064 5717
rect 4006 5657 4064 5683
rect 4106 5717 4164 5743
rect 4106 5683 4112 5717
rect 4152 5683 4164 5717
rect 4106 5657 4164 5683
rect 4206 5717 4264 5743
rect 4206 5683 4218 5717
rect 4258 5683 4264 5717
rect 4206 5657 4264 5683
rect 4306 5717 4364 5743
rect 4306 5683 4312 5717
rect 4352 5683 4364 5717
rect 4306 5657 4364 5683
rect 4406 5717 4464 5743
rect 4406 5683 4418 5717
rect 4458 5683 4464 5717
rect 4406 5657 4464 5683
rect 4506 5717 4564 5743
rect 4506 5683 4512 5717
rect 4552 5683 4564 5717
rect 4506 5657 4564 5683
rect 4606 5717 4664 5743
rect 4606 5683 4618 5717
rect 4658 5683 4664 5717
rect 4606 5657 4664 5683
rect 4706 5717 4764 5743
rect 4706 5683 4718 5717
rect 4752 5683 4764 5717
rect 4706 5657 4764 5683
rect 4806 5717 4864 5743
rect 4806 5683 4818 5717
rect 4852 5683 4864 5717
rect 4806 5657 4864 5683
rect 4906 5717 4964 5743
rect 4906 5683 4918 5717
rect 4952 5683 4964 5717
rect 4906 5657 4964 5683
rect 5006 5717 5064 5743
rect 5006 5683 5018 5717
rect 5052 5683 5064 5717
rect 5006 5657 5064 5683
rect 5106 5717 5164 5743
rect 5106 5683 5118 5717
rect 5152 5683 5164 5717
rect 5106 5657 5164 5683
rect 5206 5717 5264 5743
rect 5206 5683 5218 5717
rect 5252 5683 5264 5717
rect 5206 5657 5264 5683
rect 5306 5717 5364 5743
rect 5306 5683 5318 5717
rect 5352 5683 5364 5717
rect 5306 5657 5364 5683
rect 5406 5717 5464 5743
rect 5406 5683 5418 5717
rect 5452 5683 5464 5717
rect 5406 5657 5464 5683
rect 5506 5717 5564 5743
rect 5506 5683 5512 5717
rect 5552 5683 5564 5717
rect 5506 5657 5564 5683
rect 5606 5717 5664 5743
rect 5606 5683 5618 5717
rect 5658 5683 5664 5717
rect 5606 5657 5664 5683
rect 5706 5717 5764 5743
rect 5706 5683 5718 5717
rect 5752 5683 5764 5717
rect 5706 5657 5764 5683
rect 5806 5717 5864 5743
rect 5806 5683 5818 5717
rect 5852 5683 5864 5717
rect 5806 5657 5864 5683
rect 5906 5717 5964 5743
rect 5906 5683 5918 5717
rect 5952 5683 5964 5717
rect 5906 5657 5964 5683
rect 6006 5717 6064 5743
rect 6006 5683 6018 5717
rect 6052 5683 6064 5717
rect 6006 5657 6064 5683
rect 6106 5717 6164 5743
rect 6106 5683 6118 5717
rect 6152 5683 6164 5717
rect 6106 5657 6164 5683
rect 6206 5717 6264 5743
rect 6206 5683 6218 5717
rect 6252 5683 6264 5717
rect 6206 5657 6264 5683
rect 6306 5717 6364 5743
rect 6306 5683 6318 5717
rect 6352 5683 6364 5717
rect 6306 5657 6364 5683
rect 6406 5717 6464 5743
rect 6618 5736 6862 5770
rect 6406 5683 6418 5717
rect 6452 5683 6464 5717
rect 6508 5698 6516 5732
rect 6558 5698 6574 5732
rect 6618 5717 6652 5736
rect 6406 5657 6464 5683
rect 6828 5717 6862 5736
rect 6618 5667 6652 5683
rect 6696 5668 6712 5702
rect 6754 5668 6762 5702
rect 6828 5667 6862 5683
rect 6928 5717 7062 5733
rect 6962 5683 7028 5717
rect 6928 5667 7062 5683
rect 7128 5717 7362 5733
rect 7162 5683 7228 5717
rect 7262 5683 7328 5717
rect 7128 5667 7362 5683
rect 7428 5717 7462 5733
rect 7428 5667 7462 5683
rect 6 5577 64 5603
rect 6 5543 18 5577
rect 52 5543 64 5577
rect 6 5517 64 5543
rect 106 5577 164 5603
rect 106 5543 118 5577
rect 152 5543 164 5577
rect 106 5517 164 5543
rect 206 5577 264 5603
rect 206 5543 218 5577
rect 252 5543 264 5577
rect 206 5517 264 5543
rect 306 5577 364 5603
rect 306 5543 318 5577
rect 352 5543 364 5577
rect 306 5517 364 5543
rect 406 5577 464 5603
rect 406 5543 418 5577
rect 452 5543 464 5577
rect 406 5517 464 5543
rect 506 5577 564 5603
rect 506 5543 518 5577
rect 552 5543 564 5577
rect 506 5517 564 5543
rect 606 5577 664 5603
rect 606 5543 618 5577
rect 652 5543 664 5577
rect 606 5517 664 5543
rect 706 5577 764 5603
rect 706 5543 718 5577
rect 752 5543 764 5577
rect 706 5517 764 5543
rect 806 5577 864 5603
rect 806 5543 818 5577
rect 852 5543 864 5577
rect 806 5517 864 5543
rect 906 5577 964 5603
rect 906 5543 918 5577
rect 952 5543 964 5577
rect 906 5517 964 5543
rect 1006 5577 1064 5603
rect 1006 5543 1018 5577
rect 1052 5543 1064 5577
rect 1006 5517 1064 5543
rect 1106 5577 1164 5603
rect 1106 5543 1112 5577
rect 1152 5543 1164 5577
rect 1106 5517 1164 5543
rect 1206 5577 1264 5603
rect 1206 5543 1218 5577
rect 1258 5543 1264 5577
rect 1206 5517 1264 5543
rect 1306 5577 1364 5603
rect 1306 5543 1312 5577
rect 1352 5543 1364 5577
rect 1306 5517 1364 5543
rect 1406 5577 1464 5603
rect 1406 5543 1418 5577
rect 1458 5543 1464 5577
rect 1406 5517 1464 5543
rect 1506 5577 1564 5603
rect 1506 5543 1518 5577
rect 1552 5543 1564 5577
rect 1506 5517 1564 5543
rect 1606 5577 1664 5603
rect 1606 5543 1618 5577
rect 1652 5543 1664 5577
rect 1606 5517 1664 5543
rect 1706 5577 1764 5603
rect 1706 5543 1718 5577
rect 1752 5543 1764 5577
rect 1706 5517 1764 5543
rect 1806 5577 1864 5603
rect 1806 5543 1818 5577
rect 1852 5543 1864 5577
rect 1806 5517 1864 5543
rect 1906 5577 1964 5603
rect 1906 5543 1912 5577
rect 1952 5543 1964 5577
rect 1906 5517 1964 5543
rect 2006 5577 2064 5603
rect 2006 5543 2018 5577
rect 2058 5543 2064 5577
rect 2006 5517 2064 5543
rect 2106 5577 2164 5603
rect 2106 5543 2118 5577
rect 2152 5543 2164 5577
rect 2106 5517 2164 5543
rect 2206 5577 2264 5603
rect 2206 5543 2212 5577
rect 2252 5543 2264 5577
rect 2206 5517 2264 5543
rect 2306 5577 2364 5603
rect 2306 5543 2318 5577
rect 2358 5543 2364 5577
rect 2306 5517 2364 5543
rect 2406 5577 2464 5603
rect 2406 5543 2418 5577
rect 2452 5543 2464 5577
rect 2406 5517 2464 5543
rect 2506 5577 2564 5603
rect 2506 5543 2518 5577
rect 2552 5543 2564 5577
rect 2506 5517 2564 5543
rect 2606 5577 2664 5603
rect 2606 5543 2618 5577
rect 2652 5543 2664 5577
rect 2606 5517 2664 5543
rect 2706 5577 2764 5603
rect 2706 5543 2718 5577
rect 2752 5543 2764 5577
rect 2706 5517 2764 5543
rect 2806 5577 2864 5603
rect 2806 5543 2818 5577
rect 2852 5543 2864 5577
rect 2806 5517 2864 5543
rect 2906 5577 2964 5603
rect 2906 5543 2918 5577
rect 2952 5543 2964 5577
rect 2906 5517 2964 5543
rect 3006 5577 3064 5603
rect 3006 5543 3018 5577
rect 3052 5543 3064 5577
rect 3006 5517 3064 5543
rect 3106 5577 3164 5603
rect 3106 5543 3118 5577
rect 3152 5543 3164 5577
rect 3106 5517 3164 5543
rect 3206 5577 3264 5603
rect 3206 5543 3218 5577
rect 3252 5543 3264 5577
rect 3206 5517 3264 5543
rect 3306 5577 3364 5603
rect 3306 5543 3318 5577
rect 3352 5543 3364 5577
rect 3306 5517 3364 5543
rect 3406 5577 3464 5603
rect 3406 5543 3418 5577
rect 3452 5543 3464 5577
rect 3406 5517 3464 5543
rect 3506 5577 3564 5603
rect 3506 5543 3518 5577
rect 3552 5543 3564 5577
rect 3506 5517 3564 5543
rect 3606 5577 3664 5603
rect 3606 5543 3618 5577
rect 3652 5543 3664 5577
rect 3606 5517 3664 5543
rect 3706 5577 3764 5603
rect 3706 5543 3718 5577
rect 3752 5543 3764 5577
rect 3706 5517 3764 5543
rect 3806 5577 3864 5603
rect 3806 5543 3818 5577
rect 3852 5543 3864 5577
rect 3806 5517 3864 5543
rect 3906 5577 3964 5603
rect 3906 5543 3918 5577
rect 3952 5543 3964 5577
rect 3906 5517 3964 5543
rect 4006 5577 4064 5603
rect 4006 5543 4012 5577
rect 4052 5543 4064 5577
rect 4006 5517 4064 5543
rect 4106 5577 4164 5603
rect 4106 5543 4118 5577
rect 4158 5543 4164 5577
rect 4106 5517 4164 5543
rect 4206 5577 4264 5603
rect 4206 5543 4218 5577
rect 4252 5543 4264 5577
rect 4206 5517 4264 5543
rect 4306 5577 4364 5603
rect 4306 5543 4318 5577
rect 4352 5543 4364 5577
rect 4306 5517 4364 5543
rect 4406 5577 4464 5603
rect 4406 5543 4418 5577
rect 4452 5543 4464 5577
rect 4406 5517 4464 5543
rect 4506 5577 4564 5603
rect 4506 5543 4518 5577
rect 4552 5543 4564 5577
rect 4506 5517 4564 5543
rect 4606 5577 4664 5603
rect 4606 5543 4618 5577
rect 4652 5543 4664 5577
rect 4606 5517 4664 5543
rect 4706 5577 4764 5603
rect 4706 5543 4718 5577
rect 4752 5543 4764 5577
rect 4706 5517 4764 5543
rect 4806 5577 4864 5603
rect 4806 5543 4818 5577
rect 4852 5543 4864 5577
rect 4806 5517 4864 5543
rect 4906 5577 4964 5603
rect 4906 5543 4918 5577
rect 4952 5543 4964 5577
rect 4906 5517 4964 5543
rect 5006 5577 5064 5603
rect 5006 5543 5018 5577
rect 5052 5543 5064 5577
rect 5006 5517 5064 5543
rect 5106 5577 5164 5603
rect 5106 5543 5118 5577
rect 5152 5543 5164 5577
rect 5106 5517 5164 5543
rect 5206 5577 5264 5603
rect 5206 5543 5218 5577
rect 5252 5543 5264 5577
rect 5206 5517 5264 5543
rect 5306 5577 5364 5603
rect 5306 5543 5318 5577
rect 5352 5543 5364 5577
rect 5306 5517 5364 5543
rect 5406 5577 5464 5603
rect 5406 5543 5418 5577
rect 5452 5543 5464 5577
rect 5406 5517 5464 5543
rect 5506 5577 5564 5603
rect 5506 5543 5518 5577
rect 5552 5543 5564 5577
rect 5506 5517 5564 5543
rect 5606 5577 5664 5603
rect 5606 5543 5618 5577
rect 5652 5543 5664 5577
rect 5606 5517 5664 5543
rect 5706 5577 5764 5603
rect 5706 5543 5718 5577
rect 5752 5543 5764 5577
rect 5706 5517 5764 5543
rect 5806 5577 5864 5603
rect 5806 5543 5818 5577
rect 5852 5543 5864 5577
rect 5806 5517 5864 5543
rect 5906 5577 5964 5603
rect 5906 5543 5918 5577
rect 5952 5543 5964 5577
rect 5906 5517 5964 5543
rect 6006 5577 6064 5603
rect 6006 5543 6018 5577
rect 6052 5543 6064 5577
rect 6006 5517 6064 5543
rect 6106 5577 6164 5603
rect 6106 5543 6118 5577
rect 6152 5543 6164 5577
rect 6106 5517 6164 5543
rect 6206 5577 6264 5603
rect 6206 5543 6218 5577
rect 6252 5543 6264 5577
rect 6206 5517 6264 5543
rect 6306 5577 6364 5603
rect 6306 5543 6318 5577
rect 6352 5543 6364 5577
rect 6306 5517 6364 5543
rect 6406 5577 6464 5603
rect 6618 5596 6862 5630
rect 6406 5543 6418 5577
rect 6452 5543 6464 5577
rect 6508 5558 6516 5592
rect 6558 5558 6574 5592
rect 6618 5577 6652 5596
rect 6406 5517 6464 5543
rect 6828 5593 6862 5596
rect 6828 5577 6962 5593
rect 6618 5527 6652 5543
rect 6696 5528 6712 5562
rect 6754 5528 6762 5562
rect 6862 5543 6928 5577
rect 6828 5527 6962 5543
rect 7028 5577 7162 5593
rect 7062 5543 7128 5577
rect 7028 5527 7162 5543
rect 7228 5577 7262 5593
rect 7228 5527 7262 5543
rect 7328 5577 7462 5593
rect 7362 5543 7428 5577
rect 7328 5527 7462 5543
rect 6 5437 64 5463
rect 6 5403 18 5437
rect 58 5403 64 5437
rect 6 5377 64 5403
rect 106 5437 164 5463
rect 106 5403 118 5437
rect 152 5403 164 5437
rect 106 5377 164 5403
rect 206 5437 264 5463
rect 206 5403 218 5437
rect 252 5403 264 5437
rect 206 5377 264 5403
rect 306 5437 364 5463
rect 306 5403 318 5437
rect 352 5403 364 5437
rect 306 5377 364 5403
rect 406 5437 464 5463
rect 406 5403 412 5437
rect 452 5403 464 5437
rect 406 5377 464 5403
rect 506 5437 564 5463
rect 506 5403 518 5437
rect 558 5403 564 5437
rect 506 5377 564 5403
rect 606 5437 664 5463
rect 606 5403 618 5437
rect 652 5403 664 5437
rect 606 5377 664 5403
rect 706 5437 764 5463
rect 706 5403 718 5437
rect 752 5403 764 5437
rect 706 5377 764 5403
rect 806 5437 864 5463
rect 806 5403 818 5437
rect 852 5403 864 5437
rect 806 5377 864 5403
rect 906 5437 964 5463
rect 906 5403 918 5437
rect 952 5403 964 5437
rect 906 5377 964 5403
rect 1006 5437 1064 5463
rect 1006 5403 1018 5437
rect 1052 5403 1064 5437
rect 1006 5377 1064 5403
rect 1106 5437 1164 5463
rect 1106 5403 1118 5437
rect 1152 5403 1164 5437
rect 1106 5377 1164 5403
rect 1206 5437 1264 5463
rect 1206 5403 1218 5437
rect 1252 5403 1264 5437
rect 1206 5377 1264 5403
rect 1306 5437 1364 5463
rect 1306 5403 1318 5437
rect 1352 5403 1364 5437
rect 1306 5377 1364 5403
rect 1406 5437 1464 5463
rect 1406 5403 1412 5437
rect 1452 5403 1464 5437
rect 1406 5377 1464 5403
rect 1506 5437 1564 5463
rect 1506 5403 1518 5437
rect 1558 5403 1564 5437
rect 1506 5377 1564 5403
rect 1606 5437 1664 5463
rect 1606 5403 1618 5437
rect 1652 5403 1664 5437
rect 1606 5377 1664 5403
rect 1706 5437 1764 5463
rect 1706 5403 1712 5437
rect 1752 5403 1764 5437
rect 1706 5377 1764 5403
rect 1806 5437 1864 5463
rect 1806 5403 1818 5437
rect 1858 5403 1864 5437
rect 1806 5377 1864 5403
rect 1906 5437 1964 5463
rect 1906 5403 1918 5437
rect 1952 5403 1964 5437
rect 1906 5377 1964 5403
rect 2006 5437 2064 5463
rect 2006 5403 2018 5437
rect 2052 5403 2064 5437
rect 2006 5377 2064 5403
rect 2106 5437 2164 5463
rect 2106 5403 2118 5437
rect 2152 5403 2164 5437
rect 2106 5377 2164 5403
rect 2206 5437 2264 5463
rect 2206 5403 2212 5437
rect 2252 5403 2264 5437
rect 2206 5377 2264 5403
rect 2306 5437 2364 5463
rect 2306 5403 2318 5437
rect 2358 5403 2364 5437
rect 2306 5377 2364 5403
rect 2406 5437 2464 5463
rect 2406 5403 2418 5437
rect 2452 5403 2464 5437
rect 2406 5377 2464 5403
rect 2506 5437 2564 5463
rect 2506 5403 2518 5437
rect 2552 5403 2564 5437
rect 2506 5377 2564 5403
rect 2606 5437 2664 5463
rect 2606 5403 2618 5437
rect 2652 5403 2664 5437
rect 2606 5377 2664 5403
rect 2706 5437 2764 5463
rect 2706 5403 2718 5437
rect 2752 5403 2764 5437
rect 2706 5377 2764 5403
rect 2806 5437 2864 5463
rect 2806 5403 2818 5437
rect 2852 5403 2864 5437
rect 2806 5377 2864 5403
rect 2906 5437 2964 5463
rect 2906 5403 2918 5437
rect 2952 5403 2964 5437
rect 2906 5377 2964 5403
rect 3006 5437 3064 5463
rect 3006 5403 3018 5437
rect 3052 5403 3064 5437
rect 3006 5377 3064 5403
rect 3106 5437 3164 5463
rect 3106 5403 3118 5437
rect 3152 5403 3164 5437
rect 3106 5377 3164 5403
rect 3206 5437 3264 5463
rect 3206 5403 3218 5437
rect 3252 5403 3264 5437
rect 3206 5377 3264 5403
rect 3306 5437 3364 5463
rect 3306 5403 3318 5437
rect 3352 5403 3364 5437
rect 3306 5377 3364 5403
rect 3406 5437 3464 5463
rect 3406 5403 3418 5437
rect 3452 5403 3464 5437
rect 3406 5377 3464 5403
rect 3506 5437 3564 5463
rect 3506 5403 3518 5437
rect 3552 5403 3564 5437
rect 3506 5377 3564 5403
rect 3606 5437 3664 5463
rect 3606 5403 3618 5437
rect 3652 5403 3664 5437
rect 3606 5377 3664 5403
rect 3706 5437 3764 5463
rect 3706 5403 3712 5437
rect 3752 5403 3764 5437
rect 3706 5377 3764 5403
rect 3806 5437 3864 5463
rect 3806 5403 3818 5437
rect 3858 5403 3864 5437
rect 3806 5377 3864 5403
rect 3906 5437 3964 5463
rect 3906 5403 3918 5437
rect 3952 5403 3964 5437
rect 3906 5377 3964 5403
rect 4006 5437 4064 5463
rect 4006 5403 4018 5437
rect 4052 5403 4064 5437
rect 4006 5377 4064 5403
rect 4106 5437 4164 5463
rect 4106 5403 4118 5437
rect 4152 5403 4164 5437
rect 4106 5377 4164 5403
rect 4206 5437 4264 5463
rect 4206 5403 4218 5437
rect 4252 5403 4264 5437
rect 4206 5377 4264 5403
rect 4306 5437 4364 5463
rect 4306 5403 4318 5437
rect 4352 5403 4364 5437
rect 4306 5377 4364 5403
rect 4406 5437 4464 5463
rect 4406 5403 4418 5437
rect 4452 5403 4464 5437
rect 4406 5377 4464 5403
rect 4506 5437 4564 5463
rect 4506 5403 4518 5437
rect 4552 5403 4564 5437
rect 4506 5377 4564 5403
rect 4606 5437 4664 5463
rect 4606 5403 4618 5437
rect 4652 5403 4664 5437
rect 4606 5377 4664 5403
rect 4706 5437 4764 5463
rect 4706 5403 4718 5437
rect 4752 5403 4764 5437
rect 4706 5377 4764 5403
rect 4806 5437 4864 5463
rect 4806 5403 4818 5437
rect 4852 5403 4864 5437
rect 4806 5377 4864 5403
rect 4906 5437 4964 5463
rect 4906 5403 4918 5437
rect 4952 5403 4964 5437
rect 4906 5377 4964 5403
rect 5006 5437 5064 5463
rect 5006 5403 5018 5437
rect 5052 5403 5064 5437
rect 5006 5377 5064 5403
rect 5106 5437 5164 5463
rect 5106 5403 5112 5437
rect 5152 5403 5164 5437
rect 5106 5377 5164 5403
rect 5206 5437 5264 5463
rect 5206 5403 5218 5437
rect 5258 5403 5264 5437
rect 5206 5377 5264 5403
rect 5306 5437 5364 5463
rect 5306 5403 5312 5437
rect 5352 5403 5364 5437
rect 5306 5377 5364 5403
rect 5406 5437 5464 5463
rect 5406 5403 5418 5437
rect 5458 5403 5464 5437
rect 5406 5377 5464 5403
rect 5506 5437 5564 5463
rect 5506 5403 5512 5437
rect 5552 5403 5564 5437
rect 5506 5377 5564 5403
rect 5606 5437 5664 5463
rect 5606 5403 5618 5437
rect 5658 5403 5664 5437
rect 5606 5377 5664 5403
rect 5706 5437 5764 5463
rect 5706 5403 5712 5437
rect 5752 5403 5764 5437
rect 5706 5377 5764 5403
rect 5806 5437 5864 5463
rect 5806 5403 5818 5437
rect 5858 5403 5864 5437
rect 5806 5377 5864 5403
rect 5906 5437 5964 5463
rect 5906 5403 5918 5437
rect 5952 5403 5964 5437
rect 5906 5377 5964 5403
rect 6006 5437 6064 5463
rect 6006 5403 6018 5437
rect 6052 5403 6064 5437
rect 6006 5377 6064 5403
rect 6106 5437 6164 5463
rect 6106 5403 6118 5437
rect 6152 5403 6164 5437
rect 6106 5377 6164 5403
rect 6206 5437 6264 5463
rect 6206 5403 6218 5437
rect 6252 5403 6264 5437
rect 6206 5377 6264 5403
rect 6306 5437 6364 5463
rect 6306 5403 6318 5437
rect 6352 5403 6364 5437
rect 6306 5377 6364 5403
rect 6406 5437 6464 5463
rect 6618 5456 6862 5490
rect 6406 5403 6418 5437
rect 6452 5403 6464 5437
rect 6508 5418 6516 5452
rect 6558 5418 6574 5452
rect 6618 5437 6652 5456
rect 6406 5377 6464 5403
rect 6828 5437 6862 5456
rect 6618 5387 6652 5403
rect 6696 5388 6712 5422
rect 6754 5388 6762 5422
rect 6828 5387 6862 5403
rect 6928 5437 7162 5453
rect 6962 5403 7028 5437
rect 7062 5403 7128 5437
rect 6928 5387 7162 5403
rect 7228 5437 7262 5453
rect 7228 5387 7262 5403
rect 7328 5437 7462 5453
rect 7362 5403 7428 5437
rect 7328 5387 7462 5403
rect 6 5297 64 5323
rect 6 5263 18 5297
rect 52 5263 64 5297
rect 6 5237 64 5263
rect 106 5297 164 5323
rect 106 5263 118 5297
rect 152 5263 164 5297
rect 106 5237 164 5263
rect 206 5297 264 5323
rect 206 5263 218 5297
rect 252 5263 264 5297
rect 206 5237 264 5263
rect 306 5297 364 5323
rect 306 5263 318 5297
rect 352 5263 364 5297
rect 306 5237 364 5263
rect 406 5297 464 5323
rect 406 5263 418 5297
rect 452 5263 464 5297
rect 406 5237 464 5263
rect 506 5297 564 5323
rect 506 5263 518 5297
rect 552 5263 564 5297
rect 506 5237 564 5263
rect 606 5297 664 5323
rect 606 5263 618 5297
rect 652 5263 664 5297
rect 606 5237 664 5263
rect 706 5297 764 5323
rect 706 5263 718 5297
rect 752 5263 764 5297
rect 706 5237 764 5263
rect 806 5297 864 5323
rect 806 5263 818 5297
rect 852 5263 864 5297
rect 806 5237 864 5263
rect 906 5297 964 5323
rect 906 5263 918 5297
rect 952 5263 964 5297
rect 906 5237 964 5263
rect 1006 5297 1064 5323
rect 1006 5263 1018 5297
rect 1052 5263 1064 5297
rect 1006 5237 1064 5263
rect 1106 5297 1164 5323
rect 1106 5263 1118 5297
rect 1152 5263 1164 5297
rect 1106 5237 1164 5263
rect 1206 5297 1264 5323
rect 1206 5263 1218 5297
rect 1252 5263 1264 5297
rect 1206 5237 1264 5263
rect 1306 5297 1364 5323
rect 1306 5263 1318 5297
rect 1352 5263 1364 5297
rect 1306 5237 1364 5263
rect 1406 5297 1464 5323
rect 1406 5263 1418 5297
rect 1452 5263 1464 5297
rect 1406 5237 1464 5263
rect 1506 5297 1564 5323
rect 1506 5263 1518 5297
rect 1552 5263 1564 5297
rect 1506 5237 1564 5263
rect 1606 5297 1664 5323
rect 1606 5263 1618 5297
rect 1652 5263 1664 5297
rect 1606 5237 1664 5263
rect 1706 5297 1764 5323
rect 1706 5263 1718 5297
rect 1752 5263 1764 5297
rect 1706 5237 1764 5263
rect 1806 5297 1864 5323
rect 1806 5263 1818 5297
rect 1852 5263 1864 5297
rect 1806 5237 1864 5263
rect 1906 5297 1964 5323
rect 1906 5263 1918 5297
rect 1952 5263 1964 5297
rect 1906 5237 1964 5263
rect 2006 5297 2064 5323
rect 2006 5263 2018 5297
rect 2052 5263 2064 5297
rect 2006 5237 2064 5263
rect 2106 5297 2164 5323
rect 2106 5263 2112 5297
rect 2152 5263 2164 5297
rect 2106 5237 2164 5263
rect 2206 5297 2264 5323
rect 2206 5263 2218 5297
rect 2258 5263 2264 5297
rect 2206 5237 2264 5263
rect 2306 5297 2364 5323
rect 2306 5263 2312 5297
rect 2352 5263 2364 5297
rect 2306 5237 2364 5263
rect 2406 5297 2464 5323
rect 2406 5263 2418 5297
rect 2458 5263 2464 5297
rect 2406 5237 2464 5263
rect 2506 5297 2564 5323
rect 2506 5263 2518 5297
rect 2552 5263 2564 5297
rect 2506 5237 2564 5263
rect 2606 5297 2664 5323
rect 2606 5263 2612 5297
rect 2652 5263 2664 5297
rect 2606 5237 2664 5263
rect 2706 5297 2764 5323
rect 2706 5263 2718 5297
rect 2758 5263 2764 5297
rect 2706 5237 2764 5263
rect 2806 5297 2864 5323
rect 2806 5263 2818 5297
rect 2852 5263 2864 5297
rect 2806 5237 2864 5263
rect 2906 5297 2964 5323
rect 2906 5263 2912 5297
rect 2952 5263 2964 5297
rect 2906 5237 2964 5263
rect 3006 5297 3064 5323
rect 3006 5263 3018 5297
rect 3058 5263 3064 5297
rect 3006 5237 3064 5263
rect 3106 5297 3164 5323
rect 3106 5263 3112 5297
rect 3152 5263 3164 5297
rect 3106 5237 3164 5263
rect 3206 5297 3264 5323
rect 3206 5263 3218 5297
rect 3258 5263 3264 5297
rect 3206 5237 3264 5263
rect 3306 5297 3364 5323
rect 3306 5263 3318 5297
rect 3352 5263 3364 5297
rect 3306 5237 3364 5263
rect 3406 5297 3464 5323
rect 3406 5263 3418 5297
rect 3452 5263 3464 5297
rect 3406 5237 3464 5263
rect 3506 5297 3564 5323
rect 3506 5263 3518 5297
rect 3552 5263 3564 5297
rect 3506 5237 3564 5263
rect 3606 5297 3664 5323
rect 3606 5263 3618 5297
rect 3652 5263 3664 5297
rect 3606 5237 3664 5263
rect 3706 5297 3764 5323
rect 3706 5263 3718 5297
rect 3752 5263 3764 5297
rect 3706 5237 3764 5263
rect 3806 5297 3864 5323
rect 3806 5263 3818 5297
rect 3852 5263 3864 5297
rect 3806 5237 3864 5263
rect 3906 5297 3964 5323
rect 3906 5263 3918 5297
rect 3952 5263 3964 5297
rect 3906 5237 3964 5263
rect 4006 5297 4064 5323
rect 4006 5263 4018 5297
rect 4052 5263 4064 5297
rect 4006 5237 4064 5263
rect 4106 5297 4164 5323
rect 4106 5263 4118 5297
rect 4152 5263 4164 5297
rect 4106 5237 4164 5263
rect 4206 5297 4264 5323
rect 4206 5263 4218 5297
rect 4252 5263 4264 5297
rect 4206 5237 4264 5263
rect 4306 5297 4364 5323
rect 4306 5263 4318 5297
rect 4352 5263 4364 5297
rect 4306 5237 4364 5263
rect 4406 5297 4464 5323
rect 4406 5263 4418 5297
rect 4452 5263 4464 5297
rect 4406 5237 4464 5263
rect 4506 5297 4564 5323
rect 4506 5263 4518 5297
rect 4552 5263 4564 5297
rect 4506 5237 4564 5263
rect 4606 5297 4664 5323
rect 4606 5263 4618 5297
rect 4652 5263 4664 5297
rect 4606 5237 4664 5263
rect 4706 5297 4764 5323
rect 4706 5263 4718 5297
rect 4752 5263 4764 5297
rect 4706 5237 4764 5263
rect 4806 5297 4864 5323
rect 4806 5263 4818 5297
rect 4852 5263 4864 5297
rect 4806 5237 4864 5263
rect 4906 5297 4964 5323
rect 4906 5263 4918 5297
rect 4952 5263 4964 5297
rect 4906 5237 4964 5263
rect 5006 5297 5064 5323
rect 5006 5263 5018 5297
rect 5052 5263 5064 5297
rect 5006 5237 5064 5263
rect 5106 5297 5164 5323
rect 5106 5263 5118 5297
rect 5152 5263 5164 5297
rect 5106 5237 5164 5263
rect 5206 5297 5264 5323
rect 5206 5263 5212 5297
rect 5252 5263 5264 5297
rect 5206 5237 5264 5263
rect 5306 5297 5364 5323
rect 5306 5263 5318 5297
rect 5358 5263 5364 5297
rect 5306 5237 5364 5263
rect 5406 5297 5464 5323
rect 5406 5263 5412 5297
rect 5452 5263 5464 5297
rect 5406 5237 5464 5263
rect 5506 5297 5564 5323
rect 5506 5263 5518 5297
rect 5558 5263 5564 5297
rect 5506 5237 5564 5263
rect 5606 5297 5664 5323
rect 5606 5263 5618 5297
rect 5652 5263 5664 5297
rect 5606 5237 5664 5263
rect 5706 5297 5764 5323
rect 5706 5263 5718 5297
rect 5752 5263 5764 5297
rect 5706 5237 5764 5263
rect 5806 5297 5864 5323
rect 5806 5263 5818 5297
rect 5852 5263 5864 5297
rect 5806 5237 5864 5263
rect 5906 5297 5964 5323
rect 5906 5263 5918 5297
rect 5952 5263 5964 5297
rect 5906 5237 5964 5263
rect 6006 5297 6064 5323
rect 6006 5263 6018 5297
rect 6052 5263 6064 5297
rect 6006 5237 6064 5263
rect 6106 5297 6164 5323
rect 6106 5263 6118 5297
rect 6152 5263 6164 5297
rect 6106 5237 6164 5263
rect 6206 5297 6264 5323
rect 6206 5263 6218 5297
rect 6252 5263 6264 5297
rect 6206 5237 6264 5263
rect 6306 5297 6364 5323
rect 6306 5263 6318 5297
rect 6352 5263 6364 5297
rect 6306 5237 6364 5263
rect 6406 5297 6464 5323
rect 6618 5316 6862 5350
rect 6406 5263 6412 5297
rect 6452 5263 6464 5297
rect 6508 5278 6516 5312
rect 6558 5278 6574 5312
rect 6618 5297 6652 5316
rect 6406 5237 6464 5263
rect 6828 5313 6862 5316
rect 6828 5297 6962 5313
rect 6618 5247 6652 5263
rect 6696 5248 6712 5282
rect 6754 5248 6762 5282
rect 6862 5263 6928 5297
rect 6828 5247 6962 5263
rect 7028 5297 7062 5313
rect 7028 5247 7062 5263
rect 7128 5297 7262 5313
rect 7162 5263 7228 5297
rect 7128 5247 7262 5263
rect 7328 5297 7462 5313
rect 7362 5263 7428 5297
rect 7328 5247 7462 5263
rect 6 5157 64 5183
rect 6 5123 18 5157
rect 52 5123 64 5157
rect 6 5097 64 5123
rect 106 5157 164 5183
rect 106 5123 118 5157
rect 152 5123 164 5157
rect 106 5097 164 5123
rect 206 5157 264 5183
rect 206 5123 218 5157
rect 252 5123 264 5157
rect 206 5097 264 5123
rect 306 5157 364 5183
rect 306 5123 318 5157
rect 352 5123 364 5157
rect 306 5097 364 5123
rect 406 5157 464 5183
rect 406 5123 418 5157
rect 452 5123 464 5157
rect 406 5097 464 5123
rect 506 5157 564 5183
rect 506 5123 518 5157
rect 552 5123 564 5157
rect 506 5097 564 5123
rect 606 5157 664 5183
rect 606 5123 618 5157
rect 652 5123 664 5157
rect 606 5097 664 5123
rect 706 5157 764 5183
rect 706 5123 718 5157
rect 752 5123 764 5157
rect 706 5097 764 5123
rect 806 5157 864 5183
rect 806 5123 818 5157
rect 852 5123 864 5157
rect 806 5097 864 5123
rect 906 5157 964 5183
rect 906 5123 918 5157
rect 952 5123 964 5157
rect 906 5097 964 5123
rect 1006 5157 1064 5183
rect 1006 5123 1018 5157
rect 1052 5123 1064 5157
rect 1006 5097 1064 5123
rect 1106 5157 1164 5183
rect 1106 5123 1118 5157
rect 1152 5123 1164 5157
rect 1106 5097 1164 5123
rect 1206 5157 1264 5183
rect 1206 5123 1218 5157
rect 1252 5123 1264 5157
rect 1206 5097 1264 5123
rect 1306 5157 1364 5183
rect 1306 5123 1312 5157
rect 1352 5123 1364 5157
rect 1306 5097 1364 5123
rect 1406 5157 1464 5183
rect 1406 5123 1418 5157
rect 1458 5123 1464 5157
rect 1406 5097 1464 5123
rect 1506 5157 1564 5183
rect 1506 5123 1518 5157
rect 1552 5123 1564 5157
rect 1506 5097 1564 5123
rect 1606 5157 1664 5183
rect 1606 5123 1618 5157
rect 1652 5123 1664 5157
rect 1606 5097 1664 5123
rect 1706 5157 1764 5183
rect 1706 5123 1718 5157
rect 1752 5123 1764 5157
rect 1706 5097 1764 5123
rect 1806 5157 1864 5183
rect 1806 5123 1818 5157
rect 1852 5123 1864 5157
rect 1806 5097 1864 5123
rect 1906 5157 1964 5183
rect 1906 5123 1918 5157
rect 1952 5123 1964 5157
rect 1906 5097 1964 5123
rect 2006 5157 2064 5183
rect 2006 5123 2018 5157
rect 2052 5123 2064 5157
rect 2006 5097 2064 5123
rect 2106 5157 2164 5183
rect 2106 5123 2112 5157
rect 2152 5123 2164 5157
rect 2106 5097 2164 5123
rect 2206 5157 2264 5183
rect 2206 5123 2218 5157
rect 2258 5123 2264 5157
rect 2206 5097 2264 5123
rect 2306 5157 2364 5183
rect 2306 5123 2318 5157
rect 2352 5123 2364 5157
rect 2306 5097 2364 5123
rect 2406 5157 2464 5183
rect 2406 5123 2418 5157
rect 2452 5123 2464 5157
rect 2406 5097 2464 5123
rect 2506 5157 2564 5183
rect 2506 5123 2518 5157
rect 2552 5123 2564 5157
rect 2506 5097 2564 5123
rect 2606 5157 2664 5183
rect 2606 5123 2618 5157
rect 2652 5123 2664 5157
rect 2606 5097 2664 5123
rect 2706 5157 2764 5183
rect 2706 5123 2718 5157
rect 2752 5123 2764 5157
rect 2706 5097 2764 5123
rect 2806 5157 2864 5183
rect 2806 5123 2818 5157
rect 2852 5123 2864 5157
rect 2806 5097 2864 5123
rect 2906 5157 2964 5183
rect 2906 5123 2918 5157
rect 2952 5123 2964 5157
rect 2906 5097 2964 5123
rect 3006 5157 3064 5183
rect 3006 5123 3018 5157
rect 3052 5123 3064 5157
rect 3006 5097 3064 5123
rect 3106 5157 3164 5183
rect 3106 5123 3118 5157
rect 3152 5123 3164 5157
rect 3106 5097 3164 5123
rect 3206 5157 3264 5183
rect 3206 5123 3218 5157
rect 3252 5123 3264 5157
rect 3206 5097 3264 5123
rect 3306 5157 3364 5183
rect 3306 5123 3318 5157
rect 3352 5123 3364 5157
rect 3306 5097 3364 5123
rect 3406 5157 3464 5183
rect 3406 5123 3418 5157
rect 3452 5123 3464 5157
rect 3406 5097 3464 5123
rect 3506 5157 3564 5183
rect 3506 5123 3518 5157
rect 3552 5123 3564 5157
rect 3506 5097 3564 5123
rect 3606 5157 3664 5183
rect 3606 5123 3618 5157
rect 3652 5123 3664 5157
rect 3606 5097 3664 5123
rect 3706 5157 3764 5183
rect 3706 5123 3718 5157
rect 3752 5123 3764 5157
rect 3706 5097 3764 5123
rect 3806 5157 3864 5183
rect 3806 5123 3818 5157
rect 3852 5123 3864 5157
rect 3806 5097 3864 5123
rect 3906 5157 3964 5183
rect 3906 5123 3918 5157
rect 3952 5123 3964 5157
rect 3906 5097 3964 5123
rect 4006 5157 4064 5183
rect 4006 5123 4018 5157
rect 4052 5123 4064 5157
rect 4006 5097 4064 5123
rect 4106 5157 4164 5183
rect 4106 5123 4118 5157
rect 4152 5123 4164 5157
rect 4106 5097 4164 5123
rect 4206 5157 4264 5183
rect 4206 5123 4218 5157
rect 4252 5123 4264 5157
rect 4206 5097 4264 5123
rect 4306 5157 4364 5183
rect 4306 5123 4312 5157
rect 4352 5123 4364 5157
rect 4306 5097 4364 5123
rect 4406 5157 4464 5183
rect 4406 5123 4418 5157
rect 4458 5123 4464 5157
rect 4406 5097 4464 5123
rect 4506 5157 4564 5183
rect 4506 5123 4518 5157
rect 4552 5123 4564 5157
rect 4506 5097 4564 5123
rect 4606 5157 4664 5183
rect 4606 5123 4618 5157
rect 4652 5123 4664 5157
rect 4606 5097 4664 5123
rect 4706 5157 4764 5183
rect 4706 5123 4712 5157
rect 4752 5123 4764 5157
rect 4706 5097 4764 5123
rect 4806 5157 4864 5183
rect 4806 5123 4818 5157
rect 4858 5123 4864 5157
rect 4806 5097 4864 5123
rect 4906 5157 4964 5183
rect 4906 5123 4918 5157
rect 4952 5123 4964 5157
rect 4906 5097 4964 5123
rect 5006 5157 5064 5183
rect 5006 5123 5018 5157
rect 5052 5123 5064 5157
rect 5006 5097 5064 5123
rect 5106 5157 5164 5183
rect 5106 5123 5118 5157
rect 5152 5123 5164 5157
rect 5106 5097 5164 5123
rect 5206 5157 5264 5183
rect 5206 5123 5218 5157
rect 5252 5123 5264 5157
rect 5206 5097 5264 5123
rect 5306 5157 5364 5183
rect 5306 5123 5318 5157
rect 5352 5123 5364 5157
rect 5306 5097 5364 5123
rect 5406 5157 5464 5183
rect 5406 5123 5418 5157
rect 5452 5123 5464 5157
rect 5406 5097 5464 5123
rect 5506 5157 5564 5183
rect 5506 5123 5518 5157
rect 5552 5123 5564 5157
rect 5506 5097 5564 5123
rect 5606 5157 5664 5183
rect 5606 5123 5618 5157
rect 5652 5123 5664 5157
rect 5606 5097 5664 5123
rect 5706 5157 5764 5183
rect 5706 5123 5712 5157
rect 5752 5123 5764 5157
rect 5706 5097 5764 5123
rect 5806 5157 5864 5183
rect 5806 5123 5818 5157
rect 5858 5123 5864 5157
rect 5806 5097 5864 5123
rect 5906 5157 5964 5183
rect 5906 5123 5918 5157
rect 5952 5123 5964 5157
rect 5906 5097 5964 5123
rect 6006 5157 6064 5183
rect 6006 5123 6018 5157
rect 6052 5123 6064 5157
rect 6006 5097 6064 5123
rect 6106 5157 6164 5183
rect 6106 5123 6118 5157
rect 6152 5123 6164 5157
rect 6106 5097 6164 5123
rect 6206 5157 6264 5183
rect 6206 5123 6218 5157
rect 6252 5123 6264 5157
rect 6206 5097 6264 5123
rect 6306 5157 6364 5183
rect 6306 5123 6318 5157
rect 6352 5123 6364 5157
rect 6306 5097 6364 5123
rect 6406 5157 6464 5183
rect 6618 5176 6862 5210
rect 6406 5123 6418 5157
rect 6452 5123 6464 5157
rect 6508 5138 6516 5172
rect 6558 5138 6574 5172
rect 6618 5157 6652 5176
rect 6406 5097 6464 5123
rect 6828 5157 6862 5176
rect 6618 5107 6652 5123
rect 6696 5108 6712 5142
rect 6754 5108 6762 5142
rect 6828 5107 6862 5123
rect 6928 5157 7062 5173
rect 6962 5123 7028 5157
rect 6928 5107 7062 5123
rect 7128 5157 7262 5173
rect 7162 5123 7228 5157
rect 7128 5107 7262 5123
rect 7328 5157 7462 5173
rect 7362 5123 7428 5157
rect 7328 5107 7462 5123
rect 106 5017 164 5043
rect 106 4983 118 5017
rect 152 4983 164 5017
rect 106 4957 164 4983
rect 306 5017 364 5043
rect 306 4983 318 5017
rect 352 4983 364 5017
rect 306 4957 364 4983
rect 506 5017 564 5043
rect 506 4983 518 5017
rect 552 4983 564 5017
rect 506 4957 564 4983
rect 706 5017 764 5043
rect 706 4983 718 5017
rect 752 4983 764 5017
rect 706 4957 764 4983
rect 906 5017 964 5043
rect 906 4983 918 5017
rect 952 4983 964 5017
rect 906 4957 964 4983
rect 1106 5017 1164 5043
rect 1106 4983 1118 5017
rect 1152 4983 1164 5017
rect 1106 4957 1164 4983
rect 1306 5017 1364 5043
rect 1306 4983 1318 5017
rect 1352 4983 1364 5017
rect 1306 4957 1364 4983
rect 1506 5017 1564 5043
rect 1506 4983 1518 5017
rect 1552 4983 1564 5017
rect 1506 4957 1564 4983
rect 1706 5017 1764 5043
rect 1706 4983 1718 5017
rect 1752 4983 1764 5017
rect 1706 4957 1764 4983
rect 1906 5017 1964 5043
rect 1906 4983 1918 5017
rect 1952 4983 1964 5017
rect 1906 4957 1964 4983
rect 2106 5017 2164 5043
rect 2106 4983 2118 5017
rect 2152 4983 2164 5017
rect 2106 4957 2164 4983
rect 2306 5017 2364 5043
rect 2306 4983 2318 5017
rect 2352 4983 2364 5017
rect 2306 4957 2364 4983
rect 2506 5017 2564 5043
rect 2506 4983 2518 5017
rect 2552 4983 2564 5017
rect 2506 4957 2564 4983
rect 2706 5017 2764 5043
rect 2706 4983 2718 5017
rect 2752 4983 2764 5017
rect 2706 4957 2764 4983
rect 2906 5017 2964 5043
rect 2906 4983 2918 5017
rect 2952 4983 2964 5017
rect 2906 4957 2964 4983
rect 3106 5017 3164 5043
rect 3106 4983 3118 5017
rect 3152 4983 3164 5017
rect 3106 4957 3164 4983
rect 3306 5017 3364 5043
rect 3306 4983 3318 5017
rect 3352 4983 3364 5017
rect 3306 4957 3364 4983
rect 3506 5017 3564 5043
rect 3506 4983 3518 5017
rect 3552 4983 3564 5017
rect 3506 4957 3564 4983
rect 3706 5017 3764 5043
rect 3706 4983 3718 5017
rect 3752 4983 3764 5017
rect 3706 4957 3764 4983
rect 3906 5017 3964 5043
rect 3906 4983 3918 5017
rect 3952 4983 3964 5017
rect 3906 4957 3964 4983
rect 4106 5017 4164 5043
rect 4106 4983 4118 5017
rect 4152 4983 4164 5017
rect 4106 4957 4164 4983
rect 4306 5017 4364 5043
rect 4306 4983 4318 5017
rect 4352 4983 4364 5017
rect 4306 4957 4364 4983
rect 4506 5017 4564 5043
rect 4506 4983 4518 5017
rect 4552 4983 4564 5017
rect 4506 4957 4564 4983
rect 4706 5017 4764 5043
rect 4706 4983 4718 5017
rect 4752 4983 4764 5017
rect 4706 4957 4764 4983
rect 4906 5017 4964 5043
rect 4906 4983 4918 5017
rect 4952 4983 4964 5017
rect 4906 4957 4964 4983
rect 5106 5017 5164 5043
rect 5106 4983 5118 5017
rect 5152 4983 5164 5017
rect 5106 4957 5164 4983
rect 5306 5017 5364 5043
rect 5306 4983 5318 5017
rect 5352 4983 5364 5017
rect 5306 4957 5364 4983
rect 5506 5017 5564 5043
rect 5506 4983 5518 5017
rect 5552 4983 5564 5017
rect 5506 4957 5564 4983
rect 5706 5017 5764 5043
rect 5706 4983 5718 5017
rect 5752 4983 5764 5017
rect 5706 4957 5764 4983
rect 5906 5017 5964 5043
rect 5906 4983 5918 5017
rect 5952 4983 5964 5017
rect 5906 4957 5964 4983
rect 6106 5017 6164 5043
rect 6106 4983 6118 5017
rect 6152 4983 6164 5017
rect 6106 4957 6164 4983
rect 6306 5017 6364 5043
rect 6306 4983 6318 5017
rect 6352 4983 6364 5017
rect 6306 4957 6364 4983
rect 8 4860 18 4894
rect 52 4860 118 4894
rect 152 4860 168 4894
rect 208 4876 218 4910
rect 252 4876 318 4910
rect 352 4876 368 4910
rect 408 4860 418 4894
rect 452 4860 518 4894
rect 552 4860 568 4894
rect 608 4876 618 4910
rect 652 4876 718 4910
rect 752 4876 768 4910
rect 808 4860 818 4894
rect 852 4860 918 4894
rect 952 4860 968 4894
rect 1008 4876 1018 4910
rect 1052 4876 1118 4910
rect 1152 4876 1168 4910
rect 1208 4860 1218 4894
rect 1252 4860 1318 4894
rect 1352 4860 1368 4894
rect 1408 4876 1418 4910
rect 1452 4876 1518 4910
rect 1552 4876 1568 4910
rect 1608 4860 1618 4894
rect 1652 4860 1718 4894
rect 1752 4860 1768 4894
rect 1808 4876 1818 4910
rect 1852 4876 1918 4910
rect 1952 4876 1968 4910
rect 2008 4860 2018 4894
rect 2052 4860 2118 4894
rect 2152 4860 2168 4894
rect 2208 4876 2218 4910
rect 2252 4876 2318 4910
rect 2352 4876 2368 4910
rect 2408 4860 2418 4894
rect 2452 4860 2518 4894
rect 2552 4860 2568 4894
rect 2608 4876 2618 4910
rect 2652 4876 2718 4910
rect 2752 4876 2768 4910
rect 2808 4860 2818 4894
rect 2852 4860 2918 4894
rect 2952 4860 2968 4894
rect 3008 4876 3018 4910
rect 3052 4876 3118 4910
rect 3152 4876 3168 4910
rect 3208 4860 3218 4894
rect 3252 4860 3318 4894
rect 3352 4860 3368 4894
rect 3408 4876 3418 4910
rect 3452 4876 3518 4910
rect 3552 4876 3568 4910
rect 3608 4860 3618 4894
rect 3652 4860 3718 4894
rect 3752 4860 3768 4894
rect 3808 4876 3818 4910
rect 3852 4876 3918 4910
rect 3952 4876 3968 4910
rect 4008 4860 4018 4894
rect 4052 4860 4118 4894
rect 4152 4860 4168 4894
rect 4208 4876 4218 4910
rect 4252 4876 4318 4910
rect 4352 4876 4368 4910
rect 4408 4860 4418 4894
rect 4452 4860 4518 4894
rect 4552 4860 4568 4894
rect 4608 4876 4618 4910
rect 4652 4876 4718 4910
rect 4752 4876 4768 4910
rect 4808 4860 4818 4894
rect 4852 4860 4918 4894
rect 4952 4860 4968 4894
rect 5008 4876 5018 4910
rect 5052 4876 5118 4910
rect 5152 4876 5168 4910
rect 5208 4860 5218 4894
rect 5252 4860 5318 4894
rect 5352 4860 5368 4894
rect 5408 4876 5418 4910
rect 5452 4876 5518 4910
rect 5552 4876 5568 4910
rect 5608 4860 5618 4894
rect 5652 4860 5718 4894
rect 5752 4860 5768 4894
rect 5808 4876 5818 4910
rect 5852 4876 5918 4910
rect 5952 4876 5968 4910
rect 6008 4860 6018 4894
rect 6052 4860 6118 4894
rect 6152 4860 6168 4894
rect 6208 4876 6218 4910
rect 6252 4876 6318 4910
rect 6352 4876 6368 4910
rect 6516 4891 6568 4908
rect 6550 4874 6568 4891
rect 6602 4874 6618 4908
rect 6652 4874 6668 4908
rect 6702 4879 6720 4908
rect 6702 4874 6754 4879
rect 6862 4874 6878 4908
rect 6912 4874 6928 4908
rect 6962 4874 6978 4908
rect 7012 4874 7028 4908
rect 7062 4874 7078 4908
rect 7112 4874 7128 4908
rect 7162 4874 7178 4908
rect 7212 4874 7228 4908
rect 7262 4874 7278 4908
rect 7312 4874 7328 4908
rect 7362 4874 7378 4908
rect 7412 4874 7428 4908
rect 6 4787 64 4813
rect 6 4753 18 4787
rect 58 4753 64 4787
rect 6 4727 64 4753
rect 106 4787 164 4813
rect 106 4753 118 4787
rect 152 4753 164 4787
rect 106 4727 164 4753
rect 206 4787 264 4813
rect 206 4753 212 4787
rect 252 4753 264 4787
rect 206 4727 264 4753
rect 306 4787 364 4813
rect 306 4753 318 4787
rect 358 4753 364 4787
rect 306 4727 364 4753
rect 406 4787 464 4813
rect 406 4753 418 4787
rect 452 4753 464 4787
rect 406 4727 464 4753
rect 506 4787 564 4813
rect 506 4753 518 4787
rect 552 4753 564 4787
rect 506 4727 564 4753
rect 606 4787 664 4813
rect 606 4753 618 4787
rect 652 4753 664 4787
rect 606 4727 664 4753
rect 706 4787 764 4813
rect 706 4753 718 4787
rect 752 4753 764 4787
rect 706 4727 764 4753
rect 806 4787 864 4813
rect 806 4753 818 4787
rect 852 4753 864 4787
rect 806 4727 864 4753
rect 906 4787 964 4813
rect 906 4753 918 4787
rect 952 4753 964 4787
rect 906 4727 964 4753
rect 1006 4787 1064 4813
rect 1006 4753 1018 4787
rect 1052 4753 1064 4787
rect 1006 4727 1064 4753
rect 1106 4787 1164 4813
rect 1106 4753 1112 4787
rect 1152 4753 1164 4787
rect 1106 4727 1164 4753
rect 1206 4787 1264 4813
rect 1206 4753 1218 4787
rect 1258 4753 1264 4787
rect 1206 4727 1264 4753
rect 1306 4787 1364 4813
rect 1306 4753 1318 4787
rect 1352 4753 1364 4787
rect 1306 4727 1364 4753
rect 1406 4787 1464 4813
rect 1406 4753 1418 4787
rect 1452 4753 1464 4787
rect 1406 4727 1464 4753
rect 1506 4787 1564 4813
rect 1506 4753 1518 4787
rect 1552 4753 1564 4787
rect 1506 4727 1564 4753
rect 1606 4787 1664 4813
rect 1606 4753 1618 4787
rect 1652 4753 1664 4787
rect 1606 4727 1664 4753
rect 1706 4787 1764 4813
rect 1706 4753 1718 4787
rect 1752 4753 1764 4787
rect 1706 4727 1764 4753
rect 1806 4787 1864 4813
rect 1806 4753 1818 4787
rect 1852 4753 1864 4787
rect 1806 4727 1864 4753
rect 1906 4787 1964 4813
rect 1906 4753 1918 4787
rect 1952 4753 1964 4787
rect 1906 4727 1964 4753
rect 2006 4787 2064 4813
rect 2006 4753 2018 4787
rect 2052 4753 2064 4787
rect 2006 4727 2064 4753
rect 2106 4787 2164 4813
rect 2106 4753 2118 4787
rect 2152 4753 2164 4787
rect 2106 4727 2164 4753
rect 2206 4787 2264 4813
rect 2206 4753 2218 4787
rect 2252 4753 2264 4787
rect 2206 4727 2264 4753
rect 2306 4787 2364 4813
rect 2306 4753 2318 4787
rect 2352 4753 2364 4787
rect 2306 4727 2364 4753
rect 2406 4787 2464 4813
rect 2406 4753 2418 4787
rect 2452 4753 2464 4787
rect 2406 4727 2464 4753
rect 2506 4787 2564 4813
rect 2506 4753 2518 4787
rect 2552 4753 2564 4787
rect 2506 4727 2564 4753
rect 2606 4787 2664 4813
rect 2606 4753 2618 4787
rect 2652 4753 2664 4787
rect 2606 4727 2664 4753
rect 2706 4787 2764 4813
rect 2706 4753 2718 4787
rect 2752 4753 2764 4787
rect 2706 4727 2764 4753
rect 2806 4787 2864 4813
rect 2806 4753 2812 4787
rect 2852 4753 2864 4787
rect 2806 4727 2864 4753
rect 2906 4787 2964 4813
rect 2906 4753 2918 4787
rect 2958 4753 2964 4787
rect 2906 4727 2964 4753
rect 3006 4787 3064 4813
rect 3006 4753 3018 4787
rect 3052 4753 3064 4787
rect 3006 4727 3064 4753
rect 3106 4787 3164 4813
rect 3106 4753 3118 4787
rect 3152 4753 3164 4787
rect 3106 4727 3164 4753
rect 3206 4787 3264 4813
rect 3206 4753 3218 4787
rect 3252 4753 3264 4787
rect 3206 4727 3264 4753
rect 3306 4787 3364 4813
rect 3306 4753 3318 4787
rect 3352 4753 3364 4787
rect 3306 4727 3364 4753
rect 3406 4787 3464 4813
rect 3406 4753 3418 4787
rect 3452 4753 3464 4787
rect 3406 4727 3464 4753
rect 3506 4787 3564 4813
rect 3506 4753 3518 4787
rect 3552 4753 3564 4787
rect 3506 4727 3564 4753
rect 3606 4787 3664 4813
rect 3606 4753 3618 4787
rect 3652 4753 3664 4787
rect 3606 4727 3664 4753
rect 3706 4787 3764 4813
rect 3706 4753 3718 4787
rect 3752 4753 3764 4787
rect 3706 4727 3764 4753
rect 3806 4787 3864 4813
rect 3806 4753 3818 4787
rect 3852 4753 3864 4787
rect 3806 4727 3864 4753
rect 3906 4787 3964 4813
rect 3906 4753 3918 4787
rect 3952 4753 3964 4787
rect 3906 4727 3964 4753
rect 4006 4787 4064 4813
rect 4006 4753 4018 4787
rect 4052 4753 4064 4787
rect 4006 4727 4064 4753
rect 4106 4787 4164 4813
rect 4106 4753 4118 4787
rect 4152 4753 4164 4787
rect 4106 4727 4164 4753
rect 4206 4787 4264 4813
rect 4206 4753 4218 4787
rect 4252 4753 4264 4787
rect 4206 4727 4264 4753
rect 4306 4787 4364 4813
rect 4306 4753 4318 4787
rect 4352 4753 4364 4787
rect 4306 4727 4364 4753
rect 4406 4787 4464 4813
rect 4406 4753 4418 4787
rect 4452 4753 4464 4787
rect 4406 4727 4464 4753
rect 4506 4787 4564 4813
rect 4506 4753 4518 4787
rect 4552 4753 4564 4787
rect 4506 4727 4564 4753
rect 4606 4787 4664 4813
rect 4606 4753 4612 4787
rect 4652 4753 4664 4787
rect 4606 4727 4664 4753
rect 4706 4787 4764 4813
rect 4706 4753 4718 4787
rect 4758 4753 4764 4787
rect 4706 4727 4764 4753
rect 4806 4787 4864 4813
rect 4806 4753 4818 4787
rect 4852 4753 4864 4787
rect 4806 4727 4864 4753
rect 4906 4787 4964 4813
rect 4906 4753 4918 4787
rect 4952 4753 4964 4787
rect 4906 4727 4964 4753
rect 5006 4787 5064 4813
rect 5006 4753 5018 4787
rect 5052 4753 5064 4787
rect 5006 4727 5064 4753
rect 5106 4787 5164 4813
rect 5106 4753 5118 4787
rect 5152 4753 5164 4787
rect 5106 4727 5164 4753
rect 5206 4787 5264 4813
rect 5206 4753 5218 4787
rect 5252 4753 5264 4787
rect 5206 4727 5264 4753
rect 5306 4787 5364 4813
rect 5306 4753 5318 4787
rect 5352 4753 5364 4787
rect 5306 4727 5364 4753
rect 5406 4787 5464 4813
rect 5406 4753 5412 4787
rect 5452 4753 5464 4787
rect 5406 4727 5464 4753
rect 5506 4787 5564 4813
rect 5506 4753 5518 4787
rect 5558 4753 5564 4787
rect 5506 4727 5564 4753
rect 5606 4787 5664 4813
rect 5606 4753 5618 4787
rect 5652 4753 5664 4787
rect 5606 4727 5664 4753
rect 5706 4787 5764 4813
rect 5706 4753 5718 4787
rect 5752 4753 5764 4787
rect 5706 4727 5764 4753
rect 5806 4787 5864 4813
rect 5806 4753 5818 4787
rect 5852 4753 5864 4787
rect 5806 4727 5864 4753
rect 5906 4787 5964 4813
rect 5906 4753 5912 4787
rect 5952 4753 5964 4787
rect 5906 4727 5964 4753
rect 6006 4787 6064 4813
rect 6006 4753 6018 4787
rect 6058 4753 6064 4787
rect 6006 4727 6064 4753
rect 6106 4787 6164 4813
rect 6106 4753 6112 4787
rect 6152 4753 6164 4787
rect 6106 4727 6164 4753
rect 6206 4787 6264 4813
rect 6206 4753 6218 4787
rect 6258 4753 6264 4787
rect 6206 4727 6264 4753
rect 6306 4787 6364 4813
rect 6306 4753 6318 4787
rect 6352 4753 6364 4787
rect 6306 4727 6364 4753
rect 6406 4787 6464 4813
rect 6618 4806 6862 4840
rect 6406 4753 6418 4787
rect 6452 4753 6464 4787
rect 6508 4768 6516 4802
rect 6558 4768 6574 4802
rect 6618 4787 6652 4806
rect 6406 4727 6464 4753
rect 6828 4803 6862 4806
rect 6828 4787 6962 4803
rect 6618 4737 6652 4753
rect 6696 4738 6712 4772
rect 6754 4738 6762 4772
rect 6862 4753 6928 4787
rect 6828 4737 6962 4753
rect 7028 4787 7162 4803
rect 7062 4753 7128 4787
rect 7028 4737 7162 4753
rect 7228 4787 7362 4803
rect 7262 4753 7328 4787
rect 7228 4737 7362 4753
rect 7428 4787 7462 4803
rect 7428 4737 7462 4753
rect 6 4647 64 4673
rect 6 4613 18 4647
rect 58 4613 64 4647
rect 6 4587 64 4613
rect 106 4647 164 4673
rect 106 4613 118 4647
rect 152 4613 164 4647
rect 106 4587 164 4613
rect 206 4647 264 4673
rect 206 4613 218 4647
rect 252 4613 264 4647
rect 206 4587 264 4613
rect 306 4647 364 4673
rect 306 4613 318 4647
rect 352 4613 364 4647
rect 306 4587 364 4613
rect 406 4647 464 4673
rect 406 4613 418 4647
rect 452 4613 464 4647
rect 406 4587 464 4613
rect 506 4647 564 4673
rect 506 4613 518 4647
rect 552 4613 564 4647
rect 506 4587 564 4613
rect 606 4647 664 4673
rect 606 4613 618 4647
rect 652 4613 664 4647
rect 606 4587 664 4613
rect 706 4647 764 4673
rect 706 4613 718 4647
rect 752 4613 764 4647
rect 706 4587 764 4613
rect 806 4647 864 4673
rect 806 4613 818 4647
rect 852 4613 864 4647
rect 806 4587 864 4613
rect 906 4647 964 4673
rect 906 4613 918 4647
rect 952 4613 964 4647
rect 906 4587 964 4613
rect 1006 4647 1064 4673
rect 1006 4613 1018 4647
rect 1052 4613 1064 4647
rect 1006 4587 1064 4613
rect 1106 4647 1164 4673
rect 1106 4613 1118 4647
rect 1152 4613 1164 4647
rect 1106 4587 1164 4613
rect 1206 4647 1264 4673
rect 1206 4613 1218 4647
rect 1252 4613 1264 4647
rect 1206 4587 1264 4613
rect 1306 4647 1364 4673
rect 1306 4613 1318 4647
rect 1352 4613 1364 4647
rect 1306 4587 1364 4613
rect 1406 4647 1464 4673
rect 1406 4613 1418 4647
rect 1452 4613 1464 4647
rect 1406 4587 1464 4613
rect 1506 4647 1564 4673
rect 1506 4613 1518 4647
rect 1552 4613 1564 4647
rect 1506 4587 1564 4613
rect 1606 4647 1664 4673
rect 1606 4613 1618 4647
rect 1652 4613 1664 4647
rect 1606 4587 1664 4613
rect 1706 4647 1764 4673
rect 1706 4613 1718 4647
rect 1752 4613 1764 4647
rect 1706 4587 1764 4613
rect 1806 4647 1864 4673
rect 1806 4613 1812 4647
rect 1852 4613 1864 4647
rect 1806 4587 1864 4613
rect 1906 4647 1964 4673
rect 1906 4613 1918 4647
rect 1958 4613 1964 4647
rect 1906 4587 1964 4613
rect 2006 4647 2064 4673
rect 2006 4613 2012 4647
rect 2052 4613 2064 4647
rect 2006 4587 2064 4613
rect 2106 4647 2164 4673
rect 2106 4613 2118 4647
rect 2158 4613 2164 4647
rect 2106 4587 2164 4613
rect 2206 4647 2264 4673
rect 2206 4613 2218 4647
rect 2252 4613 2264 4647
rect 2206 4587 2264 4613
rect 2306 4647 2364 4673
rect 2306 4613 2318 4647
rect 2352 4613 2364 4647
rect 2306 4587 2364 4613
rect 2406 4647 2464 4673
rect 2406 4613 2418 4647
rect 2452 4613 2464 4647
rect 2406 4587 2464 4613
rect 2506 4647 2564 4673
rect 2506 4613 2518 4647
rect 2552 4613 2564 4647
rect 2506 4587 2564 4613
rect 2606 4647 2664 4673
rect 2606 4613 2618 4647
rect 2652 4613 2664 4647
rect 2606 4587 2664 4613
rect 2706 4647 2764 4673
rect 2706 4613 2718 4647
rect 2752 4613 2764 4647
rect 2706 4587 2764 4613
rect 2806 4647 2864 4673
rect 2806 4613 2818 4647
rect 2852 4613 2864 4647
rect 2806 4587 2864 4613
rect 2906 4647 2964 4673
rect 2906 4613 2918 4647
rect 2952 4613 2964 4647
rect 2906 4587 2964 4613
rect 3006 4647 3064 4673
rect 3006 4613 3018 4647
rect 3052 4613 3064 4647
rect 3006 4587 3064 4613
rect 3106 4647 3164 4673
rect 3106 4613 3118 4647
rect 3152 4613 3164 4647
rect 3106 4587 3164 4613
rect 3206 4647 3264 4673
rect 3206 4613 3212 4647
rect 3252 4613 3264 4647
rect 3206 4587 3264 4613
rect 3306 4647 3364 4673
rect 3306 4613 3318 4647
rect 3358 4613 3364 4647
rect 3306 4587 3364 4613
rect 3406 4647 3464 4673
rect 3406 4613 3418 4647
rect 3452 4613 3464 4647
rect 3406 4587 3464 4613
rect 3506 4647 3564 4673
rect 3506 4613 3518 4647
rect 3552 4613 3564 4647
rect 3506 4587 3564 4613
rect 3606 4647 3664 4673
rect 3606 4613 3618 4647
rect 3652 4613 3664 4647
rect 3606 4587 3664 4613
rect 3706 4647 3764 4673
rect 3706 4613 3718 4647
rect 3752 4613 3764 4647
rect 3706 4587 3764 4613
rect 3806 4647 3864 4673
rect 3806 4613 3818 4647
rect 3852 4613 3864 4647
rect 3806 4587 3864 4613
rect 3906 4647 3964 4673
rect 3906 4613 3918 4647
rect 3952 4613 3964 4647
rect 3906 4587 3964 4613
rect 4006 4647 4064 4673
rect 4006 4613 4018 4647
rect 4052 4613 4064 4647
rect 4006 4587 4064 4613
rect 4106 4647 4164 4673
rect 4106 4613 4118 4647
rect 4152 4613 4164 4647
rect 4106 4587 4164 4613
rect 4206 4647 4264 4673
rect 4206 4613 4218 4647
rect 4252 4613 4264 4647
rect 4206 4587 4264 4613
rect 4306 4647 4364 4673
rect 4306 4613 4318 4647
rect 4352 4613 4364 4647
rect 4306 4587 4364 4613
rect 4406 4647 4464 4673
rect 4406 4613 4418 4647
rect 4452 4613 4464 4647
rect 4406 4587 4464 4613
rect 4506 4647 4564 4673
rect 4506 4613 4512 4647
rect 4552 4613 4564 4647
rect 4506 4587 4564 4613
rect 4606 4647 4664 4673
rect 4606 4613 4618 4647
rect 4658 4613 4664 4647
rect 4606 4587 4664 4613
rect 4706 4647 4764 4673
rect 4706 4613 4718 4647
rect 4752 4613 4764 4647
rect 4706 4587 4764 4613
rect 4806 4647 4864 4673
rect 4806 4613 4818 4647
rect 4852 4613 4864 4647
rect 4806 4587 4864 4613
rect 4906 4647 4964 4673
rect 4906 4613 4918 4647
rect 4952 4613 4964 4647
rect 4906 4587 4964 4613
rect 5006 4647 5064 4673
rect 5006 4613 5018 4647
rect 5052 4613 5064 4647
rect 5006 4587 5064 4613
rect 5106 4647 5164 4673
rect 5106 4613 5118 4647
rect 5152 4613 5164 4647
rect 5106 4587 5164 4613
rect 5206 4647 5264 4673
rect 5206 4613 5218 4647
rect 5252 4613 5264 4647
rect 5206 4587 5264 4613
rect 5306 4647 5364 4673
rect 5306 4613 5318 4647
rect 5352 4613 5364 4647
rect 5306 4587 5364 4613
rect 5406 4647 5464 4673
rect 5406 4613 5418 4647
rect 5452 4613 5464 4647
rect 5406 4587 5464 4613
rect 5506 4647 5564 4673
rect 5506 4613 5518 4647
rect 5552 4613 5564 4647
rect 5506 4587 5564 4613
rect 5606 4647 5664 4673
rect 5606 4613 5618 4647
rect 5652 4613 5664 4647
rect 5606 4587 5664 4613
rect 5706 4647 5764 4673
rect 5706 4613 5718 4647
rect 5752 4613 5764 4647
rect 5706 4587 5764 4613
rect 5806 4647 5864 4673
rect 5806 4613 5818 4647
rect 5852 4613 5864 4647
rect 5806 4587 5864 4613
rect 5906 4647 5964 4673
rect 5906 4613 5918 4647
rect 5952 4613 5964 4647
rect 5906 4587 5964 4613
rect 6006 4647 6064 4673
rect 6006 4613 6012 4647
rect 6052 4613 6064 4647
rect 6006 4587 6064 4613
rect 6106 4647 6164 4673
rect 6106 4613 6118 4647
rect 6158 4613 6164 4647
rect 6106 4587 6164 4613
rect 6206 4647 6264 4673
rect 6206 4613 6212 4647
rect 6252 4613 6264 4647
rect 6206 4587 6264 4613
rect 6306 4647 6364 4673
rect 6306 4613 6318 4647
rect 6358 4613 6364 4647
rect 6306 4587 6364 4613
rect 6406 4647 6464 4673
rect 6618 4666 6862 4700
rect 6406 4613 6412 4647
rect 6452 4613 6464 4647
rect 6508 4628 6516 4662
rect 6558 4628 6574 4662
rect 6618 4647 6652 4666
rect 6406 4587 6464 4613
rect 6828 4647 6862 4666
rect 6618 4597 6652 4613
rect 6696 4598 6712 4632
rect 6754 4598 6762 4632
rect 6828 4597 6862 4613
rect 6928 4647 7162 4663
rect 6962 4613 7028 4647
rect 7062 4613 7128 4647
rect 6928 4597 7162 4613
rect 7228 4647 7362 4663
rect 7262 4613 7328 4647
rect 7228 4597 7362 4613
rect 7428 4647 7462 4663
rect 7428 4597 7462 4613
rect 6 4507 64 4533
rect 6 4473 18 4507
rect 58 4473 64 4507
rect 6 4447 64 4473
rect 106 4507 164 4533
rect 106 4473 112 4507
rect 152 4473 164 4507
rect 106 4447 164 4473
rect 206 4507 264 4533
rect 206 4473 218 4507
rect 258 4473 264 4507
rect 206 4447 264 4473
rect 306 4507 364 4533
rect 306 4473 318 4507
rect 352 4473 364 4507
rect 306 4447 364 4473
rect 406 4507 464 4533
rect 406 4473 418 4507
rect 452 4473 464 4507
rect 406 4447 464 4473
rect 506 4507 564 4533
rect 506 4473 518 4507
rect 552 4473 564 4507
rect 506 4447 564 4473
rect 606 4507 664 4533
rect 606 4473 618 4507
rect 652 4473 664 4507
rect 606 4447 664 4473
rect 706 4507 764 4533
rect 706 4473 718 4507
rect 752 4473 764 4507
rect 706 4447 764 4473
rect 806 4507 864 4533
rect 806 4473 818 4507
rect 852 4473 864 4507
rect 806 4447 864 4473
rect 906 4507 964 4533
rect 906 4473 918 4507
rect 952 4473 964 4507
rect 906 4447 964 4473
rect 1006 4507 1064 4533
rect 1006 4473 1018 4507
rect 1052 4473 1064 4507
rect 1006 4447 1064 4473
rect 1106 4507 1164 4533
rect 1106 4473 1118 4507
rect 1152 4473 1164 4507
rect 1106 4447 1164 4473
rect 1206 4507 1264 4533
rect 1206 4473 1218 4507
rect 1252 4473 1264 4507
rect 1206 4447 1264 4473
rect 1306 4507 1364 4533
rect 1306 4473 1318 4507
rect 1352 4473 1364 4507
rect 1306 4447 1364 4473
rect 1406 4507 1464 4533
rect 1406 4473 1418 4507
rect 1452 4473 1464 4507
rect 1406 4447 1464 4473
rect 1506 4507 1564 4533
rect 1506 4473 1518 4507
rect 1552 4473 1564 4507
rect 1506 4447 1564 4473
rect 1606 4507 1664 4533
rect 1606 4473 1612 4507
rect 1652 4473 1664 4507
rect 1606 4447 1664 4473
rect 1706 4507 1764 4533
rect 1706 4473 1718 4507
rect 1758 4473 1764 4507
rect 1706 4447 1764 4473
rect 1806 4507 1864 4533
rect 1806 4473 1818 4507
rect 1852 4473 1864 4507
rect 1806 4447 1864 4473
rect 1906 4507 1964 4533
rect 1906 4473 1918 4507
rect 1952 4473 1964 4507
rect 1906 4447 1964 4473
rect 2006 4507 2064 4533
rect 2006 4473 2018 4507
rect 2052 4473 2064 4507
rect 2006 4447 2064 4473
rect 2106 4507 2164 4533
rect 2106 4473 2118 4507
rect 2152 4473 2164 4507
rect 2106 4447 2164 4473
rect 2206 4507 2264 4533
rect 2206 4473 2218 4507
rect 2252 4473 2264 4507
rect 2206 4447 2264 4473
rect 2306 4507 2364 4533
rect 2306 4473 2318 4507
rect 2352 4473 2364 4507
rect 2306 4447 2364 4473
rect 2406 4507 2464 4533
rect 2406 4473 2412 4507
rect 2452 4473 2464 4507
rect 2406 4447 2464 4473
rect 2506 4507 2564 4533
rect 2506 4473 2518 4507
rect 2558 4473 2564 4507
rect 2506 4447 2564 4473
rect 2606 4507 2664 4533
rect 2606 4473 2618 4507
rect 2652 4473 2664 4507
rect 2606 4447 2664 4473
rect 2706 4507 2764 4533
rect 2706 4473 2718 4507
rect 2752 4473 2764 4507
rect 2706 4447 2764 4473
rect 2806 4507 2864 4533
rect 2806 4473 2818 4507
rect 2852 4473 2864 4507
rect 2806 4447 2864 4473
rect 2906 4507 2964 4533
rect 2906 4473 2918 4507
rect 2952 4473 2964 4507
rect 2906 4447 2964 4473
rect 3006 4507 3064 4533
rect 3006 4473 3018 4507
rect 3052 4473 3064 4507
rect 3006 4447 3064 4473
rect 3106 4507 3164 4533
rect 3106 4473 3118 4507
rect 3152 4473 3164 4507
rect 3106 4447 3164 4473
rect 3206 4507 3264 4533
rect 3206 4473 3218 4507
rect 3252 4473 3264 4507
rect 3206 4447 3264 4473
rect 3306 4507 3364 4533
rect 3306 4473 3312 4507
rect 3352 4473 3364 4507
rect 3306 4447 3364 4473
rect 3406 4507 3464 4533
rect 3406 4473 3418 4507
rect 3458 4473 3464 4507
rect 3406 4447 3464 4473
rect 3506 4507 3564 4533
rect 3506 4473 3518 4507
rect 3552 4473 3564 4507
rect 3506 4447 3564 4473
rect 3606 4507 3664 4533
rect 3606 4473 3618 4507
rect 3652 4473 3664 4507
rect 3606 4447 3664 4473
rect 3706 4507 3764 4533
rect 3706 4473 3718 4507
rect 3752 4473 3764 4507
rect 3706 4447 3764 4473
rect 3806 4507 3864 4533
rect 3806 4473 3818 4507
rect 3852 4473 3864 4507
rect 3806 4447 3864 4473
rect 3906 4507 3964 4533
rect 3906 4473 3918 4507
rect 3952 4473 3964 4507
rect 3906 4447 3964 4473
rect 4006 4507 4064 4533
rect 4006 4473 4018 4507
rect 4052 4473 4064 4507
rect 4006 4447 4064 4473
rect 4106 4507 4164 4533
rect 4106 4473 4118 4507
rect 4152 4473 4164 4507
rect 4106 4447 4164 4473
rect 4206 4507 4264 4533
rect 4206 4473 4218 4507
rect 4252 4473 4264 4507
rect 4206 4447 4264 4473
rect 4306 4507 4364 4533
rect 4306 4473 4312 4507
rect 4352 4473 4364 4507
rect 4306 4447 4364 4473
rect 4406 4507 4464 4533
rect 4406 4473 4418 4507
rect 4458 4473 4464 4507
rect 4406 4447 4464 4473
rect 4506 4507 4564 4533
rect 4506 4473 4518 4507
rect 4552 4473 4564 4507
rect 4506 4447 4564 4473
rect 4606 4507 4664 4533
rect 4606 4473 4618 4507
rect 4652 4473 4664 4507
rect 4606 4447 4664 4473
rect 4706 4507 4764 4533
rect 4706 4473 4718 4507
rect 4752 4473 4764 4507
rect 4706 4447 4764 4473
rect 4806 4507 4864 4533
rect 4806 4473 4818 4507
rect 4852 4473 4864 4507
rect 4806 4447 4864 4473
rect 4906 4507 4964 4533
rect 4906 4473 4918 4507
rect 4952 4473 4964 4507
rect 4906 4447 4964 4473
rect 5006 4507 5064 4533
rect 5006 4473 5018 4507
rect 5052 4473 5064 4507
rect 5006 4447 5064 4473
rect 5106 4507 5164 4533
rect 5106 4473 5118 4507
rect 5152 4473 5164 4507
rect 5106 4447 5164 4473
rect 5206 4507 5264 4533
rect 5206 4473 5212 4507
rect 5252 4473 5264 4507
rect 5206 4447 5264 4473
rect 5306 4507 5364 4533
rect 5306 4473 5318 4507
rect 5358 4473 5364 4507
rect 5306 4447 5364 4473
rect 5406 4507 5464 4533
rect 5406 4473 5418 4507
rect 5452 4473 5464 4507
rect 5406 4447 5464 4473
rect 5506 4507 5564 4533
rect 5506 4473 5518 4507
rect 5552 4473 5564 4507
rect 5506 4447 5564 4473
rect 5606 4507 5664 4533
rect 5606 4473 5618 4507
rect 5652 4473 5664 4507
rect 5606 4447 5664 4473
rect 5706 4507 5764 4533
rect 5706 4473 5712 4507
rect 5752 4473 5764 4507
rect 5706 4447 5764 4473
rect 5806 4507 5864 4533
rect 5806 4473 5818 4507
rect 5858 4473 5864 4507
rect 5806 4447 5864 4473
rect 5906 4507 5964 4533
rect 5906 4473 5918 4507
rect 5952 4473 5964 4507
rect 5906 4447 5964 4473
rect 6006 4507 6064 4533
rect 6006 4473 6018 4507
rect 6052 4473 6064 4507
rect 6006 4447 6064 4473
rect 6106 4507 6164 4533
rect 6106 4473 6118 4507
rect 6152 4473 6164 4507
rect 6106 4447 6164 4473
rect 6206 4507 6264 4533
rect 6206 4473 6212 4507
rect 6252 4473 6264 4507
rect 6206 4447 6264 4473
rect 6306 4507 6364 4533
rect 6306 4473 6318 4507
rect 6358 4473 6364 4507
rect 6306 4447 6364 4473
rect 6406 4507 6464 4533
rect 6618 4526 6862 4560
rect 6406 4473 6412 4507
rect 6452 4473 6464 4507
rect 6508 4488 6516 4522
rect 6558 4488 6574 4522
rect 6618 4507 6652 4526
rect 6406 4447 6464 4473
rect 6828 4523 6862 4526
rect 6828 4507 6962 4523
rect 6618 4457 6652 4473
rect 6696 4458 6712 4492
rect 6754 4458 6762 4492
rect 6862 4473 6928 4507
rect 6828 4457 6962 4473
rect 7028 4507 7062 4523
rect 7028 4457 7062 4473
rect 7128 4507 7362 4523
rect 7162 4473 7228 4507
rect 7262 4473 7328 4507
rect 7128 4457 7362 4473
rect 7428 4507 7462 4523
rect 7428 4457 7462 4473
rect 6 4367 64 4393
rect 6 4333 18 4367
rect 58 4333 64 4367
rect 6 4307 64 4333
rect 106 4367 164 4393
rect 106 4333 118 4367
rect 152 4333 164 4367
rect 106 4307 164 4333
rect 206 4367 264 4393
rect 206 4333 218 4367
rect 252 4333 264 4367
rect 206 4307 264 4333
rect 306 4367 364 4393
rect 306 4333 318 4367
rect 352 4333 364 4367
rect 306 4307 364 4333
rect 406 4367 464 4393
rect 406 4333 412 4367
rect 452 4333 464 4367
rect 406 4307 464 4333
rect 506 4367 564 4393
rect 506 4333 518 4367
rect 558 4333 564 4367
rect 506 4307 564 4333
rect 606 4367 664 4393
rect 606 4333 618 4367
rect 652 4333 664 4367
rect 606 4307 664 4333
rect 706 4367 764 4393
rect 706 4333 712 4367
rect 752 4333 764 4367
rect 706 4307 764 4333
rect 806 4367 864 4393
rect 806 4333 818 4367
rect 858 4333 864 4367
rect 806 4307 864 4333
rect 906 4367 964 4393
rect 906 4333 918 4367
rect 952 4333 964 4367
rect 906 4307 964 4333
rect 1006 4367 1064 4393
rect 1006 4333 1018 4367
rect 1052 4333 1064 4367
rect 1006 4307 1064 4333
rect 1106 4367 1164 4393
rect 1106 4333 1118 4367
rect 1152 4333 1164 4367
rect 1106 4307 1164 4333
rect 1206 4367 1264 4393
rect 1206 4333 1218 4367
rect 1252 4333 1264 4367
rect 1206 4307 1264 4333
rect 1306 4367 1364 4393
rect 1306 4333 1318 4367
rect 1352 4333 1364 4367
rect 1306 4307 1364 4333
rect 1406 4367 1464 4393
rect 1406 4333 1418 4367
rect 1452 4333 1464 4367
rect 1406 4307 1464 4333
rect 1506 4367 1564 4393
rect 1506 4333 1518 4367
rect 1552 4333 1564 4367
rect 1506 4307 1564 4333
rect 1606 4367 1664 4393
rect 1606 4333 1618 4367
rect 1652 4333 1664 4367
rect 1606 4307 1664 4333
rect 1706 4367 1764 4393
rect 1706 4333 1718 4367
rect 1752 4333 1764 4367
rect 1706 4307 1764 4333
rect 1806 4367 1864 4393
rect 1806 4333 1818 4367
rect 1852 4333 1864 4367
rect 1806 4307 1864 4333
rect 1906 4367 1964 4393
rect 1906 4333 1918 4367
rect 1952 4333 1964 4367
rect 1906 4307 1964 4333
rect 2006 4367 2064 4393
rect 2006 4333 2018 4367
rect 2052 4333 2064 4367
rect 2006 4307 2064 4333
rect 2106 4367 2164 4393
rect 2106 4333 2118 4367
rect 2152 4333 2164 4367
rect 2106 4307 2164 4333
rect 2206 4367 2264 4393
rect 2206 4333 2218 4367
rect 2252 4333 2264 4367
rect 2206 4307 2264 4333
rect 2306 4367 2364 4393
rect 2306 4333 2318 4367
rect 2352 4333 2364 4367
rect 2306 4307 2364 4333
rect 2406 4367 2464 4393
rect 2406 4333 2412 4367
rect 2452 4333 2464 4367
rect 2406 4307 2464 4333
rect 2506 4367 2564 4393
rect 2506 4333 2518 4367
rect 2558 4333 2564 4367
rect 2506 4307 2564 4333
rect 2606 4367 2664 4393
rect 2606 4333 2618 4367
rect 2652 4333 2664 4367
rect 2606 4307 2664 4333
rect 2706 4367 2764 4393
rect 2706 4333 2718 4367
rect 2752 4333 2764 4367
rect 2706 4307 2764 4333
rect 2806 4367 2864 4393
rect 2806 4333 2812 4367
rect 2852 4333 2864 4367
rect 2806 4307 2864 4333
rect 2906 4367 2964 4393
rect 2906 4333 2918 4367
rect 2958 4333 2964 4367
rect 2906 4307 2964 4333
rect 3006 4367 3064 4393
rect 3006 4333 3018 4367
rect 3052 4333 3064 4367
rect 3006 4307 3064 4333
rect 3106 4367 3164 4393
rect 3106 4333 3118 4367
rect 3152 4333 3164 4367
rect 3106 4307 3164 4333
rect 3206 4367 3264 4393
rect 3206 4333 3212 4367
rect 3252 4333 3264 4367
rect 3206 4307 3264 4333
rect 3306 4367 3364 4393
rect 3306 4333 3318 4367
rect 3358 4333 3364 4367
rect 3306 4307 3364 4333
rect 3406 4367 3464 4393
rect 3406 4333 3418 4367
rect 3452 4333 3464 4367
rect 3406 4307 3464 4333
rect 3506 4367 3564 4393
rect 3506 4333 3518 4367
rect 3552 4333 3564 4367
rect 3506 4307 3564 4333
rect 3606 4367 3664 4393
rect 3606 4333 3618 4367
rect 3652 4333 3664 4367
rect 3606 4307 3664 4333
rect 3706 4367 3764 4393
rect 3706 4333 3718 4367
rect 3752 4333 3764 4367
rect 3706 4307 3764 4333
rect 3806 4367 3864 4393
rect 3806 4333 3818 4367
rect 3852 4333 3864 4367
rect 3806 4307 3864 4333
rect 3906 4367 3964 4393
rect 3906 4333 3918 4367
rect 3952 4333 3964 4367
rect 3906 4307 3964 4333
rect 4006 4367 4064 4393
rect 4006 4333 4018 4367
rect 4052 4333 4064 4367
rect 4006 4307 4064 4333
rect 4106 4367 4164 4393
rect 4106 4333 4118 4367
rect 4152 4333 4164 4367
rect 4106 4307 4164 4333
rect 4206 4367 4264 4393
rect 4206 4333 4218 4367
rect 4252 4333 4264 4367
rect 4206 4307 4264 4333
rect 4306 4367 4364 4393
rect 4306 4333 4318 4367
rect 4352 4333 4364 4367
rect 4306 4307 4364 4333
rect 4406 4367 4464 4393
rect 4406 4333 4418 4367
rect 4452 4333 4464 4367
rect 4406 4307 4464 4333
rect 4506 4367 4564 4393
rect 4506 4333 4518 4367
rect 4552 4333 4564 4367
rect 4506 4307 4564 4333
rect 4606 4367 4664 4393
rect 4606 4333 4618 4367
rect 4652 4333 4664 4367
rect 4606 4307 4664 4333
rect 4706 4367 4764 4393
rect 4706 4333 4718 4367
rect 4752 4333 4764 4367
rect 4706 4307 4764 4333
rect 4806 4367 4864 4393
rect 4806 4333 4818 4367
rect 4852 4333 4864 4367
rect 4806 4307 4864 4333
rect 4906 4367 4964 4393
rect 4906 4333 4918 4367
rect 4952 4333 4964 4367
rect 4906 4307 4964 4333
rect 5006 4367 5064 4393
rect 5006 4333 5012 4367
rect 5052 4333 5064 4367
rect 5006 4307 5064 4333
rect 5106 4367 5164 4393
rect 5106 4333 5118 4367
rect 5158 4333 5164 4367
rect 5106 4307 5164 4333
rect 5206 4367 5264 4393
rect 5206 4333 5218 4367
rect 5252 4333 5264 4367
rect 5206 4307 5264 4333
rect 5306 4367 5364 4393
rect 5306 4333 5318 4367
rect 5352 4333 5364 4367
rect 5306 4307 5364 4333
rect 5406 4367 5464 4393
rect 5406 4333 5412 4367
rect 5452 4333 5464 4367
rect 5406 4307 5464 4333
rect 5506 4367 5564 4393
rect 5506 4333 5518 4367
rect 5558 4333 5564 4367
rect 5506 4307 5564 4333
rect 5606 4367 5664 4393
rect 5606 4333 5618 4367
rect 5652 4333 5664 4367
rect 5606 4307 5664 4333
rect 5706 4367 5764 4393
rect 5706 4333 5718 4367
rect 5752 4333 5764 4367
rect 5706 4307 5764 4333
rect 5806 4367 5864 4393
rect 5806 4333 5818 4367
rect 5852 4333 5864 4367
rect 5806 4307 5864 4333
rect 5906 4367 5964 4393
rect 5906 4333 5918 4367
rect 5952 4333 5964 4367
rect 5906 4307 5964 4333
rect 6006 4367 6064 4393
rect 6006 4333 6012 4367
rect 6052 4333 6064 4367
rect 6006 4307 6064 4333
rect 6106 4367 6164 4393
rect 6106 4333 6118 4367
rect 6158 4333 6164 4367
rect 6106 4307 6164 4333
rect 6206 4367 6264 4393
rect 6206 4333 6212 4367
rect 6252 4333 6264 4367
rect 6206 4307 6264 4333
rect 6306 4367 6364 4393
rect 6306 4333 6318 4367
rect 6358 4333 6364 4367
rect 6306 4307 6364 4333
rect 6406 4367 6464 4393
rect 6618 4386 6862 4420
rect 6406 4333 6412 4367
rect 6452 4333 6464 4367
rect 6508 4348 6516 4382
rect 6558 4348 6574 4382
rect 6618 4367 6652 4386
rect 6406 4307 6464 4333
rect 6828 4367 6862 4386
rect 6618 4317 6652 4333
rect 6696 4318 6712 4352
rect 6754 4318 6762 4352
rect 6828 4317 6862 4333
rect 6928 4367 7062 4383
rect 6962 4333 7028 4367
rect 6928 4317 7062 4333
rect 7128 4367 7362 4383
rect 7162 4333 7228 4367
rect 7262 4333 7328 4367
rect 7128 4317 7362 4333
rect 7428 4367 7462 4383
rect 7428 4317 7462 4333
rect 6 4227 64 4253
rect 6 4193 18 4227
rect 58 4193 64 4227
rect 6 4167 64 4193
rect 106 4227 164 4253
rect 106 4193 112 4227
rect 152 4193 164 4227
rect 106 4167 164 4193
rect 206 4227 264 4253
rect 206 4193 218 4227
rect 258 4193 264 4227
rect 206 4167 264 4193
rect 306 4227 364 4253
rect 306 4193 312 4227
rect 352 4193 364 4227
rect 306 4167 364 4193
rect 406 4227 464 4253
rect 406 4193 418 4227
rect 458 4193 464 4227
rect 406 4167 464 4193
rect 506 4227 564 4253
rect 506 4193 518 4227
rect 552 4193 564 4227
rect 506 4167 564 4193
rect 606 4227 664 4253
rect 606 4193 618 4227
rect 652 4193 664 4227
rect 606 4167 664 4193
rect 706 4227 764 4253
rect 706 4193 718 4227
rect 752 4193 764 4227
rect 706 4167 764 4193
rect 806 4227 864 4253
rect 806 4193 818 4227
rect 852 4193 864 4227
rect 806 4167 864 4193
rect 906 4227 964 4253
rect 906 4193 918 4227
rect 952 4193 964 4227
rect 906 4167 964 4193
rect 1006 4227 1064 4253
rect 1006 4193 1018 4227
rect 1052 4193 1064 4227
rect 1006 4167 1064 4193
rect 1106 4227 1164 4253
rect 1106 4193 1118 4227
rect 1152 4193 1164 4227
rect 1106 4167 1164 4193
rect 1206 4227 1264 4253
rect 1206 4193 1218 4227
rect 1252 4193 1264 4227
rect 1206 4167 1264 4193
rect 1306 4227 1364 4253
rect 1306 4193 1318 4227
rect 1352 4193 1364 4227
rect 1306 4167 1364 4193
rect 1406 4227 1464 4253
rect 1406 4193 1412 4227
rect 1452 4193 1464 4227
rect 1406 4167 1464 4193
rect 1506 4227 1564 4253
rect 1506 4193 1518 4227
rect 1558 4193 1564 4227
rect 1506 4167 1564 4193
rect 1606 4227 1664 4253
rect 1606 4193 1618 4227
rect 1652 4193 1664 4227
rect 1606 4167 1664 4193
rect 1706 4227 1764 4253
rect 1706 4193 1718 4227
rect 1752 4193 1764 4227
rect 1706 4167 1764 4193
rect 1806 4227 1864 4253
rect 1806 4193 1818 4227
rect 1852 4193 1864 4227
rect 1806 4167 1864 4193
rect 1906 4227 1964 4253
rect 1906 4193 1918 4227
rect 1952 4193 1964 4227
rect 1906 4167 1964 4193
rect 2006 4227 2064 4253
rect 2006 4193 2018 4227
rect 2052 4193 2064 4227
rect 2006 4167 2064 4193
rect 2106 4227 2164 4253
rect 2106 4193 2118 4227
rect 2152 4193 2164 4227
rect 2106 4167 2164 4193
rect 2206 4227 2264 4253
rect 2206 4193 2218 4227
rect 2252 4193 2264 4227
rect 2206 4167 2264 4193
rect 2306 4227 2364 4253
rect 2306 4193 2318 4227
rect 2352 4193 2364 4227
rect 2306 4167 2364 4193
rect 2406 4227 2464 4253
rect 2406 4193 2418 4227
rect 2452 4193 2464 4227
rect 2406 4167 2464 4193
rect 2506 4227 2564 4253
rect 2506 4193 2518 4227
rect 2552 4193 2564 4227
rect 2506 4167 2564 4193
rect 2606 4227 2664 4253
rect 2606 4193 2618 4227
rect 2652 4193 2664 4227
rect 2606 4167 2664 4193
rect 2706 4227 2764 4253
rect 2706 4193 2718 4227
rect 2752 4193 2764 4227
rect 2706 4167 2764 4193
rect 2806 4227 2864 4253
rect 2806 4193 2818 4227
rect 2852 4193 2864 4227
rect 2806 4167 2864 4193
rect 2906 4227 2964 4253
rect 2906 4193 2918 4227
rect 2952 4193 2964 4227
rect 2906 4167 2964 4193
rect 3006 4227 3064 4253
rect 3006 4193 3018 4227
rect 3052 4193 3064 4227
rect 3006 4167 3064 4193
rect 3106 4227 3164 4253
rect 3106 4193 3118 4227
rect 3152 4193 3164 4227
rect 3106 4167 3164 4193
rect 3206 4227 3264 4253
rect 3206 4193 3218 4227
rect 3252 4193 3264 4227
rect 3206 4167 3264 4193
rect 3306 4227 3364 4253
rect 3306 4193 3318 4227
rect 3352 4193 3364 4227
rect 3306 4167 3364 4193
rect 3406 4227 3464 4253
rect 3406 4193 3412 4227
rect 3452 4193 3464 4227
rect 3406 4167 3464 4193
rect 3506 4227 3564 4253
rect 3506 4193 3518 4227
rect 3558 4193 3564 4227
rect 3506 4167 3564 4193
rect 3606 4227 3664 4253
rect 3606 4193 3612 4227
rect 3652 4193 3664 4227
rect 3606 4167 3664 4193
rect 3706 4227 3764 4253
rect 3706 4193 3718 4227
rect 3758 4193 3764 4227
rect 3706 4167 3764 4193
rect 3806 4227 3864 4253
rect 3806 4193 3818 4227
rect 3852 4193 3864 4227
rect 3806 4167 3864 4193
rect 3906 4227 3964 4253
rect 3906 4193 3918 4227
rect 3952 4193 3964 4227
rect 3906 4167 3964 4193
rect 4006 4227 4064 4253
rect 4006 4193 4018 4227
rect 4052 4193 4064 4227
rect 4006 4167 4064 4193
rect 4106 4227 4164 4253
rect 4106 4193 4118 4227
rect 4152 4193 4164 4227
rect 4106 4167 4164 4193
rect 4206 4227 4264 4253
rect 4206 4193 4218 4227
rect 4252 4193 4264 4227
rect 4206 4167 4264 4193
rect 4306 4227 4364 4253
rect 4306 4193 4318 4227
rect 4352 4193 4364 4227
rect 4306 4167 4364 4193
rect 4406 4227 4464 4253
rect 4406 4193 4412 4227
rect 4452 4193 4464 4227
rect 4406 4167 4464 4193
rect 4506 4227 4564 4253
rect 4506 4193 4518 4227
rect 4558 4193 4564 4227
rect 4506 4167 4564 4193
rect 4606 4227 4664 4253
rect 4606 4193 4618 4227
rect 4652 4193 4664 4227
rect 4606 4167 4664 4193
rect 4706 4227 4764 4253
rect 4706 4193 4718 4227
rect 4752 4193 4764 4227
rect 4706 4167 4764 4193
rect 4806 4227 4864 4253
rect 4806 4193 4818 4227
rect 4852 4193 4864 4227
rect 4806 4167 4864 4193
rect 4906 4227 4964 4253
rect 4906 4193 4918 4227
rect 4952 4193 4964 4227
rect 4906 4167 4964 4193
rect 5006 4227 5064 4253
rect 5006 4193 5012 4227
rect 5052 4193 5064 4227
rect 5006 4167 5064 4193
rect 5106 4227 5164 4253
rect 5106 4193 5118 4227
rect 5158 4193 5164 4227
rect 5106 4167 5164 4193
rect 5206 4227 5264 4253
rect 5206 4193 5218 4227
rect 5252 4193 5264 4227
rect 5206 4167 5264 4193
rect 5306 4227 5364 4253
rect 5306 4193 5318 4227
rect 5352 4193 5364 4227
rect 5306 4167 5364 4193
rect 5406 4227 5464 4253
rect 5406 4193 5412 4227
rect 5452 4193 5464 4227
rect 5406 4167 5464 4193
rect 5506 4227 5564 4253
rect 5506 4193 5518 4227
rect 5558 4193 5564 4227
rect 5506 4167 5564 4193
rect 5606 4227 5664 4253
rect 5606 4193 5618 4227
rect 5652 4193 5664 4227
rect 5606 4167 5664 4193
rect 5706 4227 5764 4253
rect 5706 4193 5718 4227
rect 5752 4193 5764 4227
rect 5706 4167 5764 4193
rect 5806 4227 5864 4253
rect 5806 4193 5812 4227
rect 5852 4193 5864 4227
rect 5806 4167 5864 4193
rect 5906 4227 5964 4253
rect 5906 4193 5918 4227
rect 5958 4193 5964 4227
rect 5906 4167 5964 4193
rect 6006 4227 6064 4253
rect 6006 4193 6018 4227
rect 6052 4193 6064 4227
rect 6006 4167 6064 4193
rect 6106 4227 6164 4253
rect 6106 4193 6118 4227
rect 6152 4193 6164 4227
rect 6106 4167 6164 4193
rect 6206 4227 6264 4253
rect 6206 4193 6218 4227
rect 6252 4193 6264 4227
rect 6206 4167 6264 4193
rect 6306 4227 6364 4253
rect 6306 4193 6318 4227
rect 6352 4193 6364 4227
rect 6306 4167 6364 4193
rect 6406 4227 6464 4253
rect 6618 4246 6862 4280
rect 6406 4193 6412 4227
rect 6452 4193 6464 4227
rect 6508 4208 6516 4242
rect 6558 4208 6574 4242
rect 6618 4227 6652 4246
rect 6406 4167 6464 4193
rect 6828 4243 6862 4246
rect 6828 4227 6962 4243
rect 6618 4177 6652 4193
rect 6696 4178 6712 4212
rect 6754 4178 6762 4212
rect 6862 4193 6928 4227
rect 6828 4177 6962 4193
rect 7028 4227 7162 4243
rect 7062 4193 7128 4227
rect 7028 4177 7162 4193
rect 7228 4227 7262 4243
rect 7228 4177 7262 4193
rect 7328 4227 7462 4243
rect 7362 4193 7428 4227
rect 7328 4177 7462 4193
rect 6 4087 64 4113
rect 6 4053 18 4087
rect 58 4053 64 4087
rect 6 4027 64 4053
rect 106 4087 164 4113
rect 106 4053 118 4087
rect 152 4053 164 4087
rect 106 4027 164 4053
rect 206 4087 264 4113
rect 206 4053 218 4087
rect 252 4053 264 4087
rect 206 4027 264 4053
rect 306 4087 364 4113
rect 306 4053 318 4087
rect 352 4053 364 4087
rect 306 4027 364 4053
rect 406 4087 464 4113
rect 406 4053 412 4087
rect 452 4053 464 4087
rect 406 4027 464 4053
rect 506 4087 564 4113
rect 506 4053 518 4087
rect 558 4053 564 4087
rect 506 4027 564 4053
rect 606 4087 664 4113
rect 606 4053 612 4087
rect 652 4053 664 4087
rect 606 4027 664 4053
rect 706 4087 764 4113
rect 706 4053 718 4087
rect 758 4053 764 4087
rect 706 4027 764 4053
rect 806 4087 864 4113
rect 806 4053 818 4087
rect 852 4053 864 4087
rect 806 4027 864 4053
rect 906 4087 964 4113
rect 906 4053 918 4087
rect 952 4053 964 4087
rect 906 4027 964 4053
rect 1006 4087 1064 4113
rect 1006 4053 1018 4087
rect 1052 4053 1064 4087
rect 1006 4027 1064 4053
rect 1106 4087 1164 4113
rect 1106 4053 1118 4087
rect 1152 4053 1164 4087
rect 1106 4027 1164 4053
rect 1206 4087 1264 4113
rect 1206 4053 1218 4087
rect 1252 4053 1264 4087
rect 1206 4027 1264 4053
rect 1306 4087 1364 4113
rect 1306 4053 1318 4087
rect 1352 4053 1364 4087
rect 1306 4027 1364 4053
rect 1406 4087 1464 4113
rect 1406 4053 1418 4087
rect 1452 4053 1464 4087
rect 1406 4027 1464 4053
rect 1506 4087 1564 4113
rect 1506 4053 1512 4087
rect 1552 4053 1564 4087
rect 1506 4027 1564 4053
rect 1606 4087 1664 4113
rect 1606 4053 1618 4087
rect 1658 4053 1664 4087
rect 1606 4027 1664 4053
rect 1706 4087 1764 4113
rect 1706 4053 1712 4087
rect 1752 4053 1764 4087
rect 1706 4027 1764 4053
rect 1806 4087 1864 4113
rect 1806 4053 1818 4087
rect 1858 4053 1864 4087
rect 1806 4027 1864 4053
rect 1906 4087 1964 4113
rect 1906 4053 1912 4087
rect 1952 4053 1964 4087
rect 1906 4027 1964 4053
rect 2006 4087 2064 4113
rect 2006 4053 2018 4087
rect 2058 4053 2064 4087
rect 2006 4027 2064 4053
rect 2106 4087 2164 4113
rect 2106 4053 2118 4087
rect 2152 4053 2164 4087
rect 2106 4027 2164 4053
rect 2206 4087 2264 4113
rect 2206 4053 2212 4087
rect 2252 4053 2264 4087
rect 2206 4027 2264 4053
rect 2306 4087 2364 4113
rect 2306 4053 2318 4087
rect 2358 4053 2364 4087
rect 2306 4027 2364 4053
rect 2406 4087 2464 4113
rect 2406 4053 2412 4087
rect 2452 4053 2464 4087
rect 2406 4027 2464 4053
rect 2506 4087 2564 4113
rect 2506 4053 2518 4087
rect 2558 4053 2564 4087
rect 2506 4027 2564 4053
rect 2606 4087 2664 4113
rect 2606 4053 2618 4087
rect 2652 4053 2664 4087
rect 2606 4027 2664 4053
rect 2706 4087 2764 4113
rect 2706 4053 2718 4087
rect 2752 4053 2764 4087
rect 2706 4027 2764 4053
rect 2806 4087 2864 4113
rect 2806 4053 2818 4087
rect 2852 4053 2864 4087
rect 2806 4027 2864 4053
rect 2906 4087 2964 4113
rect 2906 4053 2918 4087
rect 2952 4053 2964 4087
rect 2906 4027 2964 4053
rect 3006 4087 3064 4113
rect 3006 4053 3018 4087
rect 3052 4053 3064 4087
rect 3006 4027 3064 4053
rect 3106 4087 3164 4113
rect 3106 4053 3118 4087
rect 3152 4053 3164 4087
rect 3106 4027 3164 4053
rect 3206 4087 3264 4113
rect 3206 4053 3212 4087
rect 3252 4053 3264 4087
rect 3206 4027 3264 4053
rect 3306 4087 3364 4113
rect 3306 4053 3318 4087
rect 3358 4053 3364 4087
rect 3306 4027 3364 4053
rect 3406 4087 3464 4113
rect 3406 4053 3412 4087
rect 3452 4053 3464 4087
rect 3406 4027 3464 4053
rect 3506 4087 3564 4113
rect 3506 4053 3518 4087
rect 3558 4053 3564 4087
rect 3506 4027 3564 4053
rect 3606 4087 3664 4113
rect 3606 4053 3618 4087
rect 3652 4053 3664 4087
rect 3606 4027 3664 4053
rect 3706 4087 3764 4113
rect 3706 4053 3718 4087
rect 3752 4053 3764 4087
rect 3706 4027 3764 4053
rect 3806 4087 3864 4113
rect 3806 4053 3818 4087
rect 3852 4053 3864 4087
rect 3806 4027 3864 4053
rect 3906 4087 3964 4113
rect 3906 4053 3918 4087
rect 3952 4053 3964 4087
rect 3906 4027 3964 4053
rect 4006 4087 4064 4113
rect 4006 4053 4018 4087
rect 4052 4053 4064 4087
rect 4006 4027 4064 4053
rect 4106 4087 4164 4113
rect 4106 4053 4118 4087
rect 4152 4053 4164 4087
rect 4106 4027 4164 4053
rect 4206 4087 4264 4113
rect 4206 4053 4218 4087
rect 4252 4053 4264 4087
rect 4206 4027 4264 4053
rect 4306 4087 4364 4113
rect 4306 4053 4318 4087
rect 4352 4053 4364 4087
rect 4306 4027 4364 4053
rect 4406 4087 4464 4113
rect 4406 4053 4418 4087
rect 4452 4053 4464 4087
rect 4406 4027 4464 4053
rect 4506 4087 4564 4113
rect 4506 4053 4518 4087
rect 4552 4053 4564 4087
rect 4506 4027 4564 4053
rect 4606 4087 4664 4113
rect 4606 4053 4618 4087
rect 4652 4053 4664 4087
rect 4606 4027 4664 4053
rect 4706 4087 4764 4113
rect 4706 4053 4712 4087
rect 4752 4053 4764 4087
rect 4706 4027 4764 4053
rect 4806 4087 4864 4113
rect 4806 4053 4818 4087
rect 4858 4053 4864 4087
rect 4806 4027 4864 4053
rect 4906 4087 4964 4113
rect 4906 4053 4918 4087
rect 4952 4053 4964 4087
rect 4906 4027 4964 4053
rect 5006 4087 5064 4113
rect 5006 4053 5018 4087
rect 5052 4053 5064 4087
rect 5006 4027 5064 4053
rect 5106 4087 5164 4113
rect 5106 4053 5118 4087
rect 5152 4053 5164 4087
rect 5106 4027 5164 4053
rect 5206 4087 5264 4113
rect 5206 4053 5218 4087
rect 5252 4053 5264 4087
rect 5206 4027 5264 4053
rect 5306 4087 5364 4113
rect 5306 4053 5318 4087
rect 5352 4053 5364 4087
rect 5306 4027 5364 4053
rect 5406 4087 5464 4113
rect 5406 4053 5418 4087
rect 5452 4053 5464 4087
rect 5406 4027 5464 4053
rect 5506 4087 5564 4113
rect 5506 4053 5518 4087
rect 5552 4053 5564 4087
rect 5506 4027 5564 4053
rect 5606 4087 5664 4113
rect 5606 4053 5612 4087
rect 5652 4053 5664 4087
rect 5606 4027 5664 4053
rect 5706 4087 5764 4113
rect 5706 4053 5718 4087
rect 5758 4053 5764 4087
rect 5706 4027 5764 4053
rect 5806 4087 5864 4113
rect 5806 4053 5818 4087
rect 5852 4053 5864 4087
rect 5806 4027 5864 4053
rect 5906 4087 5964 4113
rect 5906 4053 5918 4087
rect 5952 4053 5964 4087
rect 5906 4027 5964 4053
rect 6006 4087 6064 4113
rect 6006 4053 6018 4087
rect 6052 4053 6064 4087
rect 6006 4027 6064 4053
rect 6106 4087 6164 4113
rect 6106 4053 6118 4087
rect 6152 4053 6164 4087
rect 6106 4027 6164 4053
rect 6206 4087 6264 4113
rect 6206 4053 6218 4087
rect 6252 4053 6264 4087
rect 6206 4027 6264 4053
rect 6306 4087 6364 4113
rect 6306 4053 6318 4087
rect 6352 4053 6364 4087
rect 6306 4027 6364 4053
rect 6406 4087 6464 4113
rect 6618 4106 6862 4140
rect 6406 4053 6412 4087
rect 6452 4053 6464 4087
rect 6508 4068 6516 4102
rect 6558 4068 6574 4102
rect 6618 4087 6652 4106
rect 6406 4027 6464 4053
rect 6828 4087 6862 4106
rect 6618 4037 6652 4053
rect 6696 4038 6712 4072
rect 6754 4038 6762 4072
rect 6828 4037 6862 4053
rect 6928 4087 7162 4103
rect 6962 4053 7028 4087
rect 7062 4053 7128 4087
rect 6928 4037 7162 4053
rect 7228 4087 7262 4103
rect 7228 4037 7262 4053
rect 7328 4087 7462 4103
rect 7362 4053 7428 4087
rect 7328 4037 7462 4053
rect 6 3947 64 3973
rect 6 3913 18 3947
rect 52 3913 64 3947
rect 6 3887 64 3913
rect 106 3947 164 3973
rect 106 3913 118 3947
rect 152 3913 164 3947
rect 106 3887 164 3913
rect 206 3947 264 3973
rect 206 3913 218 3947
rect 252 3913 264 3947
rect 206 3887 264 3913
rect 306 3947 364 3973
rect 306 3913 318 3947
rect 352 3913 364 3947
rect 306 3887 364 3913
rect 406 3947 464 3973
rect 406 3913 418 3947
rect 452 3913 464 3947
rect 406 3887 464 3913
rect 506 3947 564 3973
rect 506 3913 512 3947
rect 552 3913 564 3947
rect 506 3887 564 3913
rect 606 3947 664 3973
rect 606 3913 618 3947
rect 658 3913 664 3947
rect 606 3887 664 3913
rect 706 3947 764 3973
rect 706 3913 718 3947
rect 752 3913 764 3947
rect 706 3887 764 3913
rect 806 3947 864 3973
rect 806 3913 818 3947
rect 852 3913 864 3947
rect 806 3887 864 3913
rect 906 3947 964 3973
rect 906 3913 918 3947
rect 952 3913 964 3947
rect 906 3887 964 3913
rect 1006 3947 1064 3973
rect 1006 3913 1018 3947
rect 1052 3913 1064 3947
rect 1006 3887 1064 3913
rect 1106 3947 1164 3973
rect 1106 3913 1118 3947
rect 1152 3913 1164 3947
rect 1106 3887 1164 3913
rect 1206 3947 1264 3973
rect 1206 3913 1218 3947
rect 1252 3913 1264 3947
rect 1206 3887 1264 3913
rect 1306 3947 1364 3973
rect 1306 3913 1318 3947
rect 1352 3913 1364 3947
rect 1306 3887 1364 3913
rect 1406 3947 1464 3973
rect 1406 3913 1418 3947
rect 1452 3913 1464 3947
rect 1406 3887 1464 3913
rect 1506 3947 1564 3973
rect 1506 3913 1518 3947
rect 1552 3913 1564 3947
rect 1506 3887 1564 3913
rect 1606 3947 1664 3973
rect 1606 3913 1618 3947
rect 1652 3913 1664 3947
rect 1606 3887 1664 3913
rect 1706 3947 1764 3973
rect 1706 3913 1718 3947
rect 1752 3913 1764 3947
rect 1706 3887 1764 3913
rect 1806 3947 1864 3973
rect 1806 3913 1818 3947
rect 1852 3913 1864 3947
rect 1806 3887 1864 3913
rect 1906 3947 1964 3973
rect 1906 3913 1918 3947
rect 1952 3913 1964 3947
rect 1906 3887 1964 3913
rect 2006 3947 2064 3973
rect 2006 3913 2018 3947
rect 2052 3913 2064 3947
rect 2006 3887 2064 3913
rect 2106 3947 2164 3973
rect 2106 3913 2112 3947
rect 2152 3913 2164 3947
rect 2106 3887 2164 3913
rect 2206 3947 2264 3973
rect 2206 3913 2218 3947
rect 2258 3913 2264 3947
rect 2206 3887 2264 3913
rect 2306 3947 2364 3973
rect 2306 3913 2318 3947
rect 2352 3913 2364 3947
rect 2306 3887 2364 3913
rect 2406 3947 2464 3973
rect 2406 3913 2418 3947
rect 2452 3913 2464 3947
rect 2406 3887 2464 3913
rect 2506 3947 2564 3973
rect 2506 3913 2518 3947
rect 2552 3913 2564 3947
rect 2506 3887 2564 3913
rect 2606 3947 2664 3973
rect 2606 3913 2618 3947
rect 2652 3913 2664 3947
rect 2606 3887 2664 3913
rect 2706 3947 2764 3973
rect 2706 3913 2718 3947
rect 2752 3913 2764 3947
rect 2706 3887 2764 3913
rect 2806 3947 2864 3973
rect 2806 3913 2818 3947
rect 2852 3913 2864 3947
rect 2806 3887 2864 3913
rect 2906 3947 2964 3973
rect 2906 3913 2918 3947
rect 2952 3913 2964 3947
rect 2906 3887 2964 3913
rect 3006 3947 3064 3973
rect 3006 3913 3018 3947
rect 3052 3913 3064 3947
rect 3006 3887 3064 3913
rect 3106 3947 3164 3973
rect 3106 3913 3118 3947
rect 3152 3913 3164 3947
rect 3106 3887 3164 3913
rect 3206 3947 3264 3973
rect 3206 3913 3212 3947
rect 3252 3913 3264 3947
rect 3206 3887 3264 3913
rect 3306 3947 3364 3973
rect 3306 3913 3318 3947
rect 3358 3913 3364 3947
rect 3306 3887 3364 3913
rect 3406 3947 3464 3973
rect 3406 3913 3418 3947
rect 3452 3913 3464 3947
rect 3406 3887 3464 3913
rect 3506 3947 3564 3973
rect 3506 3913 3518 3947
rect 3552 3913 3564 3947
rect 3506 3887 3564 3913
rect 3606 3947 3664 3973
rect 3606 3913 3618 3947
rect 3652 3913 3664 3947
rect 3606 3887 3664 3913
rect 3706 3947 3764 3973
rect 3706 3913 3718 3947
rect 3752 3913 3764 3947
rect 3706 3887 3764 3913
rect 3806 3947 3864 3973
rect 3806 3913 3818 3947
rect 3852 3913 3864 3947
rect 3806 3887 3864 3913
rect 3906 3947 3964 3973
rect 3906 3913 3918 3947
rect 3952 3913 3964 3947
rect 3906 3887 3964 3913
rect 4006 3947 4064 3973
rect 4006 3913 4018 3947
rect 4052 3913 4064 3947
rect 4006 3887 4064 3913
rect 4106 3947 4164 3973
rect 4106 3913 4112 3947
rect 4152 3913 4164 3947
rect 4106 3887 4164 3913
rect 4206 3947 4264 3973
rect 4206 3913 4218 3947
rect 4258 3913 4264 3947
rect 4206 3887 4264 3913
rect 4306 3947 4364 3973
rect 4306 3913 4318 3947
rect 4352 3913 4364 3947
rect 4306 3887 4364 3913
rect 4406 3947 4464 3973
rect 4406 3913 4418 3947
rect 4452 3913 4464 3947
rect 4406 3887 4464 3913
rect 4506 3947 4564 3973
rect 4506 3913 4512 3947
rect 4552 3913 4564 3947
rect 4506 3887 4564 3913
rect 4606 3947 4664 3973
rect 4606 3913 4618 3947
rect 4658 3913 4664 3947
rect 4606 3887 4664 3913
rect 4706 3947 4764 3973
rect 4706 3913 4718 3947
rect 4752 3913 4764 3947
rect 4706 3887 4764 3913
rect 4806 3947 4864 3973
rect 4806 3913 4818 3947
rect 4852 3913 4864 3947
rect 4806 3887 4864 3913
rect 4906 3947 4964 3973
rect 4906 3913 4918 3947
rect 4952 3913 4964 3947
rect 4906 3887 4964 3913
rect 5006 3947 5064 3973
rect 5006 3913 5018 3947
rect 5052 3913 5064 3947
rect 5006 3887 5064 3913
rect 5106 3947 5164 3973
rect 5106 3913 5118 3947
rect 5152 3913 5164 3947
rect 5106 3887 5164 3913
rect 5206 3947 5264 3973
rect 5206 3913 5218 3947
rect 5252 3913 5264 3947
rect 5206 3887 5264 3913
rect 5306 3947 5364 3973
rect 5306 3913 5318 3947
rect 5352 3913 5364 3947
rect 5306 3887 5364 3913
rect 5406 3947 5464 3973
rect 5406 3913 5418 3947
rect 5452 3913 5464 3947
rect 5406 3887 5464 3913
rect 5506 3947 5564 3973
rect 5506 3913 5518 3947
rect 5552 3913 5564 3947
rect 5506 3887 5564 3913
rect 5606 3947 5664 3973
rect 5606 3913 5618 3947
rect 5652 3913 5664 3947
rect 5606 3887 5664 3913
rect 5706 3947 5764 3973
rect 5706 3913 5718 3947
rect 5752 3913 5764 3947
rect 5706 3887 5764 3913
rect 5806 3947 5864 3973
rect 5806 3913 5818 3947
rect 5852 3913 5864 3947
rect 5806 3887 5864 3913
rect 5906 3947 5964 3973
rect 5906 3913 5918 3947
rect 5952 3913 5964 3947
rect 5906 3887 5964 3913
rect 6006 3947 6064 3973
rect 6006 3913 6012 3947
rect 6052 3913 6064 3947
rect 6006 3887 6064 3913
rect 6106 3947 6164 3973
rect 6106 3913 6118 3947
rect 6158 3913 6164 3947
rect 6106 3887 6164 3913
rect 6206 3947 6264 3973
rect 6206 3913 6218 3947
rect 6252 3913 6264 3947
rect 6206 3887 6264 3913
rect 6306 3947 6364 3973
rect 6306 3913 6318 3947
rect 6352 3913 6364 3947
rect 6306 3887 6364 3913
rect 6406 3947 6464 3973
rect 6618 3966 6862 4000
rect 6406 3913 6418 3947
rect 6452 3913 6464 3947
rect 6508 3928 6516 3962
rect 6558 3928 6574 3962
rect 6618 3947 6652 3966
rect 6406 3887 6464 3913
rect 6828 3963 6862 3966
rect 6828 3947 6962 3963
rect 6618 3897 6652 3913
rect 6696 3898 6712 3932
rect 6754 3898 6762 3932
rect 6862 3913 6928 3947
rect 6828 3897 6962 3913
rect 7028 3947 7062 3963
rect 7028 3897 7062 3913
rect 7128 3947 7262 3963
rect 7162 3913 7228 3947
rect 7128 3897 7262 3913
rect 7328 3947 7462 3963
rect 7362 3913 7428 3947
rect 7328 3897 7462 3913
rect 6 3807 64 3833
rect 6 3773 18 3807
rect 52 3773 64 3807
rect 6 3747 64 3773
rect 106 3807 164 3833
rect 106 3773 118 3807
rect 152 3773 164 3807
rect 106 3747 164 3773
rect 206 3807 264 3833
rect 206 3773 218 3807
rect 252 3773 264 3807
rect 206 3747 264 3773
rect 306 3807 364 3833
rect 306 3773 318 3807
rect 352 3773 364 3807
rect 306 3747 364 3773
rect 406 3807 464 3833
rect 406 3773 418 3807
rect 452 3773 464 3807
rect 406 3747 464 3773
rect 506 3807 564 3833
rect 506 3773 518 3807
rect 552 3773 564 3807
rect 506 3747 564 3773
rect 606 3807 664 3833
rect 606 3773 618 3807
rect 652 3773 664 3807
rect 606 3747 664 3773
rect 706 3807 764 3833
rect 706 3773 718 3807
rect 752 3773 764 3807
rect 706 3747 764 3773
rect 806 3807 864 3833
rect 806 3773 818 3807
rect 852 3773 864 3807
rect 806 3747 864 3773
rect 906 3807 964 3833
rect 906 3773 918 3807
rect 952 3773 964 3807
rect 906 3747 964 3773
rect 1006 3807 1064 3833
rect 1006 3773 1018 3807
rect 1052 3773 1064 3807
rect 1006 3747 1064 3773
rect 1106 3807 1164 3833
rect 1106 3773 1118 3807
rect 1152 3773 1164 3807
rect 1106 3747 1164 3773
rect 1206 3807 1264 3833
rect 1206 3773 1212 3807
rect 1252 3773 1264 3807
rect 1206 3747 1264 3773
rect 1306 3807 1364 3833
rect 1306 3773 1318 3807
rect 1358 3773 1364 3807
rect 1306 3747 1364 3773
rect 1406 3807 1464 3833
rect 1406 3773 1412 3807
rect 1452 3773 1464 3807
rect 1406 3747 1464 3773
rect 1506 3807 1564 3833
rect 1506 3773 1518 3807
rect 1558 3773 1564 3807
rect 1506 3747 1564 3773
rect 1606 3807 1664 3833
rect 1606 3773 1618 3807
rect 1652 3773 1664 3807
rect 1606 3747 1664 3773
rect 1706 3807 1764 3833
rect 1706 3773 1712 3807
rect 1752 3773 1764 3807
rect 1706 3747 1764 3773
rect 1806 3807 1864 3833
rect 1806 3773 1818 3807
rect 1858 3773 1864 3807
rect 1806 3747 1864 3773
rect 1906 3807 1964 3833
rect 1906 3773 1918 3807
rect 1952 3773 1964 3807
rect 1906 3747 1964 3773
rect 2006 3807 2064 3833
rect 2006 3773 2018 3807
rect 2052 3773 2064 3807
rect 2006 3747 2064 3773
rect 2106 3807 2164 3833
rect 2106 3773 2118 3807
rect 2152 3773 2164 3807
rect 2106 3747 2164 3773
rect 2206 3807 2264 3833
rect 2206 3773 2218 3807
rect 2252 3773 2264 3807
rect 2206 3747 2264 3773
rect 2306 3807 2364 3833
rect 2306 3773 2318 3807
rect 2352 3773 2364 3807
rect 2306 3747 2364 3773
rect 2406 3807 2464 3833
rect 2406 3773 2418 3807
rect 2452 3773 2464 3807
rect 2406 3747 2464 3773
rect 2506 3807 2564 3833
rect 2506 3773 2518 3807
rect 2552 3773 2564 3807
rect 2506 3747 2564 3773
rect 2606 3807 2664 3833
rect 2606 3773 2618 3807
rect 2652 3773 2664 3807
rect 2606 3747 2664 3773
rect 2706 3807 2764 3833
rect 2706 3773 2718 3807
rect 2752 3773 2764 3807
rect 2706 3747 2764 3773
rect 2806 3807 2864 3833
rect 2806 3773 2818 3807
rect 2852 3773 2864 3807
rect 2806 3747 2864 3773
rect 2906 3807 2964 3833
rect 2906 3773 2918 3807
rect 2952 3773 2964 3807
rect 2906 3747 2964 3773
rect 3006 3807 3064 3833
rect 3006 3773 3018 3807
rect 3052 3773 3064 3807
rect 3006 3747 3064 3773
rect 3106 3807 3164 3833
rect 3106 3773 3118 3807
rect 3152 3773 3164 3807
rect 3106 3747 3164 3773
rect 3206 3807 3264 3833
rect 3206 3773 3218 3807
rect 3252 3773 3264 3807
rect 3206 3747 3264 3773
rect 3306 3807 3364 3833
rect 3306 3773 3318 3807
rect 3352 3773 3364 3807
rect 3306 3747 3364 3773
rect 3406 3807 3464 3833
rect 3406 3773 3412 3807
rect 3452 3773 3464 3807
rect 3406 3747 3464 3773
rect 3506 3807 3564 3833
rect 3506 3773 3518 3807
rect 3558 3773 3564 3807
rect 3506 3747 3564 3773
rect 3606 3807 3664 3833
rect 3606 3773 3618 3807
rect 3652 3773 3664 3807
rect 3606 3747 3664 3773
rect 3706 3807 3764 3833
rect 3706 3773 3718 3807
rect 3752 3773 3764 3807
rect 3706 3747 3764 3773
rect 3806 3807 3864 3833
rect 3806 3773 3818 3807
rect 3852 3773 3864 3807
rect 3806 3747 3864 3773
rect 3906 3807 3964 3833
rect 3906 3773 3918 3807
rect 3952 3773 3964 3807
rect 3906 3747 3964 3773
rect 4006 3807 4064 3833
rect 4006 3773 4018 3807
rect 4052 3773 4064 3807
rect 4006 3747 4064 3773
rect 4106 3807 4164 3833
rect 4106 3773 4118 3807
rect 4152 3773 4164 3807
rect 4106 3747 4164 3773
rect 4206 3807 4264 3833
rect 4206 3773 4218 3807
rect 4252 3773 4264 3807
rect 4206 3747 4264 3773
rect 4306 3807 4364 3833
rect 4306 3773 4318 3807
rect 4352 3773 4364 3807
rect 4306 3747 4364 3773
rect 4406 3807 4464 3833
rect 4406 3773 4418 3807
rect 4452 3773 4464 3807
rect 4406 3747 4464 3773
rect 4506 3807 4564 3833
rect 4506 3773 4518 3807
rect 4552 3773 4564 3807
rect 4506 3747 4564 3773
rect 4606 3807 4664 3833
rect 4606 3773 4618 3807
rect 4652 3773 4664 3807
rect 4606 3747 4664 3773
rect 4706 3807 4764 3833
rect 4706 3773 4712 3807
rect 4752 3773 4764 3807
rect 4706 3747 4764 3773
rect 4806 3807 4864 3833
rect 4806 3773 4818 3807
rect 4858 3773 4864 3807
rect 4806 3747 4864 3773
rect 4906 3807 4964 3833
rect 4906 3773 4918 3807
rect 4952 3773 4964 3807
rect 4906 3747 4964 3773
rect 5006 3807 5064 3833
rect 5006 3773 5018 3807
rect 5052 3773 5064 3807
rect 5006 3747 5064 3773
rect 5106 3807 5164 3833
rect 5106 3773 5118 3807
rect 5152 3773 5164 3807
rect 5106 3747 5164 3773
rect 5206 3807 5264 3833
rect 5206 3773 5218 3807
rect 5252 3773 5264 3807
rect 5206 3747 5264 3773
rect 5306 3807 5364 3833
rect 5306 3773 5318 3807
rect 5352 3773 5364 3807
rect 5306 3747 5364 3773
rect 5406 3807 5464 3833
rect 5406 3773 5418 3807
rect 5452 3773 5464 3807
rect 5406 3747 5464 3773
rect 5506 3807 5564 3833
rect 5506 3773 5518 3807
rect 5552 3773 5564 3807
rect 5506 3747 5564 3773
rect 5606 3807 5664 3833
rect 5606 3773 5612 3807
rect 5652 3773 5664 3807
rect 5606 3747 5664 3773
rect 5706 3807 5764 3833
rect 5706 3773 5718 3807
rect 5758 3773 5764 3807
rect 5706 3747 5764 3773
rect 5806 3807 5864 3833
rect 5806 3773 5818 3807
rect 5852 3773 5864 3807
rect 5806 3747 5864 3773
rect 5906 3807 5964 3833
rect 5906 3773 5918 3807
rect 5952 3773 5964 3807
rect 5906 3747 5964 3773
rect 6006 3807 6064 3833
rect 6006 3773 6018 3807
rect 6052 3773 6064 3807
rect 6006 3747 6064 3773
rect 6106 3807 6164 3833
rect 6106 3773 6118 3807
rect 6152 3773 6164 3807
rect 6106 3747 6164 3773
rect 6206 3807 6264 3833
rect 6206 3773 6218 3807
rect 6252 3773 6264 3807
rect 6206 3747 6264 3773
rect 6306 3807 6364 3833
rect 6306 3773 6318 3807
rect 6352 3773 6364 3807
rect 6306 3747 6364 3773
rect 6406 3807 6464 3833
rect 6618 3826 6862 3860
rect 6406 3773 6418 3807
rect 6452 3773 6464 3807
rect 6508 3788 6516 3822
rect 6558 3788 6574 3822
rect 6618 3807 6652 3826
rect 6406 3747 6464 3773
rect 6828 3807 6862 3826
rect 6618 3757 6652 3773
rect 6696 3758 6712 3792
rect 6754 3758 6762 3792
rect 6828 3757 6862 3773
rect 6928 3807 7062 3823
rect 6962 3773 7028 3807
rect 6928 3757 7062 3773
rect 7128 3807 7262 3823
rect 7162 3773 7228 3807
rect 7128 3757 7262 3773
rect 7328 3807 7462 3823
rect 7362 3773 7428 3807
rect 7328 3757 7462 3773
rect 8 3650 18 3684
rect 52 3650 118 3684
rect 152 3650 168 3684
rect 208 3666 218 3700
rect 252 3666 318 3700
rect 352 3666 368 3700
rect 408 3650 418 3684
rect 452 3650 518 3684
rect 552 3650 568 3684
rect 608 3666 618 3700
rect 652 3666 718 3700
rect 752 3666 768 3700
rect 808 3650 818 3684
rect 852 3650 918 3684
rect 952 3650 968 3684
rect 1008 3666 1018 3700
rect 1052 3666 1118 3700
rect 1152 3666 1168 3700
rect 1208 3650 1218 3684
rect 1252 3650 1318 3684
rect 1352 3650 1368 3684
rect 1408 3666 1418 3700
rect 1452 3666 1518 3700
rect 1552 3666 1568 3700
rect 1608 3650 1618 3684
rect 1652 3650 1718 3684
rect 1752 3650 1768 3684
rect 1808 3666 1818 3700
rect 1852 3666 1918 3700
rect 1952 3666 1968 3700
rect 2008 3650 2018 3684
rect 2052 3650 2118 3684
rect 2152 3650 2168 3684
rect 2208 3666 2218 3700
rect 2252 3666 2318 3700
rect 2352 3666 2368 3700
rect 2408 3650 2418 3684
rect 2452 3650 2518 3684
rect 2552 3650 2568 3684
rect 2608 3666 2618 3700
rect 2652 3666 2718 3700
rect 2752 3666 2768 3700
rect 2808 3650 2818 3684
rect 2852 3650 2918 3684
rect 2952 3650 2968 3684
rect 3008 3666 3018 3700
rect 3052 3666 3118 3700
rect 3152 3666 3168 3700
rect 3208 3650 3218 3684
rect 3252 3650 3318 3684
rect 3352 3650 3368 3684
rect 3408 3666 3418 3700
rect 3452 3666 3518 3700
rect 3552 3666 3568 3700
rect 3608 3650 3618 3684
rect 3652 3650 3718 3684
rect 3752 3650 3768 3684
rect 3808 3666 3818 3700
rect 3852 3666 3918 3700
rect 3952 3666 3968 3700
rect 4008 3650 4018 3684
rect 4052 3650 4118 3684
rect 4152 3650 4168 3684
rect 4208 3666 4218 3700
rect 4252 3666 4318 3700
rect 4352 3666 4368 3700
rect 4408 3650 4418 3684
rect 4452 3650 4518 3684
rect 4552 3650 4568 3684
rect 4608 3666 4618 3700
rect 4652 3666 4718 3700
rect 4752 3666 4768 3700
rect 4808 3650 4818 3684
rect 4852 3650 4918 3684
rect 4952 3650 4968 3684
rect 5008 3666 5018 3700
rect 5052 3666 5118 3700
rect 5152 3666 5168 3700
rect 5208 3650 5218 3684
rect 5252 3650 5318 3684
rect 5352 3650 5368 3684
rect 5408 3666 5418 3700
rect 5452 3666 5518 3700
rect 5552 3666 5568 3700
rect 5608 3650 5618 3684
rect 5652 3650 5718 3684
rect 5752 3650 5768 3684
rect 5808 3666 5818 3700
rect 5852 3666 5918 3700
rect 5952 3666 5968 3700
rect 6008 3650 6018 3684
rect 6052 3650 6118 3684
rect 6152 3650 6168 3684
rect 6208 3666 6218 3700
rect 6252 3666 6318 3700
rect 6352 3666 6368 3700
rect 6516 3681 6568 3698
rect 6550 3664 6568 3681
rect 6602 3664 6618 3698
rect 6652 3664 6668 3698
rect 6702 3669 6720 3698
rect 6702 3664 6754 3669
rect 6862 3664 6878 3698
rect 6912 3664 6928 3698
rect 6962 3664 6978 3698
rect 7012 3664 7028 3698
rect 7062 3664 7078 3698
rect 7112 3664 7128 3698
rect 7162 3664 7178 3698
rect 7212 3664 7228 3698
rect 7262 3664 7278 3698
rect 7312 3664 7328 3698
rect 7362 3664 7378 3698
rect 7412 3664 7428 3698
rect 6 3577 64 3603
rect 6 3543 18 3577
rect 52 3543 64 3577
rect 6 3517 64 3543
rect 106 3577 164 3603
rect 106 3543 118 3577
rect 152 3543 164 3577
rect 106 3517 164 3543
rect 206 3577 264 3603
rect 206 3543 212 3577
rect 252 3543 264 3577
rect 206 3517 264 3543
rect 306 3577 364 3603
rect 306 3543 318 3577
rect 358 3543 364 3577
rect 306 3517 364 3543
rect 406 3577 464 3603
rect 406 3543 418 3577
rect 452 3543 464 3577
rect 406 3517 464 3543
rect 506 3577 564 3603
rect 506 3543 518 3577
rect 552 3543 564 3577
rect 506 3517 564 3543
rect 606 3577 664 3603
rect 606 3543 618 3577
rect 652 3543 664 3577
rect 606 3517 664 3543
rect 706 3577 764 3603
rect 706 3543 718 3577
rect 752 3543 764 3577
rect 706 3517 764 3543
rect 806 3577 864 3603
rect 806 3543 818 3577
rect 852 3543 864 3577
rect 806 3517 864 3543
rect 906 3577 964 3603
rect 906 3543 918 3577
rect 952 3543 964 3577
rect 906 3517 964 3543
rect 1006 3577 1064 3603
rect 1006 3543 1018 3577
rect 1052 3543 1064 3577
rect 1006 3517 1064 3543
rect 1106 3577 1164 3603
rect 1106 3543 1118 3577
rect 1152 3543 1164 3577
rect 1106 3517 1164 3543
rect 1206 3577 1264 3603
rect 1206 3543 1218 3577
rect 1252 3543 1264 3577
rect 1206 3517 1264 3543
rect 1306 3577 1364 3603
rect 1306 3543 1312 3577
rect 1352 3543 1364 3577
rect 1306 3517 1364 3543
rect 1406 3577 1464 3603
rect 1406 3543 1418 3577
rect 1458 3543 1464 3577
rect 1406 3517 1464 3543
rect 1506 3577 1564 3603
rect 1506 3543 1512 3577
rect 1552 3543 1564 3577
rect 1506 3517 1564 3543
rect 1606 3577 1664 3603
rect 1606 3543 1618 3577
rect 1658 3543 1664 3577
rect 1606 3517 1664 3543
rect 1706 3577 1764 3603
rect 1706 3543 1718 3577
rect 1752 3543 1764 3577
rect 1706 3517 1764 3543
rect 1806 3577 1864 3603
rect 1806 3543 1818 3577
rect 1852 3543 1864 3577
rect 1806 3517 1864 3543
rect 1906 3577 1964 3603
rect 1906 3543 1918 3577
rect 1952 3543 1964 3577
rect 1906 3517 1964 3543
rect 2006 3577 2064 3603
rect 2006 3543 2018 3577
rect 2052 3543 2064 3577
rect 2006 3517 2064 3543
rect 2106 3577 2164 3603
rect 2106 3543 2118 3577
rect 2152 3543 2164 3577
rect 2106 3517 2164 3543
rect 2206 3577 2264 3603
rect 2206 3543 2212 3577
rect 2252 3543 2264 3577
rect 2206 3517 2264 3543
rect 2306 3577 2364 3603
rect 2306 3543 2318 3577
rect 2358 3543 2364 3577
rect 2306 3517 2364 3543
rect 2406 3577 2464 3603
rect 2406 3543 2418 3577
rect 2452 3543 2464 3577
rect 2406 3517 2464 3543
rect 2506 3577 2564 3603
rect 2506 3543 2518 3577
rect 2552 3543 2564 3577
rect 2506 3517 2564 3543
rect 2606 3577 2664 3603
rect 2606 3543 2618 3577
rect 2652 3543 2664 3577
rect 2606 3517 2664 3543
rect 2706 3577 2764 3603
rect 2706 3543 2718 3577
rect 2752 3543 2764 3577
rect 2706 3517 2764 3543
rect 2806 3577 2864 3603
rect 2806 3543 2818 3577
rect 2852 3543 2864 3577
rect 2806 3517 2864 3543
rect 2906 3577 2964 3603
rect 2906 3543 2918 3577
rect 2952 3543 2964 3577
rect 2906 3517 2964 3543
rect 3006 3577 3064 3603
rect 3006 3543 3018 3577
rect 3052 3543 3064 3577
rect 3006 3517 3064 3543
rect 3106 3577 3164 3603
rect 3106 3543 3118 3577
rect 3152 3543 3164 3577
rect 3106 3517 3164 3543
rect 3206 3577 3264 3603
rect 3206 3543 3218 3577
rect 3252 3543 3264 3577
rect 3206 3517 3264 3543
rect 3306 3577 3364 3603
rect 3306 3543 3318 3577
rect 3352 3543 3364 3577
rect 3306 3517 3364 3543
rect 3406 3577 3464 3603
rect 3406 3543 3418 3577
rect 3452 3543 3464 3577
rect 3406 3517 3464 3543
rect 3506 3577 3564 3603
rect 3506 3543 3512 3577
rect 3552 3543 3564 3577
rect 3506 3517 3564 3543
rect 3606 3577 3664 3603
rect 3606 3543 3618 3577
rect 3658 3543 3664 3577
rect 3606 3517 3664 3543
rect 3706 3577 3764 3603
rect 3706 3543 3712 3577
rect 3752 3543 3764 3577
rect 3706 3517 3764 3543
rect 3806 3577 3864 3603
rect 3806 3543 3818 3577
rect 3858 3543 3864 3577
rect 3806 3517 3864 3543
rect 3906 3577 3964 3603
rect 3906 3543 3918 3577
rect 3952 3543 3964 3577
rect 3906 3517 3964 3543
rect 4006 3577 4064 3603
rect 4006 3543 4018 3577
rect 4052 3543 4064 3577
rect 4006 3517 4064 3543
rect 4106 3577 4164 3603
rect 4106 3543 4118 3577
rect 4152 3543 4164 3577
rect 4106 3517 4164 3543
rect 4206 3577 4264 3603
rect 4206 3543 4212 3577
rect 4252 3543 4264 3577
rect 4206 3517 4264 3543
rect 4306 3577 4364 3603
rect 4306 3543 4318 3577
rect 4358 3543 4364 3577
rect 4306 3517 4364 3543
rect 4406 3577 4464 3603
rect 4406 3543 4418 3577
rect 4452 3543 4464 3577
rect 4406 3517 4464 3543
rect 4506 3577 4564 3603
rect 4506 3543 4518 3577
rect 4552 3543 4564 3577
rect 4506 3517 4564 3543
rect 4606 3577 4664 3603
rect 4606 3543 4618 3577
rect 4652 3543 4664 3577
rect 4606 3517 4664 3543
rect 4706 3577 4764 3603
rect 4706 3543 4712 3577
rect 4752 3543 4764 3577
rect 4706 3517 4764 3543
rect 4806 3577 4864 3603
rect 4806 3543 4818 3577
rect 4858 3543 4864 3577
rect 4806 3517 4864 3543
rect 4906 3577 4964 3603
rect 4906 3543 4918 3577
rect 4952 3543 4964 3577
rect 4906 3517 4964 3543
rect 5006 3577 5064 3603
rect 5006 3543 5018 3577
rect 5052 3543 5064 3577
rect 5006 3517 5064 3543
rect 5106 3577 5164 3603
rect 5106 3543 5118 3577
rect 5152 3543 5164 3577
rect 5106 3517 5164 3543
rect 5206 3577 5264 3603
rect 5206 3543 5212 3577
rect 5252 3543 5264 3577
rect 5206 3517 5264 3543
rect 5306 3577 5364 3603
rect 5306 3543 5318 3577
rect 5358 3543 5364 3577
rect 5306 3517 5364 3543
rect 5406 3577 5464 3603
rect 5406 3543 5418 3577
rect 5452 3543 5464 3577
rect 5406 3517 5464 3543
rect 5506 3577 5564 3603
rect 5506 3543 5518 3577
rect 5552 3543 5564 3577
rect 5506 3517 5564 3543
rect 5606 3577 5664 3603
rect 5606 3543 5618 3577
rect 5652 3543 5664 3577
rect 5606 3517 5664 3543
rect 5706 3577 5764 3603
rect 5706 3543 5718 3577
rect 5752 3543 5764 3577
rect 5706 3517 5764 3543
rect 5806 3577 5864 3603
rect 5806 3543 5818 3577
rect 5852 3543 5864 3577
rect 5806 3517 5864 3543
rect 5906 3577 5964 3603
rect 5906 3543 5918 3577
rect 5952 3543 5964 3577
rect 5906 3517 5964 3543
rect 6006 3577 6064 3603
rect 6006 3543 6018 3577
rect 6052 3543 6064 3577
rect 6006 3517 6064 3543
rect 6106 3577 6164 3603
rect 6106 3543 6118 3577
rect 6152 3543 6164 3577
rect 6106 3517 6164 3543
rect 6206 3577 6264 3603
rect 6206 3543 6218 3577
rect 6252 3543 6264 3577
rect 6206 3517 6264 3543
rect 6306 3577 6364 3603
rect 6306 3543 6318 3577
rect 6352 3543 6364 3577
rect 6306 3517 6364 3543
rect 6406 3577 6464 3603
rect 6618 3596 6862 3630
rect 6406 3543 6412 3577
rect 6452 3543 6464 3577
rect 6508 3558 6516 3592
rect 6558 3558 6574 3592
rect 6618 3577 6652 3596
rect 6406 3517 6464 3543
rect 6828 3593 6862 3596
rect 6828 3577 6962 3593
rect 6618 3527 6652 3543
rect 6696 3528 6712 3562
rect 6754 3528 6762 3562
rect 6862 3543 6928 3577
rect 6828 3527 6962 3543
rect 7028 3577 7162 3593
rect 7062 3543 7128 3577
rect 7028 3527 7162 3543
rect 7228 3577 7362 3593
rect 7262 3543 7328 3577
rect 7228 3527 7362 3543
rect 7428 3577 7462 3593
rect 7428 3527 7462 3543
rect 6 3437 64 3463
rect 6 3403 18 3437
rect 52 3403 64 3437
rect 6 3377 64 3403
rect 106 3437 164 3463
rect 106 3403 118 3437
rect 152 3403 164 3437
rect 106 3377 164 3403
rect 206 3437 264 3463
rect 206 3403 218 3437
rect 252 3403 264 3437
rect 206 3377 264 3403
rect 306 3437 364 3463
rect 306 3403 318 3437
rect 352 3403 364 3437
rect 306 3377 364 3403
rect 406 3437 464 3463
rect 406 3403 418 3437
rect 452 3403 464 3437
rect 406 3377 464 3403
rect 506 3437 564 3463
rect 506 3403 512 3437
rect 552 3403 564 3437
rect 506 3377 564 3403
rect 606 3437 664 3463
rect 606 3403 618 3437
rect 658 3403 664 3437
rect 606 3377 664 3403
rect 706 3437 764 3463
rect 706 3403 712 3437
rect 752 3403 764 3437
rect 706 3377 764 3403
rect 806 3437 864 3463
rect 806 3403 818 3437
rect 858 3403 864 3437
rect 806 3377 864 3403
rect 906 3437 964 3463
rect 906 3403 918 3437
rect 952 3403 964 3437
rect 906 3377 964 3403
rect 1006 3437 1064 3463
rect 1006 3403 1018 3437
rect 1052 3403 1064 3437
rect 1006 3377 1064 3403
rect 1106 3437 1164 3463
rect 1106 3403 1118 3437
rect 1152 3403 1164 3437
rect 1106 3377 1164 3403
rect 1206 3437 1264 3463
rect 1206 3403 1218 3437
rect 1252 3403 1264 3437
rect 1206 3377 1264 3403
rect 1306 3437 1364 3463
rect 1306 3403 1318 3437
rect 1352 3403 1364 3437
rect 1306 3377 1364 3403
rect 1406 3437 1464 3463
rect 1406 3403 1418 3437
rect 1452 3403 1464 3437
rect 1406 3377 1464 3403
rect 1506 3437 1564 3463
rect 1506 3403 1518 3437
rect 1552 3403 1564 3437
rect 1506 3377 1564 3403
rect 1606 3437 1664 3463
rect 1606 3403 1618 3437
rect 1652 3403 1664 3437
rect 1606 3377 1664 3403
rect 1706 3437 1764 3463
rect 1706 3403 1718 3437
rect 1752 3403 1764 3437
rect 1706 3377 1764 3403
rect 1806 3437 1864 3463
rect 1806 3403 1818 3437
rect 1852 3403 1864 3437
rect 1806 3377 1864 3403
rect 1906 3437 1964 3463
rect 1906 3403 1912 3437
rect 1952 3403 1964 3437
rect 1906 3377 1964 3403
rect 2006 3437 2064 3463
rect 2006 3403 2018 3437
rect 2058 3403 2064 3437
rect 2006 3377 2064 3403
rect 2106 3437 2164 3463
rect 2106 3403 2118 3437
rect 2152 3403 2164 3437
rect 2106 3377 2164 3403
rect 2206 3437 2264 3463
rect 2206 3403 2218 3437
rect 2252 3403 2264 3437
rect 2206 3377 2264 3403
rect 2306 3437 2364 3463
rect 2306 3403 2318 3437
rect 2352 3403 2364 3437
rect 2306 3377 2364 3403
rect 2406 3437 2464 3463
rect 2406 3403 2418 3437
rect 2452 3403 2464 3437
rect 2406 3377 2464 3403
rect 2506 3437 2564 3463
rect 2506 3403 2518 3437
rect 2552 3403 2564 3437
rect 2506 3377 2564 3403
rect 2606 3437 2664 3463
rect 2606 3403 2618 3437
rect 2652 3403 2664 3437
rect 2606 3377 2664 3403
rect 2706 3437 2764 3463
rect 2706 3403 2718 3437
rect 2752 3403 2764 3437
rect 2706 3377 2764 3403
rect 2806 3437 2864 3463
rect 2806 3403 2812 3437
rect 2852 3403 2864 3437
rect 2806 3377 2864 3403
rect 2906 3437 2964 3463
rect 2906 3403 2918 3437
rect 2958 3403 2964 3437
rect 2906 3377 2964 3403
rect 3006 3437 3064 3463
rect 3006 3403 3018 3437
rect 3052 3403 3064 3437
rect 3006 3377 3064 3403
rect 3106 3437 3164 3463
rect 3106 3403 3118 3437
rect 3152 3403 3164 3437
rect 3106 3377 3164 3403
rect 3206 3437 3264 3463
rect 3206 3403 3218 3437
rect 3252 3403 3264 3437
rect 3206 3377 3264 3403
rect 3306 3437 3364 3463
rect 3306 3403 3318 3437
rect 3352 3403 3364 3437
rect 3306 3377 3364 3403
rect 3406 3437 3464 3463
rect 3406 3403 3418 3437
rect 3452 3403 3464 3437
rect 3406 3377 3464 3403
rect 3506 3437 3564 3463
rect 3506 3403 3518 3437
rect 3552 3403 3564 3437
rect 3506 3377 3564 3403
rect 3606 3437 3664 3463
rect 3606 3403 3618 3437
rect 3652 3403 3664 3437
rect 3606 3377 3664 3403
rect 3706 3437 3764 3463
rect 3706 3403 3718 3437
rect 3752 3403 3764 3437
rect 3706 3377 3764 3403
rect 3806 3437 3864 3463
rect 3806 3403 3818 3437
rect 3852 3403 3864 3437
rect 3806 3377 3864 3403
rect 3906 3437 3964 3463
rect 3906 3403 3918 3437
rect 3952 3403 3964 3437
rect 3906 3377 3964 3403
rect 4006 3437 4064 3463
rect 4006 3403 4018 3437
rect 4052 3403 4064 3437
rect 4006 3377 4064 3403
rect 4106 3437 4164 3463
rect 4106 3403 4118 3437
rect 4152 3403 4164 3437
rect 4106 3377 4164 3403
rect 4206 3437 4264 3463
rect 4206 3403 4218 3437
rect 4252 3403 4264 3437
rect 4206 3377 4264 3403
rect 4306 3437 4364 3463
rect 4306 3403 4318 3437
rect 4352 3403 4364 3437
rect 4306 3377 4364 3403
rect 4406 3437 4464 3463
rect 4406 3403 4418 3437
rect 4452 3403 4464 3437
rect 4406 3377 4464 3403
rect 4506 3437 4564 3463
rect 4506 3403 4518 3437
rect 4552 3403 4564 3437
rect 4506 3377 4564 3403
rect 4606 3437 4664 3463
rect 4606 3403 4618 3437
rect 4652 3403 4664 3437
rect 4606 3377 4664 3403
rect 4706 3437 4764 3463
rect 4706 3403 4718 3437
rect 4752 3403 4764 3437
rect 4706 3377 4764 3403
rect 4806 3437 4864 3463
rect 4806 3403 4818 3437
rect 4852 3403 4864 3437
rect 4806 3377 4864 3403
rect 4906 3437 4964 3463
rect 4906 3403 4918 3437
rect 4952 3403 4964 3437
rect 4906 3377 4964 3403
rect 5006 3437 5064 3463
rect 5006 3403 5018 3437
rect 5052 3403 5064 3437
rect 5006 3377 5064 3403
rect 5106 3437 5164 3463
rect 5106 3403 5118 3437
rect 5152 3403 5164 3437
rect 5106 3377 5164 3403
rect 5206 3437 5264 3463
rect 5206 3403 5218 3437
rect 5252 3403 5264 3437
rect 5206 3377 5264 3403
rect 5306 3437 5364 3463
rect 5306 3403 5318 3437
rect 5352 3403 5364 3437
rect 5306 3377 5364 3403
rect 5406 3437 5464 3463
rect 5406 3403 5418 3437
rect 5452 3403 5464 3437
rect 5406 3377 5464 3403
rect 5506 3437 5564 3463
rect 5506 3403 5518 3437
rect 5552 3403 5564 3437
rect 5506 3377 5564 3403
rect 5606 3437 5664 3463
rect 5606 3403 5618 3437
rect 5652 3403 5664 3437
rect 5606 3377 5664 3403
rect 5706 3437 5764 3463
rect 5706 3403 5718 3437
rect 5752 3403 5764 3437
rect 5706 3377 5764 3403
rect 5806 3437 5864 3463
rect 5806 3403 5818 3437
rect 5852 3403 5864 3437
rect 5806 3377 5864 3403
rect 5906 3437 5964 3463
rect 5906 3403 5912 3437
rect 5952 3403 5964 3437
rect 5906 3377 5964 3403
rect 6006 3437 6064 3463
rect 6006 3403 6018 3437
rect 6058 3403 6064 3437
rect 6006 3377 6064 3403
rect 6106 3437 6164 3463
rect 6106 3403 6118 3437
rect 6152 3403 6164 3437
rect 6106 3377 6164 3403
rect 6206 3437 6264 3463
rect 6206 3403 6218 3437
rect 6252 3403 6264 3437
rect 6206 3377 6264 3403
rect 6306 3437 6364 3463
rect 6306 3403 6318 3437
rect 6352 3403 6364 3437
rect 6306 3377 6364 3403
rect 6406 3437 6464 3463
rect 6618 3456 6862 3490
rect 6406 3403 6418 3437
rect 6452 3403 6464 3437
rect 6508 3418 6516 3452
rect 6558 3418 6574 3452
rect 6618 3437 6652 3456
rect 6406 3377 6464 3403
rect 6828 3437 6862 3456
rect 6618 3387 6652 3403
rect 6696 3388 6712 3422
rect 6754 3388 6762 3422
rect 6828 3387 6862 3403
rect 6928 3437 7162 3453
rect 6962 3403 7028 3437
rect 7062 3403 7128 3437
rect 6928 3387 7162 3403
rect 7228 3437 7362 3453
rect 7262 3403 7328 3437
rect 7228 3387 7362 3403
rect 7428 3437 7462 3453
rect 7428 3387 7462 3403
rect 6 3297 64 3323
rect 6 3263 18 3297
rect 58 3263 64 3297
rect 6 3237 64 3263
rect 106 3297 164 3323
rect 106 3263 118 3297
rect 152 3263 164 3297
rect 106 3237 164 3263
rect 206 3297 264 3323
rect 206 3263 218 3297
rect 252 3263 264 3297
rect 206 3237 264 3263
rect 306 3297 364 3323
rect 306 3263 318 3297
rect 352 3263 364 3297
rect 306 3237 364 3263
rect 406 3297 464 3323
rect 406 3263 418 3297
rect 452 3263 464 3297
rect 406 3237 464 3263
rect 506 3297 564 3323
rect 506 3263 518 3297
rect 552 3263 564 3297
rect 506 3237 564 3263
rect 606 3297 664 3323
rect 606 3263 618 3297
rect 652 3263 664 3297
rect 606 3237 664 3263
rect 706 3297 764 3323
rect 706 3263 718 3297
rect 752 3263 764 3297
rect 706 3237 764 3263
rect 806 3297 864 3323
rect 806 3263 818 3297
rect 852 3263 864 3297
rect 806 3237 864 3263
rect 906 3297 964 3323
rect 906 3263 918 3297
rect 952 3263 964 3297
rect 906 3237 964 3263
rect 1006 3297 1064 3323
rect 1006 3263 1018 3297
rect 1052 3263 1064 3297
rect 1006 3237 1064 3263
rect 1106 3297 1164 3323
rect 1106 3263 1118 3297
rect 1152 3263 1164 3297
rect 1106 3237 1164 3263
rect 1206 3297 1264 3323
rect 1206 3263 1212 3297
rect 1252 3263 1264 3297
rect 1206 3237 1264 3263
rect 1306 3297 1364 3323
rect 1306 3263 1318 3297
rect 1358 3263 1364 3297
rect 1306 3237 1364 3263
rect 1406 3297 1464 3323
rect 1406 3263 1418 3297
rect 1452 3263 1464 3297
rect 1406 3237 1464 3263
rect 1506 3297 1564 3323
rect 1506 3263 1518 3297
rect 1552 3263 1564 3297
rect 1506 3237 1564 3263
rect 1606 3297 1664 3323
rect 1606 3263 1618 3297
rect 1652 3263 1664 3297
rect 1606 3237 1664 3263
rect 1706 3297 1764 3323
rect 1706 3263 1718 3297
rect 1752 3263 1764 3297
rect 1706 3237 1764 3263
rect 1806 3297 1864 3323
rect 1806 3263 1818 3297
rect 1852 3263 1864 3297
rect 1806 3237 1864 3263
rect 1906 3297 1964 3323
rect 1906 3263 1918 3297
rect 1952 3263 1964 3297
rect 1906 3237 1964 3263
rect 2006 3297 2064 3323
rect 2006 3263 2018 3297
rect 2052 3263 2064 3297
rect 2006 3237 2064 3263
rect 2106 3297 2164 3323
rect 2106 3263 2118 3297
rect 2152 3263 2164 3297
rect 2106 3237 2164 3263
rect 2206 3297 2264 3323
rect 2206 3263 2218 3297
rect 2252 3263 2264 3297
rect 2206 3237 2264 3263
rect 2306 3297 2364 3323
rect 2306 3263 2318 3297
rect 2352 3263 2364 3297
rect 2306 3237 2364 3263
rect 2406 3297 2464 3323
rect 2406 3263 2418 3297
rect 2452 3263 2464 3297
rect 2406 3237 2464 3263
rect 2506 3297 2564 3323
rect 2506 3263 2518 3297
rect 2552 3263 2564 3297
rect 2506 3237 2564 3263
rect 2606 3297 2664 3323
rect 2606 3263 2618 3297
rect 2652 3263 2664 3297
rect 2606 3237 2664 3263
rect 2706 3297 2764 3323
rect 2706 3263 2712 3297
rect 2752 3263 2764 3297
rect 2706 3237 2764 3263
rect 2806 3297 2864 3323
rect 2806 3263 2818 3297
rect 2858 3263 2864 3297
rect 2806 3237 2864 3263
rect 2906 3297 2964 3323
rect 2906 3263 2912 3297
rect 2952 3263 2964 3297
rect 2906 3237 2964 3263
rect 3006 3297 3064 3323
rect 3006 3263 3018 3297
rect 3058 3263 3064 3297
rect 3006 3237 3064 3263
rect 3106 3297 3164 3323
rect 3106 3263 3118 3297
rect 3152 3263 3164 3297
rect 3106 3237 3164 3263
rect 3206 3297 3264 3323
rect 3206 3263 3218 3297
rect 3252 3263 3264 3297
rect 3206 3237 3264 3263
rect 3306 3297 3364 3323
rect 3306 3263 3318 3297
rect 3352 3263 3364 3297
rect 3306 3237 3364 3263
rect 3406 3297 3464 3323
rect 3406 3263 3418 3297
rect 3452 3263 3464 3297
rect 3406 3237 3464 3263
rect 3506 3297 3564 3323
rect 3506 3263 3518 3297
rect 3552 3263 3564 3297
rect 3506 3237 3564 3263
rect 3606 3297 3664 3323
rect 3606 3263 3618 3297
rect 3652 3263 3664 3297
rect 3606 3237 3664 3263
rect 3706 3297 3764 3323
rect 3706 3263 3718 3297
rect 3752 3263 3764 3297
rect 3706 3237 3764 3263
rect 3806 3297 3864 3323
rect 3806 3263 3818 3297
rect 3852 3263 3864 3297
rect 3806 3237 3864 3263
rect 3906 3297 3964 3323
rect 3906 3263 3918 3297
rect 3952 3263 3964 3297
rect 3906 3237 3964 3263
rect 4006 3297 4064 3323
rect 4006 3263 4018 3297
rect 4052 3263 4064 3297
rect 4006 3237 4064 3263
rect 4106 3297 4164 3323
rect 4106 3263 4118 3297
rect 4152 3263 4164 3297
rect 4106 3237 4164 3263
rect 4206 3297 4264 3323
rect 4206 3263 4218 3297
rect 4252 3263 4264 3297
rect 4206 3237 4264 3263
rect 4306 3297 4364 3323
rect 4306 3263 4312 3297
rect 4352 3263 4364 3297
rect 4306 3237 4364 3263
rect 4406 3297 4464 3323
rect 4406 3263 4418 3297
rect 4458 3263 4464 3297
rect 4406 3237 4464 3263
rect 4506 3297 4564 3323
rect 4506 3263 4518 3297
rect 4552 3263 4564 3297
rect 4506 3237 4564 3263
rect 4606 3297 4664 3323
rect 4606 3263 4618 3297
rect 4652 3263 4664 3297
rect 4606 3237 4664 3263
rect 4706 3297 4764 3323
rect 4706 3263 4718 3297
rect 4752 3263 4764 3297
rect 4706 3237 4764 3263
rect 4806 3297 4864 3323
rect 4806 3263 4812 3297
rect 4852 3263 4864 3297
rect 4806 3237 4864 3263
rect 4906 3297 4964 3323
rect 4906 3263 4918 3297
rect 4958 3263 4964 3297
rect 4906 3237 4964 3263
rect 5006 3297 5064 3323
rect 5006 3263 5018 3297
rect 5052 3263 5064 3297
rect 5006 3237 5064 3263
rect 5106 3297 5164 3323
rect 5106 3263 5118 3297
rect 5152 3263 5164 3297
rect 5106 3237 5164 3263
rect 5206 3297 5264 3323
rect 5206 3263 5218 3297
rect 5252 3263 5264 3297
rect 5206 3237 5264 3263
rect 5306 3297 5364 3323
rect 5306 3263 5318 3297
rect 5352 3263 5364 3297
rect 5306 3237 5364 3263
rect 5406 3297 5464 3323
rect 5406 3263 5418 3297
rect 5452 3263 5464 3297
rect 5406 3237 5464 3263
rect 5506 3297 5564 3323
rect 5506 3263 5512 3297
rect 5552 3263 5564 3297
rect 5506 3237 5564 3263
rect 5606 3297 5664 3323
rect 5606 3263 5618 3297
rect 5658 3263 5664 3297
rect 5606 3237 5664 3263
rect 5706 3297 5764 3323
rect 5706 3263 5718 3297
rect 5752 3263 5764 3297
rect 5706 3237 5764 3263
rect 5806 3297 5864 3323
rect 5806 3263 5818 3297
rect 5852 3263 5864 3297
rect 5806 3237 5864 3263
rect 5906 3297 5964 3323
rect 5906 3263 5918 3297
rect 5952 3263 5964 3297
rect 5906 3237 5964 3263
rect 6006 3297 6064 3323
rect 6006 3263 6018 3297
rect 6052 3263 6064 3297
rect 6006 3237 6064 3263
rect 6106 3297 6164 3323
rect 6106 3263 6118 3297
rect 6152 3263 6164 3297
rect 6106 3237 6164 3263
rect 6206 3297 6264 3323
rect 6206 3263 6218 3297
rect 6252 3263 6264 3297
rect 6206 3237 6264 3263
rect 6306 3297 6364 3323
rect 6306 3263 6318 3297
rect 6352 3263 6364 3297
rect 6306 3237 6364 3263
rect 6406 3297 6464 3323
rect 6618 3316 6862 3350
rect 6406 3263 6418 3297
rect 6452 3263 6464 3297
rect 6508 3278 6516 3312
rect 6558 3278 6574 3312
rect 6618 3297 6652 3316
rect 6406 3237 6464 3263
rect 6828 3313 6862 3316
rect 6828 3297 6962 3313
rect 6618 3247 6652 3263
rect 6696 3248 6712 3282
rect 6754 3248 6762 3282
rect 6862 3263 6928 3297
rect 6828 3247 6962 3263
rect 7028 3297 7062 3313
rect 7028 3247 7062 3263
rect 7128 3297 7362 3313
rect 7162 3263 7228 3297
rect 7262 3263 7328 3297
rect 7128 3247 7362 3263
rect 7428 3297 7462 3313
rect 7428 3247 7462 3263
rect 6 3157 64 3183
rect 6 3123 18 3157
rect 52 3123 64 3157
rect 6 3097 64 3123
rect 106 3157 164 3183
rect 106 3123 118 3157
rect 152 3123 164 3157
rect 106 3097 164 3123
rect 206 3157 264 3183
rect 206 3123 218 3157
rect 252 3123 264 3157
rect 206 3097 264 3123
rect 306 3157 364 3183
rect 306 3123 318 3157
rect 352 3123 364 3157
rect 306 3097 364 3123
rect 406 3157 464 3183
rect 406 3123 412 3157
rect 452 3123 464 3157
rect 406 3097 464 3123
rect 506 3157 564 3183
rect 506 3123 518 3157
rect 558 3123 564 3157
rect 506 3097 564 3123
rect 606 3157 664 3183
rect 606 3123 618 3157
rect 652 3123 664 3157
rect 606 3097 664 3123
rect 706 3157 764 3183
rect 706 3123 718 3157
rect 752 3123 764 3157
rect 706 3097 764 3123
rect 806 3157 864 3183
rect 806 3123 818 3157
rect 852 3123 864 3157
rect 806 3097 864 3123
rect 906 3157 964 3183
rect 906 3123 918 3157
rect 952 3123 964 3157
rect 906 3097 964 3123
rect 1006 3157 1064 3183
rect 1006 3123 1018 3157
rect 1052 3123 1064 3157
rect 1006 3097 1064 3123
rect 1106 3157 1164 3183
rect 1106 3123 1112 3157
rect 1152 3123 1164 3157
rect 1106 3097 1164 3123
rect 1206 3157 1264 3183
rect 1206 3123 1218 3157
rect 1258 3123 1264 3157
rect 1206 3097 1264 3123
rect 1306 3157 1364 3183
rect 1306 3123 1318 3157
rect 1352 3123 1364 3157
rect 1306 3097 1364 3123
rect 1406 3157 1464 3183
rect 1406 3123 1418 3157
rect 1452 3123 1464 3157
rect 1406 3097 1464 3123
rect 1506 3157 1564 3183
rect 1506 3123 1518 3157
rect 1552 3123 1564 3157
rect 1506 3097 1564 3123
rect 1606 3157 1664 3183
rect 1606 3123 1618 3157
rect 1652 3123 1664 3157
rect 1606 3097 1664 3123
rect 1706 3157 1764 3183
rect 1706 3123 1718 3157
rect 1752 3123 1764 3157
rect 1706 3097 1764 3123
rect 1806 3157 1864 3183
rect 1806 3123 1818 3157
rect 1852 3123 1864 3157
rect 1806 3097 1864 3123
rect 1906 3157 1964 3183
rect 1906 3123 1918 3157
rect 1952 3123 1964 3157
rect 1906 3097 1964 3123
rect 2006 3157 2064 3183
rect 2006 3123 2018 3157
rect 2052 3123 2064 3157
rect 2006 3097 2064 3123
rect 2106 3157 2164 3183
rect 2106 3123 2118 3157
rect 2152 3123 2164 3157
rect 2106 3097 2164 3123
rect 2206 3157 2264 3183
rect 2206 3123 2218 3157
rect 2252 3123 2264 3157
rect 2206 3097 2264 3123
rect 2306 3157 2364 3183
rect 2306 3123 2318 3157
rect 2352 3123 2364 3157
rect 2306 3097 2364 3123
rect 2406 3157 2464 3183
rect 2406 3123 2412 3157
rect 2452 3123 2464 3157
rect 2406 3097 2464 3123
rect 2506 3157 2564 3183
rect 2506 3123 2518 3157
rect 2558 3123 2564 3157
rect 2506 3097 2564 3123
rect 2606 3157 2664 3183
rect 2606 3123 2618 3157
rect 2652 3123 2664 3157
rect 2606 3097 2664 3123
rect 2706 3157 2764 3183
rect 2706 3123 2718 3157
rect 2752 3123 2764 3157
rect 2706 3097 2764 3123
rect 2806 3157 2864 3183
rect 2806 3123 2818 3157
rect 2852 3123 2864 3157
rect 2806 3097 2864 3123
rect 2906 3157 2964 3183
rect 2906 3123 2918 3157
rect 2952 3123 2964 3157
rect 2906 3097 2964 3123
rect 3006 3157 3064 3183
rect 3006 3123 3018 3157
rect 3052 3123 3064 3157
rect 3006 3097 3064 3123
rect 3106 3157 3164 3183
rect 3106 3123 3118 3157
rect 3152 3123 3164 3157
rect 3106 3097 3164 3123
rect 3206 3157 3264 3183
rect 3206 3123 3212 3157
rect 3252 3123 3264 3157
rect 3206 3097 3264 3123
rect 3306 3157 3364 3183
rect 3306 3123 3318 3157
rect 3358 3123 3364 3157
rect 3306 3097 3364 3123
rect 3406 3157 3464 3183
rect 3406 3123 3418 3157
rect 3452 3123 3464 3157
rect 3406 3097 3464 3123
rect 3506 3157 3564 3183
rect 3506 3123 3518 3157
rect 3552 3123 3564 3157
rect 3506 3097 3564 3123
rect 3606 3157 3664 3183
rect 3606 3123 3612 3157
rect 3652 3123 3664 3157
rect 3606 3097 3664 3123
rect 3706 3157 3764 3183
rect 3706 3123 3718 3157
rect 3758 3123 3764 3157
rect 3706 3097 3764 3123
rect 3806 3157 3864 3183
rect 3806 3123 3818 3157
rect 3852 3123 3864 3157
rect 3806 3097 3864 3123
rect 3906 3157 3964 3183
rect 3906 3123 3918 3157
rect 3952 3123 3964 3157
rect 3906 3097 3964 3123
rect 4006 3157 4064 3183
rect 4006 3123 4018 3157
rect 4052 3123 4064 3157
rect 4006 3097 4064 3123
rect 4106 3157 4164 3183
rect 4106 3123 4118 3157
rect 4152 3123 4164 3157
rect 4106 3097 4164 3123
rect 4206 3157 4264 3183
rect 4206 3123 4212 3157
rect 4252 3123 4264 3157
rect 4206 3097 4264 3123
rect 4306 3157 4364 3183
rect 4306 3123 4318 3157
rect 4358 3123 4364 3157
rect 4306 3097 4364 3123
rect 4406 3157 4464 3183
rect 4406 3123 4418 3157
rect 4452 3123 4464 3157
rect 4406 3097 4464 3123
rect 4506 3157 4564 3183
rect 4506 3123 4512 3157
rect 4552 3123 4564 3157
rect 4506 3097 4564 3123
rect 4606 3157 4664 3183
rect 4606 3123 4618 3157
rect 4658 3123 4664 3157
rect 4606 3097 4664 3123
rect 4706 3157 4764 3183
rect 4706 3123 4712 3157
rect 4752 3123 4764 3157
rect 4706 3097 4764 3123
rect 4806 3157 4864 3183
rect 4806 3123 4818 3157
rect 4858 3123 4864 3157
rect 4806 3097 4864 3123
rect 4906 3157 4964 3183
rect 4906 3123 4918 3157
rect 4952 3123 4964 3157
rect 4906 3097 4964 3123
rect 5006 3157 5064 3183
rect 5006 3123 5012 3157
rect 5052 3123 5064 3157
rect 5006 3097 5064 3123
rect 5106 3157 5164 3183
rect 5106 3123 5118 3157
rect 5158 3123 5164 3157
rect 5106 3097 5164 3123
rect 5206 3157 5264 3183
rect 5206 3123 5218 3157
rect 5252 3123 5264 3157
rect 5206 3097 5264 3123
rect 5306 3157 5364 3183
rect 5306 3123 5318 3157
rect 5352 3123 5364 3157
rect 5306 3097 5364 3123
rect 5406 3157 5464 3183
rect 5406 3123 5418 3157
rect 5452 3123 5464 3157
rect 5406 3097 5464 3123
rect 5506 3157 5564 3183
rect 5506 3123 5512 3157
rect 5552 3123 5564 3157
rect 5506 3097 5564 3123
rect 5606 3157 5664 3183
rect 5606 3123 5618 3157
rect 5658 3123 5664 3157
rect 5606 3097 5664 3123
rect 5706 3157 5764 3183
rect 5706 3123 5712 3157
rect 5752 3123 5764 3157
rect 5706 3097 5764 3123
rect 5806 3157 5864 3183
rect 5806 3123 5818 3157
rect 5858 3123 5864 3157
rect 5806 3097 5864 3123
rect 5906 3157 5964 3183
rect 5906 3123 5918 3157
rect 5952 3123 5964 3157
rect 5906 3097 5964 3123
rect 6006 3157 6064 3183
rect 6006 3123 6018 3157
rect 6052 3123 6064 3157
rect 6006 3097 6064 3123
rect 6106 3157 6164 3183
rect 6106 3123 6118 3157
rect 6152 3123 6164 3157
rect 6106 3097 6164 3123
rect 6206 3157 6264 3183
rect 6206 3123 6218 3157
rect 6252 3123 6264 3157
rect 6206 3097 6264 3123
rect 6306 3157 6364 3183
rect 6306 3123 6318 3157
rect 6352 3123 6364 3157
rect 6306 3097 6364 3123
rect 6406 3157 6464 3183
rect 6618 3176 6862 3210
rect 6406 3123 6418 3157
rect 6452 3123 6464 3157
rect 6508 3138 6516 3172
rect 6558 3138 6574 3172
rect 6618 3157 6652 3176
rect 6406 3097 6464 3123
rect 6828 3157 6862 3176
rect 6618 3107 6652 3123
rect 6696 3108 6712 3142
rect 6754 3108 6762 3142
rect 6828 3107 6862 3123
rect 6928 3157 7062 3173
rect 6962 3123 7028 3157
rect 6928 3107 7062 3123
rect 7128 3157 7362 3173
rect 7162 3123 7228 3157
rect 7262 3123 7328 3157
rect 7128 3107 7362 3123
rect 7428 3157 7462 3173
rect 7428 3107 7462 3123
rect 6 3017 64 3043
rect 6 2983 18 3017
rect 52 2983 64 3017
rect 6 2957 64 2983
rect 106 3017 164 3043
rect 106 2983 118 3017
rect 152 2983 164 3017
rect 106 2957 164 2983
rect 206 3017 264 3043
rect 206 2983 218 3017
rect 252 2983 264 3017
rect 206 2957 264 2983
rect 306 3017 364 3043
rect 306 2983 318 3017
rect 352 2983 364 3017
rect 306 2957 364 2983
rect 406 3017 464 3043
rect 406 2983 418 3017
rect 452 2983 464 3017
rect 406 2957 464 2983
rect 506 3017 564 3043
rect 506 2983 518 3017
rect 552 2983 564 3017
rect 506 2957 564 2983
rect 606 3017 664 3043
rect 606 2983 618 3017
rect 652 2983 664 3017
rect 606 2957 664 2983
rect 706 3017 764 3043
rect 706 2983 718 3017
rect 752 2983 764 3017
rect 706 2957 764 2983
rect 806 3017 864 3043
rect 806 2983 818 3017
rect 852 2983 864 3017
rect 806 2957 864 2983
rect 906 3017 964 3043
rect 906 2983 918 3017
rect 952 2983 964 3017
rect 906 2957 964 2983
rect 1006 3017 1064 3043
rect 1006 2983 1018 3017
rect 1052 2983 1064 3017
rect 1006 2957 1064 2983
rect 1106 3017 1164 3043
rect 1106 2983 1118 3017
rect 1152 2983 1164 3017
rect 1106 2957 1164 2983
rect 1206 3017 1264 3043
rect 1206 2983 1218 3017
rect 1252 2983 1264 3017
rect 1206 2957 1264 2983
rect 1306 3017 1364 3043
rect 1306 2983 1318 3017
rect 1352 2983 1364 3017
rect 1306 2957 1364 2983
rect 1406 3017 1464 3043
rect 1406 2983 1418 3017
rect 1452 2983 1464 3017
rect 1406 2957 1464 2983
rect 1506 3017 1564 3043
rect 1506 2983 1518 3017
rect 1552 2983 1564 3017
rect 1506 2957 1564 2983
rect 1606 3017 1664 3043
rect 1606 2983 1618 3017
rect 1652 2983 1664 3017
rect 1606 2957 1664 2983
rect 1706 3017 1764 3043
rect 1706 2983 1718 3017
rect 1752 2983 1764 3017
rect 1706 2957 1764 2983
rect 1806 3017 1864 3043
rect 1806 2983 1818 3017
rect 1852 2983 1864 3017
rect 1806 2957 1864 2983
rect 1906 3017 1964 3043
rect 1906 2983 1918 3017
rect 1952 2983 1964 3017
rect 1906 2957 1964 2983
rect 2006 3017 2064 3043
rect 2006 2983 2018 3017
rect 2052 2983 2064 3017
rect 2006 2957 2064 2983
rect 2106 3017 2164 3043
rect 2106 2983 2118 3017
rect 2152 2983 2164 3017
rect 2106 2957 2164 2983
rect 2206 3017 2264 3043
rect 2206 2983 2218 3017
rect 2252 2983 2264 3017
rect 2206 2957 2264 2983
rect 2306 3017 2364 3043
rect 2306 2983 2318 3017
rect 2352 2983 2364 3017
rect 2306 2957 2364 2983
rect 2406 3017 2464 3043
rect 2406 2983 2418 3017
rect 2452 2983 2464 3017
rect 2406 2957 2464 2983
rect 2506 3017 2564 3043
rect 2506 2983 2518 3017
rect 2552 2983 2564 3017
rect 2506 2957 2564 2983
rect 2606 3017 2664 3043
rect 2606 2983 2618 3017
rect 2652 2983 2664 3017
rect 2606 2957 2664 2983
rect 2706 3017 2764 3043
rect 2706 2983 2718 3017
rect 2752 2983 2764 3017
rect 2706 2957 2764 2983
rect 2806 3017 2864 3043
rect 2806 2983 2818 3017
rect 2852 2983 2864 3017
rect 2806 2957 2864 2983
rect 2906 3017 2964 3043
rect 2906 2983 2918 3017
rect 2952 2983 2964 3017
rect 2906 2957 2964 2983
rect 3006 3017 3064 3043
rect 3006 2983 3018 3017
rect 3052 2983 3064 3017
rect 3006 2957 3064 2983
rect 3106 3017 3164 3043
rect 3106 2983 3118 3017
rect 3152 2983 3164 3017
rect 3106 2957 3164 2983
rect 3206 3017 3264 3043
rect 3206 2983 3218 3017
rect 3252 2983 3264 3017
rect 3206 2957 3264 2983
rect 3306 3017 3364 3043
rect 3306 2983 3312 3017
rect 3352 2983 3364 3017
rect 3306 2957 3364 2983
rect 3406 3017 3464 3043
rect 3406 2983 3418 3017
rect 3458 2983 3464 3017
rect 3406 2957 3464 2983
rect 3506 3017 3564 3043
rect 3506 2983 3518 3017
rect 3552 2983 3564 3017
rect 3506 2957 3564 2983
rect 3606 3017 3664 3043
rect 3606 2983 3618 3017
rect 3652 2983 3664 3017
rect 3606 2957 3664 2983
rect 3706 3017 3764 3043
rect 3706 2983 3718 3017
rect 3752 2983 3764 3017
rect 3706 2957 3764 2983
rect 3806 3017 3864 3043
rect 3806 2983 3812 3017
rect 3852 2983 3864 3017
rect 3806 2957 3864 2983
rect 3906 3017 3964 3043
rect 3906 2983 3918 3017
rect 3958 2983 3964 3017
rect 3906 2957 3964 2983
rect 4006 3017 4064 3043
rect 4006 2983 4012 3017
rect 4052 2983 4064 3017
rect 4006 2957 4064 2983
rect 4106 3017 4164 3043
rect 4106 2983 4118 3017
rect 4158 2983 4164 3017
rect 4106 2957 4164 2983
rect 4206 3017 4264 3043
rect 4206 2983 4218 3017
rect 4252 2983 4264 3017
rect 4206 2957 4264 2983
rect 4306 3017 4364 3043
rect 4306 2983 4318 3017
rect 4352 2983 4364 3017
rect 4306 2957 4364 2983
rect 4406 3017 4464 3043
rect 4406 2983 4418 3017
rect 4452 2983 4464 3017
rect 4406 2957 4464 2983
rect 4506 3017 4564 3043
rect 4506 2983 4512 3017
rect 4552 2983 4564 3017
rect 4506 2957 4564 2983
rect 4606 3017 4664 3043
rect 4606 2983 4618 3017
rect 4658 2983 4664 3017
rect 4606 2957 4664 2983
rect 4706 3017 4764 3043
rect 4706 2983 4718 3017
rect 4752 2983 4764 3017
rect 4706 2957 4764 2983
rect 4806 3017 4864 3043
rect 4806 2983 4818 3017
rect 4852 2983 4864 3017
rect 4806 2957 4864 2983
rect 4906 3017 4964 3043
rect 4906 2983 4918 3017
rect 4952 2983 4964 3017
rect 4906 2957 4964 2983
rect 5006 3017 5064 3043
rect 5006 2983 5018 3017
rect 5052 2983 5064 3017
rect 5006 2957 5064 2983
rect 5106 3017 5164 3043
rect 5106 2983 5118 3017
rect 5152 2983 5164 3017
rect 5106 2957 5164 2983
rect 5206 3017 5264 3043
rect 5206 2983 5218 3017
rect 5252 2983 5264 3017
rect 5206 2957 5264 2983
rect 5306 3017 5364 3043
rect 5306 2983 5318 3017
rect 5352 2983 5364 3017
rect 5306 2957 5364 2983
rect 5406 3017 5464 3043
rect 5406 2983 5418 3017
rect 5452 2983 5464 3017
rect 5406 2957 5464 2983
rect 5506 3017 5564 3043
rect 5506 2983 5518 3017
rect 5552 2983 5564 3017
rect 5506 2957 5564 2983
rect 5606 3017 5664 3043
rect 5606 2983 5618 3017
rect 5652 2983 5664 3017
rect 5606 2957 5664 2983
rect 5706 3017 5764 3043
rect 5706 2983 5718 3017
rect 5752 2983 5764 3017
rect 5706 2957 5764 2983
rect 5806 3017 5864 3043
rect 5806 2983 5818 3017
rect 5852 2983 5864 3017
rect 5806 2957 5864 2983
rect 5906 3017 5964 3043
rect 5906 2983 5912 3017
rect 5952 2983 5964 3017
rect 5906 2957 5964 2983
rect 6006 3017 6064 3043
rect 6006 2983 6018 3017
rect 6058 2983 6064 3017
rect 6006 2957 6064 2983
rect 6106 3017 6164 3043
rect 6106 2983 6118 3017
rect 6152 2983 6164 3017
rect 6106 2957 6164 2983
rect 6206 3017 6264 3043
rect 6206 2983 6218 3017
rect 6252 2983 6264 3017
rect 6206 2957 6264 2983
rect 6306 3017 6364 3043
rect 6306 2983 6318 3017
rect 6352 2983 6364 3017
rect 6306 2957 6364 2983
rect 6406 3017 6464 3043
rect 6618 3036 6862 3070
rect 6406 2983 6418 3017
rect 6452 2983 6464 3017
rect 6508 2998 6516 3032
rect 6558 2998 6574 3032
rect 6618 3017 6652 3036
rect 6406 2957 6464 2983
rect 6828 3033 6862 3036
rect 6828 3017 6962 3033
rect 6618 2967 6652 2983
rect 6696 2968 6712 3002
rect 6754 2968 6762 3002
rect 6862 2983 6928 3017
rect 6828 2967 6962 2983
rect 7028 3017 7162 3033
rect 7062 2983 7128 3017
rect 7028 2967 7162 2983
rect 7228 3017 7262 3033
rect 7228 2967 7262 2983
rect 7328 3017 7462 3033
rect 7362 2983 7428 3017
rect 7328 2967 7462 2983
rect 6 2877 64 2903
rect 6 2843 18 2877
rect 52 2843 64 2877
rect 6 2817 64 2843
rect 106 2877 164 2903
rect 106 2843 118 2877
rect 152 2843 164 2877
rect 106 2817 164 2843
rect 206 2877 264 2903
rect 206 2843 218 2877
rect 252 2843 264 2877
rect 206 2817 264 2843
rect 306 2877 364 2903
rect 306 2843 312 2877
rect 352 2843 364 2877
rect 306 2817 364 2843
rect 406 2877 464 2903
rect 406 2843 418 2877
rect 458 2843 464 2877
rect 406 2817 464 2843
rect 506 2877 564 2903
rect 506 2843 518 2877
rect 552 2843 564 2877
rect 506 2817 564 2843
rect 606 2877 664 2903
rect 606 2843 618 2877
rect 652 2843 664 2877
rect 606 2817 664 2843
rect 706 2877 764 2903
rect 706 2843 712 2877
rect 752 2843 764 2877
rect 706 2817 764 2843
rect 806 2877 864 2903
rect 806 2843 818 2877
rect 858 2843 864 2877
rect 806 2817 864 2843
rect 906 2877 964 2903
rect 906 2843 918 2877
rect 952 2843 964 2877
rect 906 2817 964 2843
rect 1006 2877 1064 2903
rect 1006 2843 1018 2877
rect 1052 2843 1064 2877
rect 1006 2817 1064 2843
rect 1106 2877 1164 2903
rect 1106 2843 1118 2877
rect 1152 2843 1164 2877
rect 1106 2817 1164 2843
rect 1206 2877 1264 2903
rect 1206 2843 1218 2877
rect 1252 2843 1264 2877
rect 1206 2817 1264 2843
rect 1306 2877 1364 2903
rect 1306 2843 1318 2877
rect 1352 2843 1364 2877
rect 1306 2817 1364 2843
rect 1406 2877 1464 2903
rect 1406 2843 1412 2877
rect 1452 2843 1464 2877
rect 1406 2817 1464 2843
rect 1506 2877 1564 2903
rect 1506 2843 1518 2877
rect 1558 2843 1564 2877
rect 1506 2817 1564 2843
rect 1606 2877 1664 2903
rect 1606 2843 1618 2877
rect 1652 2843 1664 2877
rect 1606 2817 1664 2843
rect 1706 2877 1764 2903
rect 1706 2843 1718 2877
rect 1752 2843 1764 2877
rect 1706 2817 1764 2843
rect 1806 2877 1864 2903
rect 1806 2843 1818 2877
rect 1852 2843 1864 2877
rect 1806 2817 1864 2843
rect 1906 2877 1964 2903
rect 1906 2843 1918 2877
rect 1952 2843 1964 2877
rect 1906 2817 1964 2843
rect 2006 2877 2064 2903
rect 2006 2843 2018 2877
rect 2052 2843 2064 2877
rect 2006 2817 2064 2843
rect 2106 2877 2164 2903
rect 2106 2843 2112 2877
rect 2152 2843 2164 2877
rect 2106 2817 2164 2843
rect 2206 2877 2264 2903
rect 2206 2843 2218 2877
rect 2258 2843 2264 2877
rect 2206 2817 2264 2843
rect 2306 2877 2364 2903
rect 2306 2843 2312 2877
rect 2352 2843 2364 2877
rect 2306 2817 2364 2843
rect 2406 2877 2464 2903
rect 2406 2843 2418 2877
rect 2458 2843 2464 2877
rect 2406 2817 2464 2843
rect 2506 2877 2564 2903
rect 2506 2843 2512 2877
rect 2552 2843 2564 2877
rect 2506 2817 2564 2843
rect 2606 2877 2664 2903
rect 2606 2843 2618 2877
rect 2658 2843 2664 2877
rect 2606 2817 2664 2843
rect 2706 2877 2764 2903
rect 2706 2843 2718 2877
rect 2752 2843 2764 2877
rect 2706 2817 2764 2843
rect 2806 2877 2864 2903
rect 2806 2843 2818 2877
rect 2852 2843 2864 2877
rect 2806 2817 2864 2843
rect 2906 2877 2964 2903
rect 2906 2843 2918 2877
rect 2952 2843 2964 2877
rect 2906 2817 2964 2843
rect 3006 2877 3064 2903
rect 3006 2843 3012 2877
rect 3052 2843 3064 2877
rect 3006 2817 3064 2843
rect 3106 2877 3164 2903
rect 3106 2843 3118 2877
rect 3158 2843 3164 2877
rect 3106 2817 3164 2843
rect 3206 2877 3264 2903
rect 3206 2843 3218 2877
rect 3252 2843 3264 2877
rect 3206 2817 3264 2843
rect 3306 2877 3364 2903
rect 3306 2843 3318 2877
rect 3352 2843 3364 2877
rect 3306 2817 3364 2843
rect 3406 2877 3464 2903
rect 3406 2843 3418 2877
rect 3452 2843 3464 2877
rect 3406 2817 3464 2843
rect 3506 2877 3564 2903
rect 3506 2843 3518 2877
rect 3552 2843 3564 2877
rect 3506 2817 3564 2843
rect 3606 2877 3664 2903
rect 3606 2843 3618 2877
rect 3652 2843 3664 2877
rect 3606 2817 3664 2843
rect 3706 2877 3764 2903
rect 3706 2843 3718 2877
rect 3752 2843 3764 2877
rect 3706 2817 3764 2843
rect 3806 2877 3864 2903
rect 3806 2843 3818 2877
rect 3852 2843 3864 2877
rect 3806 2817 3864 2843
rect 3906 2877 3964 2903
rect 3906 2843 3918 2877
rect 3952 2843 3964 2877
rect 3906 2817 3964 2843
rect 4006 2877 4064 2903
rect 4006 2843 4018 2877
rect 4052 2843 4064 2877
rect 4006 2817 4064 2843
rect 4106 2877 4164 2903
rect 4106 2843 4118 2877
rect 4152 2843 4164 2877
rect 4106 2817 4164 2843
rect 4206 2877 4264 2903
rect 4206 2843 4218 2877
rect 4252 2843 4264 2877
rect 4206 2817 4264 2843
rect 4306 2877 4364 2903
rect 4306 2843 4318 2877
rect 4352 2843 4364 2877
rect 4306 2817 4364 2843
rect 4406 2877 4464 2903
rect 4406 2843 4418 2877
rect 4452 2843 4464 2877
rect 4406 2817 4464 2843
rect 4506 2877 4564 2903
rect 4506 2843 4518 2877
rect 4552 2843 4564 2877
rect 4506 2817 4564 2843
rect 4606 2877 4664 2903
rect 4606 2843 4618 2877
rect 4652 2843 4664 2877
rect 4606 2817 4664 2843
rect 4706 2877 4764 2903
rect 4706 2843 4718 2877
rect 4752 2843 4764 2877
rect 4706 2817 4764 2843
rect 4806 2877 4864 2903
rect 4806 2843 4818 2877
rect 4852 2843 4864 2877
rect 4806 2817 4864 2843
rect 4906 2877 4964 2903
rect 4906 2843 4918 2877
rect 4952 2843 4964 2877
rect 4906 2817 4964 2843
rect 5006 2877 5064 2903
rect 5006 2843 5018 2877
rect 5052 2843 5064 2877
rect 5006 2817 5064 2843
rect 5106 2877 5164 2903
rect 5106 2843 5118 2877
rect 5152 2843 5164 2877
rect 5106 2817 5164 2843
rect 5206 2877 5264 2903
rect 5206 2843 5218 2877
rect 5252 2843 5264 2877
rect 5206 2817 5264 2843
rect 5306 2877 5364 2903
rect 5306 2843 5318 2877
rect 5352 2843 5364 2877
rect 5306 2817 5364 2843
rect 5406 2877 5464 2903
rect 5406 2843 5418 2877
rect 5452 2843 5464 2877
rect 5406 2817 5464 2843
rect 5506 2877 5564 2903
rect 5506 2843 5518 2877
rect 5552 2843 5564 2877
rect 5506 2817 5564 2843
rect 5606 2877 5664 2903
rect 5606 2843 5618 2877
rect 5652 2843 5664 2877
rect 5606 2817 5664 2843
rect 5706 2877 5764 2903
rect 5706 2843 5718 2877
rect 5752 2843 5764 2877
rect 5706 2817 5764 2843
rect 5806 2877 5864 2903
rect 5806 2843 5818 2877
rect 5852 2843 5864 2877
rect 5806 2817 5864 2843
rect 5906 2877 5964 2903
rect 5906 2843 5918 2877
rect 5952 2843 5964 2877
rect 5906 2817 5964 2843
rect 6006 2877 6064 2903
rect 6006 2843 6012 2877
rect 6052 2843 6064 2877
rect 6006 2817 6064 2843
rect 6106 2877 6164 2903
rect 6106 2843 6118 2877
rect 6158 2843 6164 2877
rect 6106 2817 6164 2843
rect 6206 2877 6264 2903
rect 6206 2843 6218 2877
rect 6252 2843 6264 2877
rect 6206 2817 6264 2843
rect 6306 2877 6364 2903
rect 6306 2843 6318 2877
rect 6352 2843 6364 2877
rect 6306 2817 6364 2843
rect 6406 2877 6464 2903
rect 6618 2896 6862 2930
rect 6406 2843 6412 2877
rect 6452 2843 6464 2877
rect 6508 2858 6516 2892
rect 6558 2858 6574 2892
rect 6618 2877 6652 2896
rect 6406 2817 6464 2843
rect 6828 2877 6862 2896
rect 6618 2827 6652 2843
rect 6696 2828 6712 2862
rect 6754 2828 6762 2862
rect 6828 2827 6862 2843
rect 6928 2877 7162 2893
rect 6962 2843 7028 2877
rect 7062 2843 7128 2877
rect 6928 2827 7162 2843
rect 7228 2877 7262 2893
rect 7228 2827 7262 2843
rect 7328 2877 7462 2893
rect 7362 2843 7428 2877
rect 7328 2827 7462 2843
rect 6 2737 64 2763
rect 6 2703 18 2737
rect 52 2703 64 2737
rect 6 2677 64 2703
rect 106 2737 164 2763
rect 106 2703 118 2737
rect 152 2703 164 2737
rect 106 2677 164 2703
rect 206 2737 264 2763
rect 206 2703 218 2737
rect 252 2703 264 2737
rect 206 2677 264 2703
rect 306 2737 364 2763
rect 306 2703 318 2737
rect 352 2703 364 2737
rect 306 2677 364 2703
rect 406 2737 464 2763
rect 406 2703 418 2737
rect 452 2703 464 2737
rect 406 2677 464 2703
rect 506 2737 564 2763
rect 506 2703 518 2737
rect 552 2703 564 2737
rect 506 2677 564 2703
rect 606 2737 664 2763
rect 606 2703 618 2737
rect 652 2703 664 2737
rect 606 2677 664 2703
rect 706 2737 764 2763
rect 706 2703 718 2737
rect 752 2703 764 2737
rect 706 2677 764 2703
rect 806 2737 864 2763
rect 806 2703 818 2737
rect 852 2703 864 2737
rect 806 2677 864 2703
rect 906 2737 964 2763
rect 906 2703 918 2737
rect 952 2703 964 2737
rect 906 2677 964 2703
rect 1006 2737 1064 2763
rect 1006 2703 1018 2737
rect 1052 2703 1064 2737
rect 1006 2677 1064 2703
rect 1106 2737 1164 2763
rect 1106 2703 1118 2737
rect 1152 2703 1164 2737
rect 1106 2677 1164 2703
rect 1206 2737 1264 2763
rect 1206 2703 1218 2737
rect 1252 2703 1264 2737
rect 1206 2677 1264 2703
rect 1306 2737 1364 2763
rect 1306 2703 1312 2737
rect 1352 2703 1364 2737
rect 1306 2677 1364 2703
rect 1406 2737 1464 2763
rect 1406 2703 1418 2737
rect 1458 2703 1464 2737
rect 1406 2677 1464 2703
rect 1506 2737 1564 2763
rect 1506 2703 1512 2737
rect 1552 2703 1564 2737
rect 1506 2677 1564 2703
rect 1606 2737 1664 2763
rect 1606 2703 1618 2737
rect 1658 2703 1664 2737
rect 1606 2677 1664 2703
rect 1706 2737 1764 2763
rect 1706 2703 1718 2737
rect 1752 2703 1764 2737
rect 1706 2677 1764 2703
rect 1806 2737 1864 2763
rect 1806 2703 1818 2737
rect 1852 2703 1864 2737
rect 1806 2677 1864 2703
rect 1906 2737 1964 2763
rect 1906 2703 1918 2737
rect 1952 2703 1964 2737
rect 1906 2677 1964 2703
rect 2006 2737 2064 2763
rect 2006 2703 2012 2737
rect 2052 2703 2064 2737
rect 2006 2677 2064 2703
rect 2106 2737 2164 2763
rect 2106 2703 2118 2737
rect 2158 2703 2164 2737
rect 2106 2677 2164 2703
rect 2206 2737 2264 2763
rect 2206 2703 2218 2737
rect 2252 2703 2264 2737
rect 2206 2677 2264 2703
rect 2306 2737 2364 2763
rect 2306 2703 2318 2737
rect 2352 2703 2364 2737
rect 2306 2677 2364 2703
rect 2406 2737 2464 2763
rect 2406 2703 2418 2737
rect 2452 2703 2464 2737
rect 2406 2677 2464 2703
rect 2506 2737 2564 2763
rect 2506 2703 2518 2737
rect 2552 2703 2564 2737
rect 2506 2677 2564 2703
rect 2606 2737 2664 2763
rect 2606 2703 2618 2737
rect 2652 2703 2664 2737
rect 2606 2677 2664 2703
rect 2706 2737 2764 2763
rect 2706 2703 2718 2737
rect 2752 2703 2764 2737
rect 2706 2677 2764 2703
rect 2806 2737 2864 2763
rect 2806 2703 2812 2737
rect 2852 2703 2864 2737
rect 2806 2677 2864 2703
rect 2906 2737 2964 2763
rect 2906 2703 2918 2737
rect 2958 2703 2964 2737
rect 2906 2677 2964 2703
rect 3006 2737 3064 2763
rect 3006 2703 3018 2737
rect 3052 2703 3064 2737
rect 3006 2677 3064 2703
rect 3106 2737 3164 2763
rect 3106 2703 3112 2737
rect 3152 2703 3164 2737
rect 3106 2677 3164 2703
rect 3206 2737 3264 2763
rect 3206 2703 3218 2737
rect 3258 2703 3264 2737
rect 3206 2677 3264 2703
rect 3306 2737 3364 2763
rect 3306 2703 3318 2737
rect 3352 2703 3364 2737
rect 3306 2677 3364 2703
rect 3406 2737 3464 2763
rect 3406 2703 3418 2737
rect 3452 2703 3464 2737
rect 3406 2677 3464 2703
rect 3506 2737 3564 2763
rect 3506 2703 3518 2737
rect 3552 2703 3564 2737
rect 3506 2677 3564 2703
rect 3606 2737 3664 2763
rect 3606 2703 3618 2737
rect 3652 2703 3664 2737
rect 3606 2677 3664 2703
rect 3706 2737 3764 2763
rect 3706 2703 3718 2737
rect 3752 2703 3764 2737
rect 3706 2677 3764 2703
rect 3806 2737 3864 2763
rect 3806 2703 3818 2737
rect 3852 2703 3864 2737
rect 3806 2677 3864 2703
rect 3906 2737 3964 2763
rect 3906 2703 3918 2737
rect 3952 2703 3964 2737
rect 3906 2677 3964 2703
rect 4006 2737 4064 2763
rect 4006 2703 4018 2737
rect 4052 2703 4064 2737
rect 4006 2677 4064 2703
rect 4106 2737 4164 2763
rect 4106 2703 4118 2737
rect 4152 2703 4164 2737
rect 4106 2677 4164 2703
rect 4206 2737 4264 2763
rect 4206 2703 4218 2737
rect 4252 2703 4264 2737
rect 4206 2677 4264 2703
rect 4306 2737 4364 2763
rect 4306 2703 4318 2737
rect 4352 2703 4364 2737
rect 4306 2677 4364 2703
rect 4406 2737 4464 2763
rect 4406 2703 4412 2737
rect 4452 2703 4464 2737
rect 4406 2677 4464 2703
rect 4506 2737 4564 2763
rect 4506 2703 4518 2737
rect 4558 2703 4564 2737
rect 4506 2677 4564 2703
rect 4606 2737 4664 2763
rect 4606 2703 4612 2737
rect 4652 2703 4664 2737
rect 4606 2677 4664 2703
rect 4706 2737 4764 2763
rect 4706 2703 4718 2737
rect 4758 2703 4764 2737
rect 4706 2677 4764 2703
rect 4806 2737 4864 2763
rect 4806 2703 4818 2737
rect 4852 2703 4864 2737
rect 4806 2677 4864 2703
rect 4906 2737 4964 2763
rect 4906 2703 4918 2737
rect 4952 2703 4964 2737
rect 4906 2677 4964 2703
rect 5006 2737 5064 2763
rect 5006 2703 5018 2737
rect 5052 2703 5064 2737
rect 5006 2677 5064 2703
rect 5106 2737 5164 2763
rect 5106 2703 5118 2737
rect 5152 2703 5164 2737
rect 5106 2677 5164 2703
rect 5206 2737 5264 2763
rect 5206 2703 5218 2737
rect 5252 2703 5264 2737
rect 5206 2677 5264 2703
rect 5306 2737 5364 2763
rect 5306 2703 5318 2737
rect 5352 2703 5364 2737
rect 5306 2677 5364 2703
rect 5406 2737 5464 2763
rect 5406 2703 5412 2737
rect 5452 2703 5464 2737
rect 5406 2677 5464 2703
rect 5506 2737 5564 2763
rect 5506 2703 5518 2737
rect 5558 2703 5564 2737
rect 5506 2677 5564 2703
rect 5606 2737 5664 2763
rect 5606 2703 5618 2737
rect 5652 2703 5664 2737
rect 5606 2677 5664 2703
rect 5706 2737 5764 2763
rect 5706 2703 5718 2737
rect 5752 2703 5764 2737
rect 5706 2677 5764 2703
rect 5806 2737 5864 2763
rect 5806 2703 5818 2737
rect 5852 2703 5864 2737
rect 5806 2677 5864 2703
rect 5906 2737 5964 2763
rect 5906 2703 5918 2737
rect 5952 2703 5964 2737
rect 5906 2677 5964 2703
rect 6006 2737 6064 2763
rect 6006 2703 6018 2737
rect 6052 2703 6064 2737
rect 6006 2677 6064 2703
rect 6106 2737 6164 2763
rect 6106 2703 6118 2737
rect 6152 2703 6164 2737
rect 6106 2677 6164 2703
rect 6206 2737 6264 2763
rect 6206 2703 6218 2737
rect 6252 2703 6264 2737
rect 6206 2677 6264 2703
rect 6306 2737 6364 2763
rect 6306 2703 6318 2737
rect 6352 2703 6364 2737
rect 6306 2677 6364 2703
rect 6406 2737 6464 2763
rect 6618 2756 6862 2790
rect 6406 2703 6418 2737
rect 6452 2703 6464 2737
rect 6508 2718 6516 2752
rect 6558 2718 6574 2752
rect 6618 2737 6652 2756
rect 6406 2677 6464 2703
rect 6828 2753 6862 2756
rect 6828 2737 6962 2753
rect 6618 2687 6652 2703
rect 6696 2688 6712 2722
rect 6754 2688 6762 2722
rect 6862 2703 6928 2737
rect 6828 2687 6962 2703
rect 7028 2737 7062 2753
rect 7028 2687 7062 2703
rect 7128 2737 7262 2753
rect 7162 2703 7228 2737
rect 7128 2687 7262 2703
rect 7328 2737 7462 2753
rect 7362 2703 7428 2737
rect 7328 2687 7462 2703
rect 6 2597 64 2623
rect 6 2563 18 2597
rect 52 2563 64 2597
rect 6 2537 64 2563
rect 106 2597 164 2623
rect 106 2563 118 2597
rect 152 2563 164 2597
rect 106 2537 164 2563
rect 206 2597 264 2623
rect 206 2563 218 2597
rect 252 2563 264 2597
rect 206 2537 264 2563
rect 306 2597 364 2623
rect 306 2563 318 2597
rect 352 2563 364 2597
rect 306 2537 364 2563
rect 406 2597 464 2623
rect 406 2563 418 2597
rect 452 2563 464 2597
rect 406 2537 464 2563
rect 506 2597 564 2623
rect 506 2563 518 2597
rect 552 2563 564 2597
rect 506 2537 564 2563
rect 606 2597 664 2623
rect 606 2563 618 2597
rect 652 2563 664 2597
rect 606 2537 664 2563
rect 706 2597 764 2623
rect 706 2563 718 2597
rect 752 2563 764 2597
rect 706 2537 764 2563
rect 806 2597 864 2623
rect 806 2563 818 2597
rect 852 2563 864 2597
rect 806 2537 864 2563
rect 906 2597 964 2623
rect 906 2563 918 2597
rect 952 2563 964 2597
rect 906 2537 964 2563
rect 1006 2597 1064 2623
rect 1006 2563 1018 2597
rect 1052 2563 1064 2597
rect 1006 2537 1064 2563
rect 1106 2597 1164 2623
rect 1106 2563 1118 2597
rect 1152 2563 1164 2597
rect 1106 2537 1164 2563
rect 1206 2597 1264 2623
rect 1206 2563 1218 2597
rect 1252 2563 1264 2597
rect 1206 2537 1264 2563
rect 1306 2597 1364 2623
rect 1306 2563 1318 2597
rect 1352 2563 1364 2597
rect 1306 2537 1364 2563
rect 1406 2597 1464 2623
rect 1406 2563 1418 2597
rect 1452 2563 1464 2597
rect 1406 2537 1464 2563
rect 1506 2597 1564 2623
rect 1506 2563 1512 2597
rect 1552 2563 1564 2597
rect 1506 2537 1564 2563
rect 1606 2597 1664 2623
rect 1606 2563 1618 2597
rect 1658 2563 1664 2597
rect 1606 2537 1664 2563
rect 1706 2597 1764 2623
rect 1706 2563 1718 2597
rect 1752 2563 1764 2597
rect 1706 2537 1764 2563
rect 1806 2597 1864 2623
rect 1806 2563 1818 2597
rect 1852 2563 1864 2597
rect 1806 2537 1864 2563
rect 1906 2597 1964 2623
rect 1906 2563 1918 2597
rect 1952 2563 1964 2597
rect 1906 2537 1964 2563
rect 2006 2597 2064 2623
rect 2006 2563 2018 2597
rect 2052 2563 2064 2597
rect 2006 2537 2064 2563
rect 2106 2597 2164 2623
rect 2106 2563 2112 2597
rect 2152 2563 2164 2597
rect 2106 2537 2164 2563
rect 2206 2597 2264 2623
rect 2206 2563 2218 2597
rect 2258 2563 2264 2597
rect 2206 2537 2264 2563
rect 2306 2597 2364 2623
rect 2306 2563 2318 2597
rect 2352 2563 2364 2597
rect 2306 2537 2364 2563
rect 2406 2597 2464 2623
rect 2406 2563 2412 2597
rect 2452 2563 2464 2597
rect 2406 2537 2464 2563
rect 2506 2597 2564 2623
rect 2506 2563 2518 2597
rect 2558 2563 2564 2597
rect 2506 2537 2564 2563
rect 2606 2597 2664 2623
rect 2606 2563 2612 2597
rect 2652 2563 2664 2597
rect 2606 2537 2664 2563
rect 2706 2597 2764 2623
rect 2706 2563 2718 2597
rect 2758 2563 2764 2597
rect 2706 2537 2764 2563
rect 2806 2597 2864 2623
rect 2806 2563 2818 2597
rect 2852 2563 2864 2597
rect 2806 2537 2864 2563
rect 2906 2597 2964 2623
rect 2906 2563 2918 2597
rect 2952 2563 2964 2597
rect 2906 2537 2964 2563
rect 3006 2597 3064 2623
rect 3006 2563 3018 2597
rect 3052 2563 3064 2597
rect 3006 2537 3064 2563
rect 3106 2597 3164 2623
rect 3106 2563 3118 2597
rect 3152 2563 3164 2597
rect 3106 2537 3164 2563
rect 3206 2597 3264 2623
rect 3206 2563 3212 2597
rect 3252 2563 3264 2597
rect 3206 2537 3264 2563
rect 3306 2597 3364 2623
rect 3306 2563 3318 2597
rect 3358 2563 3364 2597
rect 3306 2537 3364 2563
rect 3406 2597 3464 2623
rect 3406 2563 3412 2597
rect 3452 2563 3464 2597
rect 3406 2537 3464 2563
rect 3506 2597 3564 2623
rect 3506 2563 3518 2597
rect 3558 2563 3564 2597
rect 3506 2537 3564 2563
rect 3606 2597 3664 2623
rect 3606 2563 3618 2597
rect 3652 2563 3664 2597
rect 3606 2537 3664 2563
rect 3706 2597 3764 2623
rect 3706 2563 3718 2597
rect 3752 2563 3764 2597
rect 3706 2537 3764 2563
rect 3806 2597 3864 2623
rect 3806 2563 3818 2597
rect 3852 2563 3864 2597
rect 3806 2537 3864 2563
rect 3906 2597 3964 2623
rect 3906 2563 3918 2597
rect 3952 2563 3964 2597
rect 3906 2537 3964 2563
rect 4006 2597 4064 2623
rect 4006 2563 4018 2597
rect 4052 2563 4064 2597
rect 4006 2537 4064 2563
rect 4106 2597 4164 2623
rect 4106 2563 4118 2597
rect 4152 2563 4164 2597
rect 4106 2537 4164 2563
rect 4206 2597 4264 2623
rect 4206 2563 4218 2597
rect 4252 2563 4264 2597
rect 4206 2537 4264 2563
rect 4306 2597 4364 2623
rect 4306 2563 4318 2597
rect 4352 2563 4364 2597
rect 4306 2537 4364 2563
rect 4406 2597 4464 2623
rect 4406 2563 4418 2597
rect 4452 2563 4464 2597
rect 4406 2537 4464 2563
rect 4506 2597 4564 2623
rect 4506 2563 4518 2597
rect 4552 2563 4564 2597
rect 4506 2537 4564 2563
rect 4606 2597 4664 2623
rect 4606 2563 4618 2597
rect 4652 2563 4664 2597
rect 4606 2537 4664 2563
rect 4706 2597 4764 2623
rect 4706 2563 4718 2597
rect 4752 2563 4764 2597
rect 4706 2537 4764 2563
rect 4806 2597 4864 2623
rect 4806 2563 4818 2597
rect 4852 2563 4864 2597
rect 4806 2537 4864 2563
rect 4906 2597 4964 2623
rect 4906 2563 4918 2597
rect 4952 2563 4964 2597
rect 4906 2537 4964 2563
rect 5006 2597 5064 2623
rect 5006 2563 5018 2597
rect 5052 2563 5064 2597
rect 5006 2537 5064 2563
rect 5106 2597 5164 2623
rect 5106 2563 5118 2597
rect 5152 2563 5164 2597
rect 5106 2537 5164 2563
rect 5206 2597 5264 2623
rect 5206 2563 5218 2597
rect 5252 2563 5264 2597
rect 5206 2537 5264 2563
rect 5306 2597 5364 2623
rect 5306 2563 5318 2597
rect 5352 2563 5364 2597
rect 5306 2537 5364 2563
rect 5406 2597 5464 2623
rect 5406 2563 5418 2597
rect 5452 2563 5464 2597
rect 5406 2537 5464 2563
rect 5506 2597 5564 2623
rect 5506 2563 5512 2597
rect 5552 2563 5564 2597
rect 5506 2537 5564 2563
rect 5606 2597 5664 2623
rect 5606 2563 5618 2597
rect 5658 2563 5664 2597
rect 5606 2537 5664 2563
rect 5706 2597 5764 2623
rect 5706 2563 5718 2597
rect 5752 2563 5764 2597
rect 5706 2537 5764 2563
rect 5806 2597 5864 2623
rect 5806 2563 5818 2597
rect 5852 2563 5864 2597
rect 5806 2537 5864 2563
rect 5906 2597 5964 2623
rect 5906 2563 5918 2597
rect 5952 2563 5964 2597
rect 5906 2537 5964 2563
rect 6006 2597 6064 2623
rect 6006 2563 6018 2597
rect 6052 2563 6064 2597
rect 6006 2537 6064 2563
rect 6106 2597 6164 2623
rect 6106 2563 6118 2597
rect 6152 2563 6164 2597
rect 6106 2537 6164 2563
rect 6206 2597 6264 2623
rect 6206 2563 6218 2597
rect 6252 2563 6264 2597
rect 6206 2537 6264 2563
rect 6306 2597 6364 2623
rect 6306 2563 6318 2597
rect 6352 2563 6364 2597
rect 6306 2537 6364 2563
rect 6406 2597 6464 2623
rect 6618 2616 6862 2650
rect 6406 2563 6418 2597
rect 6452 2563 6464 2597
rect 6508 2578 6516 2612
rect 6558 2578 6574 2612
rect 6618 2597 6652 2616
rect 6406 2537 6464 2563
rect 6828 2597 6862 2616
rect 6618 2547 6652 2563
rect 6696 2548 6712 2582
rect 6754 2548 6762 2582
rect 6828 2547 6862 2563
rect 6928 2597 7062 2613
rect 6962 2563 7028 2597
rect 6928 2547 7062 2563
rect 7128 2597 7262 2613
rect 7162 2563 7228 2597
rect 7128 2547 7262 2563
rect 7328 2597 7462 2613
rect 7362 2563 7428 2597
rect 7328 2547 7462 2563
rect 8 2440 18 2474
rect 52 2440 118 2474
rect 152 2440 168 2474
rect 208 2456 218 2490
rect 252 2456 318 2490
rect 352 2456 368 2490
rect 408 2440 418 2474
rect 452 2440 518 2474
rect 552 2440 568 2474
rect 608 2456 618 2490
rect 652 2456 718 2490
rect 752 2456 768 2490
rect 808 2440 818 2474
rect 852 2440 918 2474
rect 952 2440 968 2474
rect 1008 2456 1018 2490
rect 1052 2456 1118 2490
rect 1152 2456 1168 2490
rect 1208 2440 1218 2474
rect 1252 2440 1318 2474
rect 1352 2440 1368 2474
rect 1408 2456 1418 2490
rect 1452 2456 1518 2490
rect 1552 2456 1568 2490
rect 1608 2440 1618 2474
rect 1652 2440 1718 2474
rect 1752 2440 1768 2474
rect 1808 2456 1818 2490
rect 1852 2456 1918 2490
rect 1952 2456 1968 2490
rect 2008 2440 2018 2474
rect 2052 2440 2118 2474
rect 2152 2440 2168 2474
rect 2208 2456 2218 2490
rect 2252 2456 2318 2490
rect 2352 2456 2368 2490
rect 2408 2440 2418 2474
rect 2452 2440 2518 2474
rect 2552 2440 2568 2474
rect 2608 2456 2618 2490
rect 2652 2456 2718 2490
rect 2752 2456 2768 2490
rect 2808 2440 2818 2474
rect 2852 2440 2918 2474
rect 2952 2440 2968 2474
rect 3008 2456 3018 2490
rect 3052 2456 3118 2490
rect 3152 2456 3168 2490
rect 3208 2440 3218 2474
rect 3252 2440 3318 2474
rect 3352 2440 3368 2474
rect 3408 2456 3418 2490
rect 3452 2456 3518 2490
rect 3552 2456 3568 2490
rect 3608 2440 3618 2474
rect 3652 2440 3718 2474
rect 3752 2440 3768 2474
rect 3808 2456 3818 2490
rect 3852 2456 3918 2490
rect 3952 2456 3968 2490
rect 4008 2440 4018 2474
rect 4052 2440 4118 2474
rect 4152 2440 4168 2474
rect 4208 2456 4218 2490
rect 4252 2456 4318 2490
rect 4352 2456 4368 2490
rect 4408 2440 4418 2474
rect 4452 2440 4518 2474
rect 4552 2440 4568 2474
rect 4608 2456 4618 2490
rect 4652 2456 4718 2490
rect 4752 2456 4768 2490
rect 4808 2440 4818 2474
rect 4852 2440 4918 2474
rect 4952 2440 4968 2474
rect 5008 2456 5018 2490
rect 5052 2456 5118 2490
rect 5152 2456 5168 2490
rect 5208 2440 5218 2474
rect 5252 2440 5318 2474
rect 5352 2440 5368 2474
rect 5408 2456 5418 2490
rect 5452 2456 5518 2490
rect 5552 2456 5568 2490
rect 5608 2440 5618 2474
rect 5652 2440 5718 2474
rect 5752 2440 5768 2474
rect 5808 2456 5818 2490
rect 5852 2456 5918 2490
rect 5952 2456 5968 2490
rect 6008 2440 6018 2474
rect 6052 2440 6118 2474
rect 6152 2440 6168 2474
rect 6208 2456 6218 2490
rect 6252 2456 6318 2490
rect 6352 2456 6368 2490
rect 6516 2471 6568 2488
rect 6550 2454 6568 2471
rect 6602 2454 6618 2488
rect 6652 2454 6668 2488
rect 6702 2459 6720 2488
rect 6702 2454 6754 2459
rect 6862 2454 6878 2488
rect 6912 2454 6928 2488
rect 6962 2454 6978 2488
rect 7012 2454 7028 2488
rect 7062 2454 7078 2488
rect 7112 2454 7128 2488
rect 7162 2454 7178 2488
rect 7212 2454 7228 2488
rect 7262 2454 7278 2488
rect 7312 2454 7328 2488
rect 7362 2454 7378 2488
rect 7412 2454 7428 2488
rect 6 2367 64 2393
rect 6 2333 18 2367
rect 52 2333 64 2367
rect 6 2307 64 2333
rect 106 2367 164 2393
rect 106 2333 118 2367
rect 152 2333 164 2367
rect 106 2307 164 2333
rect 206 2367 264 2393
rect 206 2333 218 2367
rect 252 2333 264 2367
rect 206 2307 264 2333
rect 306 2367 364 2393
rect 306 2333 318 2367
rect 352 2333 364 2367
rect 306 2307 364 2333
rect 406 2367 464 2393
rect 406 2333 418 2367
rect 452 2333 464 2367
rect 406 2307 464 2333
rect 506 2367 564 2393
rect 506 2333 518 2367
rect 552 2333 564 2367
rect 506 2307 564 2333
rect 606 2367 664 2393
rect 606 2333 618 2367
rect 652 2333 664 2367
rect 606 2307 664 2333
rect 706 2367 764 2393
rect 706 2333 718 2367
rect 752 2333 764 2367
rect 706 2307 764 2333
rect 806 2367 864 2393
rect 806 2333 818 2367
rect 852 2333 864 2367
rect 806 2307 864 2333
rect 906 2367 964 2393
rect 906 2333 918 2367
rect 952 2333 964 2367
rect 906 2307 964 2333
rect 1006 2367 1064 2393
rect 1006 2333 1018 2367
rect 1052 2333 1064 2367
rect 1006 2307 1064 2333
rect 1106 2367 1164 2393
rect 1106 2333 1118 2367
rect 1152 2333 1164 2367
rect 1106 2307 1164 2333
rect 1206 2367 1264 2393
rect 1206 2333 1218 2367
rect 1252 2333 1264 2367
rect 1206 2307 1264 2333
rect 1306 2367 1364 2393
rect 1306 2333 1318 2367
rect 1352 2333 1364 2367
rect 1306 2307 1364 2333
rect 1406 2367 1464 2393
rect 1406 2333 1418 2367
rect 1452 2333 1464 2367
rect 1406 2307 1464 2333
rect 1506 2367 1564 2393
rect 1506 2333 1518 2367
rect 1552 2333 1564 2367
rect 1506 2307 1564 2333
rect 1606 2367 1664 2393
rect 1606 2333 1618 2367
rect 1652 2333 1664 2367
rect 1606 2307 1664 2333
rect 1706 2367 1764 2393
rect 1706 2333 1718 2367
rect 1752 2333 1764 2367
rect 1706 2307 1764 2333
rect 1806 2367 1864 2393
rect 1806 2333 1818 2367
rect 1852 2333 1864 2367
rect 1806 2307 1864 2333
rect 1906 2367 1964 2393
rect 1906 2333 1918 2367
rect 1952 2333 1964 2367
rect 1906 2307 1964 2333
rect 2006 2367 2064 2393
rect 2006 2333 2018 2367
rect 2052 2333 2064 2367
rect 2006 2307 2064 2333
rect 2106 2367 2164 2393
rect 2106 2333 2118 2367
rect 2152 2333 2164 2367
rect 2106 2307 2164 2333
rect 2206 2367 2264 2393
rect 2206 2333 2218 2367
rect 2252 2333 2264 2367
rect 2206 2307 2264 2333
rect 2306 2367 2364 2393
rect 2306 2333 2318 2367
rect 2352 2333 2364 2367
rect 2306 2307 2364 2333
rect 2406 2367 2464 2393
rect 2406 2333 2418 2367
rect 2452 2333 2464 2367
rect 2406 2307 2464 2333
rect 2506 2367 2564 2393
rect 2506 2333 2518 2367
rect 2552 2333 2564 2367
rect 2506 2307 2564 2333
rect 2606 2367 2664 2393
rect 2606 2333 2618 2367
rect 2652 2333 2664 2367
rect 2606 2307 2664 2333
rect 2706 2367 2764 2393
rect 2706 2333 2718 2367
rect 2752 2333 2764 2367
rect 2706 2307 2764 2333
rect 2806 2367 2864 2393
rect 2806 2333 2818 2367
rect 2852 2333 2864 2367
rect 2806 2307 2864 2333
rect 2906 2367 2964 2393
rect 2906 2333 2918 2367
rect 2952 2333 2964 2367
rect 2906 2307 2964 2333
rect 3006 2367 3064 2393
rect 3006 2333 3018 2367
rect 3052 2333 3064 2367
rect 3006 2307 3064 2333
rect 3106 2367 3164 2393
rect 3106 2333 3118 2367
rect 3152 2333 3164 2367
rect 3106 2307 3164 2333
rect 3206 2367 3264 2393
rect 3206 2333 3218 2367
rect 3252 2333 3264 2367
rect 3206 2307 3264 2333
rect 3306 2367 3364 2393
rect 3306 2333 3318 2367
rect 3352 2333 3364 2367
rect 3306 2307 3364 2333
rect 3406 2367 3464 2393
rect 3406 2333 3418 2367
rect 3452 2333 3464 2367
rect 3406 2307 3464 2333
rect 3506 2367 3564 2393
rect 3506 2333 3518 2367
rect 3552 2333 3564 2367
rect 3506 2307 3564 2333
rect 3606 2367 3664 2393
rect 3606 2333 3618 2367
rect 3652 2333 3664 2367
rect 3606 2307 3664 2333
rect 3706 2367 3764 2393
rect 3706 2333 3718 2367
rect 3752 2333 3764 2367
rect 3706 2307 3764 2333
rect 3806 2367 3864 2393
rect 3806 2333 3818 2367
rect 3852 2333 3864 2367
rect 3806 2307 3864 2333
rect 3906 2367 3964 2393
rect 3906 2333 3918 2367
rect 3952 2333 3964 2367
rect 3906 2307 3964 2333
rect 4006 2367 4064 2393
rect 4006 2333 4018 2367
rect 4052 2333 4064 2367
rect 4006 2307 4064 2333
rect 4106 2367 4164 2393
rect 4106 2333 4118 2367
rect 4152 2333 4164 2367
rect 4106 2307 4164 2333
rect 4206 2367 4264 2393
rect 4206 2333 4218 2367
rect 4252 2333 4264 2367
rect 4206 2307 4264 2333
rect 4306 2367 4364 2393
rect 4306 2333 4318 2367
rect 4352 2333 4364 2367
rect 4306 2307 4364 2333
rect 4406 2367 4464 2393
rect 4406 2333 4418 2367
rect 4452 2333 4464 2367
rect 4406 2307 4464 2333
rect 4506 2367 4564 2393
rect 4506 2333 4518 2367
rect 4552 2333 4564 2367
rect 4506 2307 4564 2333
rect 4606 2367 4664 2393
rect 4606 2333 4618 2367
rect 4652 2333 4664 2367
rect 4606 2307 4664 2333
rect 4706 2367 4764 2393
rect 4706 2333 4718 2367
rect 4752 2333 4764 2367
rect 4706 2307 4764 2333
rect 4806 2367 4864 2393
rect 4806 2333 4818 2367
rect 4852 2333 4864 2367
rect 4806 2307 4864 2333
rect 4906 2367 4964 2393
rect 4906 2333 4918 2367
rect 4952 2333 4964 2367
rect 4906 2307 4964 2333
rect 5006 2367 5064 2393
rect 5006 2333 5018 2367
rect 5052 2333 5064 2367
rect 5006 2307 5064 2333
rect 5106 2367 5164 2393
rect 5106 2333 5118 2367
rect 5152 2333 5164 2367
rect 5106 2307 5164 2333
rect 5206 2367 5264 2393
rect 5206 2333 5218 2367
rect 5252 2333 5264 2367
rect 5206 2307 5264 2333
rect 5306 2367 5364 2393
rect 5306 2333 5318 2367
rect 5352 2333 5364 2367
rect 5306 2307 5364 2333
rect 5406 2367 5464 2393
rect 5406 2333 5412 2367
rect 5452 2333 5464 2367
rect 5406 2307 5464 2333
rect 5506 2367 5564 2393
rect 5506 2333 5518 2367
rect 5558 2333 5564 2367
rect 5506 2307 5564 2333
rect 5606 2367 5664 2393
rect 5606 2333 5618 2367
rect 5652 2333 5664 2367
rect 5606 2307 5664 2333
rect 5706 2367 5764 2393
rect 5706 2333 5718 2367
rect 5752 2333 5764 2367
rect 5706 2307 5764 2333
rect 5806 2367 5864 2393
rect 5806 2333 5818 2367
rect 5852 2333 5864 2367
rect 5806 2307 5864 2333
rect 5906 2367 5964 2393
rect 5906 2333 5918 2367
rect 5952 2333 5964 2367
rect 5906 2307 5964 2333
rect 6006 2367 6064 2393
rect 6006 2333 6018 2367
rect 6052 2333 6064 2367
rect 6006 2307 6064 2333
rect 6106 2367 6164 2393
rect 6106 2333 6118 2367
rect 6152 2333 6164 2367
rect 6106 2307 6164 2333
rect 6206 2367 6264 2393
rect 6206 2333 6218 2367
rect 6252 2333 6264 2367
rect 6206 2307 6264 2333
rect 6306 2367 6364 2393
rect 6306 2333 6318 2367
rect 6352 2333 6364 2367
rect 6306 2307 6364 2333
rect 6406 2367 6464 2393
rect 6618 2386 6862 2420
rect 6406 2333 6412 2367
rect 6452 2333 6464 2367
rect 6508 2348 6516 2382
rect 6558 2348 6574 2382
rect 6618 2367 6652 2386
rect 6406 2307 6464 2333
rect 6828 2383 6862 2386
rect 6828 2367 6962 2383
rect 6618 2317 6652 2333
rect 6696 2318 6712 2352
rect 6754 2318 6762 2352
rect 6862 2333 6928 2367
rect 6828 2317 6962 2333
rect 7028 2367 7162 2383
rect 7062 2333 7128 2367
rect 7028 2317 7162 2333
rect 7228 2367 7362 2383
rect 7262 2333 7328 2367
rect 7228 2317 7362 2333
rect 7428 2367 7462 2383
rect 7428 2317 7462 2333
rect 6 2227 64 2253
rect 6 2193 18 2227
rect 58 2193 64 2227
rect 6 2167 64 2193
rect 106 2227 164 2253
rect 106 2193 118 2227
rect 152 2193 164 2227
rect 106 2167 164 2193
rect 206 2227 264 2253
rect 206 2193 212 2227
rect 252 2193 264 2227
rect 206 2167 264 2193
rect 306 2227 364 2253
rect 306 2193 318 2227
rect 358 2193 364 2227
rect 306 2167 364 2193
rect 406 2227 464 2253
rect 406 2193 418 2227
rect 452 2193 464 2227
rect 406 2167 464 2193
rect 506 2227 564 2253
rect 506 2193 518 2227
rect 552 2193 564 2227
rect 506 2167 564 2193
rect 606 2227 664 2253
rect 606 2193 618 2227
rect 652 2193 664 2227
rect 606 2167 664 2193
rect 706 2227 764 2253
rect 706 2193 718 2227
rect 752 2193 764 2227
rect 706 2167 764 2193
rect 806 2227 864 2253
rect 806 2193 818 2227
rect 852 2193 864 2227
rect 806 2167 864 2193
rect 906 2227 964 2253
rect 906 2193 918 2227
rect 952 2193 964 2227
rect 906 2167 964 2193
rect 1006 2227 1064 2253
rect 1006 2193 1018 2227
rect 1052 2193 1064 2227
rect 1006 2167 1064 2193
rect 1106 2227 1164 2253
rect 1106 2193 1118 2227
rect 1152 2193 1164 2227
rect 1106 2167 1164 2193
rect 1206 2227 1264 2253
rect 1206 2193 1218 2227
rect 1252 2193 1264 2227
rect 1206 2167 1264 2193
rect 1306 2227 1364 2253
rect 1306 2193 1312 2227
rect 1352 2193 1364 2227
rect 1306 2167 1364 2193
rect 1406 2227 1464 2253
rect 1406 2193 1418 2227
rect 1458 2193 1464 2227
rect 1406 2167 1464 2193
rect 1506 2227 1564 2253
rect 1506 2193 1512 2227
rect 1552 2193 1564 2227
rect 1506 2167 1564 2193
rect 1606 2227 1664 2253
rect 1606 2193 1618 2227
rect 1658 2193 1664 2227
rect 1606 2167 1664 2193
rect 1706 2227 1764 2253
rect 1706 2193 1718 2227
rect 1752 2193 1764 2227
rect 1706 2167 1764 2193
rect 1806 2227 1864 2253
rect 1806 2193 1812 2227
rect 1852 2193 1864 2227
rect 1806 2167 1864 2193
rect 1906 2227 1964 2253
rect 1906 2193 1918 2227
rect 1958 2193 1964 2227
rect 1906 2167 1964 2193
rect 2006 2227 2064 2253
rect 2006 2193 2018 2227
rect 2052 2193 2064 2227
rect 2006 2167 2064 2193
rect 2106 2227 2164 2253
rect 2106 2193 2118 2227
rect 2152 2193 2164 2227
rect 2106 2167 2164 2193
rect 2206 2227 2264 2253
rect 2206 2193 2212 2227
rect 2252 2193 2264 2227
rect 2206 2167 2264 2193
rect 2306 2227 2364 2253
rect 2306 2193 2318 2227
rect 2358 2193 2364 2227
rect 2306 2167 2364 2193
rect 2406 2227 2464 2253
rect 2406 2193 2418 2227
rect 2452 2193 2464 2227
rect 2406 2167 2464 2193
rect 2506 2227 2564 2253
rect 2506 2193 2518 2227
rect 2552 2193 2564 2227
rect 2506 2167 2564 2193
rect 2606 2227 2664 2253
rect 2606 2193 2618 2227
rect 2652 2193 2664 2227
rect 2606 2167 2664 2193
rect 2706 2227 2764 2253
rect 2706 2193 2718 2227
rect 2752 2193 2764 2227
rect 2706 2167 2764 2193
rect 2806 2227 2864 2253
rect 2806 2193 2812 2227
rect 2852 2193 2864 2227
rect 2806 2167 2864 2193
rect 2906 2227 2964 2253
rect 2906 2193 2918 2227
rect 2958 2193 2964 2227
rect 2906 2167 2964 2193
rect 3006 2227 3064 2253
rect 3006 2193 3018 2227
rect 3052 2193 3064 2227
rect 3006 2167 3064 2193
rect 3106 2227 3164 2253
rect 3106 2193 3118 2227
rect 3152 2193 3164 2227
rect 3106 2167 3164 2193
rect 3206 2227 3264 2253
rect 3206 2193 3218 2227
rect 3252 2193 3264 2227
rect 3206 2167 3264 2193
rect 3306 2227 3364 2253
rect 3306 2193 3318 2227
rect 3352 2193 3364 2227
rect 3306 2167 3364 2193
rect 3406 2227 3464 2253
rect 3406 2193 3418 2227
rect 3452 2193 3464 2227
rect 3406 2167 3464 2193
rect 3506 2227 3564 2253
rect 3506 2193 3512 2227
rect 3552 2193 3564 2227
rect 3506 2167 3564 2193
rect 3606 2227 3664 2253
rect 3606 2193 3618 2227
rect 3658 2193 3664 2227
rect 3606 2167 3664 2193
rect 3706 2227 3764 2253
rect 3706 2193 3718 2227
rect 3752 2193 3764 2227
rect 3706 2167 3764 2193
rect 3806 2227 3864 2253
rect 3806 2193 3818 2227
rect 3852 2193 3864 2227
rect 3806 2167 3864 2193
rect 3906 2227 3964 2253
rect 3906 2193 3918 2227
rect 3952 2193 3964 2227
rect 3906 2167 3964 2193
rect 4006 2227 4064 2253
rect 4006 2193 4018 2227
rect 4052 2193 4064 2227
rect 4006 2167 4064 2193
rect 4106 2227 4164 2253
rect 4106 2193 4118 2227
rect 4152 2193 4164 2227
rect 4106 2167 4164 2193
rect 4206 2227 4264 2253
rect 4206 2193 4212 2227
rect 4252 2193 4264 2227
rect 4206 2167 4264 2193
rect 4306 2227 4364 2253
rect 4306 2193 4318 2227
rect 4358 2193 4364 2227
rect 4306 2167 4364 2193
rect 4406 2227 4464 2253
rect 4406 2193 4412 2227
rect 4452 2193 4464 2227
rect 4406 2167 4464 2193
rect 4506 2227 4564 2253
rect 4506 2193 4518 2227
rect 4558 2193 4564 2227
rect 4506 2167 4564 2193
rect 4606 2227 4664 2253
rect 4606 2193 4618 2227
rect 4652 2193 4664 2227
rect 4606 2167 4664 2193
rect 4706 2227 4764 2253
rect 4706 2193 4718 2227
rect 4752 2193 4764 2227
rect 4706 2167 4764 2193
rect 4806 2227 4864 2253
rect 4806 2193 4818 2227
rect 4852 2193 4864 2227
rect 4806 2167 4864 2193
rect 4906 2227 4964 2253
rect 4906 2193 4918 2227
rect 4952 2193 4964 2227
rect 4906 2167 4964 2193
rect 5006 2227 5064 2253
rect 5006 2193 5018 2227
rect 5052 2193 5064 2227
rect 5006 2167 5064 2193
rect 5106 2227 5164 2253
rect 5106 2193 5118 2227
rect 5152 2193 5164 2227
rect 5106 2167 5164 2193
rect 5206 2227 5264 2253
rect 5206 2193 5218 2227
rect 5252 2193 5264 2227
rect 5206 2167 5264 2193
rect 5306 2227 5364 2253
rect 5306 2193 5318 2227
rect 5352 2193 5364 2227
rect 5306 2167 5364 2193
rect 5406 2227 5464 2253
rect 5406 2193 5418 2227
rect 5452 2193 5464 2227
rect 5406 2167 5464 2193
rect 5506 2227 5564 2253
rect 5506 2193 5518 2227
rect 5552 2193 5564 2227
rect 5506 2167 5564 2193
rect 5606 2227 5664 2253
rect 5606 2193 5618 2227
rect 5652 2193 5664 2227
rect 5606 2167 5664 2193
rect 5706 2227 5764 2253
rect 5706 2193 5718 2227
rect 5752 2193 5764 2227
rect 5706 2167 5764 2193
rect 5806 2227 5864 2253
rect 5806 2193 5818 2227
rect 5852 2193 5864 2227
rect 5806 2167 5864 2193
rect 5906 2227 5964 2253
rect 5906 2193 5918 2227
rect 5952 2193 5964 2227
rect 5906 2167 5964 2193
rect 6006 2227 6064 2253
rect 6006 2193 6018 2227
rect 6052 2193 6064 2227
rect 6006 2167 6064 2193
rect 6106 2227 6164 2253
rect 6106 2193 6118 2227
rect 6152 2193 6164 2227
rect 6106 2167 6164 2193
rect 6206 2227 6264 2253
rect 6206 2193 6218 2227
rect 6252 2193 6264 2227
rect 6206 2167 6264 2193
rect 6306 2227 6364 2253
rect 6306 2193 6318 2227
rect 6352 2193 6364 2227
rect 6306 2167 6364 2193
rect 6406 2227 6464 2253
rect 6618 2246 6862 2280
rect 6406 2193 6412 2227
rect 6452 2193 6464 2227
rect 6508 2208 6516 2242
rect 6558 2208 6574 2242
rect 6618 2227 6652 2246
rect 6406 2167 6464 2193
rect 6828 2227 6862 2246
rect 6618 2177 6652 2193
rect 6696 2178 6712 2212
rect 6754 2178 6762 2212
rect 6828 2177 6862 2193
rect 6928 2227 7162 2243
rect 6962 2193 7028 2227
rect 7062 2193 7128 2227
rect 6928 2177 7162 2193
rect 7228 2227 7362 2243
rect 7262 2193 7328 2227
rect 7228 2177 7362 2193
rect 7428 2227 7462 2243
rect 7428 2177 7462 2193
rect 6 2087 64 2113
rect 6 2053 18 2087
rect 58 2053 64 2087
rect 6 2027 64 2053
rect 106 2087 164 2113
rect 106 2053 118 2087
rect 152 2053 164 2087
rect 106 2027 164 2053
rect 206 2087 264 2113
rect 206 2053 218 2087
rect 252 2053 264 2087
rect 206 2027 264 2053
rect 306 2087 364 2113
rect 306 2053 312 2087
rect 352 2053 364 2087
rect 306 2027 364 2053
rect 406 2087 464 2113
rect 406 2053 418 2087
rect 458 2053 464 2087
rect 406 2027 464 2053
rect 506 2087 564 2113
rect 506 2053 518 2087
rect 552 2053 564 2087
rect 506 2027 564 2053
rect 606 2087 664 2113
rect 606 2053 618 2087
rect 652 2053 664 2087
rect 606 2027 664 2053
rect 706 2087 764 2113
rect 706 2053 718 2087
rect 752 2053 764 2087
rect 706 2027 764 2053
rect 806 2087 864 2113
rect 806 2053 818 2087
rect 852 2053 864 2087
rect 806 2027 864 2053
rect 906 2087 964 2113
rect 906 2053 918 2087
rect 952 2053 964 2087
rect 906 2027 964 2053
rect 1006 2087 1064 2113
rect 1006 2053 1018 2087
rect 1052 2053 1064 2087
rect 1006 2027 1064 2053
rect 1106 2087 1164 2113
rect 1106 2053 1118 2087
rect 1152 2053 1164 2087
rect 1106 2027 1164 2053
rect 1206 2087 1264 2113
rect 1206 2053 1218 2087
rect 1252 2053 1264 2087
rect 1206 2027 1264 2053
rect 1306 2087 1364 2113
rect 1306 2053 1312 2087
rect 1352 2053 1364 2087
rect 1306 2027 1364 2053
rect 1406 2087 1464 2113
rect 1406 2053 1418 2087
rect 1458 2053 1464 2087
rect 1406 2027 1464 2053
rect 1506 2087 1564 2113
rect 1506 2053 1512 2087
rect 1552 2053 1564 2087
rect 1506 2027 1564 2053
rect 1606 2087 1664 2113
rect 1606 2053 1618 2087
rect 1658 2053 1664 2087
rect 1606 2027 1664 2053
rect 1706 2087 1764 2113
rect 1706 2053 1718 2087
rect 1752 2053 1764 2087
rect 1706 2027 1764 2053
rect 1806 2087 1864 2113
rect 1806 2053 1812 2087
rect 1852 2053 1864 2087
rect 1806 2027 1864 2053
rect 1906 2087 1964 2113
rect 1906 2053 1918 2087
rect 1958 2053 1964 2087
rect 1906 2027 1964 2053
rect 2006 2087 2064 2113
rect 2006 2053 2018 2087
rect 2052 2053 2064 2087
rect 2006 2027 2064 2053
rect 2106 2087 2164 2113
rect 2106 2053 2118 2087
rect 2152 2053 2164 2087
rect 2106 2027 2164 2053
rect 2206 2087 2264 2113
rect 2206 2053 2212 2087
rect 2252 2053 2264 2087
rect 2206 2027 2264 2053
rect 2306 2087 2364 2113
rect 2306 2053 2318 2087
rect 2358 2053 2364 2087
rect 2306 2027 2364 2053
rect 2406 2087 2464 2113
rect 2406 2053 2412 2087
rect 2452 2053 2464 2087
rect 2406 2027 2464 2053
rect 2506 2087 2564 2113
rect 2506 2053 2518 2087
rect 2558 2053 2564 2087
rect 2506 2027 2564 2053
rect 2606 2087 2664 2113
rect 2606 2053 2618 2087
rect 2652 2053 2664 2087
rect 2606 2027 2664 2053
rect 2706 2087 2764 2113
rect 2706 2053 2718 2087
rect 2752 2053 2764 2087
rect 2706 2027 2764 2053
rect 2806 2087 2864 2113
rect 2806 2053 2818 2087
rect 2852 2053 2864 2087
rect 2806 2027 2864 2053
rect 2906 2087 2964 2113
rect 2906 2053 2918 2087
rect 2952 2053 2964 2087
rect 2906 2027 2964 2053
rect 3006 2087 3064 2113
rect 3006 2053 3018 2087
rect 3052 2053 3064 2087
rect 3006 2027 3064 2053
rect 3106 2087 3164 2113
rect 3106 2053 3118 2087
rect 3152 2053 3164 2087
rect 3106 2027 3164 2053
rect 3206 2087 3264 2113
rect 3206 2053 3218 2087
rect 3252 2053 3264 2087
rect 3206 2027 3264 2053
rect 3306 2087 3364 2113
rect 3306 2053 3312 2087
rect 3352 2053 3364 2087
rect 3306 2027 3364 2053
rect 3406 2087 3464 2113
rect 3406 2053 3418 2087
rect 3458 2053 3464 2087
rect 3406 2027 3464 2053
rect 3506 2087 3564 2113
rect 3506 2053 3518 2087
rect 3552 2053 3564 2087
rect 3506 2027 3564 2053
rect 3606 2087 3664 2113
rect 3606 2053 3612 2087
rect 3652 2053 3664 2087
rect 3606 2027 3664 2053
rect 3706 2087 3764 2113
rect 3706 2053 3718 2087
rect 3758 2053 3764 2087
rect 3706 2027 3764 2053
rect 3806 2087 3864 2113
rect 3806 2053 3818 2087
rect 3852 2053 3864 2087
rect 3806 2027 3864 2053
rect 3906 2087 3964 2113
rect 3906 2053 3912 2087
rect 3952 2053 3964 2087
rect 3906 2027 3964 2053
rect 4006 2087 4064 2113
rect 4006 2053 4018 2087
rect 4058 2053 4064 2087
rect 4006 2027 4064 2053
rect 4106 2087 4164 2113
rect 4106 2053 4118 2087
rect 4152 2053 4164 2087
rect 4106 2027 4164 2053
rect 4206 2087 4264 2113
rect 4206 2053 4218 2087
rect 4252 2053 4264 2087
rect 4206 2027 4264 2053
rect 4306 2087 4364 2113
rect 4306 2053 4318 2087
rect 4352 2053 4364 2087
rect 4306 2027 4364 2053
rect 4406 2087 4464 2113
rect 4406 2053 4412 2087
rect 4452 2053 4464 2087
rect 4406 2027 4464 2053
rect 4506 2087 4564 2113
rect 4506 2053 4518 2087
rect 4558 2053 4564 2087
rect 4506 2027 4564 2053
rect 4606 2087 4664 2113
rect 4606 2053 4618 2087
rect 4652 2053 4664 2087
rect 4606 2027 4664 2053
rect 4706 2087 4764 2113
rect 4706 2053 4718 2087
rect 4752 2053 4764 2087
rect 4706 2027 4764 2053
rect 4806 2087 4864 2113
rect 4806 2053 4818 2087
rect 4852 2053 4864 2087
rect 4806 2027 4864 2053
rect 4906 2087 4964 2113
rect 4906 2053 4918 2087
rect 4952 2053 4964 2087
rect 4906 2027 4964 2053
rect 5006 2087 5064 2113
rect 5006 2053 5018 2087
rect 5052 2053 5064 2087
rect 5006 2027 5064 2053
rect 5106 2087 5164 2113
rect 5106 2053 5118 2087
rect 5152 2053 5164 2087
rect 5106 2027 5164 2053
rect 5206 2087 5264 2113
rect 5206 2053 5218 2087
rect 5252 2053 5264 2087
rect 5206 2027 5264 2053
rect 5306 2087 5364 2113
rect 5306 2053 5318 2087
rect 5352 2053 5364 2087
rect 5306 2027 5364 2053
rect 5406 2087 5464 2113
rect 5406 2053 5418 2087
rect 5452 2053 5464 2087
rect 5406 2027 5464 2053
rect 5506 2087 5564 2113
rect 5506 2053 5518 2087
rect 5552 2053 5564 2087
rect 5506 2027 5564 2053
rect 5606 2087 5664 2113
rect 5606 2053 5618 2087
rect 5652 2053 5664 2087
rect 5606 2027 5664 2053
rect 5706 2087 5764 2113
rect 5706 2053 5718 2087
rect 5752 2053 5764 2087
rect 5706 2027 5764 2053
rect 5806 2087 5864 2113
rect 5806 2053 5818 2087
rect 5852 2053 5864 2087
rect 5806 2027 5864 2053
rect 5906 2087 5964 2113
rect 5906 2053 5918 2087
rect 5952 2053 5964 2087
rect 5906 2027 5964 2053
rect 6006 2087 6064 2113
rect 6006 2053 6018 2087
rect 6052 2053 6064 2087
rect 6006 2027 6064 2053
rect 6106 2087 6164 2113
rect 6106 2053 6118 2087
rect 6152 2053 6164 2087
rect 6106 2027 6164 2053
rect 6206 2087 6264 2113
rect 6206 2053 6218 2087
rect 6252 2053 6264 2087
rect 6206 2027 6264 2053
rect 6306 2087 6364 2113
rect 6306 2053 6318 2087
rect 6352 2053 6364 2087
rect 6306 2027 6364 2053
rect 6406 2087 6464 2113
rect 6618 2106 6862 2140
rect 6406 2053 6418 2087
rect 6452 2053 6464 2087
rect 6508 2068 6516 2102
rect 6558 2068 6574 2102
rect 6618 2087 6652 2106
rect 6406 2027 6464 2053
rect 6828 2103 6862 2106
rect 6828 2087 6962 2103
rect 6618 2037 6652 2053
rect 6696 2038 6712 2072
rect 6754 2038 6762 2072
rect 6862 2053 6928 2087
rect 6828 2037 6962 2053
rect 7028 2087 7062 2103
rect 7028 2037 7062 2053
rect 7128 2087 7362 2103
rect 7162 2053 7228 2087
rect 7262 2053 7328 2087
rect 7128 2037 7362 2053
rect 7428 2087 7462 2103
rect 7428 2037 7462 2053
rect 6 1947 64 1973
rect 6 1913 18 1947
rect 52 1913 64 1947
rect 6 1887 64 1913
rect 106 1947 164 1973
rect 106 1913 118 1947
rect 152 1913 164 1947
rect 106 1887 164 1913
rect 206 1947 264 1973
rect 206 1913 218 1947
rect 252 1913 264 1947
rect 206 1887 264 1913
rect 306 1947 364 1973
rect 306 1913 312 1947
rect 352 1913 364 1947
rect 306 1887 364 1913
rect 406 1947 464 1973
rect 406 1913 418 1947
rect 458 1913 464 1947
rect 406 1887 464 1913
rect 506 1947 564 1973
rect 506 1913 518 1947
rect 552 1913 564 1947
rect 506 1887 564 1913
rect 606 1947 664 1973
rect 606 1913 618 1947
rect 652 1913 664 1947
rect 606 1887 664 1913
rect 706 1947 764 1973
rect 706 1913 718 1947
rect 752 1913 764 1947
rect 706 1887 764 1913
rect 806 1947 864 1973
rect 806 1913 818 1947
rect 852 1913 864 1947
rect 806 1887 864 1913
rect 906 1947 964 1973
rect 906 1913 918 1947
rect 952 1913 964 1947
rect 906 1887 964 1913
rect 1006 1947 1064 1973
rect 1006 1913 1018 1947
rect 1052 1913 1064 1947
rect 1006 1887 1064 1913
rect 1106 1947 1164 1973
rect 1106 1913 1118 1947
rect 1152 1913 1164 1947
rect 1106 1887 1164 1913
rect 1206 1947 1264 1973
rect 1206 1913 1218 1947
rect 1252 1913 1264 1947
rect 1206 1887 1264 1913
rect 1306 1947 1364 1973
rect 1306 1913 1318 1947
rect 1352 1913 1364 1947
rect 1306 1887 1364 1913
rect 1406 1947 1464 1973
rect 1406 1913 1412 1947
rect 1452 1913 1464 1947
rect 1406 1887 1464 1913
rect 1506 1947 1564 1973
rect 1506 1913 1518 1947
rect 1558 1913 1564 1947
rect 1506 1887 1564 1913
rect 1606 1947 1664 1973
rect 1606 1913 1618 1947
rect 1652 1913 1664 1947
rect 1606 1887 1664 1913
rect 1706 1947 1764 1973
rect 1706 1913 1718 1947
rect 1752 1913 1764 1947
rect 1706 1887 1764 1913
rect 1806 1947 1864 1973
rect 1806 1913 1818 1947
rect 1852 1913 1864 1947
rect 1806 1887 1864 1913
rect 1906 1947 1964 1973
rect 1906 1913 1918 1947
rect 1952 1913 1964 1947
rect 1906 1887 1964 1913
rect 2006 1947 2064 1973
rect 2006 1913 2018 1947
rect 2052 1913 2064 1947
rect 2006 1887 2064 1913
rect 2106 1947 2164 1973
rect 2106 1913 2118 1947
rect 2152 1913 2164 1947
rect 2106 1887 2164 1913
rect 2206 1947 2264 1973
rect 2206 1913 2218 1947
rect 2252 1913 2264 1947
rect 2206 1887 2264 1913
rect 2306 1947 2364 1973
rect 2306 1913 2318 1947
rect 2352 1913 2364 1947
rect 2306 1887 2364 1913
rect 2406 1947 2464 1973
rect 2406 1913 2412 1947
rect 2452 1913 2464 1947
rect 2406 1887 2464 1913
rect 2506 1947 2564 1973
rect 2506 1913 2518 1947
rect 2558 1913 2564 1947
rect 2506 1887 2564 1913
rect 2606 1947 2664 1973
rect 2606 1913 2618 1947
rect 2652 1913 2664 1947
rect 2606 1887 2664 1913
rect 2706 1947 2764 1973
rect 2706 1913 2718 1947
rect 2752 1913 2764 1947
rect 2706 1887 2764 1913
rect 2806 1947 2864 1973
rect 2806 1913 2818 1947
rect 2852 1913 2864 1947
rect 2806 1887 2864 1913
rect 2906 1947 2964 1973
rect 2906 1913 2918 1947
rect 2952 1913 2964 1947
rect 2906 1887 2964 1913
rect 3006 1947 3064 1973
rect 3006 1913 3012 1947
rect 3052 1913 3064 1947
rect 3006 1887 3064 1913
rect 3106 1947 3164 1973
rect 3106 1913 3118 1947
rect 3158 1913 3164 1947
rect 3106 1887 3164 1913
rect 3206 1947 3264 1973
rect 3206 1913 3218 1947
rect 3252 1913 3264 1947
rect 3206 1887 3264 1913
rect 3306 1947 3364 1973
rect 3306 1913 3318 1947
rect 3352 1913 3364 1947
rect 3306 1887 3364 1913
rect 3406 1947 3464 1973
rect 3406 1913 3418 1947
rect 3452 1913 3464 1947
rect 3406 1887 3464 1913
rect 3506 1947 3564 1973
rect 3506 1913 3518 1947
rect 3552 1913 3564 1947
rect 3506 1887 3564 1913
rect 3606 1947 3664 1973
rect 3606 1913 3618 1947
rect 3652 1913 3664 1947
rect 3606 1887 3664 1913
rect 3706 1947 3764 1973
rect 3706 1913 3718 1947
rect 3752 1913 3764 1947
rect 3706 1887 3764 1913
rect 3806 1947 3864 1973
rect 3806 1913 3812 1947
rect 3852 1913 3864 1947
rect 3806 1887 3864 1913
rect 3906 1947 3964 1973
rect 3906 1913 3918 1947
rect 3958 1913 3964 1947
rect 3906 1887 3964 1913
rect 4006 1947 4064 1973
rect 4006 1913 4018 1947
rect 4052 1913 4064 1947
rect 4006 1887 4064 1913
rect 4106 1947 4164 1973
rect 4106 1913 4118 1947
rect 4152 1913 4164 1947
rect 4106 1887 4164 1913
rect 4206 1947 4264 1973
rect 4206 1913 4218 1947
rect 4252 1913 4264 1947
rect 4206 1887 4264 1913
rect 4306 1947 4364 1973
rect 4306 1913 4318 1947
rect 4352 1913 4364 1947
rect 4306 1887 4364 1913
rect 4406 1947 4464 1973
rect 4406 1913 4412 1947
rect 4452 1913 4464 1947
rect 4406 1887 4464 1913
rect 4506 1947 4564 1973
rect 4506 1913 4518 1947
rect 4558 1913 4564 1947
rect 4506 1887 4564 1913
rect 4606 1947 4664 1973
rect 4606 1913 4618 1947
rect 4652 1913 4664 1947
rect 4606 1887 4664 1913
rect 4706 1947 4764 1973
rect 4706 1913 4718 1947
rect 4752 1913 4764 1947
rect 4706 1887 4764 1913
rect 4806 1947 4864 1973
rect 4806 1913 4818 1947
rect 4852 1913 4864 1947
rect 4806 1887 4864 1913
rect 4906 1947 4964 1973
rect 4906 1913 4912 1947
rect 4952 1913 4964 1947
rect 4906 1887 4964 1913
rect 5006 1947 5064 1973
rect 5006 1913 5018 1947
rect 5058 1913 5064 1947
rect 5006 1887 5064 1913
rect 5106 1947 5164 1973
rect 5106 1913 5112 1947
rect 5152 1913 5164 1947
rect 5106 1887 5164 1913
rect 5206 1947 5264 1973
rect 5206 1913 5218 1947
rect 5258 1913 5264 1947
rect 5206 1887 5264 1913
rect 5306 1947 5364 1973
rect 5306 1913 5312 1947
rect 5352 1913 5364 1947
rect 5306 1887 5364 1913
rect 5406 1947 5464 1973
rect 5406 1913 5418 1947
rect 5458 1913 5464 1947
rect 5406 1887 5464 1913
rect 5506 1947 5564 1973
rect 5506 1913 5518 1947
rect 5552 1913 5564 1947
rect 5506 1887 5564 1913
rect 5606 1947 5664 1973
rect 5606 1913 5618 1947
rect 5652 1913 5664 1947
rect 5606 1887 5664 1913
rect 5706 1947 5764 1973
rect 5706 1913 5712 1947
rect 5752 1913 5764 1947
rect 5706 1887 5764 1913
rect 5806 1947 5864 1973
rect 5806 1913 5818 1947
rect 5858 1913 5864 1947
rect 5806 1887 5864 1913
rect 5906 1947 5964 1973
rect 5906 1913 5918 1947
rect 5952 1913 5964 1947
rect 5906 1887 5964 1913
rect 6006 1947 6064 1973
rect 6006 1913 6012 1947
rect 6052 1913 6064 1947
rect 6006 1887 6064 1913
rect 6106 1947 6164 1973
rect 6106 1913 6118 1947
rect 6158 1913 6164 1947
rect 6106 1887 6164 1913
rect 6206 1947 6264 1973
rect 6206 1913 6218 1947
rect 6252 1913 6264 1947
rect 6206 1887 6264 1913
rect 6306 1947 6364 1973
rect 6306 1913 6318 1947
rect 6352 1913 6364 1947
rect 6306 1887 6364 1913
rect 6406 1947 6464 1973
rect 6618 1966 6862 2000
rect 6406 1913 6418 1947
rect 6452 1913 6464 1947
rect 6508 1928 6516 1962
rect 6558 1928 6574 1962
rect 6618 1947 6652 1966
rect 6406 1887 6464 1913
rect 6828 1947 6862 1966
rect 6618 1897 6652 1913
rect 6696 1898 6712 1932
rect 6754 1898 6762 1932
rect 6828 1897 6862 1913
rect 6928 1947 7062 1963
rect 6962 1913 7028 1947
rect 6928 1897 7062 1913
rect 7128 1947 7362 1963
rect 7162 1913 7228 1947
rect 7262 1913 7328 1947
rect 7128 1897 7362 1913
rect 7428 1947 7462 1963
rect 7428 1897 7462 1913
rect 6 1807 64 1833
rect 6 1773 18 1807
rect 52 1773 64 1807
rect 6 1747 64 1773
rect 106 1807 164 1833
rect 106 1773 118 1807
rect 152 1773 164 1807
rect 106 1747 164 1773
rect 206 1807 264 1833
rect 206 1773 218 1807
rect 252 1773 264 1807
rect 206 1747 264 1773
rect 306 1807 364 1833
rect 306 1773 318 1807
rect 352 1773 364 1807
rect 306 1747 364 1773
rect 406 1807 464 1833
rect 406 1773 418 1807
rect 452 1773 464 1807
rect 406 1747 464 1773
rect 506 1807 564 1833
rect 506 1773 518 1807
rect 552 1773 564 1807
rect 506 1747 564 1773
rect 606 1807 664 1833
rect 606 1773 618 1807
rect 652 1773 664 1807
rect 606 1747 664 1773
rect 706 1807 764 1833
rect 706 1773 718 1807
rect 752 1773 764 1807
rect 706 1747 764 1773
rect 806 1807 864 1833
rect 806 1773 818 1807
rect 852 1773 864 1807
rect 806 1747 864 1773
rect 906 1807 964 1833
rect 906 1773 912 1807
rect 952 1773 964 1807
rect 906 1747 964 1773
rect 1006 1807 1064 1833
rect 1006 1773 1018 1807
rect 1058 1773 1064 1807
rect 1006 1747 1064 1773
rect 1106 1807 1164 1833
rect 1106 1773 1118 1807
rect 1152 1773 1164 1807
rect 1106 1747 1164 1773
rect 1206 1807 1264 1833
rect 1206 1773 1218 1807
rect 1252 1773 1264 1807
rect 1206 1747 1264 1773
rect 1306 1807 1364 1833
rect 1306 1773 1318 1807
rect 1352 1773 1364 1807
rect 1306 1747 1364 1773
rect 1406 1807 1464 1833
rect 1406 1773 1418 1807
rect 1452 1773 1464 1807
rect 1406 1747 1464 1773
rect 1506 1807 1564 1833
rect 1506 1773 1518 1807
rect 1552 1773 1564 1807
rect 1506 1747 1564 1773
rect 1606 1807 1664 1833
rect 1606 1773 1618 1807
rect 1652 1773 1664 1807
rect 1606 1747 1664 1773
rect 1706 1807 1764 1833
rect 1706 1773 1718 1807
rect 1752 1773 1764 1807
rect 1706 1747 1764 1773
rect 1806 1807 1864 1833
rect 1806 1773 1812 1807
rect 1852 1773 1864 1807
rect 1806 1747 1864 1773
rect 1906 1807 1964 1833
rect 1906 1773 1918 1807
rect 1958 1773 1964 1807
rect 1906 1747 1964 1773
rect 2006 1807 2064 1833
rect 2006 1773 2018 1807
rect 2052 1773 2064 1807
rect 2006 1747 2064 1773
rect 2106 1807 2164 1833
rect 2106 1773 2118 1807
rect 2152 1773 2164 1807
rect 2106 1747 2164 1773
rect 2206 1807 2264 1833
rect 2206 1773 2218 1807
rect 2252 1773 2264 1807
rect 2206 1747 2264 1773
rect 2306 1807 2364 1833
rect 2306 1773 2318 1807
rect 2352 1773 2364 1807
rect 2306 1747 2364 1773
rect 2406 1807 2464 1833
rect 2406 1773 2418 1807
rect 2452 1773 2464 1807
rect 2406 1747 2464 1773
rect 2506 1807 2564 1833
rect 2506 1773 2518 1807
rect 2552 1773 2564 1807
rect 2506 1747 2564 1773
rect 2606 1807 2664 1833
rect 2606 1773 2618 1807
rect 2652 1773 2664 1807
rect 2606 1747 2664 1773
rect 2706 1807 2764 1833
rect 2706 1773 2718 1807
rect 2752 1773 2764 1807
rect 2706 1747 2764 1773
rect 2806 1807 2864 1833
rect 2806 1773 2818 1807
rect 2852 1773 2864 1807
rect 2806 1747 2864 1773
rect 2906 1807 2964 1833
rect 2906 1773 2918 1807
rect 2952 1773 2964 1807
rect 2906 1747 2964 1773
rect 3006 1807 3064 1833
rect 3006 1773 3018 1807
rect 3052 1773 3064 1807
rect 3006 1747 3064 1773
rect 3106 1807 3164 1833
rect 3106 1773 3118 1807
rect 3152 1773 3164 1807
rect 3106 1747 3164 1773
rect 3206 1807 3264 1833
rect 3206 1773 3218 1807
rect 3252 1773 3264 1807
rect 3206 1747 3264 1773
rect 3306 1807 3364 1833
rect 3306 1773 3318 1807
rect 3352 1773 3364 1807
rect 3306 1747 3364 1773
rect 3406 1807 3464 1833
rect 3406 1773 3412 1807
rect 3452 1773 3464 1807
rect 3406 1747 3464 1773
rect 3506 1807 3564 1833
rect 3506 1773 3518 1807
rect 3558 1773 3564 1807
rect 3506 1747 3564 1773
rect 3606 1807 3664 1833
rect 3606 1773 3612 1807
rect 3652 1773 3664 1807
rect 3606 1747 3664 1773
rect 3706 1807 3764 1833
rect 3706 1773 3718 1807
rect 3758 1773 3764 1807
rect 3706 1747 3764 1773
rect 3806 1807 3864 1833
rect 3806 1773 3818 1807
rect 3852 1773 3864 1807
rect 3806 1747 3864 1773
rect 3906 1807 3964 1833
rect 3906 1773 3912 1807
rect 3952 1773 3964 1807
rect 3906 1747 3964 1773
rect 4006 1807 4064 1833
rect 4006 1773 4018 1807
rect 4058 1773 4064 1807
rect 4006 1747 4064 1773
rect 4106 1807 4164 1833
rect 4106 1773 4118 1807
rect 4152 1773 4164 1807
rect 4106 1747 4164 1773
rect 4206 1807 4264 1833
rect 4206 1773 4218 1807
rect 4252 1773 4264 1807
rect 4206 1747 4264 1773
rect 4306 1807 4364 1833
rect 4306 1773 4318 1807
rect 4352 1773 4364 1807
rect 4306 1747 4364 1773
rect 4406 1807 4464 1833
rect 4406 1773 4418 1807
rect 4452 1773 4464 1807
rect 4406 1747 4464 1773
rect 4506 1807 4564 1833
rect 4506 1773 4518 1807
rect 4552 1773 4564 1807
rect 4506 1747 4564 1773
rect 4606 1807 4664 1833
rect 4606 1773 4618 1807
rect 4652 1773 4664 1807
rect 4606 1747 4664 1773
rect 4706 1807 4764 1833
rect 4706 1773 4718 1807
rect 4752 1773 4764 1807
rect 4706 1747 4764 1773
rect 4806 1807 4864 1833
rect 4806 1773 4812 1807
rect 4852 1773 4864 1807
rect 4806 1747 4864 1773
rect 4906 1807 4964 1833
rect 4906 1773 4918 1807
rect 4958 1773 4964 1807
rect 4906 1747 4964 1773
rect 5006 1807 5064 1833
rect 5006 1773 5018 1807
rect 5052 1773 5064 1807
rect 5006 1747 5064 1773
rect 5106 1807 5164 1833
rect 5106 1773 5118 1807
rect 5152 1773 5164 1807
rect 5106 1747 5164 1773
rect 5206 1807 5264 1833
rect 5206 1773 5218 1807
rect 5252 1773 5264 1807
rect 5206 1747 5264 1773
rect 5306 1807 5364 1833
rect 5306 1773 5318 1807
rect 5352 1773 5364 1807
rect 5306 1747 5364 1773
rect 5406 1807 5464 1833
rect 5406 1773 5418 1807
rect 5452 1773 5464 1807
rect 5406 1747 5464 1773
rect 5506 1807 5564 1833
rect 5506 1773 5518 1807
rect 5552 1773 5564 1807
rect 5506 1747 5564 1773
rect 5606 1807 5664 1833
rect 5606 1773 5618 1807
rect 5652 1773 5664 1807
rect 5606 1747 5664 1773
rect 5706 1807 5764 1833
rect 5706 1773 5718 1807
rect 5752 1773 5764 1807
rect 5706 1747 5764 1773
rect 5806 1807 5864 1833
rect 5806 1773 5818 1807
rect 5852 1773 5864 1807
rect 5806 1747 5864 1773
rect 5906 1807 5964 1833
rect 5906 1773 5918 1807
rect 5952 1773 5964 1807
rect 5906 1747 5964 1773
rect 6006 1807 6064 1833
rect 6006 1773 6018 1807
rect 6052 1773 6064 1807
rect 6006 1747 6064 1773
rect 6106 1807 6164 1833
rect 6106 1773 6118 1807
rect 6152 1773 6164 1807
rect 6106 1747 6164 1773
rect 6206 1807 6264 1833
rect 6206 1773 6218 1807
rect 6252 1773 6264 1807
rect 6206 1747 6264 1773
rect 6306 1807 6364 1833
rect 6306 1773 6318 1807
rect 6352 1773 6364 1807
rect 6306 1747 6364 1773
rect 6406 1807 6464 1833
rect 6618 1826 6862 1860
rect 6406 1773 6418 1807
rect 6452 1773 6464 1807
rect 6508 1788 6516 1822
rect 6558 1788 6574 1822
rect 6618 1807 6652 1826
rect 6406 1747 6464 1773
rect 6828 1823 6862 1826
rect 6828 1807 6962 1823
rect 6618 1757 6652 1773
rect 6696 1758 6712 1792
rect 6754 1758 6762 1792
rect 6862 1773 6928 1807
rect 6828 1757 6962 1773
rect 7028 1807 7162 1823
rect 7062 1773 7128 1807
rect 7028 1757 7162 1773
rect 7228 1807 7262 1823
rect 7228 1757 7262 1773
rect 7328 1807 7462 1823
rect 7362 1773 7428 1807
rect 7328 1757 7462 1773
rect 6 1667 64 1693
rect 6 1633 18 1667
rect 58 1633 64 1667
rect 6 1607 64 1633
rect 106 1667 164 1693
rect 106 1633 112 1667
rect 152 1633 164 1667
rect 106 1607 164 1633
rect 206 1667 264 1693
rect 206 1633 218 1667
rect 258 1633 264 1667
rect 206 1607 264 1633
rect 306 1667 364 1693
rect 306 1633 318 1667
rect 352 1633 364 1667
rect 306 1607 364 1633
rect 406 1667 464 1693
rect 406 1633 418 1667
rect 452 1633 464 1667
rect 406 1607 464 1633
rect 506 1667 564 1693
rect 506 1633 518 1667
rect 552 1633 564 1667
rect 506 1607 564 1633
rect 606 1667 664 1693
rect 606 1633 618 1667
rect 652 1633 664 1667
rect 606 1607 664 1633
rect 706 1667 764 1693
rect 706 1633 712 1667
rect 752 1633 764 1667
rect 706 1607 764 1633
rect 806 1667 864 1693
rect 806 1633 818 1667
rect 858 1633 864 1667
rect 806 1607 864 1633
rect 906 1667 964 1693
rect 906 1633 912 1667
rect 952 1633 964 1667
rect 906 1607 964 1633
rect 1006 1667 1064 1693
rect 1006 1633 1018 1667
rect 1058 1633 1064 1667
rect 1006 1607 1064 1633
rect 1106 1667 1164 1693
rect 1106 1633 1118 1667
rect 1152 1633 1164 1667
rect 1106 1607 1164 1633
rect 1206 1667 1264 1693
rect 1206 1633 1218 1667
rect 1252 1633 1264 1667
rect 1206 1607 1264 1633
rect 1306 1667 1364 1693
rect 1306 1633 1318 1667
rect 1352 1633 1364 1667
rect 1306 1607 1364 1633
rect 1406 1667 1464 1693
rect 1406 1633 1418 1667
rect 1452 1633 1464 1667
rect 1406 1607 1464 1633
rect 1506 1667 1564 1693
rect 1506 1633 1512 1667
rect 1552 1633 1564 1667
rect 1506 1607 1564 1633
rect 1606 1667 1664 1693
rect 1606 1633 1618 1667
rect 1658 1633 1664 1667
rect 1606 1607 1664 1633
rect 1706 1667 1764 1693
rect 1706 1633 1712 1667
rect 1752 1633 1764 1667
rect 1706 1607 1764 1633
rect 1806 1667 1864 1693
rect 1806 1633 1818 1667
rect 1858 1633 1864 1667
rect 1806 1607 1864 1633
rect 1906 1667 1964 1693
rect 1906 1633 1912 1667
rect 1952 1633 1964 1667
rect 1906 1607 1964 1633
rect 2006 1667 2064 1693
rect 2006 1633 2018 1667
rect 2058 1633 2064 1667
rect 2006 1607 2064 1633
rect 2106 1667 2164 1693
rect 2106 1633 2118 1667
rect 2152 1633 2164 1667
rect 2106 1607 2164 1633
rect 2206 1667 2264 1693
rect 2206 1633 2218 1667
rect 2252 1633 2264 1667
rect 2206 1607 2264 1633
rect 2306 1667 2364 1693
rect 2306 1633 2318 1667
rect 2352 1633 2364 1667
rect 2306 1607 2364 1633
rect 2406 1667 2464 1693
rect 2406 1633 2418 1667
rect 2452 1633 2464 1667
rect 2406 1607 2464 1633
rect 2506 1667 2564 1693
rect 2506 1633 2518 1667
rect 2552 1633 2564 1667
rect 2506 1607 2564 1633
rect 2606 1667 2664 1693
rect 2606 1633 2612 1667
rect 2652 1633 2664 1667
rect 2606 1607 2664 1633
rect 2706 1667 2764 1693
rect 2706 1633 2718 1667
rect 2758 1633 2764 1667
rect 2706 1607 2764 1633
rect 2806 1667 2864 1693
rect 2806 1633 2818 1667
rect 2852 1633 2864 1667
rect 2806 1607 2864 1633
rect 2906 1667 2964 1693
rect 2906 1633 2918 1667
rect 2952 1633 2964 1667
rect 2906 1607 2964 1633
rect 3006 1667 3064 1693
rect 3006 1633 3018 1667
rect 3052 1633 3064 1667
rect 3006 1607 3064 1633
rect 3106 1667 3164 1693
rect 3106 1633 3118 1667
rect 3152 1633 3164 1667
rect 3106 1607 3164 1633
rect 3206 1667 3264 1693
rect 3206 1633 3218 1667
rect 3252 1633 3264 1667
rect 3206 1607 3264 1633
rect 3306 1667 3364 1693
rect 3306 1633 3318 1667
rect 3352 1633 3364 1667
rect 3306 1607 3364 1633
rect 3406 1667 3464 1693
rect 3406 1633 3412 1667
rect 3452 1633 3464 1667
rect 3406 1607 3464 1633
rect 3506 1667 3564 1693
rect 3506 1633 3518 1667
rect 3558 1633 3564 1667
rect 3506 1607 3564 1633
rect 3606 1667 3664 1693
rect 3606 1633 3618 1667
rect 3652 1633 3664 1667
rect 3606 1607 3664 1633
rect 3706 1667 3764 1693
rect 3706 1633 3712 1667
rect 3752 1633 3764 1667
rect 3706 1607 3764 1633
rect 3806 1667 3864 1693
rect 3806 1633 3818 1667
rect 3858 1633 3864 1667
rect 3806 1607 3864 1633
rect 3906 1667 3964 1693
rect 3906 1633 3918 1667
rect 3952 1633 3964 1667
rect 3906 1607 3964 1633
rect 4006 1667 4064 1693
rect 4006 1633 4018 1667
rect 4052 1633 4064 1667
rect 4006 1607 4064 1633
rect 4106 1667 4164 1693
rect 4106 1633 4118 1667
rect 4152 1633 4164 1667
rect 4106 1607 4164 1633
rect 4206 1667 4264 1693
rect 4206 1633 4218 1667
rect 4252 1633 4264 1667
rect 4206 1607 4264 1633
rect 4306 1667 4364 1693
rect 4306 1633 4318 1667
rect 4352 1633 4364 1667
rect 4306 1607 4364 1633
rect 4406 1667 4464 1693
rect 4406 1633 4412 1667
rect 4452 1633 4464 1667
rect 4406 1607 4464 1633
rect 4506 1667 4564 1693
rect 4506 1633 4518 1667
rect 4558 1633 4564 1667
rect 4506 1607 4564 1633
rect 4606 1667 4664 1693
rect 4606 1633 4618 1667
rect 4652 1633 4664 1667
rect 4606 1607 4664 1633
rect 4706 1667 4764 1693
rect 4706 1633 4718 1667
rect 4752 1633 4764 1667
rect 4706 1607 4764 1633
rect 4806 1667 4864 1693
rect 4806 1633 4818 1667
rect 4852 1633 4864 1667
rect 4806 1607 4864 1633
rect 4906 1667 4964 1693
rect 4906 1633 4918 1667
rect 4952 1633 4964 1667
rect 4906 1607 4964 1633
rect 5006 1667 5064 1693
rect 5006 1633 5018 1667
rect 5052 1633 5064 1667
rect 5006 1607 5064 1633
rect 5106 1667 5164 1693
rect 5106 1633 5118 1667
rect 5152 1633 5164 1667
rect 5106 1607 5164 1633
rect 5206 1667 5264 1693
rect 5206 1633 5218 1667
rect 5252 1633 5264 1667
rect 5206 1607 5264 1633
rect 5306 1667 5364 1693
rect 5306 1633 5312 1667
rect 5352 1633 5364 1667
rect 5306 1607 5364 1633
rect 5406 1667 5464 1693
rect 5406 1633 5418 1667
rect 5458 1633 5464 1667
rect 5406 1607 5464 1633
rect 5506 1667 5564 1693
rect 5506 1633 5518 1667
rect 5552 1633 5564 1667
rect 5506 1607 5564 1633
rect 5606 1667 5664 1693
rect 5606 1633 5618 1667
rect 5652 1633 5664 1667
rect 5606 1607 5664 1633
rect 5706 1667 5764 1693
rect 5706 1633 5712 1667
rect 5752 1633 5764 1667
rect 5706 1607 5764 1633
rect 5806 1667 5864 1693
rect 5806 1633 5818 1667
rect 5858 1633 5864 1667
rect 5806 1607 5864 1633
rect 5906 1667 5964 1693
rect 5906 1633 5912 1667
rect 5952 1633 5964 1667
rect 5906 1607 5964 1633
rect 6006 1667 6064 1693
rect 6006 1633 6018 1667
rect 6058 1633 6064 1667
rect 6006 1607 6064 1633
rect 6106 1667 6164 1693
rect 6106 1633 6118 1667
rect 6152 1633 6164 1667
rect 6106 1607 6164 1633
rect 6206 1667 6264 1693
rect 6206 1633 6218 1667
rect 6252 1633 6264 1667
rect 6206 1607 6264 1633
rect 6306 1667 6364 1693
rect 6306 1633 6318 1667
rect 6352 1633 6364 1667
rect 6306 1607 6364 1633
rect 6406 1667 6464 1693
rect 6618 1686 6862 1720
rect 6406 1633 6418 1667
rect 6452 1633 6464 1667
rect 6508 1648 6516 1682
rect 6558 1648 6574 1682
rect 6618 1667 6652 1686
rect 6406 1607 6464 1633
rect 6828 1667 6862 1686
rect 6618 1617 6652 1633
rect 6696 1618 6712 1652
rect 6754 1618 6762 1652
rect 6828 1617 6862 1633
rect 6928 1667 7162 1683
rect 6962 1633 7028 1667
rect 7062 1633 7128 1667
rect 6928 1617 7162 1633
rect 7228 1667 7262 1683
rect 7228 1617 7262 1633
rect 7328 1667 7462 1683
rect 7362 1633 7428 1667
rect 7328 1617 7462 1633
rect 6 1527 64 1553
rect 6 1493 18 1527
rect 58 1493 64 1527
rect 6 1467 64 1493
rect 106 1527 164 1553
rect 106 1493 112 1527
rect 152 1493 164 1527
rect 106 1467 164 1493
rect 206 1527 264 1553
rect 206 1493 218 1527
rect 258 1493 264 1527
rect 206 1467 264 1493
rect 306 1527 364 1553
rect 306 1493 318 1527
rect 352 1493 364 1527
rect 306 1467 364 1493
rect 406 1527 464 1553
rect 406 1493 412 1527
rect 452 1493 464 1527
rect 406 1467 464 1493
rect 506 1527 564 1553
rect 506 1493 518 1527
rect 558 1493 564 1527
rect 506 1467 564 1493
rect 606 1527 664 1553
rect 606 1493 618 1527
rect 652 1493 664 1527
rect 606 1467 664 1493
rect 706 1527 764 1553
rect 706 1493 718 1527
rect 752 1493 764 1527
rect 706 1467 764 1493
rect 806 1527 864 1553
rect 806 1493 818 1527
rect 852 1493 864 1527
rect 806 1467 864 1493
rect 906 1527 964 1553
rect 906 1493 918 1527
rect 952 1493 964 1527
rect 906 1467 964 1493
rect 1006 1527 1064 1553
rect 1006 1493 1018 1527
rect 1052 1493 1064 1527
rect 1006 1467 1064 1493
rect 1106 1527 1164 1553
rect 1106 1493 1118 1527
rect 1152 1493 1164 1527
rect 1106 1467 1164 1493
rect 1206 1527 1264 1553
rect 1206 1493 1218 1527
rect 1252 1493 1264 1527
rect 1206 1467 1264 1493
rect 1306 1527 1364 1553
rect 1306 1493 1318 1527
rect 1352 1493 1364 1527
rect 1306 1467 1364 1493
rect 1406 1527 1464 1553
rect 1406 1493 1418 1527
rect 1452 1493 1464 1527
rect 1406 1467 1464 1493
rect 1506 1527 1564 1553
rect 1506 1493 1518 1527
rect 1552 1493 1564 1527
rect 1506 1467 1564 1493
rect 1606 1527 1664 1553
rect 1606 1493 1612 1527
rect 1652 1493 1664 1527
rect 1606 1467 1664 1493
rect 1706 1527 1764 1553
rect 1706 1493 1718 1527
rect 1758 1493 1764 1527
rect 1706 1467 1764 1493
rect 1806 1527 1864 1553
rect 1806 1493 1818 1527
rect 1852 1493 1864 1527
rect 1806 1467 1864 1493
rect 1906 1527 1964 1553
rect 1906 1493 1918 1527
rect 1952 1493 1964 1527
rect 1906 1467 1964 1493
rect 2006 1527 2064 1553
rect 2006 1493 2018 1527
rect 2052 1493 2064 1527
rect 2006 1467 2064 1493
rect 2106 1527 2164 1553
rect 2106 1493 2118 1527
rect 2152 1493 2164 1527
rect 2106 1467 2164 1493
rect 2206 1527 2264 1553
rect 2206 1493 2218 1527
rect 2252 1493 2264 1527
rect 2206 1467 2264 1493
rect 2306 1527 2364 1553
rect 2306 1493 2318 1527
rect 2352 1493 2364 1527
rect 2306 1467 2364 1493
rect 2406 1527 2464 1553
rect 2406 1493 2418 1527
rect 2452 1493 2464 1527
rect 2406 1467 2464 1493
rect 2506 1527 2564 1553
rect 2506 1493 2518 1527
rect 2552 1493 2564 1527
rect 2506 1467 2564 1493
rect 2606 1527 2664 1553
rect 2606 1493 2618 1527
rect 2652 1493 2664 1527
rect 2606 1467 2664 1493
rect 2706 1527 2764 1553
rect 2706 1493 2718 1527
rect 2752 1493 2764 1527
rect 2706 1467 2764 1493
rect 2806 1527 2864 1553
rect 2806 1493 2818 1527
rect 2852 1493 2864 1527
rect 2806 1467 2864 1493
rect 2906 1527 2964 1553
rect 2906 1493 2918 1527
rect 2952 1493 2964 1527
rect 2906 1467 2964 1493
rect 3006 1527 3064 1553
rect 3006 1493 3018 1527
rect 3052 1493 3064 1527
rect 3006 1467 3064 1493
rect 3106 1527 3164 1553
rect 3106 1493 3118 1527
rect 3152 1493 3164 1527
rect 3106 1467 3164 1493
rect 3206 1527 3264 1553
rect 3206 1493 3218 1527
rect 3252 1493 3264 1527
rect 3206 1467 3264 1493
rect 3306 1527 3364 1553
rect 3306 1493 3318 1527
rect 3352 1493 3364 1527
rect 3306 1467 3364 1493
rect 3406 1527 3464 1553
rect 3406 1493 3418 1527
rect 3452 1493 3464 1527
rect 3406 1467 3464 1493
rect 3506 1527 3564 1553
rect 3506 1493 3518 1527
rect 3552 1493 3564 1527
rect 3506 1467 3564 1493
rect 3606 1527 3664 1553
rect 3606 1493 3618 1527
rect 3652 1493 3664 1527
rect 3606 1467 3664 1493
rect 3706 1527 3764 1553
rect 3706 1493 3718 1527
rect 3752 1493 3764 1527
rect 3706 1467 3764 1493
rect 3806 1527 3864 1553
rect 3806 1493 3818 1527
rect 3852 1493 3864 1527
rect 3806 1467 3864 1493
rect 3906 1527 3964 1553
rect 3906 1493 3918 1527
rect 3952 1493 3964 1527
rect 3906 1467 3964 1493
rect 4006 1527 4064 1553
rect 4006 1493 4018 1527
rect 4052 1493 4064 1527
rect 4006 1467 4064 1493
rect 4106 1527 4164 1553
rect 4106 1493 4112 1527
rect 4152 1493 4164 1527
rect 4106 1467 4164 1493
rect 4206 1527 4264 1553
rect 4206 1493 4218 1527
rect 4258 1493 4264 1527
rect 4206 1467 4264 1493
rect 4306 1527 4364 1553
rect 4306 1493 4318 1527
rect 4352 1493 4364 1527
rect 4306 1467 4364 1493
rect 4406 1527 4464 1553
rect 4406 1493 4412 1527
rect 4452 1493 4464 1527
rect 4406 1467 4464 1493
rect 4506 1527 4564 1553
rect 4506 1493 4518 1527
rect 4558 1493 4564 1527
rect 4506 1467 4564 1493
rect 4606 1527 4664 1553
rect 4606 1493 4618 1527
rect 4652 1493 4664 1527
rect 4606 1467 4664 1493
rect 4706 1527 4764 1553
rect 4706 1493 4718 1527
rect 4752 1493 4764 1527
rect 4706 1467 4764 1493
rect 4806 1527 4864 1553
rect 4806 1493 4818 1527
rect 4852 1493 4864 1527
rect 4806 1467 4864 1493
rect 4906 1527 4964 1553
rect 4906 1493 4918 1527
rect 4952 1493 4964 1527
rect 4906 1467 4964 1493
rect 5006 1527 5064 1553
rect 5006 1493 5012 1527
rect 5052 1493 5064 1527
rect 5006 1467 5064 1493
rect 5106 1527 5164 1553
rect 5106 1493 5118 1527
rect 5158 1493 5164 1527
rect 5106 1467 5164 1493
rect 5206 1527 5264 1553
rect 5206 1493 5212 1527
rect 5252 1493 5264 1527
rect 5206 1467 5264 1493
rect 5306 1527 5364 1553
rect 5306 1493 5318 1527
rect 5358 1493 5364 1527
rect 5306 1467 5364 1493
rect 5406 1527 5464 1553
rect 5406 1493 5412 1527
rect 5452 1493 5464 1527
rect 5406 1467 5464 1493
rect 5506 1527 5564 1553
rect 5506 1493 5518 1527
rect 5558 1493 5564 1527
rect 5506 1467 5564 1493
rect 5606 1527 5664 1553
rect 5606 1493 5618 1527
rect 5652 1493 5664 1527
rect 5606 1467 5664 1493
rect 5706 1527 5764 1553
rect 5706 1493 5712 1527
rect 5752 1493 5764 1527
rect 5706 1467 5764 1493
rect 5806 1527 5864 1553
rect 5806 1493 5818 1527
rect 5858 1493 5864 1527
rect 5806 1467 5864 1493
rect 5906 1527 5964 1553
rect 5906 1493 5912 1527
rect 5952 1493 5964 1527
rect 5906 1467 5964 1493
rect 6006 1527 6064 1553
rect 6006 1493 6018 1527
rect 6058 1493 6064 1527
rect 6006 1467 6064 1493
rect 6106 1527 6164 1553
rect 6106 1493 6118 1527
rect 6152 1493 6164 1527
rect 6106 1467 6164 1493
rect 6206 1527 6264 1553
rect 6206 1493 6212 1527
rect 6252 1493 6264 1527
rect 6206 1467 6264 1493
rect 6306 1527 6364 1553
rect 6306 1493 6318 1527
rect 6358 1493 6364 1527
rect 6306 1467 6364 1493
rect 6406 1527 6464 1553
rect 6618 1546 6862 1580
rect 6406 1493 6412 1527
rect 6452 1493 6464 1527
rect 6508 1508 6516 1542
rect 6558 1508 6574 1542
rect 6618 1527 6652 1546
rect 6406 1467 6464 1493
rect 6828 1543 6862 1546
rect 6828 1527 6962 1543
rect 6618 1477 6652 1493
rect 6696 1478 6712 1512
rect 6754 1478 6762 1512
rect 6862 1493 6928 1527
rect 6828 1477 6962 1493
rect 7028 1527 7062 1543
rect 7028 1477 7062 1493
rect 7128 1527 7262 1543
rect 7162 1493 7228 1527
rect 7128 1477 7262 1493
rect 7328 1527 7462 1543
rect 7362 1493 7428 1527
rect 7328 1477 7462 1493
rect 6 1387 64 1413
rect 6 1353 18 1387
rect 52 1353 64 1387
rect 6 1327 64 1353
rect 106 1387 164 1413
rect 106 1353 118 1387
rect 152 1353 164 1387
rect 106 1327 164 1353
rect 206 1387 264 1413
rect 206 1353 212 1387
rect 252 1353 264 1387
rect 206 1327 264 1353
rect 306 1387 364 1413
rect 306 1353 318 1387
rect 358 1353 364 1387
rect 306 1327 364 1353
rect 406 1387 464 1413
rect 406 1353 418 1387
rect 452 1353 464 1387
rect 406 1327 464 1353
rect 506 1387 564 1413
rect 506 1353 512 1387
rect 552 1353 564 1387
rect 506 1327 564 1353
rect 606 1387 664 1413
rect 606 1353 618 1387
rect 658 1353 664 1387
rect 606 1327 664 1353
rect 706 1387 764 1413
rect 706 1353 718 1387
rect 752 1353 764 1387
rect 706 1327 764 1353
rect 806 1387 864 1413
rect 806 1353 818 1387
rect 852 1353 864 1387
rect 806 1327 864 1353
rect 906 1387 964 1413
rect 906 1353 918 1387
rect 952 1353 964 1387
rect 906 1327 964 1353
rect 1006 1387 1064 1413
rect 1006 1353 1018 1387
rect 1052 1353 1064 1387
rect 1006 1327 1064 1353
rect 1106 1387 1164 1413
rect 1106 1353 1118 1387
rect 1152 1353 1164 1387
rect 1106 1327 1164 1353
rect 1206 1387 1264 1413
rect 1206 1353 1218 1387
rect 1252 1353 1264 1387
rect 1206 1327 1264 1353
rect 1306 1387 1364 1413
rect 1306 1353 1318 1387
rect 1352 1353 1364 1387
rect 1306 1327 1364 1353
rect 1406 1387 1464 1413
rect 1406 1353 1418 1387
rect 1452 1353 1464 1387
rect 1406 1327 1464 1353
rect 1506 1387 1564 1413
rect 1506 1353 1512 1387
rect 1552 1353 1564 1387
rect 1506 1327 1564 1353
rect 1606 1387 1664 1413
rect 1606 1353 1618 1387
rect 1658 1353 1664 1387
rect 1606 1327 1664 1353
rect 1706 1387 1764 1413
rect 1706 1353 1712 1387
rect 1752 1353 1764 1387
rect 1706 1327 1764 1353
rect 1806 1387 1864 1413
rect 1806 1353 1818 1387
rect 1858 1353 1864 1387
rect 1806 1327 1864 1353
rect 1906 1387 1964 1413
rect 1906 1353 1918 1387
rect 1952 1353 1964 1387
rect 1906 1327 1964 1353
rect 2006 1387 2064 1413
rect 2006 1353 2018 1387
rect 2052 1353 2064 1387
rect 2006 1327 2064 1353
rect 2106 1387 2164 1413
rect 2106 1353 2118 1387
rect 2152 1353 2164 1387
rect 2106 1327 2164 1353
rect 2206 1387 2264 1413
rect 2206 1353 2218 1387
rect 2252 1353 2264 1387
rect 2206 1327 2264 1353
rect 2306 1387 2364 1413
rect 2306 1353 2318 1387
rect 2352 1353 2364 1387
rect 2306 1327 2364 1353
rect 2406 1387 2464 1413
rect 2406 1353 2418 1387
rect 2452 1353 2464 1387
rect 2406 1327 2464 1353
rect 2506 1387 2564 1413
rect 2506 1353 2518 1387
rect 2552 1353 2564 1387
rect 2506 1327 2564 1353
rect 2606 1387 2664 1413
rect 2606 1353 2618 1387
rect 2652 1353 2664 1387
rect 2606 1327 2664 1353
rect 2706 1387 2764 1413
rect 2706 1353 2718 1387
rect 2752 1353 2764 1387
rect 2706 1327 2764 1353
rect 2806 1387 2864 1413
rect 2806 1353 2818 1387
rect 2852 1353 2864 1387
rect 2806 1327 2864 1353
rect 2906 1387 2964 1413
rect 2906 1353 2912 1387
rect 2952 1353 2964 1387
rect 2906 1327 2964 1353
rect 3006 1387 3064 1413
rect 3006 1353 3018 1387
rect 3058 1353 3064 1387
rect 3006 1327 3064 1353
rect 3106 1387 3164 1413
rect 3106 1353 3118 1387
rect 3152 1353 3164 1387
rect 3106 1327 3164 1353
rect 3206 1387 3264 1413
rect 3206 1353 3218 1387
rect 3252 1353 3264 1387
rect 3206 1327 3264 1353
rect 3306 1387 3364 1413
rect 3306 1353 3318 1387
rect 3352 1353 3364 1387
rect 3306 1327 3364 1353
rect 3406 1387 3464 1413
rect 3406 1353 3418 1387
rect 3452 1353 3464 1387
rect 3406 1327 3464 1353
rect 3506 1387 3564 1413
rect 3506 1353 3512 1387
rect 3552 1353 3564 1387
rect 3506 1327 3564 1353
rect 3606 1387 3664 1413
rect 3606 1353 3618 1387
rect 3658 1353 3664 1387
rect 3606 1327 3664 1353
rect 3706 1387 3764 1413
rect 3706 1353 3718 1387
rect 3752 1353 3764 1387
rect 3706 1327 3764 1353
rect 3806 1387 3864 1413
rect 3806 1353 3812 1387
rect 3852 1353 3864 1387
rect 3806 1327 3864 1353
rect 3906 1387 3964 1413
rect 3906 1353 3918 1387
rect 3958 1353 3964 1387
rect 3906 1327 3964 1353
rect 4006 1387 4064 1413
rect 4006 1353 4018 1387
rect 4052 1353 4064 1387
rect 4006 1327 4064 1353
rect 4106 1387 4164 1413
rect 4106 1353 4118 1387
rect 4152 1353 4164 1387
rect 4106 1327 4164 1353
rect 4206 1387 4264 1413
rect 4206 1353 4218 1387
rect 4252 1353 4264 1387
rect 4206 1327 4264 1353
rect 4306 1387 4364 1413
rect 4306 1353 4318 1387
rect 4352 1353 4364 1387
rect 4306 1327 4364 1353
rect 4406 1387 4464 1413
rect 4406 1353 4418 1387
rect 4452 1353 4464 1387
rect 4406 1327 4464 1353
rect 4506 1387 4564 1413
rect 4506 1353 4518 1387
rect 4552 1353 4564 1387
rect 4506 1327 4564 1353
rect 4606 1387 4664 1413
rect 4606 1353 4618 1387
rect 4652 1353 4664 1387
rect 4606 1327 4664 1353
rect 4706 1387 4764 1413
rect 4706 1353 4718 1387
rect 4752 1353 4764 1387
rect 4706 1327 4764 1353
rect 4806 1387 4864 1413
rect 4806 1353 4812 1387
rect 4852 1353 4864 1387
rect 4806 1327 4864 1353
rect 4906 1387 4964 1413
rect 4906 1353 4918 1387
rect 4958 1353 4964 1387
rect 4906 1327 4964 1353
rect 5006 1387 5064 1413
rect 5006 1353 5012 1387
rect 5052 1353 5064 1387
rect 5006 1327 5064 1353
rect 5106 1387 5164 1413
rect 5106 1353 5118 1387
rect 5158 1353 5164 1387
rect 5106 1327 5164 1353
rect 5206 1387 5264 1413
rect 5206 1353 5218 1387
rect 5252 1353 5264 1387
rect 5206 1327 5264 1353
rect 5306 1387 5364 1413
rect 5306 1353 5318 1387
rect 5352 1353 5364 1387
rect 5306 1327 5364 1353
rect 5406 1387 5464 1413
rect 5406 1353 5418 1387
rect 5452 1353 5464 1387
rect 5406 1327 5464 1353
rect 5506 1387 5564 1413
rect 5506 1353 5518 1387
rect 5552 1353 5564 1387
rect 5506 1327 5564 1353
rect 5606 1387 5664 1413
rect 5606 1353 5618 1387
rect 5652 1353 5664 1387
rect 5606 1327 5664 1353
rect 5706 1387 5764 1413
rect 5706 1353 5718 1387
rect 5752 1353 5764 1387
rect 5706 1327 5764 1353
rect 5806 1387 5864 1413
rect 5806 1353 5818 1387
rect 5852 1353 5864 1387
rect 5806 1327 5864 1353
rect 5906 1387 5964 1413
rect 5906 1353 5918 1387
rect 5952 1353 5964 1387
rect 5906 1327 5964 1353
rect 6006 1387 6064 1413
rect 6006 1353 6018 1387
rect 6052 1353 6064 1387
rect 6006 1327 6064 1353
rect 6106 1387 6164 1413
rect 6106 1353 6112 1387
rect 6152 1353 6164 1387
rect 6106 1327 6164 1353
rect 6206 1387 6264 1413
rect 6206 1353 6218 1387
rect 6258 1353 6264 1387
rect 6206 1327 6264 1353
rect 6306 1387 6364 1413
rect 6306 1353 6318 1387
rect 6352 1353 6364 1387
rect 6306 1327 6364 1353
rect 6406 1387 6464 1413
rect 6618 1406 6862 1440
rect 6406 1353 6418 1387
rect 6452 1353 6464 1387
rect 6508 1368 6516 1402
rect 6558 1368 6574 1402
rect 6618 1387 6652 1406
rect 6406 1327 6464 1353
rect 6828 1387 6862 1406
rect 6618 1337 6652 1353
rect 6696 1338 6712 1372
rect 6754 1338 6762 1372
rect 6828 1337 6862 1353
rect 6928 1387 7062 1403
rect 6962 1353 7028 1387
rect 6928 1337 7062 1353
rect 7128 1387 7262 1403
rect 7162 1353 7228 1387
rect 7128 1337 7262 1353
rect 7328 1387 7462 1403
rect 7362 1353 7428 1387
rect 7328 1337 7462 1353
rect 8 1230 18 1264
rect 52 1230 118 1264
rect 152 1230 168 1264
rect 208 1246 218 1280
rect 252 1246 318 1280
rect 352 1246 368 1280
rect 408 1230 418 1264
rect 452 1230 518 1264
rect 552 1230 568 1264
rect 608 1246 618 1280
rect 652 1246 718 1280
rect 752 1246 768 1280
rect 808 1230 818 1264
rect 852 1230 918 1264
rect 952 1230 968 1264
rect 1008 1246 1018 1280
rect 1052 1246 1118 1280
rect 1152 1246 1168 1280
rect 1208 1230 1218 1264
rect 1252 1230 1318 1264
rect 1352 1230 1368 1264
rect 1408 1246 1418 1280
rect 1452 1246 1518 1280
rect 1552 1246 1568 1280
rect 1608 1230 1618 1264
rect 1652 1230 1718 1264
rect 1752 1230 1768 1264
rect 1808 1246 1818 1280
rect 1852 1246 1918 1280
rect 1952 1246 1968 1280
rect 2008 1230 2018 1264
rect 2052 1230 2118 1264
rect 2152 1230 2168 1264
rect 2208 1246 2218 1280
rect 2252 1246 2318 1280
rect 2352 1246 2368 1280
rect 2408 1230 2418 1264
rect 2452 1230 2518 1264
rect 2552 1230 2568 1264
rect 2608 1246 2618 1280
rect 2652 1246 2718 1280
rect 2752 1246 2768 1280
rect 2808 1230 2818 1264
rect 2852 1230 2918 1264
rect 2952 1230 2968 1264
rect 3008 1246 3018 1280
rect 3052 1246 3118 1280
rect 3152 1246 3168 1280
rect 3208 1230 3218 1264
rect 3252 1230 3318 1264
rect 3352 1230 3368 1264
rect 3408 1246 3418 1280
rect 3452 1246 3518 1280
rect 3552 1246 3568 1280
rect 3608 1230 3618 1264
rect 3652 1230 3718 1264
rect 3752 1230 3768 1264
rect 3808 1246 3818 1280
rect 3852 1246 3918 1280
rect 3952 1246 3968 1280
rect 4008 1230 4018 1264
rect 4052 1230 4118 1264
rect 4152 1230 4168 1264
rect 4208 1246 4218 1280
rect 4252 1246 4318 1280
rect 4352 1246 4368 1280
rect 4408 1230 4418 1264
rect 4452 1230 4518 1264
rect 4552 1230 4568 1264
rect 4608 1246 4618 1280
rect 4652 1246 4718 1280
rect 4752 1246 4768 1280
rect 4808 1230 4818 1264
rect 4852 1230 4918 1264
rect 4952 1230 4968 1264
rect 5008 1246 5018 1280
rect 5052 1246 5118 1280
rect 5152 1246 5168 1280
rect 5208 1230 5218 1264
rect 5252 1230 5318 1264
rect 5352 1230 5368 1264
rect 5408 1246 5418 1280
rect 5452 1246 5518 1280
rect 5552 1246 5568 1280
rect 5608 1230 5618 1264
rect 5652 1230 5718 1264
rect 5752 1230 5768 1264
rect 5808 1246 5818 1280
rect 5852 1246 5918 1280
rect 5952 1246 5968 1280
rect 6008 1230 6018 1264
rect 6052 1230 6118 1264
rect 6152 1230 6168 1264
rect 6208 1246 6218 1280
rect 6252 1246 6318 1280
rect 6352 1246 6368 1280
rect 6516 1261 6568 1278
rect 6550 1244 6568 1261
rect 6602 1244 6618 1278
rect 6652 1244 6668 1278
rect 6702 1249 6720 1278
rect 6702 1244 6754 1249
rect 6862 1244 6878 1278
rect 6912 1244 6928 1278
rect 6962 1244 6978 1278
rect 7012 1244 7028 1278
rect 7062 1244 7078 1278
rect 7112 1244 7128 1278
rect 7162 1244 7178 1278
rect 7212 1244 7228 1278
rect 7262 1244 7278 1278
rect 7312 1244 7328 1278
rect 7362 1244 7378 1278
rect 7412 1244 7428 1278
rect 6 1157 64 1183
rect 6 1123 18 1157
rect 52 1123 64 1157
rect 6 1097 64 1123
rect 106 1157 164 1183
rect 106 1123 118 1157
rect 152 1123 164 1157
rect 106 1097 164 1123
rect 206 1157 264 1183
rect 206 1123 218 1157
rect 252 1123 264 1157
rect 206 1097 264 1123
rect 306 1157 364 1183
rect 306 1123 312 1157
rect 352 1123 364 1157
rect 306 1097 364 1123
rect 406 1157 464 1183
rect 406 1123 418 1157
rect 458 1123 464 1157
rect 406 1097 464 1123
rect 506 1157 564 1183
rect 506 1123 512 1157
rect 552 1123 564 1157
rect 506 1097 564 1123
rect 606 1157 664 1183
rect 606 1123 618 1157
rect 658 1123 664 1157
rect 606 1097 664 1123
rect 706 1157 764 1183
rect 706 1123 712 1157
rect 752 1123 764 1157
rect 706 1097 764 1123
rect 806 1157 864 1183
rect 806 1123 818 1157
rect 858 1123 864 1157
rect 806 1097 864 1123
rect 906 1157 964 1183
rect 906 1123 918 1157
rect 952 1123 964 1157
rect 906 1097 964 1123
rect 1006 1157 1064 1183
rect 1006 1123 1018 1157
rect 1052 1123 1064 1157
rect 1006 1097 1064 1123
rect 1106 1157 1164 1183
rect 1106 1123 1118 1157
rect 1152 1123 1164 1157
rect 1106 1097 1164 1123
rect 1206 1157 1264 1183
rect 1206 1123 1212 1157
rect 1252 1123 1264 1157
rect 1206 1097 1264 1123
rect 1306 1157 1364 1183
rect 1306 1123 1318 1157
rect 1358 1123 1364 1157
rect 1306 1097 1364 1123
rect 1406 1157 1464 1183
rect 1406 1123 1418 1157
rect 1452 1123 1464 1157
rect 1406 1097 1464 1123
rect 1506 1157 1564 1183
rect 1506 1123 1518 1157
rect 1552 1123 1564 1157
rect 1506 1097 1564 1123
rect 1606 1157 1664 1183
rect 1606 1123 1618 1157
rect 1652 1123 1664 1157
rect 1606 1097 1664 1123
rect 1706 1157 1764 1183
rect 1706 1123 1718 1157
rect 1752 1123 1764 1157
rect 1706 1097 1764 1123
rect 1806 1157 1864 1183
rect 1806 1123 1818 1157
rect 1852 1123 1864 1157
rect 1806 1097 1864 1123
rect 1906 1157 1964 1183
rect 1906 1123 1918 1157
rect 1952 1123 1964 1157
rect 1906 1097 1964 1123
rect 2006 1157 2064 1183
rect 2006 1123 2018 1157
rect 2052 1123 2064 1157
rect 2006 1097 2064 1123
rect 2106 1157 2164 1183
rect 2106 1123 2118 1157
rect 2152 1123 2164 1157
rect 2106 1097 2164 1123
rect 2206 1157 2264 1183
rect 2206 1123 2218 1157
rect 2252 1123 2264 1157
rect 2206 1097 2264 1123
rect 2306 1157 2364 1183
rect 2306 1123 2318 1157
rect 2352 1123 2364 1157
rect 2306 1097 2364 1123
rect 2406 1157 2464 1183
rect 2406 1123 2418 1157
rect 2452 1123 2464 1157
rect 2406 1097 2464 1123
rect 2506 1157 2564 1183
rect 2506 1123 2512 1157
rect 2552 1123 2564 1157
rect 2506 1097 2564 1123
rect 2606 1157 2664 1183
rect 2606 1123 2618 1157
rect 2658 1123 2664 1157
rect 2606 1097 2664 1123
rect 2706 1157 2764 1183
rect 2706 1123 2712 1157
rect 2752 1123 2764 1157
rect 2706 1097 2764 1123
rect 2806 1157 2864 1183
rect 2806 1123 2818 1157
rect 2858 1123 2864 1157
rect 2806 1097 2864 1123
rect 2906 1157 2964 1183
rect 2906 1123 2918 1157
rect 2952 1123 2964 1157
rect 2906 1097 2964 1123
rect 3006 1157 3064 1183
rect 3006 1123 3018 1157
rect 3052 1123 3064 1157
rect 3006 1097 3064 1123
rect 3106 1157 3164 1183
rect 3106 1123 3118 1157
rect 3152 1123 3164 1157
rect 3106 1097 3164 1123
rect 3206 1157 3264 1183
rect 3206 1123 3218 1157
rect 3252 1123 3264 1157
rect 3206 1097 3264 1123
rect 3306 1157 3364 1183
rect 3306 1123 3318 1157
rect 3352 1123 3364 1157
rect 3306 1097 3364 1123
rect 3406 1157 3464 1183
rect 3406 1123 3418 1157
rect 3452 1123 3464 1157
rect 3406 1097 3464 1123
rect 3506 1157 3564 1183
rect 3506 1123 3518 1157
rect 3552 1123 3564 1157
rect 3506 1097 3564 1123
rect 3606 1157 3664 1183
rect 3606 1123 3618 1157
rect 3652 1123 3664 1157
rect 3606 1097 3664 1123
rect 3706 1157 3764 1183
rect 3706 1123 3718 1157
rect 3752 1123 3764 1157
rect 3706 1097 3764 1123
rect 3806 1157 3864 1183
rect 3806 1123 3818 1157
rect 3852 1123 3864 1157
rect 3806 1097 3864 1123
rect 3906 1157 3964 1183
rect 3906 1123 3918 1157
rect 3952 1123 3964 1157
rect 3906 1097 3964 1123
rect 4006 1157 4064 1183
rect 4006 1123 4018 1157
rect 4052 1123 4064 1157
rect 4006 1097 4064 1123
rect 4106 1157 4164 1183
rect 4106 1123 4118 1157
rect 4152 1123 4164 1157
rect 4106 1097 4164 1123
rect 4206 1157 4264 1183
rect 4206 1123 4212 1157
rect 4252 1123 4264 1157
rect 4206 1097 4264 1123
rect 4306 1157 4364 1183
rect 4306 1123 4318 1157
rect 4358 1123 4364 1157
rect 4306 1097 4364 1123
rect 4406 1157 4464 1183
rect 4406 1123 4418 1157
rect 4452 1123 4464 1157
rect 4406 1097 4464 1123
rect 4506 1157 4564 1183
rect 4506 1123 4518 1157
rect 4552 1123 4564 1157
rect 4506 1097 4564 1123
rect 4606 1157 4664 1183
rect 4606 1123 4618 1157
rect 4652 1123 4664 1157
rect 4606 1097 4664 1123
rect 4706 1157 4764 1183
rect 4706 1123 4718 1157
rect 4752 1123 4764 1157
rect 4706 1097 4764 1123
rect 4806 1157 4864 1183
rect 4806 1123 4818 1157
rect 4852 1123 4864 1157
rect 4806 1097 4864 1123
rect 4906 1157 4964 1183
rect 4906 1123 4918 1157
rect 4952 1123 4964 1157
rect 4906 1097 4964 1123
rect 5006 1157 5064 1183
rect 5006 1123 5018 1157
rect 5052 1123 5064 1157
rect 5006 1097 5064 1123
rect 5106 1157 5164 1183
rect 5106 1123 5118 1157
rect 5152 1123 5164 1157
rect 5106 1097 5164 1123
rect 5206 1157 5264 1183
rect 5206 1123 5218 1157
rect 5252 1123 5264 1157
rect 5206 1097 5264 1123
rect 5306 1157 5364 1183
rect 5306 1123 5318 1157
rect 5352 1123 5364 1157
rect 5306 1097 5364 1123
rect 5406 1157 5464 1183
rect 5406 1123 5412 1157
rect 5452 1123 5464 1157
rect 5406 1097 5464 1123
rect 5506 1157 5564 1183
rect 5506 1123 5518 1157
rect 5558 1123 5564 1157
rect 5506 1097 5564 1123
rect 5606 1157 5664 1183
rect 5606 1123 5618 1157
rect 5652 1123 5664 1157
rect 5606 1097 5664 1123
rect 5706 1157 5764 1183
rect 5706 1123 5718 1157
rect 5752 1123 5764 1157
rect 5706 1097 5764 1123
rect 5806 1157 5864 1183
rect 5806 1123 5818 1157
rect 5852 1123 5864 1157
rect 5806 1097 5864 1123
rect 5906 1157 5964 1183
rect 5906 1123 5912 1157
rect 5952 1123 5964 1157
rect 5906 1097 5964 1123
rect 6006 1157 6064 1183
rect 6006 1123 6018 1157
rect 6058 1123 6064 1157
rect 6006 1097 6064 1123
rect 6106 1157 6164 1183
rect 6106 1123 6118 1157
rect 6152 1123 6164 1157
rect 6106 1097 6164 1123
rect 6206 1157 6264 1183
rect 6206 1123 6218 1157
rect 6252 1123 6264 1157
rect 6206 1097 6264 1123
rect 6306 1157 6364 1183
rect 6306 1123 6318 1157
rect 6352 1123 6364 1157
rect 6306 1097 6364 1123
rect 6406 1157 6464 1183
rect 6618 1176 6862 1210
rect 6406 1123 6412 1157
rect 6452 1123 6464 1157
rect 6508 1138 6516 1172
rect 6558 1138 6574 1172
rect 6618 1157 6652 1176
rect 6406 1097 6464 1123
rect 6828 1173 6862 1176
rect 6828 1157 6962 1173
rect 6618 1107 6652 1123
rect 6696 1108 6712 1142
rect 6754 1108 6762 1142
rect 6862 1123 6928 1157
rect 6828 1107 6962 1123
rect 7028 1157 7162 1173
rect 7062 1123 7128 1157
rect 7028 1107 7162 1123
rect 7228 1157 7362 1173
rect 7262 1123 7328 1157
rect 7228 1107 7362 1123
rect 7428 1157 7462 1173
rect 7428 1107 7462 1123
rect 6 1017 64 1043
rect 6 983 18 1017
rect 52 983 64 1017
rect 6 957 64 983
rect 106 1017 164 1043
rect 106 983 118 1017
rect 152 983 164 1017
rect 106 957 164 983
rect 206 1017 264 1043
rect 206 983 218 1017
rect 252 983 264 1017
rect 206 957 264 983
rect 306 1017 364 1043
rect 306 983 318 1017
rect 352 983 364 1017
rect 306 957 364 983
rect 406 1017 464 1043
rect 406 983 418 1017
rect 452 983 464 1017
rect 406 957 464 983
rect 506 1017 564 1043
rect 506 983 518 1017
rect 552 983 564 1017
rect 506 957 564 983
rect 606 1017 664 1043
rect 606 983 618 1017
rect 652 983 664 1017
rect 606 957 664 983
rect 706 1017 764 1043
rect 706 983 718 1017
rect 752 983 764 1017
rect 706 957 764 983
rect 806 1017 864 1043
rect 806 983 818 1017
rect 852 983 864 1017
rect 806 957 864 983
rect 906 1017 964 1043
rect 906 983 912 1017
rect 952 983 964 1017
rect 906 957 964 983
rect 1006 1017 1064 1043
rect 1006 983 1018 1017
rect 1058 983 1064 1017
rect 1006 957 1064 983
rect 1106 1017 1164 1043
rect 1106 983 1112 1017
rect 1152 983 1164 1017
rect 1106 957 1164 983
rect 1206 1017 1264 1043
rect 1206 983 1218 1017
rect 1258 983 1264 1017
rect 1206 957 1264 983
rect 1306 1017 1364 1043
rect 1306 983 1318 1017
rect 1352 983 1364 1017
rect 1306 957 1364 983
rect 1406 1017 1464 1043
rect 1406 983 1418 1017
rect 1452 983 1464 1017
rect 1406 957 1464 983
rect 1506 1017 1564 1043
rect 1506 983 1518 1017
rect 1552 983 1564 1017
rect 1506 957 1564 983
rect 1606 1017 1664 1043
rect 1606 983 1618 1017
rect 1652 983 1664 1017
rect 1606 957 1664 983
rect 1706 1017 1764 1043
rect 1706 983 1718 1017
rect 1752 983 1764 1017
rect 1706 957 1764 983
rect 1806 1017 1864 1043
rect 1806 983 1818 1017
rect 1852 983 1864 1017
rect 1806 957 1864 983
rect 1906 1017 1964 1043
rect 1906 983 1918 1017
rect 1952 983 1964 1017
rect 1906 957 1964 983
rect 2006 1017 2064 1043
rect 2006 983 2018 1017
rect 2052 983 2064 1017
rect 2006 957 2064 983
rect 2106 1017 2164 1043
rect 2106 983 2112 1017
rect 2152 983 2164 1017
rect 2106 957 2164 983
rect 2206 1017 2264 1043
rect 2206 983 2218 1017
rect 2258 983 2264 1017
rect 2206 957 2264 983
rect 2306 1017 2364 1043
rect 2306 983 2318 1017
rect 2352 983 2364 1017
rect 2306 957 2364 983
rect 2406 1017 2464 1043
rect 2406 983 2412 1017
rect 2452 983 2464 1017
rect 2406 957 2464 983
rect 2506 1017 2564 1043
rect 2506 983 2518 1017
rect 2558 983 2564 1017
rect 2506 957 2564 983
rect 2606 1017 2664 1043
rect 2606 983 2618 1017
rect 2652 983 2664 1017
rect 2606 957 2664 983
rect 2706 1017 2764 1043
rect 2706 983 2718 1017
rect 2752 983 2764 1017
rect 2706 957 2764 983
rect 2806 1017 2864 1043
rect 2806 983 2818 1017
rect 2852 983 2864 1017
rect 2806 957 2864 983
rect 2906 1017 2964 1043
rect 2906 983 2918 1017
rect 2952 983 2964 1017
rect 2906 957 2964 983
rect 3006 1017 3064 1043
rect 3006 983 3018 1017
rect 3052 983 3064 1017
rect 3006 957 3064 983
rect 3106 1017 3164 1043
rect 3106 983 3118 1017
rect 3152 983 3164 1017
rect 3106 957 3164 983
rect 3206 1017 3264 1043
rect 3206 983 3218 1017
rect 3252 983 3264 1017
rect 3206 957 3264 983
rect 3306 1017 3364 1043
rect 3306 983 3318 1017
rect 3352 983 3364 1017
rect 3306 957 3364 983
rect 3406 1017 3464 1043
rect 3406 983 3418 1017
rect 3452 983 3464 1017
rect 3406 957 3464 983
rect 3506 1017 3564 1043
rect 3506 983 3518 1017
rect 3552 983 3564 1017
rect 3506 957 3564 983
rect 3606 1017 3664 1043
rect 3606 983 3618 1017
rect 3652 983 3664 1017
rect 3606 957 3664 983
rect 3706 1017 3764 1043
rect 3706 983 3718 1017
rect 3752 983 3764 1017
rect 3706 957 3764 983
rect 3806 1017 3864 1043
rect 3806 983 3818 1017
rect 3852 983 3864 1017
rect 3806 957 3864 983
rect 3906 1017 3964 1043
rect 3906 983 3918 1017
rect 3952 983 3964 1017
rect 3906 957 3964 983
rect 4006 1017 4064 1043
rect 4006 983 4018 1017
rect 4052 983 4064 1017
rect 4006 957 4064 983
rect 4106 1017 4164 1043
rect 4106 983 4118 1017
rect 4152 983 4164 1017
rect 4106 957 4164 983
rect 4206 1017 4264 1043
rect 4206 983 4212 1017
rect 4252 983 4264 1017
rect 4206 957 4264 983
rect 4306 1017 4364 1043
rect 4306 983 4318 1017
rect 4358 983 4364 1017
rect 4306 957 4364 983
rect 4406 1017 4464 1043
rect 4406 983 4418 1017
rect 4452 983 4464 1017
rect 4406 957 4464 983
rect 4506 1017 4564 1043
rect 4506 983 4518 1017
rect 4552 983 4564 1017
rect 4506 957 4564 983
rect 4606 1017 4664 1043
rect 4606 983 4618 1017
rect 4652 983 4664 1017
rect 4606 957 4664 983
rect 4706 1017 4764 1043
rect 4706 983 4718 1017
rect 4752 983 4764 1017
rect 4706 957 4764 983
rect 4806 1017 4864 1043
rect 4806 983 4812 1017
rect 4852 983 4864 1017
rect 4806 957 4864 983
rect 4906 1017 4964 1043
rect 4906 983 4918 1017
rect 4958 983 4964 1017
rect 4906 957 4964 983
rect 5006 1017 5064 1043
rect 5006 983 5012 1017
rect 5052 983 5064 1017
rect 5006 957 5064 983
rect 5106 1017 5164 1043
rect 5106 983 5118 1017
rect 5158 983 5164 1017
rect 5106 957 5164 983
rect 5206 1017 5264 1043
rect 5206 983 5218 1017
rect 5252 983 5264 1017
rect 5206 957 5264 983
rect 5306 1017 5364 1043
rect 5306 983 5318 1017
rect 5352 983 5364 1017
rect 5306 957 5364 983
rect 5406 1017 5464 1043
rect 5406 983 5418 1017
rect 5452 983 5464 1017
rect 5406 957 5464 983
rect 5506 1017 5564 1043
rect 5506 983 5518 1017
rect 5552 983 5564 1017
rect 5506 957 5564 983
rect 5606 1017 5664 1043
rect 5606 983 5618 1017
rect 5652 983 5664 1017
rect 5606 957 5664 983
rect 5706 1017 5764 1043
rect 5706 983 5718 1017
rect 5752 983 5764 1017
rect 5706 957 5764 983
rect 5806 1017 5864 1043
rect 5806 983 5818 1017
rect 5852 983 5864 1017
rect 5806 957 5864 983
rect 5906 1017 5964 1043
rect 5906 983 5918 1017
rect 5952 983 5964 1017
rect 5906 957 5964 983
rect 6006 1017 6064 1043
rect 6006 983 6018 1017
rect 6052 983 6064 1017
rect 6006 957 6064 983
rect 6106 1017 6164 1043
rect 6106 983 6118 1017
rect 6152 983 6164 1017
rect 6106 957 6164 983
rect 6206 1017 6264 1043
rect 6206 983 6212 1017
rect 6252 983 6264 1017
rect 6206 957 6264 983
rect 6306 1017 6364 1043
rect 6306 983 6318 1017
rect 6358 983 6364 1017
rect 6306 957 6364 983
rect 6406 1017 6464 1043
rect 6618 1036 6862 1070
rect 6406 983 6412 1017
rect 6452 983 6464 1017
rect 6508 998 6516 1032
rect 6558 998 6574 1032
rect 6618 1017 6652 1036
rect 6406 957 6464 983
rect 6828 1017 6862 1036
rect 6618 967 6652 983
rect 6696 968 6712 1002
rect 6754 968 6762 1002
rect 6828 967 6862 983
rect 6928 1017 7162 1033
rect 6962 983 7028 1017
rect 7062 983 7128 1017
rect 6928 967 7162 983
rect 7228 1017 7362 1033
rect 7262 983 7328 1017
rect 7228 967 7362 983
rect 7428 1017 7462 1033
rect 7428 967 7462 983
rect 6 877 64 903
rect 6 843 18 877
rect 52 843 64 877
rect 6 817 64 843
rect 106 877 164 903
rect 106 843 118 877
rect 152 843 164 877
rect 106 817 164 843
rect 206 877 264 903
rect 206 843 218 877
rect 252 843 264 877
rect 206 817 264 843
rect 306 877 364 903
rect 306 843 318 877
rect 352 843 364 877
rect 306 817 364 843
rect 406 877 464 903
rect 406 843 418 877
rect 452 843 464 877
rect 406 817 464 843
rect 506 877 564 903
rect 506 843 518 877
rect 552 843 564 877
rect 506 817 564 843
rect 606 877 664 903
rect 606 843 618 877
rect 652 843 664 877
rect 606 817 664 843
rect 706 877 764 903
rect 706 843 718 877
rect 752 843 764 877
rect 706 817 764 843
rect 806 877 864 903
rect 806 843 818 877
rect 852 843 864 877
rect 806 817 864 843
rect 906 877 964 903
rect 906 843 918 877
rect 952 843 964 877
rect 906 817 964 843
rect 1006 877 1064 903
rect 1006 843 1012 877
rect 1052 843 1064 877
rect 1006 817 1064 843
rect 1106 877 1164 903
rect 1106 843 1118 877
rect 1158 843 1164 877
rect 1106 817 1164 843
rect 1206 877 1264 903
rect 1206 843 1218 877
rect 1252 843 1264 877
rect 1206 817 1264 843
rect 1306 877 1364 903
rect 1306 843 1318 877
rect 1352 843 1364 877
rect 1306 817 1364 843
rect 1406 877 1464 903
rect 1406 843 1418 877
rect 1452 843 1464 877
rect 1406 817 1464 843
rect 1506 877 1564 903
rect 1506 843 1518 877
rect 1552 843 1564 877
rect 1506 817 1564 843
rect 1606 877 1664 903
rect 1606 843 1618 877
rect 1652 843 1664 877
rect 1606 817 1664 843
rect 1706 877 1764 903
rect 1706 843 1712 877
rect 1752 843 1764 877
rect 1706 817 1764 843
rect 1806 877 1864 903
rect 1806 843 1818 877
rect 1858 843 1864 877
rect 1806 817 1864 843
rect 1906 877 1964 903
rect 1906 843 1918 877
rect 1952 843 1964 877
rect 1906 817 1964 843
rect 2006 877 2064 903
rect 2006 843 2018 877
rect 2052 843 2064 877
rect 2006 817 2064 843
rect 2106 877 2164 903
rect 2106 843 2118 877
rect 2152 843 2164 877
rect 2106 817 2164 843
rect 2206 877 2264 903
rect 2206 843 2218 877
rect 2252 843 2264 877
rect 2206 817 2264 843
rect 2306 877 2364 903
rect 2306 843 2318 877
rect 2352 843 2364 877
rect 2306 817 2364 843
rect 2406 877 2464 903
rect 2406 843 2418 877
rect 2452 843 2464 877
rect 2406 817 2464 843
rect 2506 877 2564 903
rect 2506 843 2518 877
rect 2552 843 2564 877
rect 2506 817 2564 843
rect 2606 877 2664 903
rect 2606 843 2618 877
rect 2652 843 2664 877
rect 2606 817 2664 843
rect 2706 877 2764 903
rect 2706 843 2718 877
rect 2752 843 2764 877
rect 2706 817 2764 843
rect 2806 877 2864 903
rect 2806 843 2818 877
rect 2852 843 2864 877
rect 2806 817 2864 843
rect 2906 877 2964 903
rect 2906 843 2918 877
rect 2952 843 2964 877
rect 2906 817 2964 843
rect 3006 877 3064 903
rect 3006 843 3018 877
rect 3052 843 3064 877
rect 3006 817 3064 843
rect 3106 877 3164 903
rect 3106 843 3118 877
rect 3152 843 3164 877
rect 3106 817 3164 843
rect 3206 877 3264 903
rect 3206 843 3218 877
rect 3252 843 3264 877
rect 3206 817 3264 843
rect 3306 877 3364 903
rect 3306 843 3318 877
rect 3352 843 3364 877
rect 3306 817 3364 843
rect 3406 877 3464 903
rect 3406 843 3418 877
rect 3452 843 3464 877
rect 3406 817 3464 843
rect 3506 877 3564 903
rect 3506 843 3518 877
rect 3552 843 3564 877
rect 3506 817 3564 843
rect 3606 877 3664 903
rect 3606 843 3618 877
rect 3652 843 3664 877
rect 3606 817 3664 843
rect 3706 877 3764 903
rect 3706 843 3718 877
rect 3752 843 3764 877
rect 3706 817 3764 843
rect 3806 877 3864 903
rect 3806 843 3818 877
rect 3852 843 3864 877
rect 3806 817 3864 843
rect 3906 877 3964 903
rect 3906 843 3918 877
rect 3952 843 3964 877
rect 3906 817 3964 843
rect 4006 877 4064 903
rect 4006 843 4018 877
rect 4052 843 4064 877
rect 4006 817 4064 843
rect 4106 877 4164 903
rect 4106 843 4118 877
rect 4152 843 4164 877
rect 4106 817 4164 843
rect 4206 877 4264 903
rect 4206 843 4218 877
rect 4252 843 4264 877
rect 4206 817 4264 843
rect 4306 877 4364 903
rect 4306 843 4312 877
rect 4352 843 4364 877
rect 4306 817 4364 843
rect 4406 877 4464 903
rect 4406 843 4418 877
rect 4458 843 4464 877
rect 4406 817 4464 843
rect 4506 877 4564 903
rect 4506 843 4512 877
rect 4552 843 4564 877
rect 4506 817 4564 843
rect 4606 877 4664 903
rect 4606 843 4618 877
rect 4658 843 4664 877
rect 4606 817 4664 843
rect 4706 877 4764 903
rect 4706 843 4718 877
rect 4752 843 4764 877
rect 4706 817 4764 843
rect 4806 877 4864 903
rect 4806 843 4818 877
rect 4852 843 4864 877
rect 4806 817 4864 843
rect 4906 877 4964 903
rect 4906 843 4918 877
rect 4952 843 4964 877
rect 4906 817 4964 843
rect 5006 877 5064 903
rect 5006 843 5018 877
rect 5052 843 5064 877
rect 5006 817 5064 843
rect 5106 877 5164 903
rect 5106 843 5118 877
rect 5152 843 5164 877
rect 5106 817 5164 843
rect 5206 877 5264 903
rect 5206 843 5218 877
rect 5252 843 5264 877
rect 5206 817 5264 843
rect 5306 877 5364 903
rect 5306 843 5318 877
rect 5352 843 5364 877
rect 5306 817 5364 843
rect 5406 877 5464 903
rect 5406 843 5418 877
rect 5452 843 5464 877
rect 5406 817 5464 843
rect 5506 877 5564 903
rect 5506 843 5518 877
rect 5552 843 5564 877
rect 5506 817 5564 843
rect 5606 877 5664 903
rect 5606 843 5618 877
rect 5652 843 5664 877
rect 5606 817 5664 843
rect 5706 877 5764 903
rect 5706 843 5718 877
rect 5752 843 5764 877
rect 5706 817 5764 843
rect 5806 877 5864 903
rect 5806 843 5818 877
rect 5852 843 5864 877
rect 5806 817 5864 843
rect 5906 877 5964 903
rect 5906 843 5918 877
rect 5952 843 5964 877
rect 5906 817 5964 843
rect 6006 877 6064 903
rect 6006 843 6018 877
rect 6052 843 6064 877
rect 6006 817 6064 843
rect 6106 877 6164 903
rect 6106 843 6118 877
rect 6152 843 6164 877
rect 6106 817 6164 843
rect 6206 877 6264 903
rect 6206 843 6218 877
rect 6252 843 6264 877
rect 6206 817 6264 843
rect 6306 877 6364 903
rect 6306 843 6318 877
rect 6352 843 6364 877
rect 6306 817 6364 843
rect 6406 877 6464 903
rect 6618 896 6862 930
rect 6406 843 6418 877
rect 6452 843 6464 877
rect 6508 858 6516 892
rect 6558 858 6574 892
rect 6618 877 6652 896
rect 6406 817 6464 843
rect 6828 893 6862 896
rect 6828 877 6962 893
rect 6618 827 6652 843
rect 6696 828 6712 862
rect 6754 828 6762 862
rect 6862 843 6928 877
rect 6828 827 6962 843
rect 7028 877 7062 893
rect 7028 827 7062 843
rect 7128 877 7362 893
rect 7162 843 7228 877
rect 7262 843 7328 877
rect 7128 827 7362 843
rect 7428 877 7462 893
rect 7428 827 7462 843
rect 6 737 64 763
rect 6 703 18 737
rect 58 703 64 737
rect 6 677 64 703
rect 106 737 164 763
rect 106 703 118 737
rect 152 703 164 737
rect 106 677 164 703
rect 206 737 264 763
rect 206 703 218 737
rect 252 703 264 737
rect 206 677 264 703
rect 306 737 364 763
rect 306 703 318 737
rect 352 703 364 737
rect 306 677 364 703
rect 406 737 464 763
rect 406 703 418 737
rect 452 703 464 737
rect 406 677 464 703
rect 506 737 564 763
rect 506 703 518 737
rect 552 703 564 737
rect 506 677 564 703
rect 606 737 664 763
rect 606 703 618 737
rect 652 703 664 737
rect 606 677 664 703
rect 706 737 764 763
rect 706 703 718 737
rect 752 703 764 737
rect 706 677 764 703
rect 806 737 864 763
rect 806 703 818 737
rect 852 703 864 737
rect 806 677 864 703
rect 906 737 964 763
rect 906 703 912 737
rect 952 703 964 737
rect 906 677 964 703
rect 1006 737 1064 763
rect 1006 703 1018 737
rect 1058 703 1064 737
rect 1006 677 1064 703
rect 1106 737 1164 763
rect 1106 703 1118 737
rect 1152 703 1164 737
rect 1106 677 1164 703
rect 1206 737 1264 763
rect 1206 703 1218 737
rect 1252 703 1264 737
rect 1206 677 1264 703
rect 1306 737 1364 763
rect 1306 703 1318 737
rect 1352 703 1364 737
rect 1306 677 1364 703
rect 1406 737 1464 763
rect 1406 703 1418 737
rect 1452 703 1464 737
rect 1406 677 1464 703
rect 1506 737 1564 763
rect 1506 703 1518 737
rect 1552 703 1564 737
rect 1506 677 1564 703
rect 1606 737 1664 763
rect 1606 703 1618 737
rect 1652 703 1664 737
rect 1606 677 1664 703
rect 1706 737 1764 763
rect 1706 703 1718 737
rect 1752 703 1764 737
rect 1706 677 1764 703
rect 1806 737 1864 763
rect 1806 703 1818 737
rect 1852 703 1864 737
rect 1806 677 1864 703
rect 1906 737 1964 763
rect 1906 703 1918 737
rect 1952 703 1964 737
rect 1906 677 1964 703
rect 2006 737 2064 763
rect 2006 703 2012 737
rect 2052 703 2064 737
rect 2006 677 2064 703
rect 2106 737 2164 763
rect 2106 703 2118 737
rect 2158 703 2164 737
rect 2106 677 2164 703
rect 2206 737 2264 763
rect 2206 703 2212 737
rect 2252 703 2264 737
rect 2206 677 2264 703
rect 2306 737 2364 763
rect 2306 703 2318 737
rect 2358 703 2364 737
rect 2306 677 2364 703
rect 2406 737 2464 763
rect 2406 703 2418 737
rect 2452 703 2464 737
rect 2406 677 2464 703
rect 2506 737 2564 763
rect 2506 703 2518 737
rect 2552 703 2564 737
rect 2506 677 2564 703
rect 2606 737 2664 763
rect 2606 703 2618 737
rect 2652 703 2664 737
rect 2606 677 2664 703
rect 2706 737 2764 763
rect 2706 703 2718 737
rect 2752 703 2764 737
rect 2706 677 2764 703
rect 2806 737 2864 763
rect 2806 703 2818 737
rect 2852 703 2864 737
rect 2806 677 2864 703
rect 2906 737 2964 763
rect 2906 703 2918 737
rect 2952 703 2964 737
rect 2906 677 2964 703
rect 3006 737 3064 763
rect 3006 703 3018 737
rect 3052 703 3064 737
rect 3006 677 3064 703
rect 3106 737 3164 763
rect 3106 703 3118 737
rect 3152 703 3164 737
rect 3106 677 3164 703
rect 3206 737 3264 763
rect 3206 703 3218 737
rect 3252 703 3264 737
rect 3206 677 3264 703
rect 3306 737 3364 763
rect 3306 703 3318 737
rect 3352 703 3364 737
rect 3306 677 3364 703
rect 3406 737 3464 763
rect 3406 703 3418 737
rect 3452 703 3464 737
rect 3406 677 3464 703
rect 3506 737 3564 763
rect 3506 703 3518 737
rect 3552 703 3564 737
rect 3506 677 3564 703
rect 3606 737 3664 763
rect 3606 703 3618 737
rect 3652 703 3664 737
rect 3606 677 3664 703
rect 3706 737 3764 763
rect 3706 703 3718 737
rect 3752 703 3764 737
rect 3706 677 3764 703
rect 3806 737 3864 763
rect 3806 703 3818 737
rect 3852 703 3864 737
rect 3806 677 3864 703
rect 3906 737 3964 763
rect 3906 703 3918 737
rect 3952 703 3964 737
rect 3906 677 3964 703
rect 4006 737 4064 763
rect 4006 703 4018 737
rect 4052 703 4064 737
rect 4006 677 4064 703
rect 4106 737 4164 763
rect 4106 703 4118 737
rect 4152 703 4164 737
rect 4106 677 4164 703
rect 4206 737 4264 763
rect 4206 703 4218 737
rect 4252 703 4264 737
rect 4206 677 4264 703
rect 4306 737 4364 763
rect 4306 703 4318 737
rect 4352 703 4364 737
rect 4306 677 4364 703
rect 4406 737 4464 763
rect 4406 703 4412 737
rect 4452 703 4464 737
rect 4406 677 4464 703
rect 4506 737 4564 763
rect 4506 703 4518 737
rect 4558 703 4564 737
rect 4506 677 4564 703
rect 4606 737 4664 763
rect 4606 703 4618 737
rect 4652 703 4664 737
rect 4606 677 4664 703
rect 4706 737 4764 763
rect 4706 703 4718 737
rect 4752 703 4764 737
rect 4706 677 4764 703
rect 4806 737 4864 763
rect 4806 703 4818 737
rect 4852 703 4864 737
rect 4806 677 4864 703
rect 4906 737 4964 763
rect 4906 703 4918 737
rect 4952 703 4964 737
rect 4906 677 4964 703
rect 5006 737 5064 763
rect 5006 703 5018 737
rect 5052 703 5064 737
rect 5006 677 5064 703
rect 5106 737 5164 763
rect 5106 703 5118 737
rect 5152 703 5164 737
rect 5106 677 5164 703
rect 5206 737 5264 763
rect 5206 703 5218 737
rect 5252 703 5264 737
rect 5206 677 5264 703
rect 5306 737 5364 763
rect 5306 703 5318 737
rect 5352 703 5364 737
rect 5306 677 5364 703
rect 5406 737 5464 763
rect 5406 703 5418 737
rect 5452 703 5464 737
rect 5406 677 5464 703
rect 5506 737 5564 763
rect 5506 703 5512 737
rect 5552 703 5564 737
rect 5506 677 5564 703
rect 5606 737 5664 763
rect 5606 703 5618 737
rect 5658 703 5664 737
rect 5606 677 5664 703
rect 5706 737 5764 763
rect 5706 703 5712 737
rect 5752 703 5764 737
rect 5706 677 5764 703
rect 5806 737 5864 763
rect 5806 703 5818 737
rect 5858 703 5864 737
rect 5806 677 5864 703
rect 5906 737 5964 763
rect 5906 703 5918 737
rect 5952 703 5964 737
rect 5906 677 5964 703
rect 6006 737 6064 763
rect 6006 703 6018 737
rect 6052 703 6064 737
rect 6006 677 6064 703
rect 6106 737 6164 763
rect 6106 703 6118 737
rect 6152 703 6164 737
rect 6106 677 6164 703
rect 6206 737 6264 763
rect 6206 703 6218 737
rect 6252 703 6264 737
rect 6206 677 6264 703
rect 6306 737 6364 763
rect 6306 703 6318 737
rect 6352 703 6364 737
rect 6306 677 6364 703
rect 6406 737 6464 763
rect 6618 756 6862 790
rect 6406 703 6418 737
rect 6452 703 6464 737
rect 6508 718 6516 752
rect 6558 718 6574 752
rect 6618 737 6652 756
rect 6406 677 6464 703
rect 6828 737 6862 756
rect 6618 687 6652 703
rect 6696 688 6712 722
rect 6754 688 6762 722
rect 6828 687 6862 703
rect 6928 737 7062 753
rect 6962 703 7028 737
rect 6928 687 7062 703
rect 7128 737 7362 753
rect 7162 703 7228 737
rect 7262 703 7328 737
rect 7128 687 7362 703
rect 7428 737 7462 753
rect 7428 687 7462 703
rect 6 597 64 623
rect 6 563 18 597
rect 52 563 64 597
rect 6 537 64 563
rect 106 597 164 623
rect 106 563 118 597
rect 152 563 164 597
rect 106 537 164 563
rect 206 597 264 623
rect 206 563 218 597
rect 252 563 264 597
rect 206 537 264 563
rect 306 597 364 623
rect 306 563 318 597
rect 352 563 364 597
rect 306 537 364 563
rect 406 597 464 623
rect 406 563 418 597
rect 452 563 464 597
rect 406 537 464 563
rect 506 597 564 623
rect 506 563 512 597
rect 552 563 564 597
rect 506 537 564 563
rect 606 597 664 623
rect 606 563 618 597
rect 658 563 664 597
rect 606 537 664 563
rect 706 597 764 623
rect 706 563 718 597
rect 752 563 764 597
rect 706 537 764 563
rect 806 597 864 623
rect 806 563 818 597
rect 852 563 864 597
rect 806 537 864 563
rect 906 597 964 623
rect 906 563 918 597
rect 952 563 964 597
rect 906 537 964 563
rect 1006 597 1064 623
rect 1006 563 1012 597
rect 1052 563 1064 597
rect 1006 537 1064 563
rect 1106 597 1164 623
rect 1106 563 1118 597
rect 1158 563 1164 597
rect 1106 537 1164 563
rect 1206 597 1264 623
rect 1206 563 1218 597
rect 1252 563 1264 597
rect 1206 537 1264 563
rect 1306 597 1364 623
rect 1306 563 1318 597
rect 1352 563 1364 597
rect 1306 537 1364 563
rect 1406 597 1464 623
rect 1406 563 1418 597
rect 1452 563 1464 597
rect 1406 537 1464 563
rect 1506 597 1564 623
rect 1506 563 1518 597
rect 1552 563 1564 597
rect 1506 537 1564 563
rect 1606 597 1664 623
rect 1606 563 1618 597
rect 1652 563 1664 597
rect 1606 537 1664 563
rect 1706 597 1764 623
rect 1706 563 1718 597
rect 1752 563 1764 597
rect 1706 537 1764 563
rect 1806 597 1864 623
rect 1806 563 1818 597
rect 1852 563 1864 597
rect 1806 537 1864 563
rect 1906 597 1964 623
rect 1906 563 1918 597
rect 1952 563 1964 597
rect 1906 537 1964 563
rect 2006 597 2064 623
rect 2006 563 2018 597
rect 2052 563 2064 597
rect 2006 537 2064 563
rect 2106 597 2164 623
rect 2106 563 2118 597
rect 2152 563 2164 597
rect 2106 537 2164 563
rect 2206 597 2264 623
rect 2206 563 2218 597
rect 2252 563 2264 597
rect 2206 537 2264 563
rect 2306 597 2364 623
rect 2306 563 2318 597
rect 2352 563 2364 597
rect 2306 537 2364 563
rect 2406 597 2464 623
rect 2406 563 2418 597
rect 2452 563 2464 597
rect 2406 537 2464 563
rect 2506 597 2564 623
rect 2506 563 2518 597
rect 2552 563 2564 597
rect 2506 537 2564 563
rect 2606 597 2664 623
rect 2606 563 2618 597
rect 2652 563 2664 597
rect 2606 537 2664 563
rect 2706 597 2764 623
rect 2706 563 2718 597
rect 2752 563 2764 597
rect 2706 537 2764 563
rect 2806 597 2864 623
rect 2806 563 2818 597
rect 2852 563 2864 597
rect 2806 537 2864 563
rect 2906 597 2964 623
rect 2906 563 2918 597
rect 2952 563 2964 597
rect 2906 537 2964 563
rect 3006 597 3064 623
rect 3006 563 3018 597
rect 3052 563 3064 597
rect 3006 537 3064 563
rect 3106 597 3164 623
rect 3106 563 3118 597
rect 3152 563 3164 597
rect 3106 537 3164 563
rect 3206 597 3264 623
rect 3206 563 3218 597
rect 3252 563 3264 597
rect 3206 537 3264 563
rect 3306 597 3364 623
rect 3306 563 3318 597
rect 3352 563 3364 597
rect 3306 537 3364 563
rect 3406 597 3464 623
rect 3406 563 3418 597
rect 3452 563 3464 597
rect 3406 537 3464 563
rect 3506 597 3564 623
rect 3506 563 3518 597
rect 3552 563 3564 597
rect 3506 537 3564 563
rect 3606 597 3664 623
rect 3606 563 3618 597
rect 3652 563 3664 597
rect 3606 537 3664 563
rect 3706 597 3764 623
rect 3706 563 3712 597
rect 3752 563 3764 597
rect 3706 537 3764 563
rect 3806 597 3864 623
rect 3806 563 3818 597
rect 3858 563 3864 597
rect 3806 537 3864 563
rect 3906 597 3964 623
rect 3906 563 3918 597
rect 3952 563 3964 597
rect 3906 537 3964 563
rect 4006 597 4064 623
rect 4006 563 4012 597
rect 4052 563 4064 597
rect 4006 537 4064 563
rect 4106 597 4164 623
rect 4106 563 4118 597
rect 4158 563 4164 597
rect 4106 537 4164 563
rect 4206 597 4264 623
rect 4206 563 4212 597
rect 4252 563 4264 597
rect 4206 537 4264 563
rect 4306 597 4364 623
rect 4306 563 4318 597
rect 4358 563 4364 597
rect 4306 537 4364 563
rect 4406 597 4464 623
rect 4406 563 4418 597
rect 4452 563 4464 597
rect 4406 537 4464 563
rect 4506 597 4564 623
rect 4506 563 4518 597
rect 4552 563 4564 597
rect 4506 537 4564 563
rect 4606 597 4664 623
rect 4606 563 4612 597
rect 4652 563 4664 597
rect 4606 537 4664 563
rect 4706 597 4764 623
rect 4706 563 4718 597
rect 4758 563 4764 597
rect 4706 537 4764 563
rect 4806 597 4864 623
rect 4806 563 4818 597
rect 4852 563 4864 597
rect 4806 537 4864 563
rect 4906 597 4964 623
rect 4906 563 4918 597
rect 4952 563 4964 597
rect 4906 537 4964 563
rect 5006 597 5064 623
rect 5006 563 5018 597
rect 5052 563 5064 597
rect 5006 537 5064 563
rect 5106 597 5164 623
rect 5106 563 5118 597
rect 5152 563 5164 597
rect 5106 537 5164 563
rect 5206 597 5264 623
rect 5206 563 5212 597
rect 5252 563 5264 597
rect 5206 537 5264 563
rect 5306 597 5364 623
rect 5306 563 5318 597
rect 5358 563 5364 597
rect 5306 537 5364 563
rect 5406 597 5464 623
rect 5406 563 5418 597
rect 5452 563 5464 597
rect 5406 537 5464 563
rect 5506 597 5564 623
rect 5506 563 5518 597
rect 5552 563 5564 597
rect 5506 537 5564 563
rect 5606 597 5664 623
rect 5606 563 5618 597
rect 5652 563 5664 597
rect 5606 537 5664 563
rect 5706 597 5764 623
rect 5706 563 5718 597
rect 5752 563 5764 597
rect 5706 537 5764 563
rect 5806 597 5864 623
rect 5806 563 5818 597
rect 5852 563 5864 597
rect 5806 537 5864 563
rect 5906 597 5964 623
rect 5906 563 5918 597
rect 5952 563 5964 597
rect 5906 537 5964 563
rect 6006 597 6064 623
rect 6006 563 6012 597
rect 6052 563 6064 597
rect 6006 537 6064 563
rect 6106 597 6164 623
rect 6106 563 6118 597
rect 6158 563 6164 597
rect 6106 537 6164 563
rect 6206 597 6264 623
rect 6206 563 6218 597
rect 6252 563 6264 597
rect 6206 537 6264 563
rect 6306 597 6364 623
rect 6306 563 6318 597
rect 6352 563 6364 597
rect 6306 537 6364 563
rect 6406 597 6464 623
rect 6618 616 6862 650
rect 6406 563 6412 597
rect 6452 563 6464 597
rect 6508 578 6516 612
rect 6558 578 6574 612
rect 6618 597 6652 616
rect 6406 537 6464 563
rect 6828 613 6862 616
rect 6828 597 6962 613
rect 6618 547 6652 563
rect 6696 548 6712 582
rect 6754 548 6762 582
rect 6862 563 6928 597
rect 6828 547 6962 563
rect 7028 597 7162 613
rect 7062 563 7128 597
rect 7028 547 7162 563
rect 7228 597 7262 613
rect 7228 547 7262 563
rect 7328 597 7462 613
rect 7362 563 7428 597
rect 7328 547 7462 563
rect 6 457 64 483
rect 6 423 18 457
rect 52 423 64 457
rect 6 397 64 423
rect 106 457 164 483
rect 106 423 118 457
rect 152 423 164 457
rect 106 397 164 423
rect 206 457 264 483
rect 206 423 212 457
rect 252 423 264 457
rect 206 397 264 423
rect 306 457 364 483
rect 306 423 318 457
rect 358 423 364 457
rect 306 397 364 423
rect 406 457 464 483
rect 406 423 412 457
rect 452 423 464 457
rect 406 397 464 423
rect 506 457 564 483
rect 506 423 518 457
rect 558 423 564 457
rect 506 397 564 423
rect 606 457 664 483
rect 606 423 618 457
rect 652 423 664 457
rect 606 397 664 423
rect 706 457 764 483
rect 706 423 718 457
rect 752 423 764 457
rect 706 397 764 423
rect 806 457 864 483
rect 806 423 818 457
rect 852 423 864 457
rect 806 397 864 423
rect 906 457 964 483
rect 906 423 918 457
rect 952 423 964 457
rect 906 397 964 423
rect 1006 457 1064 483
rect 1006 423 1018 457
rect 1052 423 1064 457
rect 1006 397 1064 423
rect 1106 457 1164 483
rect 1106 423 1118 457
rect 1152 423 1164 457
rect 1106 397 1164 423
rect 1206 457 1264 483
rect 1206 423 1218 457
rect 1252 423 1264 457
rect 1206 397 1264 423
rect 1306 457 1364 483
rect 1306 423 1318 457
rect 1352 423 1364 457
rect 1306 397 1364 423
rect 1406 457 1464 483
rect 1406 423 1412 457
rect 1452 423 1464 457
rect 1406 397 1464 423
rect 1506 457 1564 483
rect 1506 423 1518 457
rect 1558 423 1564 457
rect 1506 397 1564 423
rect 1606 457 1664 483
rect 1606 423 1618 457
rect 1652 423 1664 457
rect 1606 397 1664 423
rect 1706 457 1764 483
rect 1706 423 1718 457
rect 1752 423 1764 457
rect 1706 397 1764 423
rect 1806 457 1864 483
rect 1806 423 1818 457
rect 1852 423 1864 457
rect 1806 397 1864 423
rect 1906 457 1964 483
rect 1906 423 1918 457
rect 1952 423 1964 457
rect 1906 397 1964 423
rect 2006 457 2064 483
rect 2006 423 2018 457
rect 2052 423 2064 457
rect 2006 397 2064 423
rect 2106 457 2164 483
rect 2106 423 2118 457
rect 2152 423 2164 457
rect 2106 397 2164 423
rect 2206 457 2264 483
rect 2206 423 2218 457
rect 2252 423 2264 457
rect 2206 397 2264 423
rect 2306 457 2364 483
rect 2306 423 2318 457
rect 2352 423 2364 457
rect 2306 397 2364 423
rect 2406 457 2464 483
rect 2406 423 2418 457
rect 2452 423 2464 457
rect 2406 397 2464 423
rect 2506 457 2564 483
rect 2506 423 2518 457
rect 2552 423 2564 457
rect 2506 397 2564 423
rect 2606 457 2664 483
rect 2606 423 2618 457
rect 2652 423 2664 457
rect 2606 397 2664 423
rect 2706 457 2764 483
rect 2706 423 2718 457
rect 2752 423 2764 457
rect 2706 397 2764 423
rect 2806 457 2864 483
rect 2806 423 2818 457
rect 2852 423 2864 457
rect 2806 397 2864 423
rect 2906 457 2964 483
rect 2906 423 2918 457
rect 2952 423 2964 457
rect 2906 397 2964 423
rect 3006 457 3064 483
rect 3006 423 3012 457
rect 3052 423 3064 457
rect 3006 397 3064 423
rect 3106 457 3164 483
rect 3106 423 3118 457
rect 3158 423 3164 457
rect 3106 397 3164 423
rect 3206 457 3264 483
rect 3206 423 3212 457
rect 3252 423 3264 457
rect 3206 397 3264 423
rect 3306 457 3364 483
rect 3306 423 3318 457
rect 3358 423 3364 457
rect 3306 397 3364 423
rect 3406 457 3464 483
rect 3406 423 3418 457
rect 3452 423 3464 457
rect 3406 397 3464 423
rect 3506 457 3564 483
rect 3506 423 3512 457
rect 3552 423 3564 457
rect 3506 397 3564 423
rect 3606 457 3664 483
rect 3606 423 3618 457
rect 3658 423 3664 457
rect 3606 397 3664 423
rect 3706 457 3764 483
rect 3706 423 3712 457
rect 3752 423 3764 457
rect 3706 397 3764 423
rect 3806 457 3864 483
rect 3806 423 3818 457
rect 3858 423 3864 457
rect 3806 397 3864 423
rect 3906 457 3964 483
rect 3906 423 3918 457
rect 3952 423 3964 457
rect 3906 397 3964 423
rect 4006 457 4064 483
rect 4006 423 4018 457
rect 4052 423 4064 457
rect 4006 397 4064 423
rect 4106 457 4164 483
rect 4106 423 4118 457
rect 4152 423 4164 457
rect 4106 397 4164 423
rect 4206 457 4264 483
rect 4206 423 4218 457
rect 4252 423 4264 457
rect 4206 397 4264 423
rect 4306 457 4364 483
rect 4306 423 4318 457
rect 4352 423 4364 457
rect 4306 397 4364 423
rect 4406 457 4464 483
rect 4406 423 4418 457
rect 4452 423 4464 457
rect 4406 397 4464 423
rect 4506 457 4564 483
rect 4506 423 4518 457
rect 4552 423 4564 457
rect 4506 397 4564 423
rect 4606 457 4664 483
rect 4606 423 4618 457
rect 4652 423 4664 457
rect 4606 397 4664 423
rect 4706 457 4764 483
rect 4706 423 4718 457
rect 4752 423 4764 457
rect 4706 397 4764 423
rect 4806 457 4864 483
rect 4806 423 4818 457
rect 4852 423 4864 457
rect 4806 397 4864 423
rect 4906 457 4964 483
rect 4906 423 4918 457
rect 4952 423 4964 457
rect 4906 397 4964 423
rect 5006 457 5064 483
rect 5006 423 5018 457
rect 5052 423 5064 457
rect 5006 397 5064 423
rect 5106 457 5164 483
rect 5106 423 5118 457
rect 5152 423 5164 457
rect 5106 397 5164 423
rect 5206 457 5264 483
rect 5206 423 5218 457
rect 5252 423 5264 457
rect 5206 397 5264 423
rect 5306 457 5364 483
rect 5306 423 5318 457
rect 5352 423 5364 457
rect 5306 397 5364 423
rect 5406 457 5464 483
rect 5406 423 5418 457
rect 5452 423 5464 457
rect 5406 397 5464 423
rect 5506 457 5564 483
rect 5506 423 5512 457
rect 5552 423 5564 457
rect 5506 397 5564 423
rect 5606 457 5664 483
rect 5606 423 5618 457
rect 5658 423 5664 457
rect 5606 397 5664 423
rect 5706 457 5764 483
rect 5706 423 5718 457
rect 5752 423 5764 457
rect 5706 397 5764 423
rect 5806 457 5864 483
rect 5806 423 5818 457
rect 5852 423 5864 457
rect 5806 397 5864 423
rect 5906 457 5964 483
rect 5906 423 5918 457
rect 5952 423 5964 457
rect 5906 397 5964 423
rect 6006 457 6064 483
rect 6006 423 6018 457
rect 6052 423 6064 457
rect 6006 397 6064 423
rect 6106 457 6164 483
rect 6106 423 6118 457
rect 6152 423 6164 457
rect 6106 397 6164 423
rect 6206 457 6264 483
rect 6206 423 6212 457
rect 6252 423 6264 457
rect 6206 397 6264 423
rect 6306 457 6364 483
rect 6306 423 6318 457
rect 6358 423 6364 457
rect 6306 397 6364 423
rect 6406 457 6464 483
rect 6618 476 6862 510
rect 6406 423 6412 457
rect 6452 423 6464 457
rect 6508 438 6516 472
rect 6558 438 6574 472
rect 6618 457 6652 476
rect 6406 397 6464 423
rect 6828 457 6862 476
rect 6618 407 6652 423
rect 6696 408 6712 442
rect 6754 408 6762 442
rect 6828 407 6862 423
rect 6928 457 7162 473
rect 6962 423 7028 457
rect 7062 423 7128 457
rect 6928 407 7162 423
rect 7228 457 7262 473
rect 7228 407 7262 423
rect 7328 457 7462 473
rect 7362 423 7428 457
rect 7328 407 7462 423
rect 6 317 64 343
rect 6 283 18 317
rect 52 283 64 317
rect 6 257 64 283
rect 106 317 164 343
rect 106 283 118 317
rect 152 283 164 317
rect 106 257 164 283
rect 206 317 264 343
rect 206 283 218 317
rect 252 283 264 317
rect 206 257 264 283
rect 306 317 364 343
rect 306 283 318 317
rect 352 283 364 317
rect 306 257 364 283
rect 406 317 464 343
rect 406 283 418 317
rect 452 283 464 317
rect 406 257 464 283
rect 506 317 564 343
rect 506 283 518 317
rect 552 283 564 317
rect 506 257 564 283
rect 606 317 664 343
rect 606 283 612 317
rect 652 283 664 317
rect 606 257 664 283
rect 706 317 764 343
rect 706 283 718 317
rect 758 283 764 317
rect 706 257 764 283
rect 806 317 864 343
rect 806 283 818 317
rect 852 283 864 317
rect 806 257 864 283
rect 906 317 964 343
rect 906 283 918 317
rect 952 283 964 317
rect 906 257 964 283
rect 1006 317 1064 343
rect 1006 283 1018 317
rect 1052 283 1064 317
rect 1006 257 1064 283
rect 1106 317 1164 343
rect 1106 283 1118 317
rect 1152 283 1164 317
rect 1106 257 1164 283
rect 1206 317 1264 343
rect 1206 283 1218 317
rect 1252 283 1264 317
rect 1206 257 1264 283
rect 1306 317 1364 343
rect 1306 283 1318 317
rect 1352 283 1364 317
rect 1306 257 1364 283
rect 1406 317 1464 343
rect 1406 283 1418 317
rect 1452 283 1464 317
rect 1406 257 1464 283
rect 1506 317 1564 343
rect 1506 283 1512 317
rect 1552 283 1564 317
rect 1506 257 1564 283
rect 1606 317 1664 343
rect 1606 283 1618 317
rect 1658 283 1664 317
rect 1606 257 1664 283
rect 1706 317 1764 343
rect 1706 283 1718 317
rect 1752 283 1764 317
rect 1706 257 1764 283
rect 1806 317 1864 343
rect 1806 283 1818 317
rect 1852 283 1864 317
rect 1806 257 1864 283
rect 1906 317 1964 343
rect 1906 283 1918 317
rect 1952 283 1964 317
rect 1906 257 1964 283
rect 2006 317 2064 343
rect 2006 283 2018 317
rect 2052 283 2064 317
rect 2006 257 2064 283
rect 2106 317 2164 343
rect 2106 283 2118 317
rect 2152 283 2164 317
rect 2106 257 2164 283
rect 2206 317 2264 343
rect 2206 283 2212 317
rect 2252 283 2264 317
rect 2206 257 2264 283
rect 2306 317 2364 343
rect 2306 283 2318 317
rect 2358 283 2364 317
rect 2306 257 2364 283
rect 2406 317 2464 343
rect 2406 283 2412 317
rect 2452 283 2464 317
rect 2406 257 2464 283
rect 2506 317 2564 343
rect 2506 283 2518 317
rect 2558 283 2564 317
rect 2506 257 2564 283
rect 2606 317 2664 343
rect 2606 283 2612 317
rect 2652 283 2664 317
rect 2606 257 2664 283
rect 2706 317 2764 343
rect 2706 283 2718 317
rect 2758 283 2764 317
rect 2706 257 2764 283
rect 2806 317 2864 343
rect 2806 283 2812 317
rect 2852 283 2864 317
rect 2806 257 2864 283
rect 2906 317 2964 343
rect 2906 283 2918 317
rect 2958 283 2964 317
rect 2906 257 2964 283
rect 3006 317 3064 343
rect 3006 283 3018 317
rect 3052 283 3064 317
rect 3006 257 3064 283
rect 3106 317 3164 343
rect 3106 283 3118 317
rect 3152 283 3164 317
rect 3106 257 3164 283
rect 3206 317 3264 343
rect 3206 283 3218 317
rect 3252 283 3264 317
rect 3206 257 3264 283
rect 3306 317 3364 343
rect 3306 283 3318 317
rect 3352 283 3364 317
rect 3306 257 3364 283
rect 3406 317 3464 343
rect 3406 283 3418 317
rect 3452 283 3464 317
rect 3406 257 3464 283
rect 3506 317 3564 343
rect 3506 283 3512 317
rect 3552 283 3564 317
rect 3506 257 3564 283
rect 3606 317 3664 343
rect 3606 283 3618 317
rect 3658 283 3664 317
rect 3606 257 3664 283
rect 3706 317 3764 343
rect 3706 283 3718 317
rect 3752 283 3764 317
rect 3706 257 3764 283
rect 3806 317 3864 343
rect 3806 283 3818 317
rect 3852 283 3864 317
rect 3806 257 3864 283
rect 3906 317 3964 343
rect 3906 283 3918 317
rect 3952 283 3964 317
rect 3906 257 3964 283
rect 4006 317 4064 343
rect 4006 283 4018 317
rect 4052 283 4064 317
rect 4006 257 4064 283
rect 4106 317 4164 343
rect 4106 283 4118 317
rect 4152 283 4164 317
rect 4106 257 4164 283
rect 4206 317 4264 343
rect 4206 283 4218 317
rect 4252 283 4264 317
rect 4206 257 4264 283
rect 4306 317 4364 343
rect 4306 283 4318 317
rect 4352 283 4364 317
rect 4306 257 4364 283
rect 4406 317 4464 343
rect 4406 283 4418 317
rect 4452 283 4464 317
rect 4406 257 4464 283
rect 4506 317 4564 343
rect 4506 283 4518 317
rect 4552 283 4564 317
rect 4506 257 4564 283
rect 4606 317 4664 343
rect 4606 283 4618 317
rect 4652 283 4664 317
rect 4606 257 4664 283
rect 4706 317 4764 343
rect 4706 283 4718 317
rect 4752 283 4764 317
rect 4706 257 4764 283
rect 4806 317 4864 343
rect 4806 283 4818 317
rect 4852 283 4864 317
rect 4806 257 4864 283
rect 4906 317 4964 343
rect 4906 283 4918 317
rect 4952 283 4964 317
rect 4906 257 4964 283
rect 5006 317 5064 343
rect 5006 283 5018 317
rect 5052 283 5064 317
rect 5006 257 5064 283
rect 5106 317 5164 343
rect 5106 283 5118 317
rect 5152 283 5164 317
rect 5106 257 5164 283
rect 5206 317 5264 343
rect 5206 283 5218 317
rect 5252 283 5264 317
rect 5206 257 5264 283
rect 5306 317 5364 343
rect 5306 283 5318 317
rect 5352 283 5364 317
rect 5306 257 5364 283
rect 5406 317 5464 343
rect 5406 283 5418 317
rect 5452 283 5464 317
rect 5406 257 5464 283
rect 5506 317 5564 343
rect 5506 283 5518 317
rect 5552 283 5564 317
rect 5506 257 5564 283
rect 5606 317 5664 343
rect 5606 283 5612 317
rect 5652 283 5664 317
rect 5606 257 5664 283
rect 5706 317 5764 343
rect 5706 283 5718 317
rect 5758 283 5764 317
rect 5706 257 5764 283
rect 5806 317 5864 343
rect 5806 283 5818 317
rect 5852 283 5864 317
rect 5806 257 5864 283
rect 5906 317 5964 343
rect 5906 283 5918 317
rect 5952 283 5964 317
rect 5906 257 5964 283
rect 6006 317 6064 343
rect 6006 283 6018 317
rect 6052 283 6064 317
rect 6006 257 6064 283
rect 6106 317 6164 343
rect 6106 283 6118 317
rect 6152 283 6164 317
rect 6106 257 6164 283
rect 6206 317 6264 343
rect 6206 283 6218 317
rect 6252 283 6264 317
rect 6206 257 6264 283
rect 6306 317 6364 343
rect 6306 283 6318 317
rect 6352 283 6364 317
rect 6306 257 6364 283
rect 6406 317 6464 343
rect 6618 336 6862 370
rect 6406 283 6412 317
rect 6452 283 6464 317
rect 6508 298 6516 332
rect 6558 298 6574 332
rect 6618 317 6652 336
rect 6406 257 6464 283
rect 6828 333 6862 336
rect 6828 317 6962 333
rect 6618 267 6652 283
rect 6696 268 6712 302
rect 6754 268 6762 302
rect 6862 283 6928 317
rect 6828 267 6962 283
rect 7028 317 7062 333
rect 7028 267 7062 283
rect 7128 317 7262 333
rect 7162 283 7228 317
rect 7128 267 7262 283
rect 7328 317 7462 333
rect 7362 283 7428 317
rect 7328 267 7462 283
rect 6 177 64 203
rect 6 143 18 177
rect 58 143 64 177
rect 6 117 64 143
rect 106 177 164 203
rect 106 143 118 177
rect 152 143 164 177
rect 106 117 164 143
rect 206 177 264 203
rect 206 143 218 177
rect 252 143 264 177
rect 206 117 264 143
rect 306 177 364 203
rect 306 143 318 177
rect 352 143 364 177
rect 306 117 364 143
rect 406 177 464 203
rect 406 143 418 177
rect 452 143 464 177
rect 406 117 464 143
rect 506 177 564 203
rect 506 143 518 177
rect 552 143 564 177
rect 506 117 564 143
rect 606 177 664 203
rect 606 143 618 177
rect 652 143 664 177
rect 606 117 664 143
rect 706 177 764 203
rect 706 143 718 177
rect 752 143 764 177
rect 706 117 764 143
rect 806 177 864 203
rect 806 143 812 177
rect 852 143 864 177
rect 806 117 864 143
rect 906 177 964 203
rect 906 143 918 177
rect 958 143 964 177
rect 906 117 964 143
rect 1006 177 1064 203
rect 1006 143 1018 177
rect 1052 143 1064 177
rect 1006 117 1064 143
rect 1106 177 1164 203
rect 1106 143 1118 177
rect 1152 143 1164 177
rect 1106 117 1164 143
rect 1206 177 1264 203
rect 1206 143 1218 177
rect 1252 143 1264 177
rect 1206 117 1264 143
rect 1306 177 1364 203
rect 1306 143 1318 177
rect 1352 143 1364 177
rect 1306 117 1364 143
rect 1406 177 1464 203
rect 1406 143 1418 177
rect 1452 143 1464 177
rect 1406 117 1464 143
rect 1506 177 1564 203
rect 1506 143 1518 177
rect 1552 143 1564 177
rect 1506 117 1564 143
rect 1606 177 1664 203
rect 1606 143 1618 177
rect 1652 143 1664 177
rect 1606 117 1664 143
rect 1706 177 1764 203
rect 1706 143 1718 177
rect 1752 143 1764 177
rect 1706 117 1764 143
rect 1806 177 1864 203
rect 1806 143 1818 177
rect 1852 143 1864 177
rect 1806 117 1864 143
rect 1906 177 1964 203
rect 1906 143 1912 177
rect 1952 143 1964 177
rect 1906 117 1964 143
rect 2006 177 2064 203
rect 2006 143 2018 177
rect 2058 143 2064 177
rect 2006 117 2064 143
rect 2106 177 2164 203
rect 2106 143 2118 177
rect 2152 143 2164 177
rect 2106 117 2164 143
rect 2206 177 2264 203
rect 2206 143 2218 177
rect 2252 143 2264 177
rect 2206 117 2264 143
rect 2306 177 2364 203
rect 2306 143 2318 177
rect 2352 143 2364 177
rect 2306 117 2364 143
rect 2406 177 2464 203
rect 2406 143 2418 177
rect 2452 143 2464 177
rect 2406 117 2464 143
rect 2506 177 2564 203
rect 2506 143 2518 177
rect 2552 143 2564 177
rect 2506 117 2564 143
rect 2606 177 2664 203
rect 2606 143 2618 177
rect 2652 143 2664 177
rect 2606 117 2664 143
rect 2706 177 2764 203
rect 2706 143 2718 177
rect 2752 143 2764 177
rect 2706 117 2764 143
rect 2806 177 2864 203
rect 2806 143 2818 177
rect 2852 143 2864 177
rect 2806 117 2864 143
rect 2906 177 2964 203
rect 2906 143 2918 177
rect 2952 143 2964 177
rect 2906 117 2964 143
rect 3006 177 3064 203
rect 3006 143 3018 177
rect 3052 143 3064 177
rect 3006 117 3064 143
rect 3106 177 3164 203
rect 3106 143 3118 177
rect 3152 143 3164 177
rect 3106 117 3164 143
rect 3206 177 3264 203
rect 3206 143 3218 177
rect 3252 143 3264 177
rect 3206 117 3264 143
rect 3306 177 3364 203
rect 3306 143 3318 177
rect 3352 143 3364 177
rect 3306 117 3364 143
rect 3406 177 3464 203
rect 3406 143 3418 177
rect 3452 143 3464 177
rect 3406 117 3464 143
rect 3506 177 3564 203
rect 3506 143 3512 177
rect 3552 143 3564 177
rect 3506 117 3564 143
rect 3606 177 3664 203
rect 3606 143 3618 177
rect 3658 143 3664 177
rect 3606 117 3664 143
rect 3706 177 3764 203
rect 3706 143 3718 177
rect 3752 143 3764 177
rect 3706 117 3764 143
rect 3806 177 3864 203
rect 3806 143 3818 177
rect 3852 143 3864 177
rect 3806 117 3864 143
rect 3906 177 3964 203
rect 3906 143 3918 177
rect 3952 143 3964 177
rect 3906 117 3964 143
rect 4006 177 4064 203
rect 4006 143 4018 177
rect 4052 143 4064 177
rect 4006 117 4064 143
rect 4106 177 4164 203
rect 4106 143 4118 177
rect 4152 143 4164 177
rect 4106 117 4164 143
rect 4206 177 4264 203
rect 4206 143 4218 177
rect 4252 143 4264 177
rect 4206 117 4264 143
rect 4306 177 4364 203
rect 4306 143 4318 177
rect 4352 143 4364 177
rect 4306 117 4364 143
rect 4406 177 4464 203
rect 4406 143 4418 177
rect 4452 143 4464 177
rect 4406 117 4464 143
rect 4506 177 4564 203
rect 4506 143 4518 177
rect 4552 143 4564 177
rect 4506 117 4564 143
rect 4606 177 4664 203
rect 4606 143 4618 177
rect 4652 143 4664 177
rect 4606 117 4664 143
rect 4706 177 4764 203
rect 4706 143 4712 177
rect 4752 143 4764 177
rect 4706 117 4764 143
rect 4806 177 4864 203
rect 4806 143 4818 177
rect 4858 143 4864 177
rect 4806 117 4864 143
rect 4906 177 4964 203
rect 4906 143 4918 177
rect 4952 143 4964 177
rect 4906 117 4964 143
rect 5006 177 5064 203
rect 5006 143 5018 177
rect 5052 143 5064 177
rect 5006 117 5064 143
rect 5106 177 5164 203
rect 5106 143 5118 177
rect 5152 143 5164 177
rect 5106 117 5164 143
rect 5206 177 5264 203
rect 5206 143 5218 177
rect 5252 143 5264 177
rect 5206 117 5264 143
rect 5306 177 5364 203
rect 5306 143 5318 177
rect 5352 143 5364 177
rect 5306 117 5364 143
rect 5406 177 5464 203
rect 5406 143 5418 177
rect 5452 143 5464 177
rect 5406 117 5464 143
rect 5506 177 5564 203
rect 5506 143 5518 177
rect 5552 143 5564 177
rect 5506 117 5564 143
rect 5606 177 5664 203
rect 5606 143 5618 177
rect 5652 143 5664 177
rect 5606 117 5664 143
rect 5706 177 5764 203
rect 5706 143 5718 177
rect 5752 143 5764 177
rect 5706 117 5764 143
rect 5806 177 5864 203
rect 5806 143 5818 177
rect 5852 143 5864 177
rect 5806 117 5864 143
rect 5906 177 5964 203
rect 5906 143 5918 177
rect 5952 143 5964 177
rect 5906 117 5964 143
rect 6006 177 6064 203
rect 6006 143 6018 177
rect 6052 143 6064 177
rect 6006 117 6064 143
rect 6106 177 6164 203
rect 6106 143 6112 177
rect 6152 143 6164 177
rect 6106 117 6164 143
rect 6206 177 6264 203
rect 6206 143 6218 177
rect 6258 143 6264 177
rect 6206 117 6264 143
rect 6306 177 6364 203
rect 6306 143 6318 177
rect 6352 143 6364 177
rect 6306 117 6364 143
rect 6406 177 6464 203
rect 6618 196 6862 230
rect 6406 143 6412 177
rect 6452 143 6464 177
rect 6508 158 6516 192
rect 6558 158 6574 192
rect 6618 177 6652 196
rect 6406 117 6464 143
rect 6828 177 6862 196
rect 6618 127 6652 143
rect 6696 128 6712 162
rect 6754 128 6762 162
rect 6828 127 6862 143
rect 6928 177 7062 193
rect 6962 143 7028 177
rect 6928 127 7062 143
rect 7128 177 7262 193
rect 7162 143 7228 177
rect 7128 127 7262 143
rect 7328 177 7462 193
rect 7362 143 7428 177
rect 7328 127 7462 143
rect 8 20 18 54
rect 52 20 118 54
rect 152 20 168 54
rect 208 36 218 70
rect 252 36 318 70
rect 352 36 368 70
rect 408 20 418 54
rect 452 20 518 54
rect 552 20 568 54
rect 608 36 618 70
rect 652 36 718 70
rect 752 36 768 70
rect 808 20 818 54
rect 852 20 918 54
rect 952 20 968 54
rect 1008 36 1018 70
rect 1052 36 1118 70
rect 1152 36 1168 70
rect 1208 20 1218 54
rect 1252 20 1318 54
rect 1352 20 1368 54
rect 1408 36 1418 70
rect 1452 36 1518 70
rect 1552 36 1568 70
rect 1608 20 1618 54
rect 1652 20 1718 54
rect 1752 20 1768 54
rect 1808 36 1818 70
rect 1852 36 1918 70
rect 1952 36 1968 70
rect 2008 20 2018 54
rect 2052 20 2118 54
rect 2152 20 2168 54
rect 2208 36 2218 70
rect 2252 36 2318 70
rect 2352 36 2368 70
rect 2408 20 2418 54
rect 2452 20 2518 54
rect 2552 20 2568 54
rect 2608 36 2618 70
rect 2652 36 2718 70
rect 2752 36 2768 70
rect 2808 20 2818 54
rect 2852 20 2918 54
rect 2952 20 2968 54
rect 3008 36 3018 70
rect 3052 36 3118 70
rect 3152 36 3168 70
rect 3208 20 3218 54
rect 3252 20 3318 54
rect 3352 20 3368 54
rect 3408 36 3418 70
rect 3452 36 3518 70
rect 3552 36 3568 70
rect 3608 20 3618 54
rect 3652 20 3718 54
rect 3752 20 3768 54
rect 3808 36 3818 70
rect 3852 36 3918 70
rect 3952 36 3968 70
rect 4008 20 4018 54
rect 4052 20 4118 54
rect 4152 20 4168 54
rect 4208 36 4218 70
rect 4252 36 4318 70
rect 4352 36 4368 70
rect 4408 20 4418 54
rect 4452 20 4518 54
rect 4552 20 4568 54
rect 4608 36 4618 70
rect 4652 36 4718 70
rect 4752 36 4768 70
rect 4808 20 4818 54
rect 4852 20 4918 54
rect 4952 20 4968 54
rect 5008 36 5018 70
rect 5052 36 5118 70
rect 5152 36 5168 70
rect 5208 20 5218 54
rect 5252 20 5318 54
rect 5352 20 5368 54
rect 5408 36 5418 70
rect 5452 36 5518 70
rect 5552 36 5568 70
rect 5608 20 5618 54
rect 5652 20 5718 54
rect 5752 20 5768 54
rect 5808 36 5818 70
rect 5852 36 5918 70
rect 5952 36 5968 70
rect 6008 20 6018 54
rect 6052 20 6118 54
rect 6152 20 6168 54
rect 6208 36 6218 70
rect 6252 36 6318 70
rect 6352 36 6368 70
rect 6516 51 6568 68
rect 6550 34 6568 51
rect 6602 34 6618 68
rect 6652 34 6668 68
rect 6702 39 6720 68
rect 6702 34 6754 39
rect 6862 34 6878 68
rect 6912 34 6928 68
rect 6962 34 6978 68
rect 7012 34 7028 68
rect 7062 34 7078 68
rect 7112 34 7128 68
rect 7162 34 7178 68
rect 7212 34 7228 68
rect 7262 34 7278 68
rect 7312 34 7328 68
rect 7362 34 7378 68
rect 7412 34 7428 68
rect 8148 51 8164 85
rect 8198 51 8232 85
rect 8266 51 8282 85
rect 8148 -8 8282 51
rect 8424 51 8447 85
rect 8481 51 8515 85
rect 8549 51 8583 85
rect 8617 51 8651 85
rect 8685 51 8708 85
rect 8424 -8 8708 51
rect 8834 51 8857 85
rect 8891 51 8925 85
rect 8959 51 8993 85
rect 9027 51 9061 85
rect 9095 51 9118 85
rect 8834 -8 9118 51
rect 9260 51 9276 85
rect 9310 51 9344 85
rect 9378 51 9394 85
rect 9260 -8 9394 51
rect -132 -61 -116 -27
rect -82 -60 -48 -27
rect -14 -61 84 -27
rect 118 -60 152 -27
rect -82 -132 -48 -94
rect 186 -61 284 -27
rect 318 -60 352 -27
rect -82 -214 -48 -183
rect 18 -133 52 -95
rect 18 -214 52 -183
rect 118 -132 152 -94
rect 386 -61 484 -27
rect 518 -60 552 -27
rect 118 -214 152 -183
rect 218 -133 252 -95
rect 218 -214 252 -183
rect 318 -132 352 -94
rect 586 -61 684 -27
rect 718 -60 752 -27
rect 318 -214 352 -183
rect 418 -133 452 -95
rect 418 -214 452 -183
rect 518 -132 552 -94
rect 786 -61 884 -27
rect 918 -60 952 -27
rect 518 -214 552 -183
rect 618 -133 652 -95
rect 618 -214 652 -183
rect 718 -132 752 -94
rect 986 -61 1084 -27
rect 1118 -60 1152 -27
rect 718 -214 752 -183
rect 818 -133 852 -95
rect 818 -214 852 -183
rect 918 -132 952 -94
rect 1186 -61 1284 -27
rect 1318 -60 1352 -27
rect 918 -214 952 -183
rect 1018 -133 1052 -95
rect 1018 -214 1052 -183
rect 1118 -132 1152 -94
rect 1386 -61 1484 -27
rect 1518 -60 1552 -27
rect 1118 -214 1152 -183
rect 1218 -133 1252 -95
rect 1218 -214 1252 -183
rect 1318 -132 1352 -94
rect 1586 -61 1684 -27
rect 1718 -60 1752 -27
rect 1318 -214 1352 -183
rect 1418 -133 1452 -95
rect 1418 -214 1452 -183
rect 1518 -132 1552 -94
rect 1786 -61 1884 -27
rect 1918 -60 1952 -27
rect 1518 -214 1552 -183
rect 1618 -133 1652 -95
rect 1618 -214 1652 -183
rect 1718 -132 1752 -94
rect 1986 -61 2084 -27
rect 2118 -60 2152 -27
rect 1718 -214 1752 -183
rect 1818 -133 1852 -95
rect 1818 -214 1852 -183
rect 1918 -132 1952 -94
rect 2186 -61 2284 -27
rect 2318 -60 2352 -27
rect 1918 -214 1952 -183
rect 2018 -133 2052 -95
rect 2018 -214 2052 -183
rect 2118 -132 2152 -94
rect 2386 -61 2484 -27
rect 2518 -60 2552 -27
rect 2118 -214 2152 -183
rect 2218 -133 2252 -95
rect 2218 -214 2252 -183
rect 2318 -132 2352 -94
rect 2586 -61 2684 -27
rect 2718 -60 2752 -27
rect 2318 -214 2352 -183
rect 2418 -133 2452 -95
rect 2418 -214 2452 -183
rect 2518 -132 2552 -94
rect 2786 -61 2884 -27
rect 2918 -60 2952 -27
rect 2518 -214 2552 -183
rect 2618 -133 2652 -95
rect 2618 -214 2652 -183
rect 2718 -132 2752 -94
rect 2986 -61 3084 -27
rect 3118 -60 3152 -27
rect 2718 -214 2752 -183
rect 2818 -133 2852 -95
rect 2818 -214 2852 -183
rect 2918 -132 2952 -94
rect 3186 -61 3284 -27
rect 3318 -60 3352 -27
rect 2918 -214 2952 -183
rect 3018 -133 3052 -95
rect 3018 -214 3052 -183
rect 3118 -132 3152 -94
rect 3386 -61 3484 -27
rect 3518 -60 3552 -27
rect 3118 -214 3152 -183
rect 3218 -133 3252 -95
rect 3218 -214 3252 -183
rect 3318 -132 3352 -94
rect 3586 -61 3684 -27
rect 3718 -60 3752 -27
rect 3318 -214 3352 -183
rect 3418 -133 3452 -95
rect 3418 -214 3452 -183
rect 3518 -132 3552 -94
rect 3786 -61 3884 -27
rect 3918 -60 3952 -27
rect 3518 -214 3552 -183
rect 3618 -133 3652 -95
rect 3618 -214 3652 -183
rect 3718 -132 3752 -94
rect 3986 -61 4084 -27
rect 4118 -60 4152 -27
rect 3718 -214 3752 -183
rect 3818 -133 3852 -95
rect 3818 -214 3852 -183
rect 3918 -132 3952 -94
rect 4186 -61 4284 -27
rect 4318 -60 4352 -27
rect 3918 -214 3952 -183
rect 4018 -133 4052 -95
rect 4018 -214 4052 -183
rect 4118 -132 4152 -94
rect 4386 -61 4484 -27
rect 4518 -60 4552 -27
rect 4118 -214 4152 -183
rect 4218 -133 4252 -95
rect 4218 -214 4252 -183
rect 4318 -132 4352 -94
rect 4586 -61 4684 -27
rect 4718 -60 4752 -27
rect 4318 -214 4352 -183
rect 4418 -133 4452 -95
rect 4418 -214 4452 -183
rect 4518 -132 4552 -94
rect 4786 -61 4884 -27
rect 4918 -60 4952 -27
rect 4518 -214 4552 -183
rect 4618 -133 4652 -95
rect 4618 -214 4652 -183
rect 4718 -132 4752 -94
rect 4986 -61 5084 -27
rect 5118 -60 5152 -27
rect 4718 -214 4752 -183
rect 4818 -133 4852 -95
rect 4818 -214 4852 -183
rect 4918 -132 4952 -94
rect 5186 -61 5284 -27
rect 5318 -60 5352 -27
rect 4918 -214 4952 -183
rect 5018 -133 5052 -95
rect 5018 -214 5052 -183
rect 5118 -132 5152 -94
rect 5386 -61 5484 -27
rect 5518 -60 5552 -27
rect 5118 -214 5152 -183
rect 5218 -133 5252 -95
rect 5218 -214 5252 -183
rect 5318 -132 5352 -94
rect 5586 -61 5684 -27
rect 5718 -60 5752 -27
rect 5318 -214 5352 -183
rect 5418 -133 5452 -95
rect 5418 -214 5452 -183
rect 5518 -132 5552 -94
rect 5786 -61 5884 -27
rect 5918 -60 5952 -27
rect 5518 -214 5552 -183
rect 5618 -133 5652 -95
rect 5618 -214 5652 -183
rect 5718 -132 5752 -94
rect 5986 -61 6084 -27
rect 6118 -60 6152 -27
rect 5718 -214 5752 -183
rect 5818 -133 5852 -95
rect 5818 -214 5852 -183
rect 5918 -132 5952 -94
rect 6186 -61 6284 -27
rect 6318 -60 6352 -27
rect 5918 -214 5952 -183
rect 6018 -133 6052 -95
rect 6018 -214 6052 -183
rect 6118 -132 6152 -94
rect 6386 -61 6402 -27
rect 8132 -42 8158 -8
rect 8196 -42 8230 -8
rect 8264 -42 8294 -8
rect 8408 -42 8442 -8
rect 8481 -42 8514 -8
rect 8549 -42 8583 -8
rect 8620 -42 8651 -8
rect 8692 -42 8724 -8
rect 8818 -42 8849 -8
rect 8891 -42 8921 -8
rect 8959 -42 8993 -8
rect 9027 -42 9061 -8
rect 9099 -42 9134 -8
rect 9248 -42 9277 -8
rect 9312 -42 9346 -8
rect 9383 -42 9410 -8
rect 6118 -214 6152 -183
rect 6218 -133 6252 -95
rect 6218 -214 6252 -183
rect 6318 -132 6352 -94
rect 8132 -142 8160 -108
rect 8196 -142 8230 -108
rect 8266 -142 8294 -108
rect 8334 -109 8368 -92
rect 6318 -214 6352 -183
rect 8408 -142 8441 -108
rect 8481 -142 8513 -108
rect 8549 -142 8583 -108
rect 8619 -142 8651 -108
rect 8691 -142 8724 -108
rect 8818 -142 8851 -108
rect 8891 -142 8923 -108
rect 8959 -142 8993 -108
rect 9029 -142 9061 -108
rect 9101 -142 9134 -108
rect 9174 -109 9208 -92
rect 8334 -208 8368 -143
rect 9248 -142 9276 -108
rect 9312 -142 9346 -108
rect 9382 -142 9410 -108
rect 9174 -208 9208 -143
rect 8132 -242 8158 -208
rect 8196 -242 8230 -208
rect 8264 -242 8294 -208
rect 8408 -242 8442 -208
rect 8481 -242 8514 -208
rect 8549 -242 8583 -208
rect 8620 -242 8651 -208
rect 8692 -242 8724 -208
rect 8818 -242 8849 -208
rect 8891 -242 8921 -208
rect 8959 -242 8993 -208
rect 9027 -242 9061 -208
rect 9099 -242 9134 -208
rect 9248 -242 9277 -208
rect 9312 -242 9346 -208
rect 9383 -242 9410 -208
rect -32 -282 18 -248
rect 52 -282 68 -248
rect 168 -282 218 -248
rect 252 -282 268 -248
rect 368 -282 418 -248
rect 452 -282 468 -248
rect 568 -282 618 -248
rect 652 -282 668 -248
rect 768 -282 818 -248
rect 852 -282 868 -248
rect 968 -282 1018 -248
rect 1052 -282 1068 -248
rect 1168 -282 1218 -248
rect 1252 -282 1268 -248
rect 1368 -282 1418 -248
rect 1452 -282 1468 -248
rect 1568 -282 1618 -248
rect 1652 -282 1668 -248
rect 1768 -282 1818 -248
rect 1852 -282 1868 -248
rect 1968 -282 2018 -248
rect 2052 -282 2068 -248
rect 2168 -282 2218 -248
rect 2252 -282 2268 -248
rect 2368 -282 2418 -248
rect 2452 -282 2468 -248
rect 2568 -282 2618 -248
rect 2652 -282 2668 -248
rect 2768 -282 2818 -248
rect 2852 -282 2868 -248
rect 2968 -282 3018 -248
rect 3052 -282 3068 -248
rect 3168 -282 3218 -248
rect 3252 -282 3268 -248
rect 3368 -282 3418 -248
rect 3452 -282 3468 -248
rect 3568 -282 3618 -248
rect 3652 -282 3668 -248
rect 3768 -282 3818 -248
rect 3852 -282 3868 -248
rect 3968 -282 4018 -248
rect 4052 -282 4068 -248
rect 4168 -282 4218 -248
rect 4252 -282 4268 -248
rect 4368 -282 4418 -248
rect 4452 -282 4468 -248
rect 4568 -282 4618 -248
rect 4652 -282 4668 -248
rect 4768 -282 4818 -248
rect 4852 -282 4868 -248
rect 4968 -282 5018 -248
rect 5052 -282 5068 -248
rect 5168 -282 5218 -248
rect 5252 -282 5268 -248
rect 5368 -282 5418 -248
rect 5452 -282 5468 -248
rect 5568 -282 5618 -248
rect 5652 -282 5668 -248
rect 5768 -282 5818 -248
rect 5852 -282 5868 -248
rect 5968 -282 6018 -248
rect 6052 -282 6068 -248
rect 6168 -282 6218 -248
rect 6252 -282 6268 -248
rect -82 -363 -48 -322
rect -82 -431 -48 -397
rect -82 -561 -48 -469
rect 18 -363 52 -322
rect 18 -431 52 -397
rect 18 -506 52 -469
rect 118 -363 152 -322
rect 118 -431 152 -397
rect -125 -595 -118 -561
rect -84 -595 -82 -561
rect -48 -595 -46 -561
rect -12 -595 -5 -561
rect 44 -577 78 -561
rect 44 -630 78 -611
rect -30 -683 4 -667
rect -30 -803 4 -717
rect 118 -683 152 -469
rect 218 -363 252 -322
rect 218 -431 252 -397
rect 218 -506 252 -469
rect 318 -363 352 -322
rect 318 -431 352 -397
rect 318 -561 352 -469
rect 418 -363 452 -322
rect 418 -431 452 -397
rect 418 -506 452 -469
rect 518 -363 552 -322
rect 518 -431 552 -397
rect 192 -577 226 -561
rect 275 -595 282 -561
rect 316 -595 318 -561
rect 352 -595 354 -561
rect 388 -595 395 -561
rect 444 -577 478 -561
rect 192 -630 226 -611
rect 444 -630 478 -611
rect 118 -733 152 -717
rect 266 -683 300 -667
rect 266 -803 300 -717
rect -30 -837 24 -803
rect 246 -837 300 -803
rect 370 -683 404 -667
rect 370 -803 404 -717
rect 518 -683 552 -469
rect 618 -363 652 -322
rect 618 -431 652 -397
rect 618 -506 652 -469
rect 718 -363 752 -322
rect 718 -431 752 -397
rect 718 -561 752 -469
rect 818 -363 852 -322
rect 818 -431 852 -397
rect 818 -506 852 -469
rect 918 -363 952 -322
rect 918 -431 952 -397
rect 592 -577 626 -561
rect 675 -595 682 -561
rect 716 -595 718 -561
rect 752 -595 754 -561
rect 788 -595 795 -561
rect 844 -577 878 -561
rect 592 -630 626 -611
rect 844 -630 878 -611
rect 518 -733 552 -717
rect 666 -683 700 -667
rect 666 -803 700 -717
rect 370 -837 424 -803
rect 646 -837 700 -803
rect 770 -683 804 -667
rect 770 -803 804 -717
rect 918 -683 952 -469
rect 1018 -363 1052 -322
rect 1018 -431 1052 -397
rect 1018 -506 1052 -469
rect 1118 -363 1152 -322
rect 1118 -431 1152 -397
rect 1118 -561 1152 -469
rect 1218 -363 1252 -322
rect 1218 -431 1252 -397
rect 1218 -506 1252 -469
rect 1318 -363 1352 -322
rect 1318 -431 1352 -397
rect 992 -577 1026 -561
rect 1075 -595 1082 -561
rect 1116 -595 1118 -561
rect 1152 -595 1154 -561
rect 1188 -595 1195 -561
rect 1244 -577 1278 -561
rect 992 -630 1026 -611
rect 1244 -630 1278 -611
rect 918 -733 952 -717
rect 1066 -683 1100 -667
rect 1066 -803 1100 -717
rect 770 -837 824 -803
rect 1046 -837 1100 -803
rect 1170 -683 1204 -667
rect 1170 -803 1204 -717
rect 1318 -683 1352 -469
rect 1418 -363 1452 -322
rect 1418 -431 1452 -397
rect 1418 -506 1452 -469
rect 1518 -363 1552 -322
rect 1518 -431 1552 -397
rect 1518 -561 1552 -469
rect 1618 -363 1652 -322
rect 1618 -431 1652 -397
rect 1618 -506 1652 -469
rect 1718 -363 1752 -322
rect 1718 -431 1752 -397
rect 1392 -577 1426 -561
rect 1475 -595 1482 -561
rect 1516 -595 1518 -561
rect 1552 -595 1554 -561
rect 1588 -595 1595 -561
rect 1644 -577 1678 -561
rect 1392 -630 1426 -611
rect 1644 -630 1678 -611
rect 1318 -733 1352 -717
rect 1466 -683 1500 -667
rect 1466 -803 1500 -717
rect 1170 -837 1224 -803
rect 1446 -837 1500 -803
rect 1570 -683 1604 -667
rect 1570 -803 1604 -717
rect 1718 -683 1752 -469
rect 1818 -363 1852 -322
rect 1818 -431 1852 -397
rect 1818 -506 1852 -469
rect 1918 -363 1952 -322
rect 1918 -431 1952 -397
rect 1918 -561 1952 -469
rect 2018 -363 2052 -322
rect 2018 -431 2052 -397
rect 2018 -506 2052 -469
rect 2118 -363 2152 -322
rect 2118 -431 2152 -397
rect 1792 -577 1826 -561
rect 1875 -595 1882 -561
rect 1916 -595 1918 -561
rect 1952 -595 1954 -561
rect 1988 -595 1995 -561
rect 2044 -577 2078 -561
rect 1792 -630 1826 -611
rect 2044 -630 2078 -611
rect 1718 -733 1752 -717
rect 1866 -683 1900 -667
rect 1866 -803 1900 -717
rect 1570 -837 1624 -803
rect 1846 -837 1900 -803
rect 1970 -683 2004 -667
rect 1970 -803 2004 -717
rect 2118 -683 2152 -469
rect 2218 -363 2252 -322
rect 2218 -431 2252 -397
rect 2218 -506 2252 -469
rect 2318 -363 2352 -322
rect 2318 -431 2352 -397
rect 2318 -561 2352 -469
rect 2418 -363 2452 -322
rect 2418 -431 2452 -397
rect 2418 -506 2452 -469
rect 2518 -363 2552 -322
rect 2518 -431 2552 -397
rect 2192 -577 2226 -561
rect 2275 -595 2282 -561
rect 2316 -595 2318 -561
rect 2352 -595 2354 -561
rect 2388 -595 2395 -561
rect 2444 -577 2478 -561
rect 2192 -630 2226 -611
rect 2444 -630 2478 -611
rect 2118 -733 2152 -717
rect 2266 -683 2300 -667
rect 2266 -803 2300 -717
rect 1970 -837 2024 -803
rect 2246 -837 2300 -803
rect 2370 -683 2404 -667
rect 2370 -803 2404 -717
rect 2518 -683 2552 -469
rect 2618 -363 2652 -322
rect 2618 -431 2652 -397
rect 2618 -506 2652 -469
rect 2718 -363 2752 -322
rect 2718 -431 2752 -397
rect 2718 -561 2752 -469
rect 2818 -363 2852 -322
rect 2818 -431 2852 -397
rect 2818 -506 2852 -469
rect 2918 -363 2952 -322
rect 2918 -431 2952 -397
rect 2592 -577 2626 -561
rect 2675 -595 2682 -561
rect 2716 -595 2718 -561
rect 2752 -595 2754 -561
rect 2788 -595 2795 -561
rect 2844 -577 2878 -561
rect 2592 -630 2626 -611
rect 2844 -630 2878 -611
rect 2518 -733 2552 -717
rect 2666 -683 2700 -667
rect 2666 -803 2700 -717
rect 2370 -837 2424 -803
rect 2646 -837 2700 -803
rect 2770 -683 2804 -667
rect 2770 -803 2804 -717
rect 2918 -683 2952 -469
rect 3018 -363 3052 -322
rect 3018 -431 3052 -397
rect 3018 -506 3052 -469
rect 3118 -363 3152 -322
rect 3118 -431 3152 -397
rect 3118 -561 3152 -469
rect 3218 -363 3252 -322
rect 3218 -431 3252 -397
rect 3218 -506 3252 -469
rect 3318 -363 3352 -322
rect 3318 -431 3352 -397
rect 2992 -577 3026 -561
rect 3075 -595 3082 -561
rect 3116 -595 3118 -561
rect 3152 -595 3154 -561
rect 3188 -595 3195 -561
rect 3244 -577 3278 -561
rect 2992 -630 3026 -611
rect 3244 -630 3278 -611
rect 2918 -733 2952 -717
rect 3066 -683 3100 -667
rect 3066 -803 3100 -717
rect 2770 -837 2824 -803
rect 3046 -837 3100 -803
rect 3170 -683 3204 -667
rect 3170 -803 3204 -717
rect 3318 -683 3352 -469
rect 3418 -363 3452 -322
rect 3418 -431 3452 -397
rect 3418 -506 3452 -469
rect 3518 -363 3552 -322
rect 3518 -431 3552 -397
rect 3518 -561 3552 -469
rect 3618 -363 3652 -322
rect 3618 -431 3652 -397
rect 3618 -506 3652 -469
rect 3718 -363 3752 -322
rect 3718 -431 3752 -397
rect 3392 -577 3426 -561
rect 3475 -595 3482 -561
rect 3516 -595 3518 -561
rect 3552 -595 3554 -561
rect 3588 -595 3595 -561
rect 3644 -577 3678 -561
rect 3392 -630 3426 -611
rect 3644 -630 3678 -611
rect 3318 -733 3352 -717
rect 3466 -683 3500 -667
rect 3466 -803 3500 -717
rect 3170 -837 3224 -803
rect 3446 -837 3500 -803
rect 3570 -683 3604 -667
rect 3570 -803 3604 -717
rect 3718 -683 3752 -469
rect 3818 -363 3852 -322
rect 3818 -431 3852 -397
rect 3818 -506 3852 -469
rect 3918 -363 3952 -322
rect 3918 -431 3952 -397
rect 3918 -561 3952 -469
rect 4018 -363 4052 -322
rect 4018 -431 4052 -397
rect 4018 -506 4052 -469
rect 4118 -363 4152 -322
rect 4118 -431 4152 -397
rect 3792 -577 3826 -561
rect 3875 -595 3882 -561
rect 3916 -595 3918 -561
rect 3952 -595 3954 -561
rect 3988 -595 3995 -561
rect 4044 -577 4078 -561
rect 3792 -630 3826 -611
rect 4044 -630 4078 -611
rect 3718 -733 3752 -717
rect 3866 -683 3900 -667
rect 3866 -803 3900 -717
rect 3570 -837 3624 -803
rect 3846 -837 3900 -803
rect 3970 -683 4004 -667
rect 3970 -803 4004 -717
rect 4118 -683 4152 -469
rect 4218 -363 4252 -322
rect 4218 -431 4252 -397
rect 4218 -506 4252 -469
rect 4318 -363 4352 -322
rect 4318 -431 4352 -397
rect 4318 -561 4352 -469
rect 4418 -363 4452 -322
rect 4418 -431 4452 -397
rect 4418 -506 4452 -469
rect 4518 -363 4552 -322
rect 4518 -431 4552 -397
rect 4192 -577 4226 -561
rect 4275 -595 4282 -561
rect 4316 -595 4318 -561
rect 4352 -595 4354 -561
rect 4388 -595 4395 -561
rect 4444 -577 4478 -561
rect 4192 -630 4226 -611
rect 4444 -630 4478 -611
rect 4118 -733 4152 -717
rect 4266 -683 4300 -667
rect 4266 -803 4300 -717
rect 3970 -837 4024 -803
rect 4246 -837 4300 -803
rect 4370 -683 4404 -667
rect 4370 -803 4404 -717
rect 4518 -683 4552 -469
rect 4618 -363 4652 -322
rect 4618 -431 4652 -397
rect 4618 -506 4652 -469
rect 4718 -363 4752 -322
rect 4718 -431 4752 -397
rect 4718 -561 4752 -469
rect 4818 -363 4852 -322
rect 4818 -431 4852 -397
rect 4818 -506 4852 -469
rect 4918 -363 4952 -322
rect 4918 -431 4952 -397
rect 4592 -577 4626 -561
rect 4675 -595 4682 -561
rect 4716 -595 4718 -561
rect 4752 -595 4754 -561
rect 4788 -595 4795 -561
rect 4844 -577 4878 -561
rect 4592 -630 4626 -611
rect 4844 -630 4878 -611
rect 4518 -733 4552 -717
rect 4666 -683 4700 -667
rect 4666 -803 4700 -717
rect 4370 -837 4424 -803
rect 4646 -837 4700 -803
rect 4770 -683 4804 -667
rect 4770 -803 4804 -717
rect 4918 -683 4952 -469
rect 5018 -363 5052 -322
rect 5018 -431 5052 -397
rect 5018 -506 5052 -469
rect 5118 -363 5152 -322
rect 5118 -431 5152 -397
rect 5118 -561 5152 -469
rect 5218 -363 5252 -322
rect 5218 -431 5252 -397
rect 5218 -506 5252 -469
rect 5318 -363 5352 -322
rect 5318 -431 5352 -397
rect 4992 -577 5026 -561
rect 5075 -595 5082 -561
rect 5116 -595 5118 -561
rect 5152 -595 5154 -561
rect 5188 -595 5195 -561
rect 5244 -577 5278 -561
rect 4992 -630 5026 -611
rect 5244 -630 5278 -611
rect 4918 -733 4952 -717
rect 5066 -683 5100 -667
rect 5066 -803 5100 -717
rect 4770 -837 4824 -803
rect 5046 -837 5100 -803
rect 5170 -683 5204 -667
rect 5170 -803 5204 -717
rect 5318 -683 5352 -469
rect 5418 -363 5452 -322
rect 5418 -431 5452 -397
rect 5418 -506 5452 -469
rect 5518 -363 5552 -322
rect 5518 -431 5552 -397
rect 5518 -561 5552 -469
rect 5618 -363 5652 -322
rect 5618 -431 5652 -397
rect 5618 -506 5652 -469
rect 5718 -363 5752 -322
rect 5718 -431 5752 -397
rect 5392 -577 5426 -561
rect 5475 -595 5482 -561
rect 5516 -595 5518 -561
rect 5552 -595 5554 -561
rect 5588 -595 5595 -561
rect 5644 -577 5678 -561
rect 5392 -630 5426 -611
rect 5644 -630 5678 -611
rect 5318 -733 5352 -717
rect 5466 -683 5500 -667
rect 5466 -803 5500 -717
rect 5170 -837 5224 -803
rect 5446 -837 5500 -803
rect 5570 -683 5604 -667
rect 5570 -803 5604 -717
rect 5718 -683 5752 -469
rect 5818 -363 5852 -322
rect 5818 -431 5852 -397
rect 5818 -506 5852 -469
rect 5918 -363 5952 -322
rect 5918 -431 5952 -397
rect 5918 -561 5952 -469
rect 6018 -363 6052 -322
rect 6018 -431 6052 -397
rect 6018 -506 6052 -469
rect 6118 -363 6152 -322
rect 6118 -431 6152 -397
rect 5792 -577 5826 -561
rect 5875 -595 5882 -561
rect 5916 -595 5918 -561
rect 5952 -595 5954 -561
rect 5988 -595 5995 -561
rect 6044 -577 6078 -561
rect 5792 -630 5826 -611
rect 6044 -630 6078 -611
rect 5718 -733 5752 -717
rect 5866 -683 5900 -667
rect 5866 -803 5900 -717
rect 5570 -837 5624 -803
rect 5846 -837 5900 -803
rect 5970 -683 6004 -667
rect 5970 -803 6004 -717
rect 6118 -683 6152 -469
rect 6218 -363 6252 -322
rect 6218 -431 6252 -397
rect 6218 -506 6252 -469
rect 6318 -363 6352 -322
rect 8132 -342 8160 -308
rect 8196 -342 8230 -308
rect 8266 -342 8294 -308
rect 8334 -309 8368 -292
rect 6318 -431 6352 -397
rect 8408 -342 8441 -308
rect 8481 -342 8513 -308
rect 8549 -342 8583 -308
rect 8619 -342 8651 -308
rect 8691 -342 8724 -308
rect 8818 -342 8851 -308
rect 8891 -342 8923 -308
rect 8959 -342 8993 -308
rect 9029 -342 9061 -308
rect 9101 -342 9134 -308
rect 9174 -309 9208 -292
rect 8334 -408 8368 -343
rect 9248 -342 9276 -308
rect 9312 -342 9346 -308
rect 9382 -342 9410 -308
rect 9174 -408 9208 -343
rect 8132 -442 8158 -408
rect 8196 -442 8230 -408
rect 8264 -442 8294 -408
rect 8408 -442 8442 -408
rect 8481 -442 8514 -408
rect 8549 -442 8583 -408
rect 8620 -442 8651 -408
rect 8692 -442 8724 -408
rect 8818 -442 8849 -408
rect 8891 -442 8921 -408
rect 8959 -442 8993 -408
rect 9027 -442 9061 -408
rect 9099 -442 9134 -408
rect 9248 -442 9277 -408
rect 9312 -442 9346 -408
rect 9383 -442 9410 -408
rect 6318 -561 6352 -469
rect 8132 -542 8160 -508
rect 8196 -542 8230 -508
rect 8266 -542 8294 -508
rect 8334 -509 8368 -492
rect 8408 -542 8441 -508
rect 8481 -542 8513 -508
rect 8549 -542 8583 -508
rect 8619 -542 8651 -508
rect 8691 -542 8724 -508
rect 8818 -542 8851 -508
rect 8891 -542 8923 -508
rect 8959 -542 8993 -508
rect 9029 -542 9061 -508
rect 9101 -542 9134 -508
rect 9174 -509 9208 -492
rect 6192 -577 6226 -561
rect 6275 -595 6282 -561
rect 6316 -595 6318 -561
rect 6352 -595 6354 -561
rect 6388 -595 6395 -561
rect 8334 -608 8368 -543
rect 9248 -542 9276 -508
rect 9312 -542 9346 -508
rect 9382 -542 9410 -508
rect 9174 -608 9208 -543
rect 6192 -630 6226 -611
rect 8132 -642 8158 -608
rect 8196 -642 8230 -608
rect 8264 -642 8294 -608
rect 8408 -642 8442 -608
rect 8481 -642 8514 -608
rect 8549 -642 8583 -608
rect 8620 -642 8651 -608
rect 8692 -642 8724 -608
rect 8818 -642 8849 -608
rect 8891 -642 8921 -608
rect 8959 -642 8993 -608
rect 9027 -642 9061 -608
rect 9099 -642 9134 -608
rect 9248 -642 9277 -608
rect 9312 -642 9346 -608
rect 9383 -642 9410 -608
rect 6118 -733 6152 -717
rect 6266 -683 6300 -667
rect 6266 -803 6300 -717
rect 8132 -742 8160 -708
rect 8196 -742 8230 -708
rect 8266 -742 8294 -708
rect 8334 -709 8368 -692
rect 5970 -837 6024 -803
rect 6246 -837 6300 -803
rect 8408 -742 8441 -708
rect 8481 -742 8513 -708
rect 8549 -742 8583 -708
rect 8619 -742 8651 -708
rect 8691 -742 8724 -708
rect 8818 -742 8851 -708
rect 8891 -742 8923 -708
rect 8959 -742 8993 -708
rect 9029 -742 9061 -708
rect 9101 -742 9134 -708
rect 9174 -709 9208 -692
rect 8334 -808 8368 -743
rect 9248 -742 9276 -708
rect 9312 -742 9346 -708
rect 9382 -742 9410 -708
rect 9174 -808 9208 -743
rect -10 -871 -4 -837
rect 30 -858 68 -837
rect -10 -892 -2 -871
rect 32 -892 66 -858
rect 102 -871 108 -837
rect 100 -892 108 -871
rect -82 -908 -48 -892
rect -82 -958 -48 -942
rect -10 -958 108 -892
rect 162 -871 168 -837
rect 202 -858 240 -837
rect 162 -892 170 -871
rect 204 -892 238 -858
rect 274 -871 280 -837
rect 272 -892 280 -871
rect 162 -908 280 -892
rect 390 -871 396 -837
rect 430 -858 468 -837
rect 390 -892 398 -871
rect 432 -892 466 -858
rect 502 -871 508 -837
rect 500 -892 508 -871
rect -10 -992 -2 -958
rect 32 -992 66 -958
rect 100 -992 108 -958
rect -82 -1008 -48 -992
rect -10 -1008 108 -992
rect 162 -958 280 -942
rect 162 -992 170 -958
rect 204 -992 238 -958
rect 272 -992 280 -958
rect -82 -1058 -48 -1042
rect -10 -1058 108 -1042
rect -10 -1092 -2 -1058
rect 32 -1092 66 -1058
rect 100 -1092 108 -1058
rect -82 -1108 -48 -1092
rect -82 -1158 -48 -1142
rect -10 -1158 108 -1092
rect -10 -1192 -2 -1158
rect 32 -1192 66 -1158
rect 100 -1192 108 -1158
rect -82 -1208 -48 -1192
rect -10 -1208 108 -1192
rect 162 -1058 280 -992
rect 390 -958 508 -892
rect 562 -871 568 -837
rect 602 -858 640 -837
rect 562 -892 570 -871
rect 604 -892 638 -858
rect 674 -871 680 -837
rect 672 -892 680 -871
rect 790 -871 796 -837
rect 830 -858 868 -837
rect 790 -892 798 -871
rect 832 -892 866 -858
rect 902 -871 908 -837
rect 900 -892 908 -871
rect 562 -908 680 -892
rect 718 -908 752 -892
rect 390 -992 398 -958
rect 432 -992 466 -958
rect 500 -992 508 -958
rect 390 -1008 508 -992
rect 562 -958 680 -942
rect 718 -958 752 -942
rect 790 -958 908 -892
rect 962 -871 968 -837
rect 1002 -858 1040 -837
rect 962 -892 970 -871
rect 1004 -892 1038 -858
rect 1074 -871 1080 -837
rect 1072 -892 1080 -871
rect 962 -908 1080 -892
rect 1190 -871 1196 -837
rect 1230 -858 1268 -837
rect 1190 -892 1198 -871
rect 1232 -892 1266 -858
rect 1302 -871 1308 -837
rect 1300 -892 1308 -871
rect 562 -992 570 -958
rect 604 -992 638 -958
rect 672 -992 680 -958
rect 790 -992 798 -958
rect 832 -992 866 -958
rect 900 -992 908 -958
rect 162 -1092 170 -1058
rect 204 -1092 238 -1058
rect 272 -1092 280 -1058
rect 162 -1158 280 -1092
rect 390 -1058 508 -1042
rect 390 -1092 398 -1058
rect 432 -1092 466 -1058
rect 500 -1092 508 -1058
rect 390 -1108 508 -1092
rect 562 -1058 680 -992
rect 718 -1008 752 -992
rect 790 -1008 908 -992
rect 962 -958 1080 -942
rect 962 -992 970 -958
rect 1004 -992 1038 -958
rect 1072 -992 1080 -958
rect 718 -1058 752 -1042
rect 790 -1058 908 -1042
rect 562 -1092 570 -1058
rect 604 -1092 638 -1058
rect 672 -1092 680 -1058
rect 790 -1092 798 -1058
rect 832 -1092 866 -1058
rect 900 -1092 908 -1058
rect 562 -1108 680 -1092
rect 718 -1108 752 -1092
rect 162 -1192 170 -1158
rect 204 -1192 238 -1158
rect 272 -1192 280 -1158
rect 162 -1208 280 -1192
rect 390 -1158 508 -1142
rect 390 -1192 398 -1158
rect 432 -1192 466 -1158
rect 500 -1192 508 -1158
rect -82 -1258 -48 -1242
rect -10 -1258 108 -1242
rect -10 -1292 -2 -1258
rect 32 -1292 66 -1258
rect 100 -1292 108 -1258
rect -82 -1308 -48 -1292
rect -82 -1358 -48 -1342
rect -10 -1358 108 -1292
rect -10 -1392 -2 -1358
rect 32 -1392 66 -1358
rect 100 -1392 108 -1358
rect -82 -1408 -48 -1392
rect -10 -1408 108 -1392
rect 162 -1258 280 -1242
rect 162 -1292 170 -1258
rect 204 -1292 238 -1258
rect 272 -1292 280 -1258
rect 162 -1358 280 -1292
rect 162 -1392 170 -1358
rect 204 -1392 238 -1358
rect 272 -1392 280 -1358
rect 162 -1408 280 -1392
rect 390 -1258 508 -1192
rect 390 -1292 398 -1258
rect 432 -1292 466 -1258
rect 500 -1292 508 -1258
rect 390 -1358 508 -1292
rect 390 -1392 398 -1358
rect 432 -1392 466 -1358
rect 500 -1392 508 -1358
rect 390 -1408 508 -1392
rect 562 -1158 680 -1142
rect 718 -1158 752 -1142
rect 790 -1158 908 -1092
rect 562 -1192 570 -1158
rect 604 -1192 638 -1158
rect 672 -1192 680 -1158
rect 790 -1192 798 -1158
rect 832 -1192 866 -1158
rect 900 -1192 908 -1158
rect 562 -1258 680 -1192
rect 718 -1208 752 -1192
rect 790 -1208 908 -1192
rect 962 -1058 1080 -992
rect 1190 -958 1308 -892
rect 1362 -871 1368 -837
rect 1402 -858 1440 -837
rect 1362 -892 1370 -871
rect 1404 -892 1438 -858
rect 1474 -871 1480 -837
rect 1472 -892 1480 -871
rect 1590 -871 1596 -837
rect 1630 -858 1668 -837
rect 1590 -892 1598 -871
rect 1632 -892 1666 -858
rect 1702 -871 1708 -837
rect 1700 -892 1708 -871
rect 1362 -908 1480 -892
rect 1518 -908 1552 -892
rect 1190 -992 1198 -958
rect 1232 -992 1266 -958
rect 1300 -992 1308 -958
rect 1190 -1008 1308 -992
rect 1362 -958 1480 -942
rect 1518 -958 1552 -942
rect 1590 -958 1708 -892
rect 1762 -871 1768 -837
rect 1802 -858 1840 -837
rect 1762 -892 1770 -871
rect 1804 -892 1838 -858
rect 1874 -871 1880 -837
rect 1872 -892 1880 -871
rect 1762 -908 1880 -892
rect 1990 -871 1996 -837
rect 2030 -858 2068 -837
rect 1990 -892 1998 -871
rect 2032 -892 2066 -858
rect 2102 -871 2108 -837
rect 2100 -892 2108 -871
rect 1362 -992 1370 -958
rect 1404 -992 1438 -958
rect 1472 -992 1480 -958
rect 1590 -992 1598 -958
rect 1632 -992 1666 -958
rect 1700 -992 1708 -958
rect 962 -1092 970 -1058
rect 1004 -1092 1038 -1058
rect 1072 -1092 1080 -1058
rect 962 -1158 1080 -1092
rect 1190 -1058 1308 -1042
rect 1190 -1092 1198 -1058
rect 1232 -1092 1266 -1058
rect 1300 -1092 1308 -1058
rect 1190 -1108 1308 -1092
rect 1362 -1058 1480 -992
rect 1518 -1008 1552 -992
rect 1590 -1008 1708 -992
rect 1762 -958 1880 -942
rect 1762 -992 1770 -958
rect 1804 -992 1838 -958
rect 1872 -992 1880 -958
rect 1518 -1058 1552 -1042
rect 1590 -1058 1708 -1042
rect 1362 -1092 1370 -1058
rect 1404 -1092 1438 -1058
rect 1472 -1092 1480 -1058
rect 1590 -1092 1598 -1058
rect 1632 -1092 1666 -1058
rect 1700 -1092 1708 -1058
rect 1362 -1108 1480 -1092
rect 1518 -1108 1552 -1092
rect 962 -1192 970 -1158
rect 1004 -1192 1038 -1158
rect 1072 -1192 1080 -1158
rect 962 -1208 1080 -1192
rect 1190 -1158 1308 -1142
rect 1190 -1192 1198 -1158
rect 1232 -1192 1266 -1158
rect 1300 -1192 1308 -1158
rect 718 -1258 752 -1242
rect 790 -1258 908 -1242
rect 562 -1292 570 -1258
rect 604 -1292 638 -1258
rect 672 -1292 680 -1258
rect 790 -1292 798 -1258
rect 832 -1292 866 -1258
rect 900 -1292 908 -1258
rect 562 -1358 680 -1292
rect 718 -1308 752 -1292
rect 790 -1308 908 -1292
rect 962 -1258 1080 -1242
rect 962 -1292 970 -1258
rect 1004 -1292 1038 -1258
rect 1072 -1292 1080 -1258
rect 962 -1308 1080 -1292
rect 1190 -1258 1308 -1192
rect 1190 -1292 1198 -1258
rect 1232 -1292 1266 -1258
rect 1300 -1292 1308 -1258
rect 1190 -1308 1308 -1292
rect 1362 -1158 1480 -1142
rect 1518 -1158 1552 -1142
rect 1590 -1158 1708 -1092
rect 1362 -1192 1370 -1158
rect 1404 -1192 1438 -1158
rect 1472 -1192 1480 -1158
rect 1590 -1192 1598 -1158
rect 1632 -1192 1666 -1158
rect 1700 -1192 1708 -1158
rect 1362 -1258 1480 -1192
rect 1518 -1208 1552 -1192
rect 1590 -1208 1708 -1192
rect 1762 -1058 1880 -992
rect 1990 -958 2108 -892
rect 2162 -871 2168 -837
rect 2202 -858 2240 -837
rect 2162 -892 2170 -871
rect 2204 -892 2238 -858
rect 2274 -871 2280 -837
rect 2272 -892 2280 -871
rect 2390 -871 2396 -837
rect 2430 -858 2468 -837
rect 2390 -892 2398 -871
rect 2432 -892 2466 -858
rect 2502 -871 2508 -837
rect 2500 -892 2508 -871
rect 2162 -908 2280 -892
rect 2318 -908 2352 -892
rect 1990 -992 1998 -958
rect 2032 -992 2066 -958
rect 2100 -992 2108 -958
rect 1990 -1008 2108 -992
rect 2162 -958 2280 -942
rect 2318 -958 2352 -942
rect 2390 -958 2508 -892
rect 2562 -871 2568 -837
rect 2602 -858 2640 -837
rect 2562 -892 2570 -871
rect 2604 -892 2638 -858
rect 2674 -871 2680 -837
rect 2672 -892 2680 -871
rect 2562 -908 2680 -892
rect 2790 -871 2796 -837
rect 2830 -858 2868 -837
rect 2790 -892 2798 -871
rect 2832 -892 2866 -858
rect 2902 -871 2908 -837
rect 2900 -892 2908 -871
rect 2162 -992 2170 -958
rect 2204 -992 2238 -958
rect 2272 -992 2280 -958
rect 2390 -992 2398 -958
rect 2432 -992 2466 -958
rect 2500 -992 2508 -958
rect 1762 -1092 1770 -1058
rect 1804 -1092 1838 -1058
rect 1872 -1092 1880 -1058
rect 1762 -1158 1880 -1092
rect 1990 -1058 2108 -1042
rect 1990 -1092 1998 -1058
rect 2032 -1092 2066 -1058
rect 2100 -1092 2108 -1058
rect 1990 -1108 2108 -1092
rect 2162 -1058 2280 -992
rect 2318 -1008 2352 -992
rect 2390 -1008 2508 -992
rect 2562 -958 2680 -942
rect 2562 -992 2570 -958
rect 2604 -992 2638 -958
rect 2672 -992 2680 -958
rect 2318 -1058 2352 -1042
rect 2390 -1058 2508 -1042
rect 2162 -1092 2170 -1058
rect 2204 -1092 2238 -1058
rect 2272 -1092 2280 -1058
rect 2390 -1092 2398 -1058
rect 2432 -1092 2466 -1058
rect 2500 -1092 2508 -1058
rect 2162 -1108 2280 -1092
rect 2318 -1108 2352 -1092
rect 1762 -1192 1770 -1158
rect 1804 -1192 1838 -1158
rect 1872 -1192 1880 -1158
rect 1762 -1208 1880 -1192
rect 1990 -1158 2108 -1142
rect 1990 -1192 1998 -1158
rect 2032 -1192 2066 -1158
rect 2100 -1192 2108 -1158
rect 1518 -1258 1552 -1242
rect 1590 -1258 1708 -1242
rect 1362 -1292 1370 -1258
rect 1404 -1292 1438 -1258
rect 1472 -1292 1480 -1258
rect 1590 -1292 1598 -1258
rect 1632 -1292 1666 -1258
rect 1700 -1292 1708 -1258
rect 1362 -1308 1480 -1292
rect 1518 -1308 1552 -1292
rect 718 -1358 752 -1342
rect 790 -1358 908 -1342
rect 562 -1392 570 -1358
rect 604 -1392 638 -1358
rect 672 -1392 680 -1358
rect 790 -1392 798 -1358
rect 832 -1392 866 -1358
rect 900 -1392 908 -1358
rect 562 -1408 680 -1392
rect 718 -1408 752 -1392
rect -82 -1458 -48 -1442
rect -10 -1458 108 -1442
rect -10 -1492 -2 -1458
rect 32 -1492 66 -1458
rect 100 -1492 108 -1458
rect -82 -1508 -48 -1492
rect -82 -1558 -48 -1542
rect -10 -1558 108 -1492
rect -10 -1592 -2 -1558
rect 32 -1592 66 -1558
rect 100 -1592 108 -1558
rect -82 -1608 -48 -1592
rect -10 -1608 108 -1592
rect 162 -1458 280 -1442
rect 162 -1492 170 -1458
rect 204 -1492 238 -1458
rect 272 -1492 280 -1458
rect 162 -1558 280 -1492
rect 162 -1592 170 -1558
rect 204 -1592 238 -1558
rect 272 -1592 280 -1558
rect 162 -1608 280 -1592
rect 390 -1458 508 -1442
rect 390 -1492 398 -1458
rect 432 -1492 466 -1458
rect 500 -1492 508 -1458
rect 390 -1558 508 -1492
rect 390 -1592 398 -1558
rect 432 -1592 466 -1558
rect 500 -1592 508 -1558
rect 390 -1608 508 -1592
rect 562 -1458 680 -1442
rect 718 -1458 752 -1442
rect 790 -1458 908 -1392
rect 562 -1492 570 -1458
rect 604 -1492 638 -1458
rect 672 -1492 680 -1458
rect 790 -1492 798 -1458
rect 832 -1492 866 -1458
rect 900 -1492 908 -1458
rect 562 -1558 680 -1492
rect 718 -1508 752 -1492
rect 718 -1558 752 -1542
rect 790 -1558 908 -1492
rect 562 -1592 570 -1558
rect 604 -1592 638 -1558
rect 672 -1592 680 -1558
rect 790 -1592 798 -1558
rect 832 -1592 866 -1558
rect 900 -1592 908 -1558
rect 562 -1608 680 -1592
rect 718 -1608 752 -1592
rect 790 -1608 908 -1592
rect 962 -1358 1080 -1342
rect 962 -1392 970 -1358
rect 1004 -1392 1038 -1358
rect 1072 -1392 1080 -1358
rect 962 -1458 1080 -1392
rect 962 -1492 970 -1458
rect 1004 -1492 1038 -1458
rect 1072 -1492 1080 -1458
rect 962 -1558 1080 -1492
rect 962 -1592 970 -1558
rect 1004 -1592 1038 -1558
rect 1072 -1592 1080 -1558
rect 962 -1608 1080 -1592
rect 1190 -1358 1308 -1342
rect 1190 -1392 1198 -1358
rect 1232 -1392 1266 -1358
rect 1300 -1392 1308 -1358
rect 1190 -1458 1308 -1392
rect 1190 -1492 1198 -1458
rect 1232 -1492 1266 -1458
rect 1300 -1492 1308 -1458
rect 1190 -1558 1308 -1492
rect 1190 -1592 1198 -1558
rect 1232 -1592 1266 -1558
rect 1300 -1592 1308 -1558
rect 1190 -1608 1308 -1592
rect 1362 -1358 1480 -1342
rect 1518 -1358 1552 -1342
rect 1590 -1358 1708 -1292
rect 1362 -1392 1370 -1358
rect 1404 -1392 1438 -1358
rect 1472 -1392 1480 -1358
rect 1590 -1392 1598 -1358
rect 1632 -1392 1666 -1358
rect 1700 -1392 1708 -1358
rect 1362 -1458 1480 -1392
rect 1518 -1408 1552 -1392
rect 1590 -1408 1708 -1392
rect 1762 -1258 1880 -1242
rect 1762 -1292 1770 -1258
rect 1804 -1292 1838 -1258
rect 1872 -1292 1880 -1258
rect 1762 -1358 1880 -1292
rect 1762 -1392 1770 -1358
rect 1804 -1392 1838 -1358
rect 1872 -1392 1880 -1358
rect 1762 -1408 1880 -1392
rect 1990 -1258 2108 -1192
rect 1990 -1292 1998 -1258
rect 2032 -1292 2066 -1258
rect 2100 -1292 2108 -1258
rect 1990 -1358 2108 -1292
rect 1990 -1392 1998 -1358
rect 2032 -1392 2066 -1358
rect 2100 -1392 2108 -1358
rect 1990 -1408 2108 -1392
rect 2162 -1158 2280 -1142
rect 2318 -1158 2352 -1142
rect 2390 -1158 2508 -1092
rect 2162 -1192 2170 -1158
rect 2204 -1192 2238 -1158
rect 2272 -1192 2280 -1158
rect 2390 -1192 2398 -1158
rect 2432 -1192 2466 -1158
rect 2500 -1192 2508 -1158
rect 2162 -1258 2280 -1192
rect 2318 -1208 2352 -1192
rect 2390 -1208 2508 -1192
rect 2562 -1058 2680 -992
rect 2790 -958 2908 -892
rect 2962 -871 2968 -837
rect 3002 -858 3040 -837
rect 2962 -892 2970 -871
rect 3004 -892 3038 -858
rect 3074 -871 3080 -837
rect 3072 -892 3080 -871
rect 3190 -871 3196 -837
rect 3230 -858 3268 -837
rect 3190 -892 3198 -871
rect 3232 -892 3266 -858
rect 3302 -871 3308 -837
rect 3300 -892 3308 -871
rect 2962 -908 3080 -892
rect 3118 -908 3152 -892
rect 2790 -992 2798 -958
rect 2832 -992 2866 -958
rect 2900 -992 2908 -958
rect 2790 -1008 2908 -992
rect 2962 -958 3080 -942
rect 3118 -958 3152 -942
rect 3190 -958 3308 -892
rect 3362 -871 3368 -837
rect 3402 -858 3440 -837
rect 3362 -892 3370 -871
rect 3404 -892 3438 -858
rect 3474 -871 3480 -837
rect 3472 -892 3480 -871
rect 3362 -908 3480 -892
rect 3590 -871 3596 -837
rect 3630 -858 3668 -837
rect 3590 -892 3598 -871
rect 3632 -892 3666 -858
rect 3702 -871 3708 -837
rect 3700 -892 3708 -871
rect 2962 -992 2970 -958
rect 3004 -992 3038 -958
rect 3072 -992 3080 -958
rect 3190 -992 3198 -958
rect 3232 -992 3266 -958
rect 3300 -992 3308 -958
rect 2562 -1092 2570 -1058
rect 2604 -1092 2638 -1058
rect 2672 -1092 2680 -1058
rect 2562 -1158 2680 -1092
rect 2790 -1058 2908 -1042
rect 2790 -1092 2798 -1058
rect 2832 -1092 2866 -1058
rect 2900 -1092 2908 -1058
rect 2790 -1108 2908 -1092
rect 2962 -1058 3080 -992
rect 3118 -1008 3152 -992
rect 3190 -1008 3308 -992
rect 3362 -958 3480 -942
rect 3362 -992 3370 -958
rect 3404 -992 3438 -958
rect 3472 -992 3480 -958
rect 3118 -1058 3152 -1042
rect 3190 -1058 3308 -1042
rect 2962 -1092 2970 -1058
rect 3004 -1092 3038 -1058
rect 3072 -1092 3080 -1058
rect 3190 -1092 3198 -1058
rect 3232 -1092 3266 -1058
rect 3300 -1092 3308 -1058
rect 2962 -1108 3080 -1092
rect 3118 -1108 3152 -1092
rect 2562 -1192 2570 -1158
rect 2604 -1192 2638 -1158
rect 2672 -1192 2680 -1158
rect 2562 -1208 2680 -1192
rect 2790 -1158 2908 -1142
rect 2790 -1192 2798 -1158
rect 2832 -1192 2866 -1158
rect 2900 -1192 2908 -1158
rect 2318 -1258 2352 -1242
rect 2390 -1258 2508 -1242
rect 2162 -1292 2170 -1258
rect 2204 -1292 2238 -1258
rect 2272 -1292 2280 -1258
rect 2390 -1292 2398 -1258
rect 2432 -1292 2466 -1258
rect 2500 -1292 2508 -1258
rect 2162 -1358 2280 -1292
rect 2318 -1308 2352 -1292
rect 2390 -1308 2508 -1292
rect 2562 -1258 2680 -1242
rect 2562 -1292 2570 -1258
rect 2604 -1292 2638 -1258
rect 2672 -1292 2680 -1258
rect 2562 -1308 2680 -1292
rect 2790 -1258 2908 -1192
rect 2790 -1292 2798 -1258
rect 2832 -1292 2866 -1258
rect 2900 -1292 2908 -1258
rect 2790 -1308 2908 -1292
rect 2962 -1158 3080 -1142
rect 3118 -1158 3152 -1142
rect 3190 -1158 3308 -1092
rect 2962 -1192 2970 -1158
rect 3004 -1192 3038 -1158
rect 3072 -1192 3080 -1158
rect 3190 -1192 3198 -1158
rect 3232 -1192 3266 -1158
rect 3300 -1192 3308 -1158
rect 2962 -1258 3080 -1192
rect 3118 -1208 3152 -1192
rect 3190 -1208 3308 -1192
rect 3362 -1058 3480 -992
rect 3590 -958 3708 -892
rect 3762 -871 3768 -837
rect 3802 -858 3840 -837
rect 3762 -892 3770 -871
rect 3804 -892 3838 -858
rect 3874 -871 3880 -837
rect 3872 -892 3880 -871
rect 3990 -871 3996 -837
rect 4030 -858 4068 -837
rect 3990 -892 3998 -871
rect 4032 -892 4066 -858
rect 4102 -871 4108 -837
rect 4100 -892 4108 -871
rect 3762 -908 3880 -892
rect 3918 -908 3952 -892
rect 3590 -992 3598 -958
rect 3632 -992 3666 -958
rect 3700 -992 3708 -958
rect 3590 -1008 3708 -992
rect 3762 -958 3880 -942
rect 3918 -958 3952 -942
rect 3990 -958 4108 -892
rect 4162 -871 4168 -837
rect 4202 -858 4240 -837
rect 4162 -892 4170 -871
rect 4204 -892 4238 -858
rect 4274 -871 4280 -837
rect 4272 -892 4280 -871
rect 4162 -908 4280 -892
rect 4390 -871 4396 -837
rect 4430 -858 4468 -837
rect 4390 -892 4398 -871
rect 4432 -892 4466 -858
rect 4502 -871 4508 -837
rect 4500 -892 4508 -871
rect 3762 -992 3770 -958
rect 3804 -992 3838 -958
rect 3872 -992 3880 -958
rect 3990 -992 3998 -958
rect 4032 -992 4066 -958
rect 4100 -992 4108 -958
rect 3362 -1092 3370 -1058
rect 3404 -1092 3438 -1058
rect 3472 -1092 3480 -1058
rect 3362 -1158 3480 -1092
rect 3590 -1058 3708 -1042
rect 3590 -1092 3598 -1058
rect 3632 -1092 3666 -1058
rect 3700 -1092 3708 -1058
rect 3590 -1108 3708 -1092
rect 3762 -1058 3880 -992
rect 3918 -1008 3952 -992
rect 3990 -1008 4108 -992
rect 4162 -958 4280 -942
rect 4162 -992 4170 -958
rect 4204 -992 4238 -958
rect 4272 -992 4280 -958
rect 3918 -1058 3952 -1042
rect 3990 -1058 4108 -1042
rect 3762 -1092 3770 -1058
rect 3804 -1092 3838 -1058
rect 3872 -1092 3880 -1058
rect 3990 -1092 3998 -1058
rect 4032 -1092 4066 -1058
rect 4100 -1092 4108 -1058
rect 3762 -1108 3880 -1092
rect 3918 -1108 3952 -1092
rect 3362 -1192 3370 -1158
rect 3404 -1192 3438 -1158
rect 3472 -1192 3480 -1158
rect 3362 -1208 3480 -1192
rect 3590 -1158 3708 -1142
rect 3590 -1192 3598 -1158
rect 3632 -1192 3666 -1158
rect 3700 -1192 3708 -1158
rect 3118 -1258 3152 -1242
rect 3190 -1258 3308 -1242
rect 2962 -1292 2970 -1258
rect 3004 -1292 3038 -1258
rect 3072 -1292 3080 -1258
rect 3190 -1292 3198 -1258
rect 3232 -1292 3266 -1258
rect 3300 -1292 3308 -1258
rect 2962 -1308 3080 -1292
rect 3118 -1308 3152 -1292
rect 2318 -1358 2352 -1342
rect 2390 -1358 2508 -1342
rect 2162 -1392 2170 -1358
rect 2204 -1392 2238 -1358
rect 2272 -1392 2280 -1358
rect 2390 -1392 2398 -1358
rect 2432 -1392 2466 -1358
rect 2500 -1392 2508 -1358
rect 2162 -1408 2280 -1392
rect 2318 -1408 2352 -1392
rect 1518 -1458 1552 -1442
rect 1590 -1458 1708 -1442
rect 1362 -1492 1370 -1458
rect 1404 -1492 1438 -1458
rect 1472 -1492 1480 -1458
rect 1590 -1492 1598 -1458
rect 1632 -1492 1666 -1458
rect 1700 -1492 1708 -1458
rect 1362 -1558 1480 -1492
rect 1518 -1508 1552 -1492
rect 1590 -1508 1708 -1492
rect 1762 -1458 1880 -1442
rect 1762 -1492 1770 -1458
rect 1804 -1492 1838 -1458
rect 1872 -1492 1880 -1458
rect 1762 -1508 1880 -1492
rect 1990 -1458 2108 -1442
rect 1990 -1492 1998 -1458
rect 2032 -1492 2066 -1458
rect 2100 -1492 2108 -1458
rect 1990 -1508 2108 -1492
rect 2162 -1458 2280 -1442
rect 2318 -1458 2352 -1442
rect 2390 -1458 2508 -1392
rect 2162 -1492 2170 -1458
rect 2204 -1492 2238 -1458
rect 2272 -1492 2280 -1458
rect 2390 -1492 2398 -1458
rect 2432 -1492 2466 -1458
rect 2500 -1492 2508 -1458
rect 2162 -1508 2280 -1492
rect 2318 -1508 2352 -1492
rect 2390 -1508 2508 -1492
rect 2562 -1358 2680 -1342
rect 2562 -1392 2570 -1358
rect 2604 -1392 2638 -1358
rect 2672 -1392 2680 -1358
rect 2562 -1458 2680 -1392
rect 2562 -1492 2570 -1458
rect 2604 -1492 2638 -1458
rect 2672 -1492 2680 -1458
rect 2562 -1508 2680 -1492
rect 2790 -1358 2908 -1342
rect 2790 -1392 2798 -1358
rect 2832 -1392 2866 -1358
rect 2900 -1392 2908 -1358
rect 2790 -1458 2908 -1392
rect 2790 -1492 2798 -1458
rect 2832 -1492 2866 -1458
rect 2900 -1492 2908 -1458
rect 2790 -1508 2908 -1492
rect 2962 -1358 3080 -1342
rect 3118 -1358 3152 -1342
rect 3190 -1358 3308 -1292
rect 2962 -1392 2970 -1358
rect 3004 -1392 3038 -1358
rect 3072 -1392 3080 -1358
rect 3190 -1392 3198 -1358
rect 3232 -1392 3266 -1358
rect 3300 -1392 3308 -1358
rect 2962 -1458 3080 -1392
rect 3118 -1408 3152 -1392
rect 3190 -1408 3308 -1392
rect 3362 -1258 3480 -1242
rect 3362 -1292 3370 -1258
rect 3404 -1292 3438 -1258
rect 3472 -1292 3480 -1258
rect 3362 -1358 3480 -1292
rect 3362 -1392 3370 -1358
rect 3404 -1392 3438 -1358
rect 3472 -1392 3480 -1358
rect 3362 -1408 3480 -1392
rect 3590 -1258 3708 -1192
rect 3590 -1292 3598 -1258
rect 3632 -1292 3666 -1258
rect 3700 -1292 3708 -1258
rect 3590 -1358 3708 -1292
rect 3590 -1392 3598 -1358
rect 3632 -1392 3666 -1358
rect 3700 -1392 3708 -1358
rect 3590 -1408 3708 -1392
rect 3762 -1158 3880 -1142
rect 3918 -1158 3952 -1142
rect 3990 -1158 4108 -1092
rect 3762 -1192 3770 -1158
rect 3804 -1192 3838 -1158
rect 3872 -1192 3880 -1158
rect 3990 -1192 3998 -1158
rect 4032 -1192 4066 -1158
rect 4100 -1192 4108 -1158
rect 3762 -1258 3880 -1192
rect 3918 -1208 3952 -1192
rect 3990 -1208 4108 -1192
rect 4162 -1058 4280 -992
rect 4390 -958 4508 -892
rect 4562 -871 4568 -837
rect 4602 -858 4640 -837
rect 4562 -892 4570 -871
rect 4604 -892 4638 -858
rect 4674 -871 4680 -837
rect 4672 -892 4680 -871
rect 4790 -871 4796 -837
rect 4830 -858 4868 -837
rect 4790 -892 4798 -871
rect 4832 -892 4866 -858
rect 4902 -871 4908 -837
rect 4900 -892 4908 -871
rect 4562 -908 4680 -892
rect 4718 -908 4752 -892
rect 4390 -992 4398 -958
rect 4432 -992 4466 -958
rect 4500 -992 4508 -958
rect 4390 -1008 4508 -992
rect 4562 -958 4680 -942
rect 4718 -958 4752 -942
rect 4790 -958 4908 -892
rect 4962 -871 4968 -837
rect 5002 -858 5040 -837
rect 4962 -892 4970 -871
rect 5004 -892 5038 -858
rect 5074 -871 5080 -837
rect 5072 -892 5080 -871
rect 4962 -908 5080 -892
rect 5190 -871 5196 -837
rect 5230 -858 5268 -837
rect 5190 -892 5198 -871
rect 5232 -892 5266 -858
rect 5302 -871 5308 -837
rect 5300 -892 5308 -871
rect 4562 -992 4570 -958
rect 4604 -992 4638 -958
rect 4672 -992 4680 -958
rect 4790 -992 4798 -958
rect 4832 -992 4866 -958
rect 4900 -992 4908 -958
rect 4162 -1092 4170 -1058
rect 4204 -1092 4238 -1058
rect 4272 -1092 4280 -1058
rect 4162 -1158 4280 -1092
rect 4390 -1058 4508 -1042
rect 4390 -1092 4398 -1058
rect 4432 -1092 4466 -1058
rect 4500 -1092 4508 -1058
rect 4390 -1108 4508 -1092
rect 4562 -1058 4680 -992
rect 4718 -1008 4752 -992
rect 4790 -1008 4908 -992
rect 4962 -958 5080 -942
rect 4962 -992 4970 -958
rect 5004 -992 5038 -958
rect 5072 -992 5080 -958
rect 4718 -1058 4752 -1042
rect 4790 -1058 4908 -1042
rect 4562 -1092 4570 -1058
rect 4604 -1092 4638 -1058
rect 4672 -1092 4680 -1058
rect 4790 -1092 4798 -1058
rect 4832 -1092 4866 -1058
rect 4900 -1092 4908 -1058
rect 4562 -1108 4680 -1092
rect 4718 -1108 4752 -1092
rect 4162 -1192 4170 -1158
rect 4204 -1192 4238 -1158
rect 4272 -1192 4280 -1158
rect 4162 -1208 4280 -1192
rect 4390 -1158 4508 -1142
rect 4390 -1192 4398 -1158
rect 4432 -1192 4466 -1158
rect 4500 -1192 4508 -1158
rect 3918 -1258 3952 -1242
rect 3990 -1258 4108 -1242
rect 3762 -1292 3770 -1258
rect 3804 -1292 3838 -1258
rect 3872 -1292 3880 -1258
rect 3990 -1292 3998 -1258
rect 4032 -1292 4066 -1258
rect 4100 -1292 4108 -1258
rect 3762 -1358 3880 -1292
rect 3918 -1308 3952 -1292
rect 3990 -1308 4108 -1292
rect 4162 -1258 4280 -1242
rect 4162 -1292 4170 -1258
rect 4204 -1292 4238 -1258
rect 4272 -1292 4280 -1258
rect 4162 -1308 4280 -1292
rect 4390 -1258 4508 -1192
rect 4390 -1292 4398 -1258
rect 4432 -1292 4466 -1258
rect 4500 -1292 4508 -1258
rect 4390 -1308 4508 -1292
rect 4562 -1158 4680 -1142
rect 4718 -1158 4752 -1142
rect 4790 -1158 4908 -1092
rect 4562 -1192 4570 -1158
rect 4604 -1192 4638 -1158
rect 4672 -1192 4680 -1158
rect 4790 -1192 4798 -1158
rect 4832 -1192 4866 -1158
rect 4900 -1192 4908 -1158
rect 4562 -1258 4680 -1192
rect 4718 -1208 4752 -1192
rect 4790 -1208 4908 -1192
rect 4962 -1058 5080 -992
rect 5190 -958 5308 -892
rect 5362 -871 5368 -837
rect 5402 -858 5440 -837
rect 5362 -892 5370 -871
rect 5404 -892 5438 -858
rect 5474 -871 5480 -837
rect 5472 -892 5480 -871
rect 5590 -871 5596 -837
rect 5630 -858 5668 -837
rect 5590 -892 5598 -871
rect 5632 -892 5666 -858
rect 5702 -871 5708 -837
rect 5700 -892 5708 -871
rect 5362 -908 5480 -892
rect 5518 -908 5552 -892
rect 5190 -992 5198 -958
rect 5232 -992 5266 -958
rect 5300 -992 5308 -958
rect 5190 -1008 5308 -992
rect 5362 -958 5480 -942
rect 5518 -958 5552 -942
rect 5590 -958 5708 -892
rect 5762 -871 5768 -837
rect 5802 -858 5840 -837
rect 5762 -892 5770 -871
rect 5804 -892 5838 -858
rect 5874 -871 5880 -837
rect 5872 -892 5880 -871
rect 5762 -908 5880 -892
rect 5990 -871 5996 -837
rect 6030 -858 6068 -837
rect 5990 -892 5998 -871
rect 6032 -892 6066 -858
rect 6102 -871 6108 -837
rect 6100 -892 6108 -871
rect 5362 -992 5370 -958
rect 5404 -992 5438 -958
rect 5472 -992 5480 -958
rect 5590 -992 5598 -958
rect 5632 -992 5666 -958
rect 5700 -992 5708 -958
rect 4962 -1092 4970 -1058
rect 5004 -1092 5038 -1058
rect 5072 -1092 5080 -1058
rect 4962 -1158 5080 -1092
rect 5190 -1058 5308 -1042
rect 5190 -1092 5198 -1058
rect 5232 -1092 5266 -1058
rect 5300 -1092 5308 -1058
rect 5190 -1108 5308 -1092
rect 5362 -1058 5480 -992
rect 5518 -1008 5552 -992
rect 5590 -1008 5708 -992
rect 5762 -958 5880 -942
rect 5762 -992 5770 -958
rect 5804 -992 5838 -958
rect 5872 -992 5880 -958
rect 5518 -1058 5552 -1042
rect 5590 -1058 5708 -1042
rect 5362 -1092 5370 -1058
rect 5404 -1092 5438 -1058
rect 5472 -1092 5480 -1058
rect 5590 -1092 5598 -1058
rect 5632 -1092 5666 -1058
rect 5700 -1092 5708 -1058
rect 5362 -1108 5480 -1092
rect 5518 -1108 5552 -1092
rect 4962 -1192 4970 -1158
rect 5004 -1192 5038 -1158
rect 5072 -1192 5080 -1158
rect 4962 -1208 5080 -1192
rect 5190 -1158 5308 -1142
rect 5190 -1192 5198 -1158
rect 5232 -1192 5266 -1158
rect 5300 -1192 5308 -1158
rect 4718 -1258 4752 -1242
rect 4790 -1258 4908 -1242
rect 4562 -1292 4570 -1258
rect 4604 -1292 4638 -1258
rect 4672 -1292 4680 -1258
rect 4790 -1292 4798 -1258
rect 4832 -1292 4866 -1258
rect 4900 -1292 4908 -1258
rect 4562 -1308 4680 -1292
rect 4718 -1308 4752 -1292
rect 3918 -1358 3952 -1342
rect 3990 -1358 4108 -1342
rect 3762 -1392 3770 -1358
rect 3804 -1392 3838 -1358
rect 3872 -1392 3880 -1358
rect 3990 -1392 3998 -1358
rect 4032 -1392 4066 -1358
rect 4100 -1392 4108 -1358
rect 3762 -1408 3880 -1392
rect 3918 -1408 3952 -1392
rect 3118 -1458 3152 -1442
rect 3190 -1458 3308 -1442
rect 2962 -1492 2970 -1458
rect 3004 -1492 3038 -1458
rect 3072 -1492 3080 -1458
rect 3190 -1492 3198 -1458
rect 3232 -1492 3266 -1458
rect 3300 -1492 3308 -1458
rect 2962 -1508 3080 -1492
rect 3118 -1508 3152 -1492
rect 1518 -1558 1552 -1542
rect 1590 -1558 1708 -1542
rect 1362 -1592 1370 -1558
rect 1404 -1592 1438 -1558
rect 1472 -1592 1480 -1558
rect 1590 -1592 1598 -1558
rect 1632 -1592 1666 -1558
rect 1700 -1592 1708 -1558
rect 1362 -1608 1480 -1592
rect 1518 -1608 1552 -1592
rect -82 -1658 -48 -1642
rect -10 -1658 108 -1642
rect -10 -1692 -2 -1658
rect 32 -1692 66 -1658
rect 100 -1692 108 -1658
rect -82 -1708 -48 -1692
rect -82 -1758 -48 -1742
rect -10 -1758 108 -1692
rect -10 -1792 -2 -1758
rect 32 -1792 66 -1758
rect 100 -1792 108 -1758
rect -82 -1808 -48 -1792
rect -10 -1808 108 -1792
rect 162 -1658 280 -1642
rect 162 -1692 170 -1658
rect 204 -1692 238 -1658
rect 272 -1692 280 -1658
rect 162 -1758 280 -1692
rect 162 -1792 170 -1758
rect 204 -1792 238 -1758
rect 272 -1792 280 -1758
rect 162 -1808 280 -1792
rect 390 -1658 508 -1642
rect 390 -1692 398 -1658
rect 432 -1692 466 -1658
rect 500 -1692 508 -1658
rect 390 -1758 508 -1692
rect 390 -1792 398 -1758
rect 432 -1792 466 -1758
rect 500 -1792 508 -1758
rect 390 -1808 508 -1792
rect 562 -1658 680 -1642
rect 718 -1658 752 -1642
rect 790 -1658 908 -1642
rect 562 -1692 570 -1658
rect 604 -1692 638 -1658
rect 672 -1692 680 -1658
rect 790 -1692 798 -1658
rect 832 -1692 866 -1658
rect 900 -1692 908 -1658
rect 562 -1758 680 -1692
rect 718 -1708 752 -1692
rect 718 -1758 752 -1742
rect 790 -1758 908 -1692
rect 562 -1792 570 -1758
rect 604 -1792 638 -1758
rect 672 -1792 680 -1758
rect 790 -1792 798 -1758
rect 832 -1792 866 -1758
rect 900 -1792 908 -1758
rect 562 -1808 680 -1792
rect 718 -1808 752 -1792
rect 790 -1808 908 -1792
rect 962 -1658 1080 -1642
rect 962 -1692 970 -1658
rect 1004 -1692 1038 -1658
rect 1072 -1692 1080 -1658
rect 962 -1758 1080 -1692
rect 962 -1792 970 -1758
rect 1004 -1792 1038 -1758
rect 1072 -1792 1080 -1758
rect 962 -1808 1080 -1792
rect 1190 -1658 1308 -1642
rect 1190 -1692 1198 -1658
rect 1232 -1692 1266 -1658
rect 1300 -1692 1308 -1658
rect 1190 -1758 1308 -1692
rect 1190 -1792 1198 -1758
rect 1232 -1792 1266 -1758
rect 1300 -1792 1308 -1758
rect 1190 -1808 1308 -1792
rect 1362 -1658 1480 -1642
rect 1518 -1658 1552 -1642
rect 1590 -1658 1708 -1592
rect 1362 -1692 1370 -1658
rect 1404 -1692 1438 -1658
rect 1472 -1692 1480 -1658
rect 1590 -1692 1598 -1658
rect 1632 -1692 1666 -1658
rect 1700 -1692 1708 -1658
rect 1362 -1758 1480 -1692
rect 1518 -1708 1552 -1692
rect 1518 -1758 1552 -1742
rect 1590 -1758 1708 -1692
rect 1362 -1792 1370 -1758
rect 1404 -1792 1438 -1758
rect 1472 -1792 1480 -1758
rect 1590 -1792 1598 -1758
rect 1632 -1792 1666 -1758
rect 1700 -1792 1708 -1758
rect 1362 -1808 1480 -1792
rect 1518 -1808 1552 -1792
rect 1590 -1808 1708 -1792
rect 1762 -1558 1880 -1542
rect 1762 -1592 1770 -1558
rect 1804 -1592 1838 -1558
rect 1872 -1592 1880 -1558
rect 1762 -1658 1880 -1592
rect 1762 -1692 1770 -1658
rect 1804 -1692 1838 -1658
rect 1872 -1692 1880 -1658
rect 1762 -1758 1880 -1692
rect 1762 -1792 1770 -1758
rect 1804 -1792 1838 -1758
rect 1872 -1792 1880 -1758
rect 1762 -1808 1880 -1792
rect 1990 -1558 2108 -1542
rect 1990 -1592 1998 -1558
rect 2032 -1592 2066 -1558
rect 2100 -1592 2108 -1558
rect 1990 -1658 2108 -1592
rect 1990 -1692 1998 -1658
rect 2032 -1692 2066 -1658
rect 2100 -1692 2108 -1658
rect 1990 -1758 2108 -1692
rect 1990 -1792 1998 -1758
rect 2032 -1792 2066 -1758
rect 2100 -1792 2108 -1758
rect 1990 -1808 2108 -1792
rect 2162 -1558 2280 -1542
rect 2318 -1558 2352 -1542
rect 2390 -1558 2508 -1542
rect 2162 -1592 2170 -1558
rect 2204 -1592 2238 -1558
rect 2272 -1592 2280 -1558
rect 2390 -1592 2398 -1558
rect 2432 -1592 2466 -1558
rect 2500 -1592 2508 -1558
rect 2162 -1658 2280 -1592
rect 2318 -1608 2352 -1592
rect 2318 -1658 2352 -1642
rect 2390 -1658 2508 -1592
rect 2162 -1692 2170 -1658
rect 2204 -1692 2238 -1658
rect 2272 -1692 2280 -1658
rect 2390 -1692 2398 -1658
rect 2432 -1692 2466 -1658
rect 2500 -1692 2508 -1658
rect 2162 -1758 2280 -1692
rect 2318 -1708 2352 -1692
rect 2318 -1758 2352 -1742
rect 2390 -1758 2508 -1692
rect 2162 -1792 2170 -1758
rect 2204 -1792 2238 -1758
rect 2272 -1792 2280 -1758
rect 2390 -1792 2398 -1758
rect 2432 -1792 2466 -1758
rect 2500 -1792 2508 -1758
rect 2162 -1808 2280 -1792
rect 2318 -1808 2352 -1792
rect 2390 -1808 2508 -1792
rect 2562 -1558 2680 -1542
rect 2562 -1592 2570 -1558
rect 2604 -1592 2638 -1558
rect 2672 -1592 2680 -1558
rect 2562 -1658 2680 -1592
rect 2562 -1692 2570 -1658
rect 2604 -1692 2638 -1658
rect 2672 -1692 2680 -1658
rect 2562 -1758 2680 -1692
rect 2562 -1792 2570 -1758
rect 2604 -1792 2638 -1758
rect 2672 -1792 2680 -1758
rect 2562 -1808 2680 -1792
rect 2790 -1558 2908 -1542
rect 2790 -1592 2798 -1558
rect 2832 -1592 2866 -1558
rect 2900 -1592 2908 -1558
rect 2790 -1658 2908 -1592
rect 2790 -1692 2798 -1658
rect 2832 -1692 2866 -1658
rect 2900 -1692 2908 -1658
rect 2790 -1758 2908 -1692
rect 2790 -1792 2798 -1758
rect 2832 -1792 2866 -1758
rect 2900 -1792 2908 -1758
rect 2790 -1808 2908 -1792
rect 2962 -1558 3080 -1542
rect 3118 -1558 3152 -1542
rect 3190 -1558 3308 -1492
rect 2962 -1592 2970 -1558
rect 3004 -1592 3038 -1558
rect 3072 -1592 3080 -1558
rect 3190 -1592 3198 -1558
rect 3232 -1592 3266 -1558
rect 3300 -1592 3308 -1558
rect 2962 -1658 3080 -1592
rect 3118 -1608 3152 -1592
rect 3190 -1608 3308 -1592
rect 3362 -1458 3480 -1442
rect 3362 -1492 3370 -1458
rect 3404 -1492 3438 -1458
rect 3472 -1492 3480 -1458
rect 3362 -1558 3480 -1492
rect 3362 -1592 3370 -1558
rect 3404 -1592 3438 -1558
rect 3472 -1592 3480 -1558
rect 3362 -1608 3480 -1592
rect 3590 -1458 3708 -1442
rect 3590 -1492 3598 -1458
rect 3632 -1492 3666 -1458
rect 3700 -1492 3708 -1458
rect 3590 -1558 3708 -1492
rect 3590 -1592 3598 -1558
rect 3632 -1592 3666 -1558
rect 3700 -1592 3708 -1558
rect 3590 -1608 3708 -1592
rect 3762 -1458 3880 -1442
rect 3918 -1458 3952 -1442
rect 3990 -1458 4108 -1392
rect 3762 -1492 3770 -1458
rect 3804 -1492 3838 -1458
rect 3872 -1492 3880 -1458
rect 3990 -1492 3998 -1458
rect 4032 -1492 4066 -1458
rect 4100 -1492 4108 -1458
rect 3762 -1558 3880 -1492
rect 3918 -1508 3952 -1492
rect 3918 -1558 3952 -1542
rect 3990 -1558 4108 -1492
rect 3762 -1592 3770 -1558
rect 3804 -1592 3838 -1558
rect 3872 -1592 3880 -1558
rect 3990 -1592 3998 -1558
rect 4032 -1592 4066 -1558
rect 4100 -1592 4108 -1558
rect 3762 -1608 3880 -1592
rect 3918 -1608 3952 -1592
rect 3990 -1608 4108 -1592
rect 4162 -1358 4280 -1342
rect 4162 -1392 4170 -1358
rect 4204 -1392 4238 -1358
rect 4272 -1392 4280 -1358
rect 4162 -1458 4280 -1392
rect 4162 -1492 4170 -1458
rect 4204 -1492 4238 -1458
rect 4272 -1492 4280 -1458
rect 4162 -1558 4280 -1492
rect 4162 -1592 4170 -1558
rect 4204 -1592 4238 -1558
rect 4272 -1592 4280 -1558
rect 4162 -1608 4280 -1592
rect 4390 -1358 4508 -1342
rect 4390 -1392 4398 -1358
rect 4432 -1392 4466 -1358
rect 4500 -1392 4508 -1358
rect 4390 -1458 4508 -1392
rect 4390 -1492 4398 -1458
rect 4432 -1492 4466 -1458
rect 4500 -1492 4508 -1458
rect 4390 -1558 4508 -1492
rect 4390 -1592 4398 -1558
rect 4432 -1592 4466 -1558
rect 4500 -1592 4508 -1558
rect 4390 -1608 4508 -1592
rect 4562 -1358 4680 -1342
rect 4718 -1358 4752 -1342
rect 4790 -1358 4908 -1292
rect 4562 -1392 4570 -1358
rect 4604 -1392 4638 -1358
rect 4672 -1392 4680 -1358
rect 4790 -1392 4798 -1358
rect 4832 -1392 4866 -1358
rect 4900 -1392 4908 -1358
rect 4562 -1458 4680 -1392
rect 4718 -1408 4752 -1392
rect 4790 -1408 4908 -1392
rect 4962 -1258 5080 -1242
rect 4962 -1292 4970 -1258
rect 5004 -1292 5038 -1258
rect 5072 -1292 5080 -1258
rect 4962 -1358 5080 -1292
rect 4962 -1392 4970 -1358
rect 5004 -1392 5038 -1358
rect 5072 -1392 5080 -1358
rect 4962 -1408 5080 -1392
rect 5190 -1258 5308 -1192
rect 5190 -1292 5198 -1258
rect 5232 -1292 5266 -1258
rect 5300 -1292 5308 -1258
rect 5190 -1358 5308 -1292
rect 5190 -1392 5198 -1358
rect 5232 -1392 5266 -1358
rect 5300 -1392 5308 -1358
rect 5190 -1408 5308 -1392
rect 5362 -1158 5480 -1142
rect 5518 -1158 5552 -1142
rect 5590 -1158 5708 -1092
rect 5362 -1192 5370 -1158
rect 5404 -1192 5438 -1158
rect 5472 -1192 5480 -1158
rect 5590 -1192 5598 -1158
rect 5632 -1192 5666 -1158
rect 5700 -1192 5708 -1158
rect 5362 -1258 5480 -1192
rect 5518 -1208 5552 -1192
rect 5590 -1208 5708 -1192
rect 5762 -1058 5880 -992
rect 5990 -958 6108 -892
rect 6162 -871 6168 -837
rect 6202 -858 6240 -837
rect 6162 -892 6170 -871
rect 6204 -892 6238 -858
rect 6274 -871 6280 -837
rect 8132 -842 8158 -808
rect 8196 -842 8230 -808
rect 8264 -842 8294 -808
rect 8408 -842 8442 -808
rect 8481 -842 8514 -808
rect 8549 -842 8583 -808
rect 8620 -842 8651 -808
rect 8692 -842 8724 -808
rect 8818 -842 8849 -808
rect 8891 -842 8921 -808
rect 8959 -842 8993 -808
rect 9027 -842 9061 -808
rect 9099 -842 9134 -808
rect 9248 -842 9277 -808
rect 9312 -842 9346 -808
rect 9383 -842 9410 -808
rect 6272 -892 6280 -871
rect 6162 -908 6280 -892
rect 6318 -908 6352 -892
rect 8132 -942 8160 -908
rect 8196 -942 8230 -908
rect 8266 -942 8294 -908
rect 8334 -909 8368 -892
rect 5990 -992 5998 -958
rect 6032 -992 6066 -958
rect 6100 -992 6108 -958
rect 5990 -1008 6108 -992
rect 6162 -958 6280 -942
rect 6318 -958 6352 -942
rect 8408 -942 8441 -908
rect 8481 -942 8513 -908
rect 8549 -942 8583 -908
rect 8619 -942 8651 -908
rect 8691 -942 8724 -908
rect 8818 -942 8851 -908
rect 8891 -942 8923 -908
rect 8959 -942 8993 -908
rect 9029 -942 9061 -908
rect 9101 -942 9134 -908
rect 9174 -909 9208 -892
rect 6162 -992 6170 -958
rect 6204 -992 6238 -958
rect 6272 -992 6280 -958
rect 5762 -1092 5770 -1058
rect 5804 -1092 5838 -1058
rect 5872 -1092 5880 -1058
rect 5762 -1158 5880 -1092
rect 5990 -1058 6108 -1042
rect 5990 -1092 5998 -1058
rect 6032 -1092 6066 -1058
rect 6100 -1092 6108 -1058
rect 5990 -1108 6108 -1092
rect 6162 -1058 6280 -992
rect 6318 -1008 6352 -992
rect 8334 -1008 8368 -943
rect 9248 -942 9276 -908
rect 9312 -942 9346 -908
rect 9382 -942 9410 -908
rect 9174 -1008 9208 -943
rect 8132 -1042 8158 -1008
rect 8196 -1042 8230 -1008
rect 8264 -1042 8294 -1008
rect 8408 -1042 8442 -1008
rect 8481 -1042 8514 -1008
rect 8549 -1042 8583 -1008
rect 8620 -1042 8651 -1008
rect 8692 -1042 8724 -1008
rect 8818 -1042 8849 -1008
rect 8891 -1042 8921 -1008
rect 8959 -1042 8993 -1008
rect 9027 -1042 9061 -1008
rect 9099 -1042 9134 -1008
rect 9248 -1042 9277 -1008
rect 9312 -1042 9346 -1008
rect 9383 -1042 9410 -1008
rect 6318 -1058 6352 -1042
rect 6162 -1092 6170 -1058
rect 6204 -1092 6238 -1058
rect 6272 -1092 6280 -1058
rect 6162 -1108 6280 -1092
rect 6318 -1108 6352 -1092
rect 8132 -1142 8160 -1108
rect 8196 -1142 8230 -1108
rect 8266 -1142 8294 -1108
rect 8334 -1109 8368 -1092
rect 5762 -1192 5770 -1158
rect 5804 -1192 5838 -1158
rect 5872 -1192 5880 -1158
rect 5762 -1208 5880 -1192
rect 5990 -1158 6108 -1142
rect 5990 -1192 5998 -1158
rect 6032 -1192 6066 -1158
rect 6100 -1192 6108 -1158
rect 5518 -1258 5552 -1242
rect 5590 -1258 5708 -1242
rect 5362 -1292 5370 -1258
rect 5404 -1292 5438 -1258
rect 5472 -1292 5480 -1258
rect 5590 -1292 5598 -1258
rect 5632 -1292 5666 -1258
rect 5700 -1292 5708 -1258
rect 5362 -1358 5480 -1292
rect 5518 -1308 5552 -1292
rect 5590 -1308 5708 -1292
rect 5762 -1258 5880 -1242
rect 5762 -1292 5770 -1258
rect 5804 -1292 5838 -1258
rect 5872 -1292 5880 -1258
rect 5762 -1308 5880 -1292
rect 5990 -1258 6108 -1192
rect 5990 -1292 5998 -1258
rect 6032 -1292 6066 -1258
rect 6100 -1292 6108 -1258
rect 5990 -1308 6108 -1292
rect 6162 -1158 6280 -1142
rect 6318 -1158 6352 -1142
rect 8408 -1142 8441 -1108
rect 8481 -1142 8513 -1108
rect 8549 -1142 8583 -1108
rect 8619 -1142 8651 -1108
rect 8691 -1142 8724 -1108
rect 8818 -1142 8851 -1108
rect 8891 -1142 8923 -1108
rect 8959 -1142 8993 -1108
rect 9029 -1142 9061 -1108
rect 9101 -1142 9134 -1108
rect 9174 -1109 9208 -1092
rect 6162 -1192 6170 -1158
rect 6204 -1192 6238 -1158
rect 6272 -1192 6280 -1158
rect 6162 -1258 6280 -1192
rect 6318 -1208 6352 -1192
rect 8334 -1208 8368 -1143
rect 9248 -1142 9276 -1108
rect 9312 -1142 9346 -1108
rect 9382 -1142 9410 -1108
rect 9174 -1208 9208 -1143
rect 8132 -1242 8158 -1208
rect 8196 -1242 8230 -1208
rect 8264 -1242 8294 -1208
rect 8408 -1242 8442 -1208
rect 8481 -1242 8514 -1208
rect 8549 -1242 8583 -1208
rect 8620 -1242 8651 -1208
rect 8692 -1242 8724 -1208
rect 8818 -1242 8849 -1208
rect 8891 -1242 8921 -1208
rect 8959 -1242 8993 -1208
rect 9027 -1242 9061 -1208
rect 9099 -1242 9134 -1208
rect 9248 -1242 9277 -1208
rect 9312 -1242 9346 -1208
rect 9383 -1242 9410 -1208
rect 6318 -1258 6352 -1242
rect 6162 -1292 6170 -1258
rect 6204 -1292 6238 -1258
rect 6272 -1292 6280 -1258
rect 6162 -1308 6280 -1292
rect 6318 -1308 6352 -1292
rect 8132 -1342 8160 -1308
rect 8196 -1342 8230 -1308
rect 8266 -1342 8294 -1308
rect 8334 -1309 8368 -1292
rect 5518 -1358 5552 -1342
rect 5590 -1358 5708 -1342
rect 5362 -1392 5370 -1358
rect 5404 -1392 5438 -1358
rect 5472 -1392 5480 -1358
rect 5590 -1392 5598 -1358
rect 5632 -1392 5666 -1358
rect 5700 -1392 5708 -1358
rect 5362 -1408 5480 -1392
rect 5518 -1408 5552 -1392
rect 4718 -1458 4752 -1442
rect 4790 -1458 4908 -1442
rect 4562 -1492 4570 -1458
rect 4604 -1492 4638 -1458
rect 4672 -1492 4680 -1458
rect 4790 -1492 4798 -1458
rect 4832 -1492 4866 -1458
rect 4900 -1492 4908 -1458
rect 4562 -1558 4680 -1492
rect 4718 -1508 4752 -1492
rect 4790 -1508 4908 -1492
rect 4962 -1458 5080 -1442
rect 4962 -1492 4970 -1458
rect 5004 -1492 5038 -1458
rect 5072 -1492 5080 -1458
rect 4962 -1508 5080 -1492
rect 5190 -1458 5308 -1442
rect 5190 -1492 5198 -1458
rect 5232 -1492 5266 -1458
rect 5300 -1492 5308 -1458
rect 5190 -1508 5308 -1492
rect 5362 -1458 5480 -1442
rect 5518 -1458 5552 -1442
rect 5590 -1458 5708 -1392
rect 5362 -1492 5370 -1458
rect 5404 -1492 5438 -1458
rect 5472 -1492 5480 -1458
rect 5590 -1492 5598 -1458
rect 5632 -1492 5666 -1458
rect 5700 -1492 5708 -1458
rect 5362 -1508 5480 -1492
rect 5518 -1508 5552 -1492
rect 5590 -1508 5708 -1492
rect 5762 -1358 5880 -1342
rect 5762 -1392 5770 -1358
rect 5804 -1392 5838 -1358
rect 5872 -1392 5880 -1358
rect 5762 -1458 5880 -1392
rect 5762 -1492 5770 -1458
rect 5804 -1492 5838 -1458
rect 5872 -1492 5880 -1458
rect 5762 -1508 5880 -1492
rect 5990 -1358 6108 -1342
rect 5990 -1392 5998 -1358
rect 6032 -1392 6066 -1358
rect 6100 -1392 6108 -1358
rect 5990 -1458 6108 -1392
rect 5990 -1492 5998 -1458
rect 6032 -1492 6066 -1458
rect 6100 -1492 6108 -1458
rect 5990 -1508 6108 -1492
rect 6162 -1358 6280 -1342
rect 6318 -1358 6352 -1342
rect 8408 -1342 8441 -1308
rect 8481 -1342 8513 -1308
rect 8549 -1342 8583 -1308
rect 8619 -1342 8651 -1308
rect 8691 -1342 8724 -1308
rect 8818 -1342 8851 -1308
rect 8891 -1342 8923 -1308
rect 8959 -1342 8993 -1308
rect 9029 -1342 9061 -1308
rect 9101 -1342 9134 -1308
rect 9174 -1309 9208 -1292
rect 6162 -1392 6170 -1358
rect 6204 -1392 6238 -1358
rect 6272 -1392 6280 -1358
rect 6162 -1458 6280 -1392
rect 6318 -1408 6352 -1392
rect 8334 -1408 8368 -1343
rect 9248 -1342 9276 -1308
rect 9312 -1342 9346 -1308
rect 9382 -1342 9410 -1308
rect 9174 -1408 9208 -1343
rect 8132 -1442 8158 -1408
rect 8196 -1442 8230 -1408
rect 8264 -1442 8294 -1408
rect 8408 -1442 8442 -1408
rect 8481 -1442 8514 -1408
rect 8549 -1442 8583 -1408
rect 8620 -1442 8651 -1408
rect 8692 -1442 8724 -1408
rect 8818 -1442 8849 -1408
rect 8891 -1442 8921 -1408
rect 8959 -1442 8993 -1408
rect 9027 -1442 9061 -1408
rect 9099 -1442 9134 -1408
rect 9248 -1442 9277 -1408
rect 9312 -1442 9346 -1408
rect 9383 -1442 9410 -1408
rect 6318 -1458 6352 -1442
rect 6162 -1492 6170 -1458
rect 6204 -1492 6238 -1458
rect 6272 -1492 6280 -1458
rect 6162 -1508 6280 -1492
rect 6318 -1508 6352 -1492
rect 8132 -1542 8160 -1508
rect 8196 -1542 8230 -1508
rect 8266 -1542 8294 -1508
rect 8334 -1509 8368 -1492
rect 4718 -1558 4752 -1542
rect 4790 -1558 4908 -1542
rect 4562 -1592 4570 -1558
rect 4604 -1592 4638 -1558
rect 4672 -1592 4680 -1558
rect 4790 -1592 4798 -1558
rect 4832 -1592 4866 -1558
rect 4900 -1592 4908 -1558
rect 4562 -1608 4680 -1592
rect 4718 -1608 4752 -1592
rect 3118 -1658 3152 -1642
rect 3190 -1658 3308 -1642
rect 2962 -1692 2970 -1658
rect 3004 -1692 3038 -1658
rect 3072 -1692 3080 -1658
rect 3190 -1692 3198 -1658
rect 3232 -1692 3266 -1658
rect 3300 -1692 3308 -1658
rect 2962 -1758 3080 -1692
rect 3118 -1708 3152 -1692
rect 3190 -1708 3308 -1692
rect 3362 -1658 3480 -1642
rect 3362 -1692 3370 -1658
rect 3404 -1692 3438 -1658
rect 3472 -1692 3480 -1658
rect 3362 -1708 3480 -1692
rect 3590 -1658 3708 -1642
rect 3590 -1692 3598 -1658
rect 3632 -1692 3666 -1658
rect 3700 -1692 3708 -1658
rect 3590 -1708 3708 -1692
rect 3762 -1658 3880 -1642
rect 3918 -1658 3952 -1642
rect 3990 -1658 4108 -1642
rect 3762 -1692 3770 -1658
rect 3804 -1692 3838 -1658
rect 3872 -1692 3880 -1658
rect 3990 -1692 3998 -1658
rect 4032 -1692 4066 -1658
rect 4100 -1692 4108 -1658
rect 3762 -1708 3880 -1692
rect 3918 -1708 3952 -1692
rect 3990 -1708 4108 -1692
rect 4162 -1658 4280 -1642
rect 4162 -1692 4170 -1658
rect 4204 -1692 4238 -1658
rect 4272 -1692 4280 -1658
rect 4162 -1708 4280 -1692
rect 4390 -1658 4508 -1642
rect 4390 -1692 4398 -1658
rect 4432 -1692 4466 -1658
rect 4500 -1692 4508 -1658
rect 4390 -1708 4508 -1692
rect 4562 -1658 4680 -1642
rect 4718 -1658 4752 -1642
rect 4790 -1658 4908 -1592
rect 4562 -1692 4570 -1658
rect 4604 -1692 4638 -1658
rect 4672 -1692 4680 -1658
rect 4790 -1692 4798 -1658
rect 4832 -1692 4866 -1658
rect 4900 -1692 4908 -1658
rect 4562 -1708 4680 -1692
rect 4718 -1708 4752 -1692
rect 4790 -1708 4908 -1692
rect 4962 -1558 5080 -1542
rect 4962 -1592 4970 -1558
rect 5004 -1592 5038 -1558
rect 5072 -1592 5080 -1558
rect 4962 -1658 5080 -1592
rect 4962 -1692 4970 -1658
rect 5004 -1692 5038 -1658
rect 5072 -1692 5080 -1658
rect 4962 -1708 5080 -1692
rect 5190 -1558 5308 -1542
rect 5190 -1592 5198 -1558
rect 5232 -1592 5266 -1558
rect 5300 -1592 5308 -1558
rect 5190 -1658 5308 -1592
rect 5190 -1692 5198 -1658
rect 5232 -1692 5266 -1658
rect 5300 -1692 5308 -1658
rect 5190 -1708 5308 -1692
rect 5362 -1558 5480 -1542
rect 5518 -1558 5552 -1542
rect 5590 -1558 5708 -1542
rect 5362 -1592 5370 -1558
rect 5404 -1592 5438 -1558
rect 5472 -1592 5480 -1558
rect 5590 -1592 5598 -1558
rect 5632 -1592 5666 -1558
rect 5700 -1592 5708 -1558
rect 5362 -1658 5480 -1592
rect 5518 -1608 5552 -1592
rect 5518 -1658 5552 -1642
rect 5590 -1658 5708 -1592
rect 5362 -1692 5370 -1658
rect 5404 -1692 5438 -1658
rect 5472 -1692 5480 -1658
rect 5590 -1692 5598 -1658
rect 5632 -1692 5666 -1658
rect 5700 -1692 5708 -1658
rect 5362 -1708 5480 -1692
rect 5518 -1708 5552 -1692
rect 5590 -1708 5708 -1692
rect 5762 -1558 5880 -1542
rect 5762 -1592 5770 -1558
rect 5804 -1592 5838 -1558
rect 5872 -1592 5880 -1558
rect 5762 -1658 5880 -1592
rect 5762 -1692 5770 -1658
rect 5804 -1692 5838 -1658
rect 5872 -1692 5880 -1658
rect 5762 -1708 5880 -1692
rect 5990 -1558 6108 -1542
rect 5990 -1592 5998 -1558
rect 6032 -1592 6066 -1558
rect 6100 -1592 6108 -1558
rect 5990 -1658 6108 -1592
rect 5990 -1692 5998 -1658
rect 6032 -1692 6066 -1658
rect 6100 -1692 6108 -1658
rect 5990 -1708 6108 -1692
rect 6162 -1558 6280 -1542
rect 6318 -1558 6352 -1542
rect 8408 -1542 8441 -1508
rect 8481 -1542 8513 -1508
rect 8549 -1542 8583 -1508
rect 8619 -1542 8651 -1508
rect 8691 -1542 8724 -1508
rect 8818 -1542 8851 -1508
rect 8891 -1542 8923 -1508
rect 8959 -1542 8993 -1508
rect 9029 -1542 9061 -1508
rect 9101 -1542 9134 -1508
rect 9174 -1509 9208 -1492
rect 6162 -1592 6170 -1558
rect 6204 -1592 6238 -1558
rect 6272 -1592 6280 -1558
rect 6162 -1658 6280 -1592
rect 6318 -1608 6352 -1592
rect 8334 -1608 8368 -1543
rect 9248 -1542 9276 -1508
rect 9312 -1542 9346 -1508
rect 9382 -1542 9410 -1508
rect 9174 -1608 9208 -1543
rect 8132 -1642 8158 -1608
rect 8196 -1642 8230 -1608
rect 8264 -1642 8294 -1608
rect 8408 -1642 8442 -1608
rect 8481 -1642 8514 -1608
rect 8549 -1642 8583 -1608
rect 8620 -1642 8651 -1608
rect 8692 -1642 8724 -1608
rect 8818 -1642 8849 -1608
rect 8891 -1642 8921 -1608
rect 8959 -1642 8993 -1608
rect 9027 -1642 9061 -1608
rect 9099 -1642 9134 -1608
rect 9248 -1642 9277 -1608
rect 9312 -1642 9346 -1608
rect 9383 -1642 9410 -1608
rect 6318 -1658 6352 -1642
rect 6162 -1692 6170 -1658
rect 6204 -1692 6238 -1658
rect 6272 -1692 6280 -1658
rect 6162 -1708 6280 -1692
rect 6318 -1708 6352 -1692
rect 8132 -1742 8160 -1708
rect 8196 -1742 8230 -1708
rect 8266 -1742 8294 -1708
rect 8334 -1709 8368 -1692
rect 3118 -1758 3152 -1742
rect 3190 -1758 3308 -1742
rect 2962 -1792 2970 -1758
rect 3004 -1792 3038 -1758
rect 3072 -1792 3080 -1758
rect 3190 -1792 3198 -1758
rect 3232 -1792 3266 -1758
rect 3300 -1792 3308 -1758
rect 2962 -1808 3080 -1792
rect 3118 -1808 3152 -1792
rect -82 -1858 -48 -1842
rect -10 -1858 108 -1842
rect -10 -1892 -2 -1858
rect 32 -1892 66 -1858
rect 100 -1892 108 -1858
rect -10 -1917 108 -1892
rect 162 -1858 280 -1842
rect 162 -1892 170 -1858
rect 204 -1892 238 -1858
rect 272 -1892 280 -1858
rect 162 -1917 280 -1892
rect 390 -1858 508 -1842
rect 390 -1892 398 -1858
rect 432 -1892 466 -1858
rect 500 -1892 508 -1858
rect 390 -1917 508 -1892
rect 562 -1858 680 -1842
rect 718 -1858 752 -1842
rect 790 -1858 908 -1842
rect 562 -1892 570 -1858
rect 604 -1892 638 -1858
rect 672 -1892 680 -1858
rect 562 -1917 680 -1892
rect 790 -1892 798 -1858
rect 832 -1892 866 -1858
rect 900 -1892 908 -1858
rect 790 -1917 908 -1892
rect 962 -1858 1080 -1842
rect 962 -1892 970 -1858
rect 1004 -1892 1038 -1858
rect 1072 -1892 1080 -1858
rect 962 -1917 1080 -1892
rect 1190 -1858 1308 -1842
rect 1190 -1892 1198 -1858
rect 1232 -1892 1266 -1858
rect 1300 -1892 1308 -1858
rect 1190 -1917 1308 -1892
rect 1362 -1858 1480 -1842
rect 1518 -1858 1552 -1842
rect 1590 -1858 1708 -1842
rect 1362 -1892 1370 -1858
rect 1404 -1892 1438 -1858
rect 1472 -1892 1480 -1858
rect 1362 -1917 1480 -1892
rect 1590 -1892 1598 -1858
rect 1632 -1892 1666 -1858
rect 1700 -1892 1708 -1858
rect 1590 -1917 1708 -1892
rect 1762 -1858 1880 -1842
rect 1762 -1892 1770 -1858
rect 1804 -1892 1838 -1858
rect 1872 -1892 1880 -1858
rect 1762 -1917 1880 -1892
rect 1990 -1858 2108 -1842
rect 1990 -1892 1998 -1858
rect 2032 -1892 2066 -1858
rect 2100 -1892 2108 -1858
rect 1990 -1917 2108 -1892
rect 2162 -1858 2280 -1842
rect 2318 -1858 2352 -1842
rect 2390 -1858 2508 -1842
rect 2162 -1892 2170 -1858
rect 2204 -1892 2238 -1858
rect 2272 -1892 2280 -1858
rect 2162 -1917 2280 -1892
rect 2390 -1892 2398 -1858
rect 2432 -1892 2466 -1858
rect 2500 -1892 2508 -1858
rect 2390 -1917 2508 -1892
rect 2562 -1858 2680 -1842
rect 2562 -1892 2570 -1858
rect 2604 -1892 2638 -1858
rect 2672 -1892 2680 -1858
rect 2562 -1917 2680 -1892
rect 2790 -1858 2908 -1842
rect 2790 -1892 2798 -1858
rect 2832 -1892 2866 -1858
rect 2900 -1892 2908 -1858
rect 2790 -1917 2908 -1892
rect 2962 -1858 3080 -1842
rect 3118 -1858 3152 -1842
rect 3190 -1858 3308 -1792
rect 2962 -1892 2970 -1858
rect 3004 -1892 3038 -1858
rect 3072 -1892 3080 -1858
rect 2962 -1917 3080 -1892
rect 3190 -1892 3198 -1858
rect 3232 -1892 3266 -1858
rect 3300 -1892 3308 -1858
rect 3190 -1917 3308 -1892
rect 3362 -1758 3480 -1742
rect 3362 -1792 3370 -1758
rect 3404 -1792 3438 -1758
rect 3472 -1792 3480 -1758
rect 3362 -1858 3480 -1792
rect 3362 -1892 3370 -1858
rect 3404 -1892 3438 -1858
rect 3472 -1892 3480 -1858
rect 3362 -1917 3480 -1892
rect 3590 -1758 3708 -1742
rect 3590 -1792 3598 -1758
rect 3632 -1792 3666 -1758
rect 3700 -1792 3708 -1758
rect 3590 -1858 3708 -1792
rect 3590 -1892 3598 -1858
rect 3632 -1892 3666 -1858
rect 3700 -1892 3708 -1858
rect 3590 -1917 3708 -1892
rect 3762 -1758 3880 -1742
rect 3918 -1758 3952 -1742
rect 3990 -1758 4108 -1742
rect 3762 -1792 3770 -1758
rect 3804 -1792 3838 -1758
rect 3872 -1792 3880 -1758
rect 3990 -1792 3998 -1758
rect 4032 -1792 4066 -1758
rect 4100 -1792 4108 -1758
rect 3762 -1858 3880 -1792
rect 3918 -1808 3952 -1792
rect 3918 -1858 3952 -1842
rect 3990 -1858 4108 -1792
rect 3762 -1892 3770 -1858
rect 3804 -1892 3838 -1858
rect 3872 -1892 3880 -1858
rect 3762 -1917 3880 -1892
rect 3990 -1892 3998 -1858
rect 4032 -1892 4066 -1858
rect 4100 -1892 4108 -1858
rect 3990 -1917 4108 -1892
rect 4162 -1758 4280 -1742
rect 4162 -1792 4170 -1758
rect 4204 -1792 4238 -1758
rect 4272 -1792 4280 -1758
rect 4162 -1858 4280 -1792
rect 4162 -1892 4170 -1858
rect 4204 -1892 4238 -1858
rect 4272 -1892 4280 -1858
rect 4162 -1917 4280 -1892
rect 4390 -1758 4508 -1742
rect 4390 -1792 4398 -1758
rect 4432 -1792 4466 -1758
rect 4500 -1792 4508 -1758
rect 4390 -1858 4508 -1792
rect 4390 -1892 4398 -1858
rect 4432 -1892 4466 -1858
rect 4500 -1892 4508 -1858
rect 4390 -1917 4508 -1892
rect 4562 -1758 4680 -1742
rect 4718 -1758 4752 -1742
rect 4790 -1758 4908 -1742
rect 4562 -1792 4570 -1758
rect 4604 -1792 4638 -1758
rect 4672 -1792 4680 -1758
rect 4790 -1792 4798 -1758
rect 4832 -1792 4866 -1758
rect 4900 -1792 4908 -1758
rect 4562 -1858 4680 -1792
rect 4718 -1808 4752 -1792
rect 4718 -1858 4752 -1842
rect 4790 -1858 4908 -1792
rect 4562 -1892 4570 -1858
rect 4604 -1892 4638 -1858
rect 4672 -1892 4680 -1858
rect 4562 -1917 4680 -1892
rect 4790 -1892 4798 -1858
rect 4832 -1892 4866 -1858
rect 4900 -1892 4908 -1858
rect 4790 -1917 4908 -1892
rect 4962 -1758 5080 -1742
rect 4962 -1792 4970 -1758
rect 5004 -1792 5038 -1758
rect 5072 -1792 5080 -1758
rect 4962 -1858 5080 -1792
rect 4962 -1892 4970 -1858
rect 5004 -1892 5038 -1858
rect 5072 -1892 5080 -1858
rect 4962 -1917 5080 -1892
rect 5190 -1758 5308 -1742
rect 5190 -1792 5198 -1758
rect 5232 -1792 5266 -1758
rect 5300 -1792 5308 -1758
rect 5190 -1858 5308 -1792
rect 5190 -1892 5198 -1858
rect 5232 -1892 5266 -1858
rect 5300 -1892 5308 -1858
rect 5190 -1917 5308 -1892
rect 5362 -1758 5480 -1742
rect 5518 -1758 5552 -1742
rect 5590 -1758 5708 -1742
rect 5362 -1792 5370 -1758
rect 5404 -1792 5438 -1758
rect 5472 -1792 5480 -1758
rect 5590 -1792 5598 -1758
rect 5632 -1792 5666 -1758
rect 5700 -1792 5708 -1758
rect 5362 -1858 5480 -1792
rect 5518 -1808 5552 -1792
rect 5518 -1858 5552 -1842
rect 5590 -1858 5708 -1792
rect 5362 -1892 5370 -1858
rect 5404 -1892 5438 -1858
rect 5472 -1892 5480 -1858
rect 5362 -1917 5480 -1892
rect 5590 -1892 5598 -1858
rect 5632 -1892 5666 -1858
rect 5700 -1892 5708 -1858
rect 5590 -1917 5708 -1892
rect 5762 -1758 5880 -1742
rect 5762 -1792 5770 -1758
rect 5804 -1792 5838 -1758
rect 5872 -1792 5880 -1758
rect 5762 -1858 5880 -1792
rect 5762 -1892 5770 -1858
rect 5804 -1892 5838 -1858
rect 5872 -1892 5880 -1858
rect 5762 -1917 5880 -1892
rect 5990 -1758 6108 -1742
rect 5990 -1792 5998 -1758
rect 6032 -1792 6066 -1758
rect 6100 -1792 6108 -1758
rect 5990 -1858 6108 -1792
rect 5990 -1892 5998 -1858
rect 6032 -1892 6066 -1858
rect 6100 -1892 6108 -1858
rect 5990 -1917 6108 -1892
rect 6162 -1758 6280 -1742
rect 6318 -1758 6352 -1742
rect 8408 -1742 8441 -1708
rect 8481 -1742 8513 -1708
rect 8549 -1742 8583 -1708
rect 8619 -1742 8651 -1708
rect 8691 -1742 8724 -1708
rect 8818 -1742 8851 -1708
rect 8891 -1742 8923 -1708
rect 8959 -1742 8993 -1708
rect 9029 -1742 9061 -1708
rect 9101 -1742 9134 -1708
rect 9174 -1709 9208 -1692
rect 6162 -1792 6170 -1758
rect 6204 -1792 6238 -1758
rect 6272 -1792 6280 -1758
rect 6162 -1858 6280 -1792
rect 6318 -1808 6352 -1792
rect 8334 -1808 8368 -1743
rect 9248 -1742 9276 -1708
rect 9312 -1742 9346 -1708
rect 9382 -1742 9410 -1708
rect 9174 -1808 9208 -1743
rect 8132 -1842 8158 -1808
rect 8196 -1842 8230 -1808
rect 8264 -1842 8294 -1808
rect 8408 -1842 8442 -1808
rect 8481 -1842 8514 -1808
rect 8549 -1842 8583 -1808
rect 8620 -1842 8651 -1808
rect 8692 -1842 8724 -1808
rect 8818 -1842 8849 -1808
rect 8891 -1842 8921 -1808
rect 8959 -1842 8993 -1808
rect 9027 -1842 9061 -1808
rect 9099 -1842 9134 -1808
rect 9248 -1842 9277 -1808
rect 9312 -1842 9346 -1808
rect 9383 -1842 9410 -1808
rect 6318 -1858 6352 -1842
rect 6162 -1892 6170 -1858
rect 6204 -1892 6238 -1858
rect 6272 -1892 6280 -1858
rect 6162 -1917 6280 -1892
rect 8148 -1901 8282 -1842
rect -65 -1935 6335 -1917
rect 8148 -1935 8164 -1901
rect 8198 -1935 8232 -1901
rect 8266 -1935 8282 -1901
rect 8424 -1901 8708 -1842
rect 8424 -1935 8447 -1901
rect 8481 -1935 8515 -1901
rect 8549 -1935 8583 -1901
rect 8617 -1935 8651 -1901
rect 8685 -1935 8708 -1901
rect 8834 -1901 9118 -1842
rect 8834 -1935 8857 -1901
rect 8891 -1935 8925 -1901
rect 8959 -1935 8993 -1901
rect 9027 -1935 9061 -1901
rect 9095 -1935 9118 -1901
rect 9260 -1901 9394 -1842
rect 9260 -1935 9276 -1901
rect 9310 -1935 9344 -1901
rect 9378 -1935 9394 -1901
rect -65 -1969 -4 -1935
rect 30 -1951 68 -1935
rect 30 -1969 32 -1951
rect -65 -1985 32 -1969
rect 66 -1969 68 -1951
rect 102 -1969 168 -1935
rect 202 -1951 240 -1935
rect 202 -1969 204 -1951
rect 66 -1985 204 -1969
rect 238 -1969 240 -1951
rect 274 -1969 396 -1935
rect 430 -1951 468 -1935
rect 430 -1969 432 -1951
rect 238 -1985 432 -1969
rect 466 -1969 468 -1951
rect 502 -1969 568 -1935
rect 602 -1951 640 -1935
rect 602 -1969 604 -1951
rect 466 -1985 604 -1969
rect 638 -1969 640 -1951
rect 674 -1969 796 -1935
rect 830 -1951 868 -1935
rect 830 -1969 832 -1951
rect 638 -1985 832 -1969
rect 866 -1969 868 -1951
rect 902 -1969 968 -1935
rect 1002 -1951 1040 -1935
rect 1002 -1969 1004 -1951
rect 866 -1985 1004 -1969
rect 1038 -1969 1040 -1951
rect 1074 -1969 1196 -1935
rect 1230 -1951 1268 -1935
rect 1230 -1969 1232 -1951
rect 1038 -1985 1232 -1969
rect 1266 -1969 1268 -1951
rect 1302 -1969 1368 -1935
rect 1402 -1951 1440 -1935
rect 1402 -1969 1404 -1951
rect 1266 -1985 1404 -1969
rect 1438 -1969 1440 -1951
rect 1474 -1969 1596 -1935
rect 1630 -1951 1668 -1935
rect 1630 -1969 1632 -1951
rect 1438 -1985 1632 -1969
rect 1666 -1969 1668 -1951
rect 1702 -1969 1768 -1935
rect 1802 -1951 1840 -1935
rect 1802 -1969 1804 -1951
rect 1666 -1985 1804 -1969
rect 1838 -1969 1840 -1951
rect 1874 -1969 1996 -1935
rect 2030 -1951 2068 -1935
rect 2030 -1969 2032 -1951
rect 1838 -1985 2032 -1969
rect 2066 -1969 2068 -1951
rect 2102 -1969 2168 -1935
rect 2202 -1951 2240 -1935
rect 2202 -1969 2204 -1951
rect 2066 -1985 2204 -1969
rect 2238 -1969 2240 -1951
rect 2274 -1969 2396 -1935
rect 2430 -1951 2468 -1935
rect 2430 -1969 2432 -1951
rect 2238 -1985 2432 -1969
rect 2466 -1969 2468 -1951
rect 2502 -1969 2568 -1935
rect 2602 -1951 2640 -1935
rect 2602 -1969 2604 -1951
rect 2466 -1985 2604 -1969
rect 2638 -1969 2640 -1951
rect 2674 -1969 2796 -1935
rect 2830 -1951 2868 -1935
rect 2830 -1969 2832 -1951
rect 2638 -1985 2832 -1969
rect 2866 -1969 2868 -1951
rect 2902 -1969 2968 -1935
rect 3002 -1951 3040 -1935
rect 3002 -1969 3004 -1951
rect 2866 -1985 3004 -1969
rect 3038 -1969 3040 -1951
rect 3074 -1969 3196 -1935
rect 3230 -1951 3268 -1935
rect 3230 -1969 3232 -1951
rect 3038 -1985 3232 -1969
rect 3266 -1969 3268 -1951
rect 3302 -1969 3368 -1935
rect 3402 -1951 3440 -1935
rect 3402 -1969 3404 -1951
rect 3266 -1985 3404 -1969
rect 3438 -1969 3440 -1951
rect 3474 -1969 3596 -1935
rect 3630 -1951 3668 -1935
rect 3630 -1969 3632 -1951
rect 3438 -1985 3632 -1969
rect 3666 -1969 3668 -1951
rect 3702 -1969 3768 -1935
rect 3802 -1951 3840 -1935
rect 3802 -1969 3804 -1951
rect 3666 -1985 3804 -1969
rect 3838 -1969 3840 -1951
rect 3874 -1969 3996 -1935
rect 4030 -1951 4068 -1935
rect 4030 -1969 4032 -1951
rect 3838 -1985 4032 -1969
rect 4066 -1969 4068 -1951
rect 4102 -1969 4168 -1935
rect 4202 -1951 4240 -1935
rect 4202 -1969 4204 -1951
rect 4066 -1985 4204 -1969
rect 4238 -1969 4240 -1951
rect 4274 -1969 4396 -1935
rect 4430 -1951 4468 -1935
rect 4430 -1969 4432 -1951
rect 4238 -1985 4432 -1969
rect 4466 -1969 4468 -1951
rect 4502 -1969 4568 -1935
rect 4602 -1951 4640 -1935
rect 4602 -1969 4604 -1951
rect 4466 -1985 4604 -1969
rect 4638 -1969 4640 -1951
rect 4674 -1969 4796 -1935
rect 4830 -1951 4868 -1935
rect 4830 -1969 4832 -1951
rect 4638 -1985 4832 -1969
rect 4866 -1969 4868 -1951
rect 4902 -1969 4968 -1935
rect 5002 -1951 5040 -1935
rect 5002 -1969 5004 -1951
rect 4866 -1985 5004 -1969
rect 5038 -1969 5040 -1951
rect 5074 -1969 5196 -1935
rect 5230 -1951 5268 -1935
rect 5230 -1969 5232 -1951
rect 5038 -1985 5232 -1969
rect 5266 -1969 5268 -1951
rect 5302 -1969 5368 -1935
rect 5402 -1951 5440 -1935
rect 5402 -1969 5404 -1951
rect 5266 -1985 5404 -1969
rect 5438 -1969 5440 -1951
rect 5474 -1969 5596 -1935
rect 5630 -1951 5668 -1935
rect 5630 -1969 5632 -1951
rect 5438 -1985 5632 -1969
rect 5666 -1969 5668 -1951
rect 5702 -1969 5768 -1935
rect 5802 -1951 5840 -1935
rect 5802 -1969 5804 -1951
rect 5666 -1985 5804 -1969
rect 5838 -1969 5840 -1951
rect 5874 -1969 5996 -1935
rect 6030 -1951 6068 -1935
rect 6030 -1969 6032 -1951
rect 5838 -1985 6032 -1969
rect 6066 -1969 6068 -1951
rect 6102 -1969 6168 -1935
rect 6202 -1951 6240 -1935
rect 6202 -1969 6204 -1951
rect 6066 -1985 6204 -1969
rect 6238 -1969 6240 -1951
rect 6274 -1969 6335 -1935
rect 6238 -1985 6335 -1969
rect -65 -1987 6335 -1985
<< viali >>
rect 118 9963 152 9997
rect 318 9963 352 9997
rect 518 9963 552 9997
rect 718 9963 752 9997
rect 918 9963 952 9997
rect 1118 9963 1152 9997
rect 1318 9963 1352 9997
rect 1518 9963 1552 9997
rect 1718 9963 1752 9997
rect 1918 9963 1952 9997
rect 2118 9963 2152 9997
rect 2318 9963 2352 9997
rect 2518 9963 2552 9997
rect 2718 9963 2752 9997
rect 2918 9963 2952 9997
rect 3118 9963 3152 9997
rect 3318 9963 3352 9997
rect 3518 9963 3552 9997
rect 3718 9963 3752 9997
rect 3918 9963 3952 9997
rect 4118 9963 4152 9997
rect 4318 9963 4352 9997
rect 4518 9963 4552 9997
rect 4718 9963 4752 9997
rect 4918 9963 4952 9997
rect 5118 9963 5152 9997
rect 5318 9963 5352 9997
rect 5518 9963 5552 9997
rect 5718 9963 5752 9997
rect 5918 9963 5952 9997
rect 6118 9963 6152 9997
rect 6318 9963 6352 9997
rect 18 9840 52 9874
rect 218 9856 252 9890
rect 418 9840 452 9874
rect 618 9856 652 9890
rect 818 9840 852 9874
rect 1018 9856 1052 9890
rect 1218 9840 1252 9874
rect 1418 9856 1452 9890
rect 1618 9840 1652 9874
rect 1818 9856 1852 9890
rect 2018 9840 2052 9874
rect 2218 9856 2252 9890
rect 2418 9840 2452 9874
rect 2618 9856 2652 9890
rect 2818 9840 2852 9874
rect 3018 9856 3052 9890
rect 3218 9840 3252 9874
rect 3418 9856 3452 9890
rect 3618 9840 3652 9874
rect 3818 9856 3852 9890
rect 4018 9840 4052 9874
rect 4218 9856 4252 9890
rect 4418 9840 4452 9874
rect 4618 9856 4652 9890
rect 4818 9840 4852 9874
rect 5018 9856 5052 9890
rect 5218 9840 5252 9874
rect 5418 9856 5452 9890
rect 5618 9840 5652 9874
rect 5818 9856 5852 9890
rect 6018 9840 6052 9874
rect 6218 9856 6252 9890
rect 6516 9837 6550 9871
rect 6720 9859 6754 9893
rect 6878 9854 6912 9888
rect 6978 9854 7012 9888
rect 7078 9854 7112 9888
rect 7178 9854 7212 9888
rect 7278 9854 7312 9888
rect 7378 9854 7412 9888
rect 18 9733 52 9767
rect 118 9733 152 9767
rect 218 9733 252 9767
rect 318 9733 352 9767
rect 418 9733 452 9767
rect 518 9733 552 9767
rect 618 9733 652 9767
rect 718 9733 752 9767
rect 818 9733 852 9767
rect 918 9733 952 9767
rect 1018 9733 1052 9767
rect 1118 9733 1152 9767
rect 1218 9733 1252 9767
rect 1318 9733 1352 9767
rect 1418 9733 1452 9767
rect 1518 9733 1546 9767
rect 1546 9733 1552 9767
rect 1618 9733 1624 9767
rect 1624 9733 1652 9767
rect 1718 9733 1752 9767
rect 1818 9733 1852 9767
rect 1918 9733 1952 9767
rect 2018 9733 2052 9767
rect 2118 9733 2146 9767
rect 2146 9733 2152 9767
rect 2218 9733 2224 9767
rect 2224 9733 2252 9767
rect 2318 9733 2352 9767
rect 2418 9733 2452 9767
rect 2518 9733 2552 9767
rect 2618 9733 2652 9767
rect 2718 9733 2746 9767
rect 2746 9733 2752 9767
rect 2818 9733 2824 9767
rect 2824 9733 2852 9767
rect 2918 9733 2952 9767
rect 3018 9733 3052 9767
rect 3118 9733 3152 9767
rect 3218 9733 3246 9767
rect 3246 9733 3252 9767
rect 3318 9733 3324 9767
rect 3324 9733 3352 9767
rect 3418 9733 3452 9767
rect 3518 9733 3546 9767
rect 3546 9733 3552 9767
rect 3618 9733 3624 9767
rect 3624 9733 3652 9767
rect 3718 9733 3752 9767
rect 3818 9733 3852 9767
rect 3918 9733 3952 9767
rect 4018 9733 4052 9767
rect 4118 9733 4152 9767
rect 4218 9733 4252 9767
rect 4318 9733 4352 9767
rect 4418 9733 4452 9767
rect 4518 9733 4552 9767
rect 4618 9733 4652 9767
rect 4718 9733 4752 9767
rect 4818 9733 4852 9767
rect 4918 9733 4952 9767
rect 5018 9733 5052 9767
rect 5118 9733 5152 9767
rect 5218 9733 5252 9767
rect 5318 9733 5352 9767
rect 5418 9733 5446 9767
rect 5446 9733 5452 9767
rect 5518 9733 5524 9767
rect 5524 9733 5552 9767
rect 5618 9733 5652 9767
rect 5718 9733 5746 9767
rect 5746 9733 5752 9767
rect 5818 9733 5824 9767
rect 5824 9733 5852 9767
rect 5918 9733 5946 9767
rect 5946 9733 5952 9767
rect 6018 9733 6024 9767
rect 6024 9733 6052 9767
rect 6118 9733 6152 9767
rect 6218 9733 6252 9767
rect 6318 9733 6352 9767
rect 6418 9733 6446 9767
rect 6446 9733 6452 9767
rect 6516 9748 6524 9782
rect 6524 9748 6550 9782
rect 6720 9718 6746 9752
rect 6746 9718 6754 9752
rect 18 9593 52 9627
rect 118 9593 152 9627
rect 218 9593 252 9627
rect 318 9593 352 9627
rect 418 9593 452 9627
rect 518 9593 552 9627
rect 618 9593 646 9627
rect 646 9593 652 9627
rect 718 9593 724 9627
rect 724 9593 752 9627
rect 818 9593 852 9627
rect 918 9593 952 9627
rect 1018 9593 1052 9627
rect 1118 9593 1152 9627
rect 1218 9593 1252 9627
rect 1318 9593 1352 9627
rect 1418 9593 1452 9627
rect 1518 9593 1552 9627
rect 1618 9593 1652 9627
rect 1718 9593 1752 9627
rect 1818 9593 1852 9627
rect 1918 9593 1952 9627
rect 2018 9593 2052 9627
rect 2118 9593 2146 9627
rect 2146 9593 2152 9627
rect 2218 9593 2224 9627
rect 2224 9593 2252 9627
rect 2318 9593 2346 9627
rect 2346 9593 2352 9627
rect 2418 9593 2424 9627
rect 2424 9593 2452 9627
rect 2518 9593 2552 9627
rect 2618 9593 2652 9627
rect 2718 9593 2752 9627
rect 2818 9593 2852 9627
rect 2918 9593 2946 9627
rect 2946 9593 2952 9627
rect 3018 9593 3024 9627
rect 3024 9593 3052 9627
rect 3118 9593 3152 9627
rect 3218 9593 3252 9627
rect 3318 9593 3352 9627
rect 3418 9593 3452 9627
rect 3518 9593 3552 9627
rect 3618 9593 3652 9627
rect 3718 9593 3752 9627
rect 3818 9593 3852 9627
rect 3918 9593 3952 9627
rect 4018 9593 4046 9627
rect 4046 9593 4052 9627
rect 4118 9593 4124 9627
rect 4124 9593 4152 9627
rect 4218 9593 4252 9627
rect 4318 9593 4352 9627
rect 4418 9593 4452 9627
rect 4518 9593 4552 9627
rect 4618 9593 4652 9627
rect 4718 9593 4752 9627
rect 4818 9593 4852 9627
rect 4918 9593 4952 9627
rect 5018 9593 5052 9627
rect 5118 9593 5152 9627
rect 5218 9593 5252 9627
rect 5318 9593 5352 9627
rect 5418 9593 5452 9627
rect 5518 9593 5552 9627
rect 5618 9593 5652 9627
rect 5718 9593 5752 9627
rect 5818 9593 5852 9627
rect 5918 9593 5946 9627
rect 5946 9593 5952 9627
rect 6018 9593 6024 9627
rect 6024 9593 6052 9627
rect 6118 9593 6152 9627
rect 6218 9593 6252 9627
rect 6318 9593 6352 9627
rect 6418 9593 6446 9627
rect 6446 9593 6452 9627
rect 6516 9608 6524 9642
rect 6524 9608 6550 9642
rect 6720 9578 6746 9612
rect 6746 9578 6754 9612
rect 18 9453 52 9487
rect 118 9453 152 9487
rect 218 9453 252 9487
rect 318 9453 352 9487
rect 418 9453 446 9487
rect 446 9453 452 9487
rect 518 9453 524 9487
rect 524 9453 552 9487
rect 618 9453 652 9487
rect 718 9453 752 9487
rect 818 9453 852 9487
rect 918 9453 946 9487
rect 946 9453 952 9487
rect 1018 9453 1024 9487
rect 1024 9453 1052 9487
rect 1118 9453 1146 9487
rect 1146 9453 1152 9487
rect 1218 9453 1224 9487
rect 1224 9453 1252 9487
rect 1318 9453 1352 9487
rect 1418 9453 1452 9487
rect 1518 9453 1552 9487
rect 1618 9453 1652 9487
rect 1718 9453 1746 9487
rect 1746 9453 1752 9487
rect 1818 9453 1824 9487
rect 1824 9453 1852 9487
rect 1918 9453 1952 9487
rect 2018 9453 2046 9487
rect 2046 9453 2052 9487
rect 2118 9453 2124 9487
rect 2124 9453 2152 9487
rect 2218 9453 2252 9487
rect 2318 9453 2346 9487
rect 2346 9453 2352 9487
rect 2418 9453 2424 9487
rect 2424 9453 2452 9487
rect 2518 9453 2546 9487
rect 2546 9453 2552 9487
rect 2618 9453 2624 9487
rect 2624 9453 2652 9487
rect 2718 9453 2746 9487
rect 2746 9453 2752 9487
rect 2818 9453 2824 9487
rect 2824 9453 2852 9487
rect 2918 9453 2952 9487
rect 3018 9453 3052 9487
rect 3118 9453 3152 9487
rect 3218 9453 3252 9487
rect 3318 9453 3352 9487
rect 3418 9453 3452 9487
rect 3518 9453 3552 9487
rect 3618 9453 3652 9487
rect 3718 9453 3752 9487
rect 3818 9453 3852 9487
rect 3918 9453 3952 9487
rect 4018 9453 4046 9487
rect 4046 9453 4052 9487
rect 4118 9453 4124 9487
rect 4124 9453 4152 9487
rect 4218 9453 4252 9487
rect 4318 9453 4352 9487
rect 4418 9453 4452 9487
rect 4518 9453 4546 9487
rect 4546 9453 4552 9487
rect 4618 9453 4624 9487
rect 4624 9453 4652 9487
rect 4718 9453 4752 9487
rect 4818 9453 4846 9487
rect 4846 9453 4852 9487
rect 4918 9453 4924 9487
rect 4924 9453 4952 9487
rect 5018 9453 5046 9487
rect 5046 9453 5052 9487
rect 5118 9453 5124 9487
rect 5124 9453 5152 9487
rect 5218 9453 5246 9487
rect 5246 9453 5252 9487
rect 5318 9453 5324 9487
rect 5324 9453 5352 9487
rect 5418 9453 5452 9487
rect 5518 9453 5552 9487
rect 5618 9453 5646 9487
rect 5646 9453 5652 9487
rect 5718 9453 5724 9487
rect 5724 9453 5752 9487
rect 5818 9453 5846 9487
rect 5846 9453 5852 9487
rect 5918 9453 5924 9487
rect 5924 9453 5952 9487
rect 6018 9453 6052 9487
rect 6118 9453 6146 9487
rect 6146 9453 6152 9487
rect 6218 9453 6224 9487
rect 6224 9453 6252 9487
rect 6318 9453 6352 9487
rect 6418 9453 6446 9487
rect 6446 9453 6452 9487
rect 6516 9468 6524 9502
rect 6524 9468 6550 9502
rect 6720 9438 6746 9472
rect 6746 9438 6754 9472
rect 18 9313 52 9347
rect 118 9313 152 9347
rect 218 9313 252 9347
rect 318 9313 352 9347
rect 418 9313 452 9347
rect 518 9313 552 9347
rect 618 9313 652 9347
rect 718 9313 752 9347
rect 818 9313 852 9347
rect 918 9313 952 9347
rect 1018 9313 1052 9347
rect 1118 9313 1152 9347
rect 1218 9313 1252 9347
rect 1318 9313 1352 9347
rect 1418 9313 1452 9347
rect 1518 9313 1552 9347
rect 1618 9313 1652 9347
rect 1718 9313 1746 9347
rect 1746 9313 1752 9347
rect 1818 9313 1824 9347
rect 1824 9313 1852 9347
rect 1918 9313 1952 9347
rect 2018 9313 2052 9347
rect 2118 9313 2152 9347
rect 2218 9313 2252 9347
rect 2318 9313 2352 9347
rect 2418 9313 2452 9347
rect 2518 9313 2552 9347
rect 2618 9313 2652 9347
rect 2718 9313 2752 9347
rect 2818 9313 2852 9347
rect 2918 9313 2952 9347
rect 3018 9313 3052 9347
rect 3118 9313 3152 9347
rect 3218 9313 3252 9347
rect 3318 9313 3352 9347
rect 3418 9313 3452 9347
rect 3518 9313 3552 9347
rect 3618 9313 3652 9347
rect 3718 9313 3752 9347
rect 3818 9313 3852 9347
rect 3918 9313 3952 9347
rect 4018 9313 4052 9347
rect 4118 9313 4146 9347
rect 4146 9313 4152 9347
rect 4218 9313 4224 9347
rect 4224 9313 4252 9347
rect 4318 9313 4352 9347
rect 4418 9313 4452 9347
rect 4518 9313 4552 9347
rect 4618 9313 4652 9347
rect 4718 9313 4752 9347
rect 4818 9313 4852 9347
rect 4918 9313 4952 9347
rect 5018 9313 5052 9347
rect 5118 9313 5152 9347
rect 5218 9313 5252 9347
rect 5318 9313 5352 9347
rect 5418 9313 5452 9347
rect 5518 9313 5552 9347
rect 5618 9313 5652 9347
rect 5718 9313 5752 9347
rect 5818 9313 5852 9347
rect 5918 9313 5952 9347
rect 6018 9313 6052 9347
rect 6118 9313 6152 9347
rect 6218 9313 6252 9347
rect 6318 9313 6352 9347
rect 6418 9313 6446 9347
rect 6446 9313 6452 9347
rect 6516 9328 6524 9362
rect 6524 9328 6550 9362
rect 6720 9298 6746 9332
rect 6746 9298 6754 9332
rect 18 9173 24 9207
rect 24 9173 52 9207
rect 118 9173 152 9207
rect 218 9173 252 9207
rect 318 9173 352 9207
rect 418 9173 452 9207
rect 518 9173 552 9207
rect 618 9173 652 9207
rect 718 9173 752 9207
rect 818 9173 852 9207
rect 918 9173 952 9207
rect 1018 9173 1052 9207
rect 1118 9173 1152 9207
rect 1218 9173 1252 9207
rect 1318 9173 1352 9207
rect 1418 9173 1452 9207
rect 1518 9173 1546 9207
rect 1546 9173 1552 9207
rect 1618 9173 1624 9207
rect 1624 9173 1652 9207
rect 1718 9173 1752 9207
rect 1818 9173 1852 9207
rect 1918 9173 1952 9207
rect 2018 9173 2052 9207
rect 2118 9173 2152 9207
rect 2218 9173 2252 9207
rect 2318 9173 2352 9207
rect 2418 9173 2446 9207
rect 2446 9173 2452 9207
rect 2518 9173 2524 9207
rect 2524 9173 2552 9207
rect 2618 9173 2652 9207
rect 2718 9173 2752 9207
rect 2818 9173 2852 9207
rect 2918 9173 2952 9207
rect 3018 9173 3052 9207
rect 3118 9173 3152 9207
rect 3218 9173 3252 9207
rect 3318 9173 3352 9207
rect 3418 9173 3452 9207
rect 3518 9173 3552 9207
rect 3618 9173 3652 9207
rect 3718 9173 3752 9207
rect 3818 9173 3852 9207
rect 3918 9173 3952 9207
rect 4018 9173 4046 9207
rect 4046 9173 4052 9207
rect 4118 9173 4124 9207
rect 4124 9173 4152 9207
rect 4218 9173 4252 9207
rect 4318 9173 4352 9207
rect 4418 9173 4452 9207
rect 4518 9173 4552 9207
rect 4618 9173 4652 9207
rect 4718 9173 4752 9207
rect 4818 9173 4852 9207
rect 4918 9173 4952 9207
rect 5018 9173 5046 9207
rect 5046 9173 5052 9207
rect 5118 9173 5124 9207
rect 5124 9173 5152 9207
rect 5218 9173 5252 9207
rect 5318 9173 5352 9207
rect 5418 9173 5446 9207
rect 5446 9173 5452 9207
rect 5518 9173 5524 9207
rect 5524 9173 5552 9207
rect 5618 9173 5652 9207
rect 5718 9173 5746 9207
rect 5746 9173 5752 9207
rect 5818 9173 5824 9207
rect 5824 9173 5852 9207
rect 5918 9173 5952 9207
rect 6018 9173 6052 9207
rect 6118 9173 6152 9207
rect 6218 9173 6252 9207
rect 6318 9173 6352 9207
rect 6418 9173 6452 9207
rect 6516 9188 6524 9222
rect 6524 9188 6550 9222
rect 6720 9158 6746 9192
rect 6746 9158 6754 9192
rect 18 9033 52 9067
rect 118 9033 152 9067
rect 218 9033 252 9067
rect 318 9033 352 9067
rect 418 9033 452 9067
rect 518 9033 552 9067
rect 618 9033 646 9067
rect 646 9033 652 9067
rect 718 9033 724 9067
rect 724 9033 752 9067
rect 818 9033 852 9067
rect 918 9033 952 9067
rect 1018 9033 1052 9067
rect 1118 9033 1152 9067
rect 1218 9033 1252 9067
rect 1318 9033 1352 9067
rect 1418 9033 1452 9067
rect 1518 9033 1552 9067
rect 1618 9033 1652 9067
rect 1718 9033 1746 9067
rect 1746 9033 1752 9067
rect 1818 9033 1824 9067
rect 1824 9033 1852 9067
rect 1918 9033 1946 9067
rect 1946 9033 1952 9067
rect 2018 9033 2024 9067
rect 2024 9033 2052 9067
rect 2118 9033 2152 9067
rect 2218 9033 2252 9067
rect 2318 9033 2352 9067
rect 2418 9033 2452 9067
rect 2518 9033 2552 9067
rect 2618 9033 2646 9067
rect 2646 9033 2652 9067
rect 2718 9033 2724 9067
rect 2724 9033 2752 9067
rect 2818 9033 2846 9067
rect 2846 9033 2852 9067
rect 2918 9033 2924 9067
rect 2924 9033 2952 9067
rect 3018 9033 3052 9067
rect 3118 9033 3152 9067
rect 3218 9033 3246 9067
rect 3246 9033 3252 9067
rect 3318 9033 3324 9067
rect 3324 9033 3352 9067
rect 3418 9033 3452 9067
rect 3518 9033 3552 9067
rect 3618 9033 3652 9067
rect 3718 9033 3752 9067
rect 3818 9033 3852 9067
rect 3918 9033 3952 9067
rect 4018 9033 4052 9067
rect 4118 9033 4152 9067
rect 4218 9033 4252 9067
rect 4318 9033 4352 9067
rect 4418 9033 4452 9067
rect 4518 9033 4546 9067
rect 4546 9033 4552 9067
rect 4618 9033 4624 9067
rect 4624 9033 4652 9067
rect 4718 9033 4746 9067
rect 4746 9033 4752 9067
rect 4818 9033 4824 9067
rect 4824 9033 4852 9067
rect 4918 9033 4952 9067
rect 5018 9033 5052 9067
rect 5118 9033 5152 9067
rect 5218 9033 5246 9067
rect 5246 9033 5252 9067
rect 5318 9033 5324 9067
rect 5324 9033 5352 9067
rect 5418 9033 5452 9067
rect 5518 9033 5552 9067
rect 5618 9033 5652 9067
rect 5718 9033 5752 9067
rect 5818 9033 5852 9067
rect 5918 9033 5952 9067
rect 6018 9033 6052 9067
rect 6118 9033 6152 9067
rect 6218 9033 6252 9067
rect 6318 9033 6352 9067
rect 6418 9033 6446 9067
rect 6446 9033 6452 9067
rect 6516 9048 6524 9082
rect 6524 9048 6550 9082
rect 6720 9018 6746 9052
rect 6746 9018 6754 9052
rect 18 8893 52 8927
rect 118 8893 152 8927
rect 218 8893 252 8927
rect 318 8893 352 8927
rect 418 8893 452 8927
rect 518 8893 552 8927
rect 618 8893 652 8927
rect 718 8893 752 8927
rect 818 8893 852 8927
rect 918 8893 952 8927
rect 1018 8893 1052 8927
rect 1118 8893 1152 8927
rect 1218 8893 1252 8927
rect 1318 8893 1352 8927
rect 1418 8893 1452 8927
rect 1518 8893 1552 8927
rect 1618 8893 1652 8927
rect 1718 8893 1752 8927
rect 1818 8893 1852 8927
rect 1918 8893 1952 8927
rect 2018 8893 2052 8927
rect 2118 8893 2152 8927
rect 2218 8893 2252 8927
rect 2318 8893 2352 8927
rect 2418 8893 2452 8927
rect 2518 8893 2552 8927
rect 2618 8893 2646 8927
rect 2646 8893 2652 8927
rect 2718 8893 2724 8927
rect 2724 8893 2752 8927
rect 2818 8893 2852 8927
rect 2918 8893 2952 8927
rect 3018 8893 3052 8927
rect 3118 8893 3152 8927
rect 3218 8893 3252 8927
rect 3318 8893 3352 8927
rect 3418 8893 3452 8927
rect 3518 8893 3552 8927
rect 3618 8893 3652 8927
rect 3718 8893 3752 8927
rect 3818 8893 3852 8927
rect 3918 8893 3952 8927
rect 4018 8893 4052 8927
rect 4118 8893 4152 8927
rect 4218 8893 4252 8927
rect 4318 8893 4352 8927
rect 4418 8893 4446 8927
rect 4446 8893 4452 8927
rect 4518 8893 4524 8927
rect 4524 8893 4552 8927
rect 4618 8893 4646 8927
rect 4646 8893 4652 8927
rect 4718 8893 4724 8927
rect 4724 8893 4752 8927
rect 4818 8893 4846 8927
rect 4846 8893 4852 8927
rect 4918 8893 4924 8927
rect 4924 8893 4952 8927
rect 5018 8893 5052 8927
rect 5118 8893 5152 8927
rect 5218 8893 5252 8927
rect 5318 8893 5352 8927
rect 5418 8893 5452 8927
rect 5518 8893 5552 8927
rect 5618 8893 5646 8927
rect 5646 8893 5652 8927
rect 5718 8893 5724 8927
rect 5724 8893 5752 8927
rect 5818 8893 5852 8927
rect 5918 8893 5952 8927
rect 6018 8893 6052 8927
rect 6118 8893 6146 8927
rect 6146 8893 6152 8927
rect 6218 8893 6224 8927
rect 6224 8893 6252 8927
rect 6318 8893 6352 8927
rect 6418 8893 6452 8927
rect 6516 8908 6524 8942
rect 6524 8908 6550 8942
rect 6720 8878 6746 8912
rect 6746 8878 6754 8912
rect 18 8753 24 8787
rect 24 8753 52 8787
rect 118 8753 152 8787
rect 218 8753 246 8787
rect 246 8753 252 8787
rect 318 8753 324 8787
rect 324 8753 352 8787
rect 418 8753 452 8787
rect 518 8753 552 8787
rect 618 8753 652 8787
rect 718 8753 752 8787
rect 818 8753 852 8787
rect 918 8753 952 8787
rect 1018 8753 1052 8787
rect 1118 8753 1152 8787
rect 1218 8753 1252 8787
rect 1318 8753 1352 8787
rect 1418 8753 1452 8787
rect 1518 8753 1552 8787
rect 1618 8753 1652 8787
rect 1718 8753 1752 8787
rect 1818 8753 1852 8787
rect 1918 8753 1952 8787
rect 2018 8753 2052 8787
rect 2118 8753 2152 8787
rect 2218 8753 2252 8787
rect 2318 8753 2352 8787
rect 2418 8753 2452 8787
rect 2518 8753 2552 8787
rect 2618 8753 2646 8787
rect 2646 8753 2652 8787
rect 2718 8753 2724 8787
rect 2724 8753 2752 8787
rect 2818 8753 2852 8787
rect 2918 8753 2952 8787
rect 3018 8753 3052 8787
rect 3118 8753 3146 8787
rect 3146 8753 3152 8787
rect 3218 8753 3224 8787
rect 3224 8753 3252 8787
rect 3318 8753 3352 8787
rect 3418 8753 3452 8787
rect 3518 8753 3552 8787
rect 3618 8753 3652 8787
rect 3718 8753 3752 8787
rect 3818 8753 3852 8787
rect 3918 8753 3952 8787
rect 4018 8753 4052 8787
rect 4118 8753 4152 8787
rect 4218 8753 4252 8787
rect 4318 8753 4352 8787
rect 4418 8753 4452 8787
rect 4518 8753 4552 8787
rect 4618 8753 4652 8787
rect 4718 8753 4752 8787
rect 4818 8753 4852 8787
rect 4918 8753 4952 8787
rect 5018 8753 5052 8787
rect 5118 8753 5152 8787
rect 5218 8753 5252 8787
rect 5318 8753 5352 8787
rect 5418 8753 5452 8787
rect 5518 8753 5546 8787
rect 5546 8753 5552 8787
rect 5618 8753 5624 8787
rect 5624 8753 5652 8787
rect 5718 8753 5752 8787
rect 5818 8753 5852 8787
rect 5918 8753 5946 8787
rect 5946 8753 5952 8787
rect 6018 8753 6024 8787
rect 6024 8753 6052 8787
rect 6118 8753 6152 8787
rect 6218 8753 6252 8787
rect 6318 8753 6352 8787
rect 6418 8753 6452 8787
rect 6516 8768 6524 8802
rect 6524 8768 6550 8802
rect 6720 8738 6746 8772
rect 6746 8738 6754 8772
rect 18 8630 52 8664
rect 218 8646 252 8680
rect 418 8630 452 8664
rect 618 8646 652 8680
rect 818 8630 852 8664
rect 1018 8646 1052 8680
rect 1218 8630 1252 8664
rect 1418 8646 1452 8680
rect 1618 8630 1652 8664
rect 1818 8646 1852 8680
rect 2018 8630 2052 8664
rect 2218 8646 2252 8680
rect 2418 8630 2452 8664
rect 2618 8646 2652 8680
rect 2818 8630 2852 8664
rect 3018 8646 3052 8680
rect 3218 8630 3252 8664
rect 3418 8646 3452 8680
rect 3618 8630 3652 8664
rect 3818 8646 3852 8680
rect 4018 8630 4052 8664
rect 4218 8646 4252 8680
rect 4418 8630 4452 8664
rect 4618 8646 4652 8680
rect 4818 8630 4852 8664
rect 5018 8646 5052 8680
rect 5218 8630 5252 8664
rect 5418 8646 5452 8680
rect 5618 8630 5652 8664
rect 5818 8646 5852 8680
rect 6018 8630 6052 8664
rect 6218 8646 6252 8680
rect 6516 8627 6550 8661
rect 6720 8649 6754 8683
rect 6878 8644 6912 8678
rect 6978 8644 7012 8678
rect 7078 8644 7112 8678
rect 7178 8644 7212 8678
rect 7278 8644 7312 8678
rect 7378 8644 7412 8678
rect 18 8523 52 8557
rect 118 8523 152 8557
rect 218 8523 252 8557
rect 318 8523 352 8557
rect 418 8523 452 8557
rect 518 8523 552 8557
rect 618 8523 652 8557
rect 718 8523 752 8557
rect 818 8523 846 8557
rect 846 8523 852 8557
rect 918 8523 924 8557
rect 924 8523 952 8557
rect 1018 8523 1046 8557
rect 1046 8523 1052 8557
rect 1118 8523 1124 8557
rect 1124 8523 1152 8557
rect 1218 8523 1252 8557
rect 1318 8523 1352 8557
rect 1418 8523 1452 8557
rect 1518 8523 1552 8557
rect 1618 8523 1652 8557
rect 1718 8523 1752 8557
rect 1818 8523 1852 8557
rect 1918 8523 1952 8557
rect 2018 8523 2052 8557
rect 2118 8523 2152 8557
rect 2218 8523 2252 8557
rect 2318 8523 2352 8557
rect 2418 8523 2452 8557
rect 2518 8523 2552 8557
rect 2618 8523 2652 8557
rect 2718 8523 2746 8557
rect 2746 8523 2752 8557
rect 2818 8523 2824 8557
rect 2824 8523 2852 8557
rect 2918 8523 2952 8557
rect 3018 8523 3052 8557
rect 3118 8523 3152 8557
rect 3218 8523 3252 8557
rect 3318 8523 3346 8557
rect 3346 8523 3352 8557
rect 3418 8523 3424 8557
rect 3424 8523 3452 8557
rect 3518 8523 3546 8557
rect 3546 8523 3552 8557
rect 3618 8523 3624 8557
rect 3624 8523 3652 8557
rect 3718 8523 3752 8557
rect 3818 8523 3852 8557
rect 3918 8523 3952 8557
rect 4018 8523 4046 8557
rect 4046 8523 4052 8557
rect 4118 8523 4124 8557
rect 4124 8523 4152 8557
rect 4218 8523 4252 8557
rect 4318 8523 4346 8557
rect 4346 8523 4352 8557
rect 4418 8523 4424 8557
rect 4424 8523 4452 8557
rect 4518 8523 4552 8557
rect 4618 8523 4652 8557
rect 4718 8523 4746 8557
rect 4746 8523 4752 8557
rect 4818 8523 4824 8557
rect 4824 8523 4852 8557
rect 4918 8523 4952 8557
rect 5018 8523 5052 8557
rect 5118 8523 5152 8557
rect 5218 8523 5252 8557
rect 5318 8523 5352 8557
rect 5418 8523 5452 8557
rect 5518 8523 5552 8557
rect 5618 8523 5646 8557
rect 5646 8523 5652 8557
rect 5718 8523 5724 8557
rect 5724 8523 5752 8557
rect 5818 8523 5852 8557
rect 5918 8523 5952 8557
rect 6018 8523 6052 8557
rect 6118 8523 6152 8557
rect 6218 8523 6252 8557
rect 6318 8523 6352 8557
rect 6418 8523 6452 8557
rect 6516 8538 6524 8572
rect 6524 8538 6550 8572
rect 6720 8508 6746 8542
rect 6746 8508 6754 8542
rect 18 8383 24 8417
rect 24 8383 52 8417
rect 118 8383 152 8417
rect 218 8383 252 8417
rect 318 8383 352 8417
rect 418 8383 452 8417
rect 518 8383 552 8417
rect 618 8383 652 8417
rect 718 8383 752 8417
rect 818 8383 852 8417
rect 918 8383 952 8417
rect 1018 8383 1052 8417
rect 1118 8383 1152 8417
rect 1218 8383 1252 8417
rect 1318 8383 1346 8417
rect 1346 8383 1352 8417
rect 1418 8383 1424 8417
rect 1424 8383 1452 8417
rect 1518 8383 1552 8417
rect 1618 8383 1652 8417
rect 1718 8383 1752 8417
rect 1818 8383 1846 8417
rect 1846 8383 1852 8417
rect 1918 8383 1924 8417
rect 1924 8383 1952 8417
rect 2018 8383 2046 8417
rect 2046 8383 2052 8417
rect 2118 8383 2124 8417
rect 2124 8383 2152 8417
rect 2218 8383 2252 8417
rect 2318 8383 2346 8417
rect 2346 8383 2352 8417
rect 2418 8383 2424 8417
rect 2424 8383 2452 8417
rect 2518 8383 2552 8417
rect 2618 8383 2652 8417
rect 2718 8383 2752 8417
rect 2818 8383 2852 8417
rect 2918 8383 2952 8417
rect 3018 8383 3052 8417
rect 3118 8383 3152 8417
rect 3218 8383 3252 8417
rect 3318 8383 3352 8417
rect 3418 8383 3452 8417
rect 3518 8383 3552 8417
rect 3618 8383 3652 8417
rect 3718 8383 3752 8417
rect 3818 8383 3846 8417
rect 3846 8383 3852 8417
rect 3918 8383 3924 8417
rect 3924 8383 3952 8417
rect 4018 8383 4052 8417
rect 4118 8383 4152 8417
rect 4218 8383 4252 8417
rect 4318 8383 4352 8417
rect 4418 8383 4452 8417
rect 4518 8383 4552 8417
rect 4618 8383 4652 8417
rect 4718 8383 4746 8417
rect 4746 8383 4752 8417
rect 4818 8383 4824 8417
rect 4824 8383 4852 8417
rect 4918 8383 4946 8417
rect 4946 8383 4952 8417
rect 5018 8383 5024 8417
rect 5024 8383 5052 8417
rect 5118 8383 5152 8417
rect 5218 8383 5252 8417
rect 5318 8383 5352 8417
rect 5418 8383 5452 8417
rect 5518 8383 5552 8417
rect 5618 8383 5652 8417
rect 5718 8383 5752 8417
rect 5818 8383 5846 8417
rect 5846 8383 5852 8417
rect 5918 8383 5924 8417
rect 5924 8383 5952 8417
rect 6018 8383 6052 8417
rect 6118 8383 6152 8417
rect 6218 8383 6252 8417
rect 6318 8383 6352 8417
rect 6418 8383 6446 8417
rect 6446 8383 6452 8417
rect 6516 8398 6524 8432
rect 6524 8398 6550 8432
rect 6720 8368 6746 8402
rect 6746 8368 6754 8402
rect 18 8243 52 8277
rect 118 8243 152 8277
rect 218 8243 252 8277
rect 318 8243 352 8277
rect 418 8243 452 8277
rect 518 8243 552 8277
rect 618 8243 646 8277
rect 646 8243 652 8277
rect 718 8243 724 8277
rect 724 8243 752 8277
rect 818 8243 846 8277
rect 846 8243 852 8277
rect 918 8243 924 8277
rect 924 8243 952 8277
rect 1018 8243 1052 8277
rect 1118 8243 1152 8277
rect 1218 8243 1252 8277
rect 1318 8243 1352 8277
rect 1418 8243 1452 8277
rect 1518 8243 1552 8277
rect 1618 8243 1652 8277
rect 1718 8243 1752 8277
rect 1818 8243 1852 8277
rect 1918 8243 1946 8277
rect 1946 8243 1952 8277
rect 2018 8243 2024 8277
rect 2024 8243 2052 8277
rect 2118 8243 2152 8277
rect 2218 8243 2252 8277
rect 2318 8243 2346 8277
rect 2346 8243 2352 8277
rect 2418 8243 2424 8277
rect 2424 8243 2452 8277
rect 2518 8243 2546 8277
rect 2546 8243 2552 8277
rect 2618 8243 2624 8277
rect 2624 8243 2652 8277
rect 2718 8243 2752 8277
rect 2818 8243 2852 8277
rect 2918 8243 2952 8277
rect 3018 8243 3052 8277
rect 3118 8243 3146 8277
rect 3146 8243 3152 8277
rect 3218 8243 3224 8277
rect 3224 8243 3252 8277
rect 3318 8243 3352 8277
rect 3418 8243 3452 8277
rect 3518 8243 3546 8277
rect 3546 8243 3552 8277
rect 3618 8243 3624 8277
rect 3624 8243 3652 8277
rect 3718 8243 3752 8277
rect 3818 8243 3852 8277
rect 3918 8243 3952 8277
rect 4018 8243 4052 8277
rect 4118 8243 4152 8277
rect 4218 8243 4252 8277
rect 4318 8243 4352 8277
rect 4418 8243 4452 8277
rect 4518 8243 4552 8277
rect 4618 8243 4652 8277
rect 4718 8243 4752 8277
rect 4818 8243 4852 8277
rect 4918 8243 4952 8277
rect 5018 8243 5052 8277
rect 5118 8243 5152 8277
rect 5218 8243 5252 8277
rect 5318 8243 5352 8277
rect 5418 8243 5452 8277
rect 5518 8243 5552 8277
rect 5618 8243 5652 8277
rect 5718 8243 5752 8277
rect 5818 8243 5852 8277
rect 5918 8243 5952 8277
rect 6018 8243 6052 8277
rect 6118 8243 6152 8277
rect 6218 8243 6252 8277
rect 6318 8243 6352 8277
rect 6418 8243 6446 8277
rect 6446 8243 6452 8277
rect 6516 8258 6524 8292
rect 6524 8258 6550 8292
rect 6720 8228 6746 8262
rect 6746 8228 6754 8262
rect 18 8103 52 8137
rect 118 8103 152 8137
rect 218 8103 252 8137
rect 318 8103 352 8137
rect 418 8103 452 8137
rect 518 8103 552 8137
rect 618 8103 652 8137
rect 718 8103 752 8137
rect 818 8103 852 8137
rect 918 8103 952 8137
rect 1018 8103 1052 8137
rect 1118 8103 1152 8137
rect 1218 8103 1246 8137
rect 1246 8103 1252 8137
rect 1318 8103 1324 8137
rect 1324 8103 1352 8137
rect 1418 8103 1452 8137
rect 1518 8103 1552 8137
rect 1618 8103 1652 8137
rect 1718 8103 1752 8137
rect 1818 8103 1852 8137
rect 1918 8103 1952 8137
rect 2018 8103 2052 8137
rect 2118 8103 2152 8137
rect 2218 8103 2252 8137
rect 2318 8103 2352 8137
rect 2418 8103 2452 8137
rect 2518 8103 2552 8137
rect 2618 8103 2646 8137
rect 2646 8103 2652 8137
rect 2718 8103 2724 8137
rect 2724 8103 2752 8137
rect 2818 8103 2846 8137
rect 2846 8103 2852 8137
rect 2918 8103 2924 8137
rect 2924 8103 2952 8137
rect 3018 8103 3052 8137
rect 3118 8103 3152 8137
rect 3218 8103 3252 8137
rect 3318 8103 3352 8137
rect 3418 8103 3452 8137
rect 3518 8103 3552 8137
rect 3618 8103 3652 8137
rect 3718 8103 3746 8137
rect 3746 8103 3752 8137
rect 3818 8103 3824 8137
rect 3824 8103 3852 8137
rect 3918 8103 3952 8137
rect 4018 8103 4052 8137
rect 4118 8103 4152 8137
rect 4218 8103 4252 8137
rect 4318 8103 4352 8137
rect 4418 8103 4452 8137
rect 4518 8103 4552 8137
rect 4618 8103 4652 8137
rect 4718 8103 4752 8137
rect 4818 8103 4852 8137
rect 4918 8103 4952 8137
rect 5018 8103 5052 8137
rect 5118 8103 5152 8137
rect 5218 8103 5252 8137
rect 5318 8103 5352 8137
rect 5418 8103 5452 8137
rect 5518 8103 5552 8137
rect 5618 8103 5652 8137
rect 5718 8103 5752 8137
rect 5818 8103 5852 8137
rect 5918 8103 5952 8137
rect 6018 8103 6052 8137
rect 6118 8103 6152 8137
rect 6218 8103 6252 8137
rect 6318 8103 6352 8137
rect 6418 8103 6452 8137
rect 6516 8118 6524 8152
rect 6524 8118 6550 8152
rect 6720 8088 6746 8122
rect 6746 8088 6754 8122
rect 18 7963 52 7997
rect 118 7963 152 7997
rect 218 7963 246 7997
rect 246 7963 252 7997
rect 318 7963 324 7997
rect 324 7963 352 7997
rect 418 7963 452 7997
rect 518 7963 552 7997
rect 618 7963 652 7997
rect 718 7963 752 7997
rect 818 7963 852 7997
rect 918 7963 952 7997
rect 1018 7963 1046 7997
rect 1046 7963 1052 7997
rect 1118 7963 1124 7997
rect 1124 7963 1152 7997
rect 1218 7963 1252 7997
rect 1318 7963 1346 7997
rect 1346 7963 1352 7997
rect 1418 7963 1424 7997
rect 1424 7963 1452 7997
rect 1518 7963 1552 7997
rect 1618 7963 1652 7997
rect 1718 7963 1746 7997
rect 1746 7963 1752 7997
rect 1818 7963 1824 7997
rect 1824 7963 1852 7997
rect 1918 7963 1952 7997
rect 2018 7963 2046 7997
rect 2046 7963 2052 7997
rect 2118 7963 2124 7997
rect 2124 7963 2152 7997
rect 2218 7963 2252 7997
rect 2318 7963 2352 7997
rect 2418 7963 2452 7997
rect 2518 7963 2552 7997
rect 2618 7963 2652 7997
rect 2718 7963 2746 7997
rect 2746 7963 2752 7997
rect 2818 7963 2824 7997
rect 2824 7963 2852 7997
rect 2918 7963 2946 7997
rect 2946 7963 2952 7997
rect 3018 7963 3024 7997
rect 3024 7963 3052 7997
rect 3118 7963 3152 7997
rect 3218 7963 3252 7997
rect 3318 7963 3352 7997
rect 3418 7963 3452 7997
rect 3518 7963 3552 7997
rect 3618 7963 3652 7997
rect 3718 7963 3752 7997
rect 3818 7963 3852 7997
rect 3918 7963 3952 7997
rect 4018 7963 4052 7997
rect 4118 7963 4152 7997
rect 4218 7963 4252 7997
rect 4318 7963 4352 7997
rect 4418 7963 4452 7997
rect 4518 7963 4552 7997
rect 4618 7963 4652 7997
rect 4718 7963 4752 7997
rect 4818 7963 4852 7997
rect 4918 7963 4946 7997
rect 4946 7963 4952 7997
rect 5018 7963 5024 7997
rect 5024 7963 5052 7997
rect 5118 7963 5152 7997
rect 5218 7963 5252 7997
rect 5318 7963 5352 7997
rect 5418 7963 5452 7997
rect 5518 7963 5552 7997
rect 5618 7963 5652 7997
rect 5718 7963 5752 7997
rect 5818 7963 5852 7997
rect 5918 7963 5952 7997
rect 6018 7963 6052 7997
rect 6118 7963 6152 7997
rect 6218 7963 6252 7997
rect 6318 7963 6352 7997
rect 6418 7963 6452 7997
rect 6516 7978 6524 8012
rect 6524 7978 6550 8012
rect 6720 7948 6746 7982
rect 6746 7948 6754 7982
rect 18 7823 24 7857
rect 24 7823 52 7857
rect 118 7823 152 7857
rect 218 7823 252 7857
rect 318 7823 352 7857
rect 418 7823 452 7857
rect 518 7823 552 7857
rect 618 7823 646 7857
rect 646 7823 652 7857
rect 718 7823 724 7857
rect 724 7823 752 7857
rect 818 7823 846 7857
rect 846 7823 852 7857
rect 918 7823 924 7857
rect 924 7823 952 7857
rect 1018 7823 1052 7857
rect 1118 7823 1152 7857
rect 1218 7823 1252 7857
rect 1318 7823 1352 7857
rect 1418 7823 1446 7857
rect 1446 7823 1452 7857
rect 1518 7823 1524 7857
rect 1524 7823 1552 7857
rect 1618 7823 1646 7857
rect 1646 7823 1652 7857
rect 1718 7823 1724 7857
rect 1724 7823 1752 7857
rect 1818 7823 1852 7857
rect 1918 7823 1952 7857
rect 2018 7823 2052 7857
rect 2118 7823 2152 7857
rect 2218 7823 2252 7857
rect 2318 7823 2352 7857
rect 2418 7823 2452 7857
rect 2518 7823 2546 7857
rect 2546 7823 2552 7857
rect 2618 7823 2624 7857
rect 2624 7823 2652 7857
rect 2718 7823 2752 7857
rect 2818 7823 2852 7857
rect 2918 7823 2952 7857
rect 3018 7823 3052 7857
rect 3118 7823 3152 7857
rect 3218 7823 3252 7857
rect 3318 7823 3346 7857
rect 3346 7823 3352 7857
rect 3418 7823 3424 7857
rect 3424 7823 3452 7857
rect 3518 7823 3552 7857
rect 3618 7823 3652 7857
rect 3718 7823 3746 7857
rect 3746 7823 3752 7857
rect 3818 7823 3824 7857
rect 3824 7823 3852 7857
rect 3918 7823 3946 7857
rect 3946 7823 3952 7857
rect 4018 7823 4024 7857
rect 4024 7823 4052 7857
rect 4118 7823 4146 7857
rect 4146 7823 4152 7857
rect 4218 7823 4224 7857
rect 4224 7823 4252 7857
rect 4318 7823 4352 7857
rect 4418 7823 4452 7857
rect 4518 7823 4546 7857
rect 4546 7823 4552 7857
rect 4618 7823 4624 7857
rect 4624 7823 4652 7857
rect 4718 7823 4746 7857
rect 4746 7823 4752 7857
rect 4818 7823 4824 7857
rect 4824 7823 4852 7857
rect 4918 7823 4946 7857
rect 4946 7823 4952 7857
rect 5018 7823 5024 7857
rect 5024 7823 5052 7857
rect 5118 7823 5152 7857
rect 5218 7823 5252 7857
rect 5318 7823 5352 7857
rect 5418 7823 5452 7857
rect 5518 7823 5546 7857
rect 5546 7823 5552 7857
rect 5618 7823 5624 7857
rect 5624 7823 5652 7857
rect 5718 7823 5746 7857
rect 5746 7823 5752 7857
rect 5818 7823 5824 7857
rect 5824 7823 5852 7857
rect 5918 7823 5952 7857
rect 6018 7823 6052 7857
rect 6118 7823 6152 7857
rect 6218 7823 6252 7857
rect 6318 7823 6352 7857
rect 6418 7823 6446 7857
rect 6446 7823 6452 7857
rect 6516 7838 6524 7872
rect 6524 7838 6550 7872
rect 6720 7808 6746 7842
rect 6746 7808 6754 7842
rect 18 7683 24 7717
rect 24 7683 52 7717
rect 118 7683 152 7717
rect 218 7683 252 7717
rect 318 7683 352 7717
rect 418 7683 452 7717
rect 518 7683 552 7717
rect 618 7683 652 7717
rect 718 7683 752 7717
rect 818 7683 852 7717
rect 918 7683 952 7717
rect 1018 7683 1052 7717
rect 1118 7683 1152 7717
rect 1218 7683 1252 7717
rect 1318 7683 1352 7717
rect 1418 7683 1452 7717
rect 1518 7683 1546 7717
rect 1546 7683 1552 7717
rect 1618 7683 1624 7717
rect 1624 7683 1652 7717
rect 1718 7683 1746 7717
rect 1746 7683 1752 7717
rect 1818 7683 1824 7717
rect 1824 7683 1852 7717
rect 1918 7683 1952 7717
rect 2018 7683 2052 7717
rect 2118 7683 2152 7717
rect 2218 7683 2252 7717
rect 2318 7683 2352 7717
rect 2418 7683 2452 7717
rect 2518 7683 2552 7717
rect 2618 7683 2652 7717
rect 2718 7683 2746 7717
rect 2746 7683 2752 7717
rect 2818 7683 2824 7717
rect 2824 7683 2852 7717
rect 2918 7683 2952 7717
rect 3018 7683 3052 7717
rect 3118 7683 3152 7717
rect 3218 7683 3252 7717
rect 3318 7683 3352 7717
rect 3418 7683 3452 7717
rect 3518 7683 3552 7717
rect 3618 7683 3652 7717
rect 3718 7683 3752 7717
rect 3818 7683 3852 7717
rect 3918 7683 3952 7717
rect 4018 7683 4052 7717
rect 4118 7683 4146 7717
rect 4146 7683 4152 7717
rect 4218 7683 4224 7717
rect 4224 7683 4252 7717
rect 4318 7683 4346 7717
rect 4346 7683 4352 7717
rect 4418 7683 4424 7717
rect 4424 7683 4452 7717
rect 4518 7683 4552 7717
rect 4618 7683 4652 7717
rect 4718 7683 4752 7717
rect 4818 7683 4852 7717
rect 4918 7683 4952 7717
rect 5018 7683 5052 7717
rect 5118 7683 5152 7717
rect 5218 7683 5252 7717
rect 5318 7683 5352 7717
rect 5418 7683 5452 7717
rect 5518 7683 5546 7717
rect 5546 7683 5552 7717
rect 5618 7683 5624 7717
rect 5624 7683 5652 7717
rect 5718 7683 5746 7717
rect 5746 7683 5752 7717
rect 5818 7683 5824 7717
rect 5824 7683 5852 7717
rect 5918 7683 5952 7717
rect 6018 7683 6052 7717
rect 6118 7683 6152 7717
rect 6218 7683 6252 7717
rect 6318 7683 6352 7717
rect 6418 7683 6452 7717
rect 6516 7698 6524 7732
rect 6524 7698 6550 7732
rect 6720 7668 6746 7702
rect 6746 7668 6754 7702
rect 18 7543 24 7577
rect 24 7543 52 7577
rect 118 7543 152 7577
rect 218 7543 252 7577
rect 318 7543 352 7577
rect 418 7543 452 7577
rect 518 7543 552 7577
rect 618 7543 652 7577
rect 718 7543 752 7577
rect 818 7543 852 7577
rect 918 7543 952 7577
rect 1018 7543 1046 7577
rect 1046 7543 1052 7577
rect 1118 7543 1124 7577
rect 1124 7543 1152 7577
rect 1218 7543 1252 7577
rect 1318 7543 1346 7577
rect 1346 7543 1352 7577
rect 1418 7543 1424 7577
rect 1424 7543 1452 7577
rect 1518 7543 1552 7577
rect 1618 7543 1652 7577
rect 1718 7543 1752 7577
rect 1818 7543 1852 7577
rect 1918 7543 1952 7577
rect 2018 7543 2052 7577
rect 2118 7543 2152 7577
rect 2218 7543 2252 7577
rect 2318 7543 2352 7577
rect 2418 7543 2452 7577
rect 2518 7543 2552 7577
rect 2618 7543 2652 7577
rect 2718 7543 2746 7577
rect 2746 7543 2752 7577
rect 2818 7543 2824 7577
rect 2824 7543 2852 7577
rect 2918 7543 2952 7577
rect 3018 7543 3046 7577
rect 3046 7543 3052 7577
rect 3118 7543 3124 7577
rect 3124 7543 3152 7577
rect 3218 7543 3246 7577
rect 3246 7543 3252 7577
rect 3318 7543 3324 7577
rect 3324 7543 3352 7577
rect 3418 7543 3452 7577
rect 3518 7543 3552 7577
rect 3618 7543 3652 7577
rect 3718 7543 3752 7577
rect 3818 7543 3852 7577
rect 3918 7543 3946 7577
rect 3946 7543 3952 7577
rect 4018 7543 4024 7577
rect 4024 7543 4052 7577
rect 4118 7543 4152 7577
rect 4218 7543 4252 7577
rect 4318 7543 4352 7577
rect 4418 7543 4452 7577
rect 4518 7543 4552 7577
rect 4618 7543 4652 7577
rect 4718 7543 4752 7577
rect 4818 7543 4852 7577
rect 4918 7543 4946 7577
rect 4946 7543 4952 7577
rect 5018 7543 5024 7577
rect 5024 7543 5052 7577
rect 5118 7543 5146 7577
rect 5146 7543 5152 7577
rect 5218 7543 5224 7577
rect 5224 7543 5252 7577
rect 5318 7543 5352 7577
rect 5418 7543 5452 7577
rect 5518 7543 5552 7577
rect 5618 7543 5652 7577
rect 5718 7543 5752 7577
rect 5818 7543 5852 7577
rect 5918 7543 5952 7577
rect 6018 7543 6052 7577
rect 6118 7543 6152 7577
rect 6218 7543 6252 7577
rect 6318 7543 6352 7577
rect 6418 7543 6446 7577
rect 6446 7543 6452 7577
rect 6516 7558 6524 7592
rect 6524 7558 6550 7592
rect 6720 7528 6746 7562
rect 6746 7528 6754 7562
rect 18 7420 52 7454
rect 218 7436 252 7470
rect 418 7420 452 7454
rect 618 7436 652 7470
rect 818 7420 852 7454
rect 1018 7436 1052 7470
rect 1218 7420 1252 7454
rect 1418 7436 1452 7470
rect 1618 7420 1652 7454
rect 1818 7436 1852 7470
rect 2018 7420 2052 7454
rect 2218 7436 2252 7470
rect 2418 7420 2452 7454
rect 2618 7436 2652 7470
rect 2818 7420 2852 7454
rect 3018 7436 3052 7470
rect 3218 7420 3252 7454
rect 3418 7436 3452 7470
rect 3618 7420 3652 7454
rect 3818 7436 3852 7470
rect 4018 7420 4052 7454
rect 4218 7436 4252 7470
rect 4418 7420 4452 7454
rect 4618 7436 4652 7470
rect 4818 7420 4852 7454
rect 5018 7436 5052 7470
rect 5218 7420 5252 7454
rect 5418 7436 5452 7470
rect 5618 7420 5652 7454
rect 5818 7436 5852 7470
rect 6018 7420 6052 7454
rect 6218 7436 6252 7470
rect 6516 7417 6550 7451
rect 6720 7439 6754 7473
rect 6878 7434 6912 7468
rect 6978 7434 7012 7468
rect 7078 7434 7112 7468
rect 7178 7434 7212 7468
rect 7278 7434 7312 7468
rect 7378 7434 7412 7468
rect 18 7313 52 7347
rect 118 7313 152 7347
rect 218 7313 252 7347
rect 318 7313 352 7347
rect 418 7313 452 7347
rect 518 7313 552 7347
rect 618 7313 652 7347
rect 718 7313 752 7347
rect 818 7313 852 7347
rect 918 7313 952 7347
rect 1018 7313 1052 7347
rect 1118 7313 1152 7347
rect 1218 7313 1246 7347
rect 1246 7313 1252 7347
rect 1318 7313 1324 7347
rect 1324 7313 1352 7347
rect 1418 7313 1452 7347
rect 1518 7313 1546 7347
rect 1546 7313 1552 7347
rect 1618 7313 1624 7347
rect 1624 7313 1652 7347
rect 1718 7313 1752 7347
rect 1818 7313 1852 7347
rect 1918 7313 1952 7347
rect 2018 7313 2052 7347
rect 2118 7313 2146 7347
rect 2146 7313 2152 7347
rect 2218 7313 2224 7347
rect 2224 7313 2252 7347
rect 2318 7313 2346 7347
rect 2346 7313 2352 7347
rect 2418 7313 2424 7347
rect 2424 7313 2452 7347
rect 2518 7313 2546 7347
rect 2546 7313 2552 7347
rect 2618 7313 2624 7347
rect 2624 7313 2652 7347
rect 2718 7313 2752 7347
rect 2818 7313 2852 7347
rect 2918 7313 2952 7347
rect 3018 7313 3052 7347
rect 3118 7313 3152 7347
rect 3218 7313 3252 7347
rect 3318 7313 3352 7347
rect 3418 7313 3452 7347
rect 3518 7313 3552 7347
rect 3618 7313 3652 7347
rect 3718 7313 3752 7347
rect 3818 7313 3852 7347
rect 3918 7313 3952 7347
rect 4018 7313 4052 7347
rect 4118 7313 4152 7347
rect 4218 7313 4252 7347
rect 4318 7313 4352 7347
rect 4418 7313 4452 7347
rect 4518 7313 4552 7347
rect 4618 7313 4652 7347
rect 4718 7313 4752 7347
rect 4818 7313 4852 7347
rect 4918 7313 4952 7347
rect 5018 7313 5052 7347
rect 5118 7313 5152 7347
rect 5218 7313 5252 7347
rect 5318 7313 5352 7347
rect 5418 7313 5452 7347
rect 5518 7313 5552 7347
rect 5618 7313 5652 7347
rect 5718 7313 5752 7347
rect 5818 7313 5852 7347
rect 5918 7313 5952 7347
rect 6018 7313 6052 7347
rect 6118 7313 6152 7347
rect 6218 7313 6252 7347
rect 6318 7313 6352 7347
rect 6418 7313 6452 7347
rect 6516 7328 6524 7362
rect 6524 7328 6550 7362
rect 6720 7298 6746 7332
rect 6746 7298 6754 7332
rect 18 7173 52 7207
rect 118 7173 152 7207
rect 218 7173 252 7207
rect 318 7173 346 7207
rect 346 7173 352 7207
rect 418 7173 424 7207
rect 424 7173 452 7207
rect 518 7173 552 7207
rect 618 7173 652 7207
rect 718 7173 752 7207
rect 818 7173 852 7207
rect 918 7173 952 7207
rect 1018 7173 1052 7207
rect 1118 7173 1152 7207
rect 1218 7173 1252 7207
rect 1318 7173 1352 7207
rect 1418 7173 1452 7207
rect 1518 7173 1552 7207
rect 1618 7173 1652 7207
rect 1718 7173 1752 7207
rect 1818 7173 1852 7207
rect 1918 7173 1952 7207
rect 2018 7173 2052 7207
rect 2118 7173 2152 7207
rect 2218 7173 2252 7207
rect 2318 7173 2352 7207
rect 2418 7173 2452 7207
rect 2518 7173 2546 7207
rect 2546 7173 2552 7207
rect 2618 7173 2624 7207
rect 2624 7173 2652 7207
rect 2718 7173 2752 7207
rect 2818 7173 2852 7207
rect 2918 7173 2946 7207
rect 2946 7173 2952 7207
rect 3018 7173 3024 7207
rect 3024 7173 3052 7207
rect 3118 7173 3152 7207
rect 3218 7173 3246 7207
rect 3246 7173 3252 7207
rect 3318 7173 3324 7207
rect 3324 7173 3352 7207
rect 3418 7173 3452 7207
rect 3518 7173 3552 7207
rect 3618 7173 3652 7207
rect 3718 7173 3752 7207
rect 3818 7173 3852 7207
rect 3918 7173 3952 7207
rect 4018 7173 4052 7207
rect 4118 7173 4152 7207
rect 4218 7173 4252 7207
rect 4318 7173 4346 7207
rect 4346 7173 4352 7207
rect 4418 7173 4424 7207
rect 4424 7173 4452 7207
rect 4518 7173 4552 7207
rect 4618 7173 4646 7207
rect 4646 7173 4652 7207
rect 4718 7173 4724 7207
rect 4724 7173 4752 7207
rect 4818 7173 4852 7207
rect 4918 7173 4952 7207
rect 5018 7173 5046 7207
rect 5046 7173 5052 7207
rect 5118 7173 5124 7207
rect 5124 7173 5152 7207
rect 5218 7173 5252 7207
rect 5318 7173 5352 7207
rect 5418 7173 5452 7207
rect 5518 7173 5552 7207
rect 5618 7173 5652 7207
rect 5718 7173 5752 7207
rect 5818 7173 5852 7207
rect 5918 7173 5952 7207
rect 6018 7173 6046 7207
rect 6046 7173 6052 7207
rect 6118 7173 6124 7207
rect 6124 7173 6152 7207
rect 6218 7173 6252 7207
rect 6318 7173 6352 7207
rect 6418 7173 6446 7207
rect 6446 7173 6452 7207
rect 6516 7188 6524 7222
rect 6524 7188 6550 7222
rect 6720 7158 6746 7192
rect 6746 7158 6754 7192
rect 18 7033 24 7067
rect 24 7033 52 7067
rect 118 7033 152 7067
rect 218 7033 252 7067
rect 318 7033 346 7067
rect 346 7033 352 7067
rect 418 7033 424 7067
rect 424 7033 452 7067
rect 518 7033 552 7067
rect 618 7033 652 7067
rect 718 7033 752 7067
rect 818 7033 852 7067
rect 918 7033 952 7067
rect 1018 7033 1052 7067
rect 1118 7033 1152 7067
rect 1218 7033 1246 7067
rect 1246 7033 1252 7067
rect 1318 7033 1324 7067
rect 1324 7033 1352 7067
rect 1418 7033 1452 7067
rect 1518 7033 1552 7067
rect 1618 7033 1652 7067
rect 1718 7033 1752 7067
rect 1818 7033 1852 7067
rect 1918 7033 1952 7067
rect 2018 7033 2052 7067
rect 2118 7033 2152 7067
rect 2218 7033 2246 7067
rect 2246 7033 2252 7067
rect 2318 7033 2324 7067
rect 2324 7033 2352 7067
rect 2418 7033 2452 7067
rect 2518 7033 2552 7067
rect 2618 7033 2652 7067
rect 2718 7033 2752 7067
rect 2818 7033 2852 7067
rect 2918 7033 2952 7067
rect 3018 7033 3046 7067
rect 3046 7033 3052 7067
rect 3118 7033 3124 7067
rect 3124 7033 3152 7067
rect 3218 7033 3252 7067
rect 3318 7033 3352 7067
rect 3418 7033 3446 7067
rect 3446 7033 3452 7067
rect 3518 7033 3524 7067
rect 3524 7033 3552 7067
rect 3618 7033 3652 7067
rect 3718 7033 3752 7067
rect 3818 7033 3852 7067
rect 3918 7033 3952 7067
rect 4018 7033 4046 7067
rect 4046 7033 4052 7067
rect 4118 7033 4124 7067
rect 4124 7033 4152 7067
rect 4218 7033 4252 7067
rect 4318 7033 4352 7067
rect 4418 7033 4452 7067
rect 4518 7033 4552 7067
rect 4618 7033 4652 7067
rect 4718 7033 4752 7067
rect 4818 7033 4852 7067
rect 4918 7033 4952 7067
rect 5018 7033 5052 7067
rect 5118 7033 5146 7067
rect 5146 7033 5152 7067
rect 5218 7033 5224 7067
rect 5224 7033 5252 7067
rect 5318 7033 5352 7067
rect 5418 7033 5452 7067
rect 5518 7033 5552 7067
rect 5618 7033 5652 7067
rect 5718 7033 5752 7067
rect 5818 7033 5852 7067
rect 5918 7033 5952 7067
rect 6018 7033 6052 7067
rect 6118 7033 6146 7067
rect 6146 7033 6152 7067
rect 6218 7033 6224 7067
rect 6224 7033 6252 7067
rect 6318 7033 6352 7067
rect 6418 7033 6452 7067
rect 6516 7048 6524 7082
rect 6524 7048 6550 7082
rect 6720 7018 6746 7052
rect 6746 7018 6754 7052
rect 18 6893 24 6927
rect 24 6893 52 6927
rect 118 6893 152 6927
rect 218 6893 252 6927
rect 318 6893 352 6927
rect 418 6893 452 6927
rect 518 6893 552 6927
rect 618 6893 652 6927
rect 718 6893 752 6927
rect 818 6893 852 6927
rect 918 6893 952 6927
rect 1018 6893 1052 6927
rect 1118 6893 1152 6927
rect 1218 6893 1252 6927
rect 1318 6893 1352 6927
rect 1418 6893 1446 6927
rect 1446 6893 1452 6927
rect 1518 6893 1524 6927
rect 1524 6893 1552 6927
rect 1618 6893 1652 6927
rect 1718 6893 1752 6927
rect 1818 6893 1852 6927
rect 1918 6893 1952 6927
rect 2018 6893 2046 6927
rect 2046 6893 2052 6927
rect 2118 6893 2124 6927
rect 2124 6893 2152 6927
rect 2218 6893 2252 6927
rect 2318 6893 2352 6927
rect 2418 6893 2452 6927
rect 2518 6893 2552 6927
rect 2618 6893 2652 6927
rect 2718 6893 2752 6927
rect 2818 6893 2852 6927
rect 2918 6893 2946 6927
rect 2946 6893 2952 6927
rect 3018 6893 3024 6927
rect 3024 6893 3052 6927
rect 3118 6893 3146 6927
rect 3146 6893 3152 6927
rect 3218 6893 3224 6927
rect 3224 6893 3252 6927
rect 3318 6893 3352 6927
rect 3418 6893 3446 6927
rect 3446 6893 3452 6927
rect 3518 6893 3524 6927
rect 3524 6893 3552 6927
rect 3618 6893 3652 6927
rect 3718 6893 3752 6927
rect 3818 6893 3852 6927
rect 3918 6893 3952 6927
rect 4018 6893 4052 6927
rect 4118 6893 4152 6927
rect 4218 6893 4246 6927
rect 4246 6893 4252 6927
rect 4318 6893 4324 6927
rect 4324 6893 4352 6927
rect 4418 6893 4452 6927
rect 4518 6893 4552 6927
rect 4618 6893 4652 6927
rect 4718 6893 4752 6927
rect 4818 6893 4846 6927
rect 4846 6893 4852 6927
rect 4918 6893 4924 6927
rect 4924 6893 4952 6927
rect 5018 6893 5052 6927
rect 5118 6893 5146 6927
rect 5146 6893 5152 6927
rect 5218 6893 5224 6927
rect 5224 6893 5252 6927
rect 5318 6893 5346 6927
rect 5346 6893 5352 6927
rect 5418 6893 5424 6927
rect 5424 6893 5452 6927
rect 5518 6893 5552 6927
rect 5618 6893 5652 6927
rect 5718 6893 5752 6927
rect 5818 6893 5852 6927
rect 5918 6893 5952 6927
rect 6018 6893 6052 6927
rect 6118 6893 6146 6927
rect 6146 6893 6152 6927
rect 6218 6893 6224 6927
rect 6224 6893 6252 6927
rect 6318 6893 6352 6927
rect 6418 6893 6452 6927
rect 6516 6908 6524 6942
rect 6524 6908 6550 6942
rect 6720 6878 6746 6912
rect 6746 6878 6754 6912
rect 18 6753 52 6787
rect 118 6753 152 6787
rect 218 6753 252 6787
rect 318 6753 352 6787
rect 418 6753 452 6787
rect 518 6753 552 6787
rect 618 6753 652 6787
rect 718 6753 752 6787
rect 818 6753 852 6787
rect 918 6753 952 6787
rect 1018 6753 1052 6787
rect 1118 6753 1152 6787
rect 1218 6753 1252 6787
rect 1318 6753 1346 6787
rect 1346 6753 1352 6787
rect 1418 6753 1424 6787
rect 1424 6753 1452 6787
rect 1518 6753 1546 6787
rect 1546 6753 1552 6787
rect 1618 6753 1624 6787
rect 1624 6753 1652 6787
rect 1718 6753 1752 6787
rect 1818 6753 1852 6787
rect 1918 6753 1952 6787
rect 2018 6753 2052 6787
rect 2118 6753 2146 6787
rect 2146 6753 2152 6787
rect 2218 6753 2224 6787
rect 2224 6753 2252 6787
rect 2318 6753 2352 6787
rect 2418 6753 2452 6787
rect 2518 6753 2552 6787
rect 2618 6753 2652 6787
rect 2718 6753 2752 6787
rect 2818 6753 2852 6787
rect 2918 6753 2952 6787
rect 3018 6753 3052 6787
rect 3118 6753 3152 6787
rect 3218 6753 3252 6787
rect 3318 6753 3352 6787
rect 3418 6753 3452 6787
rect 3518 6753 3552 6787
rect 3618 6753 3652 6787
rect 3718 6753 3752 6787
rect 3818 6753 3852 6787
rect 3918 6753 3952 6787
rect 4018 6753 4052 6787
rect 4118 6753 4152 6787
rect 4218 6753 4252 6787
rect 4318 6753 4352 6787
rect 4418 6753 4452 6787
rect 4518 6753 4552 6787
rect 4618 6753 4652 6787
rect 4718 6753 4752 6787
rect 4818 6753 4852 6787
rect 4918 6753 4952 6787
rect 5018 6753 5052 6787
rect 5118 6753 5152 6787
rect 5218 6753 5252 6787
rect 5318 6753 5352 6787
rect 5418 6753 5446 6787
rect 5446 6753 5452 6787
rect 5518 6753 5524 6787
rect 5524 6753 5552 6787
rect 5618 6753 5646 6787
rect 5646 6753 5652 6787
rect 5718 6753 5724 6787
rect 5724 6753 5752 6787
rect 5818 6753 5846 6787
rect 5846 6753 5852 6787
rect 5918 6753 5924 6787
rect 5924 6753 5952 6787
rect 6018 6753 6052 6787
rect 6118 6753 6152 6787
rect 6218 6753 6252 6787
rect 6318 6753 6352 6787
rect 6418 6753 6452 6787
rect 6516 6768 6524 6802
rect 6524 6768 6550 6802
rect 6720 6738 6746 6772
rect 6746 6738 6754 6772
rect 18 6613 24 6647
rect 24 6613 52 6647
rect 118 6613 152 6647
rect 218 6613 246 6647
rect 246 6613 252 6647
rect 318 6613 324 6647
rect 324 6613 352 6647
rect 418 6613 452 6647
rect 518 6613 552 6647
rect 618 6613 652 6647
rect 718 6613 752 6647
rect 818 6613 852 6647
rect 918 6613 952 6647
rect 1018 6613 1046 6647
rect 1046 6613 1052 6647
rect 1118 6613 1124 6647
rect 1124 6613 1152 6647
rect 1218 6613 1246 6647
rect 1246 6613 1252 6647
rect 1318 6613 1324 6647
rect 1324 6613 1352 6647
rect 1418 6613 1452 6647
rect 1518 6613 1552 6647
rect 1618 6613 1652 6647
rect 1718 6613 1752 6647
rect 1818 6613 1852 6647
rect 1918 6613 1952 6647
rect 2018 6613 2052 6647
rect 2118 6613 2152 6647
rect 2218 6613 2252 6647
rect 2318 6613 2352 6647
rect 2418 6613 2452 6647
rect 2518 6613 2552 6647
rect 2618 6613 2652 6647
rect 2718 6613 2752 6647
rect 2818 6613 2852 6647
rect 2918 6613 2952 6647
rect 3018 6613 3052 6647
rect 3118 6613 3152 6647
rect 3218 6613 3252 6647
rect 3318 6613 3352 6647
rect 3418 6613 3446 6647
rect 3446 6613 3452 6647
rect 3518 6613 3524 6647
rect 3524 6613 3552 6647
rect 3618 6613 3646 6647
rect 3646 6613 3652 6647
rect 3718 6613 3724 6647
rect 3724 6613 3752 6647
rect 3818 6613 3852 6647
rect 3918 6613 3952 6647
rect 4018 6613 4052 6647
rect 4118 6613 4152 6647
rect 4218 6613 4252 6647
rect 4318 6613 4352 6647
rect 4418 6613 4446 6647
rect 4446 6613 4452 6647
rect 4518 6613 4524 6647
rect 4524 6613 4552 6647
rect 4618 6613 4652 6647
rect 4718 6613 4752 6647
rect 4818 6613 4852 6647
rect 4918 6613 4952 6647
rect 5018 6613 5052 6647
rect 5118 6613 5152 6647
rect 5218 6613 5252 6647
rect 5318 6613 5352 6647
rect 5418 6613 5452 6647
rect 5518 6613 5552 6647
rect 5618 6613 5652 6647
rect 5718 6613 5752 6647
rect 5818 6613 5846 6647
rect 5846 6613 5852 6647
rect 5918 6613 5924 6647
rect 5924 6613 5952 6647
rect 6018 6613 6052 6647
rect 6118 6613 6152 6647
rect 6218 6613 6252 6647
rect 6318 6613 6352 6647
rect 6418 6613 6452 6647
rect 6516 6628 6524 6662
rect 6524 6628 6550 6662
rect 6720 6598 6746 6632
rect 6746 6598 6754 6632
rect 18 6473 52 6507
rect 118 6473 152 6507
rect 218 6473 252 6507
rect 318 6473 352 6507
rect 418 6473 452 6507
rect 518 6473 546 6507
rect 546 6473 552 6507
rect 618 6473 624 6507
rect 624 6473 652 6507
rect 718 6473 752 6507
rect 818 6473 852 6507
rect 918 6473 952 6507
rect 1018 6473 1052 6507
rect 1118 6473 1152 6507
rect 1218 6473 1252 6507
rect 1318 6473 1352 6507
rect 1418 6473 1452 6507
rect 1518 6473 1552 6507
rect 1618 6473 1646 6507
rect 1646 6473 1652 6507
rect 1718 6473 1724 6507
rect 1724 6473 1752 6507
rect 1818 6473 1852 6507
rect 1918 6473 1952 6507
rect 2018 6473 2052 6507
rect 2118 6473 2152 6507
rect 2218 6473 2252 6507
rect 2318 6473 2352 6507
rect 2418 6473 2452 6507
rect 2518 6473 2552 6507
rect 2618 6473 2652 6507
rect 2718 6473 2752 6507
rect 2818 6473 2852 6507
rect 2918 6473 2952 6507
rect 3018 6473 3052 6507
rect 3118 6473 3152 6507
rect 3218 6473 3252 6507
rect 3318 6473 3352 6507
rect 3418 6473 3452 6507
rect 3518 6473 3552 6507
rect 3618 6473 3652 6507
rect 3718 6473 3746 6507
rect 3746 6473 3752 6507
rect 3818 6473 3824 6507
rect 3824 6473 3852 6507
rect 3918 6473 3952 6507
rect 4018 6473 4052 6507
rect 4118 6473 4152 6507
rect 4218 6473 4252 6507
rect 4318 6473 4352 6507
rect 4418 6473 4452 6507
rect 4518 6473 4552 6507
rect 4618 6473 4652 6507
rect 4718 6473 4752 6507
rect 4818 6473 4852 6507
rect 4918 6473 4952 6507
rect 5018 6473 5052 6507
rect 5118 6473 5146 6507
rect 5146 6473 5152 6507
rect 5218 6473 5224 6507
rect 5224 6473 5252 6507
rect 5318 6473 5346 6507
rect 5346 6473 5352 6507
rect 5418 6473 5424 6507
rect 5424 6473 5452 6507
rect 5518 6473 5552 6507
rect 5618 6473 5652 6507
rect 5718 6473 5752 6507
rect 5818 6473 5852 6507
rect 5918 6473 5952 6507
rect 6018 6473 6052 6507
rect 6118 6473 6152 6507
rect 6218 6473 6252 6507
rect 6318 6473 6352 6507
rect 6418 6473 6452 6507
rect 6516 6488 6524 6522
rect 6524 6488 6550 6522
rect 6720 6458 6746 6492
rect 6746 6458 6754 6492
rect 18 6333 24 6367
rect 24 6333 52 6367
rect 118 6333 146 6367
rect 146 6333 152 6367
rect 218 6333 224 6367
rect 224 6333 252 6367
rect 318 6333 352 6367
rect 418 6333 452 6367
rect 518 6333 552 6367
rect 618 6333 652 6367
rect 718 6333 752 6367
rect 818 6333 846 6367
rect 846 6333 852 6367
rect 918 6333 924 6367
rect 924 6333 952 6367
rect 1018 6333 1046 6367
rect 1046 6333 1052 6367
rect 1118 6333 1124 6367
rect 1124 6333 1152 6367
rect 1218 6333 1252 6367
rect 1318 6333 1352 6367
rect 1418 6333 1452 6367
rect 1518 6333 1552 6367
rect 1618 6333 1646 6367
rect 1646 6333 1652 6367
rect 1718 6333 1724 6367
rect 1724 6333 1752 6367
rect 1818 6333 1852 6367
rect 1918 6333 1946 6367
rect 1946 6333 1952 6367
rect 2018 6333 2024 6367
rect 2024 6333 2052 6367
rect 2118 6333 2152 6367
rect 2218 6333 2252 6367
rect 2318 6333 2352 6367
rect 2418 6333 2452 6367
rect 2518 6333 2552 6367
rect 2618 6333 2652 6367
rect 2718 6333 2752 6367
rect 2818 6333 2846 6367
rect 2846 6333 2852 6367
rect 2918 6333 2924 6367
rect 2924 6333 2952 6367
rect 3018 6333 3052 6367
rect 3118 6333 3152 6367
rect 3218 6333 3252 6367
rect 3318 6333 3346 6367
rect 3346 6333 3352 6367
rect 3418 6333 3424 6367
rect 3424 6333 3452 6367
rect 3518 6333 3552 6367
rect 3618 6333 3652 6367
rect 3718 6333 3752 6367
rect 3818 6333 3852 6367
rect 3918 6333 3952 6367
rect 4018 6333 4052 6367
rect 4118 6333 4152 6367
rect 4218 6333 4252 6367
rect 4318 6333 4352 6367
rect 4418 6333 4452 6367
rect 4518 6333 4552 6367
rect 4618 6333 4652 6367
rect 4718 6333 4752 6367
rect 4818 6333 4852 6367
rect 4918 6333 4952 6367
rect 5018 6333 5046 6367
rect 5046 6333 5052 6367
rect 5118 6333 5124 6367
rect 5124 6333 5152 6367
rect 5218 6333 5252 6367
rect 5318 6333 5346 6367
rect 5346 6333 5352 6367
rect 5418 6333 5424 6367
rect 5424 6333 5452 6367
rect 5518 6333 5552 6367
rect 5618 6333 5652 6367
rect 5718 6333 5752 6367
rect 5818 6333 5852 6367
rect 5918 6333 5952 6367
rect 6018 6333 6052 6367
rect 6118 6333 6146 6367
rect 6146 6333 6152 6367
rect 6218 6333 6224 6367
rect 6224 6333 6252 6367
rect 6318 6333 6352 6367
rect 6418 6333 6446 6367
rect 6446 6333 6452 6367
rect 6516 6348 6524 6382
rect 6524 6348 6550 6382
rect 6720 6318 6746 6352
rect 6746 6318 6754 6352
rect 18 6210 52 6244
rect 218 6226 252 6260
rect 418 6210 452 6244
rect 618 6226 652 6260
rect 818 6210 852 6244
rect 1018 6226 1052 6260
rect 1218 6210 1252 6244
rect 1418 6226 1452 6260
rect 1618 6210 1652 6244
rect 1818 6226 1852 6260
rect 2018 6210 2052 6244
rect 2218 6226 2252 6260
rect 2418 6210 2452 6244
rect 2618 6226 2652 6260
rect 2818 6210 2852 6244
rect 3018 6226 3052 6260
rect 3218 6210 3252 6244
rect 3418 6226 3452 6260
rect 3618 6210 3652 6244
rect 3818 6226 3852 6260
rect 4018 6210 4052 6244
rect 4218 6226 4252 6260
rect 4418 6210 4452 6244
rect 4618 6226 4652 6260
rect 4818 6210 4852 6244
rect 5018 6226 5052 6260
rect 5218 6210 5252 6244
rect 5418 6226 5452 6260
rect 5618 6210 5652 6244
rect 5818 6226 5852 6260
rect 6018 6210 6052 6244
rect 6218 6226 6252 6260
rect 6516 6207 6550 6241
rect 6720 6229 6754 6263
rect 6878 6224 6912 6258
rect 6978 6224 7012 6258
rect 7078 6224 7112 6258
rect 7178 6224 7212 6258
rect 7278 6224 7312 6258
rect 7378 6224 7412 6258
rect 18 6103 52 6137
rect 118 6103 152 6137
rect 218 6103 252 6137
rect 318 6103 352 6137
rect 418 6103 452 6137
rect 518 6103 552 6137
rect 618 6103 652 6137
rect 718 6103 752 6137
rect 818 6103 852 6137
rect 918 6103 952 6137
rect 1018 6103 1052 6137
rect 1118 6103 1152 6137
rect 1218 6103 1252 6137
rect 1318 6103 1352 6137
rect 1418 6103 1452 6137
rect 1518 6103 1552 6137
rect 1618 6103 1652 6137
rect 1718 6103 1752 6137
rect 1818 6103 1852 6137
rect 1918 6103 1952 6137
rect 2018 6103 2052 6137
rect 2118 6103 2152 6137
rect 2218 6103 2252 6137
rect 2318 6103 2352 6137
rect 2418 6103 2446 6137
rect 2446 6103 2452 6137
rect 2518 6103 2524 6137
rect 2524 6103 2552 6137
rect 2618 6103 2652 6137
rect 2718 6103 2752 6137
rect 2818 6103 2852 6137
rect 2918 6103 2952 6137
rect 3018 6103 3052 6137
rect 3118 6103 3152 6137
rect 3218 6103 3252 6137
rect 3318 6103 3352 6137
rect 3418 6103 3452 6137
rect 3518 6103 3552 6137
rect 3618 6103 3652 6137
rect 3718 6103 3746 6137
rect 3746 6103 3752 6137
rect 3818 6103 3824 6137
rect 3824 6103 3852 6137
rect 3918 6103 3952 6137
rect 4018 6103 4046 6137
rect 4046 6103 4052 6137
rect 4118 6103 4124 6137
rect 4124 6103 4152 6137
rect 4218 6103 4252 6137
rect 4318 6103 4352 6137
rect 4418 6103 4446 6137
rect 4446 6103 4452 6137
rect 4518 6103 4524 6137
rect 4524 6103 4552 6137
rect 4618 6103 4646 6137
rect 4646 6103 4652 6137
rect 4718 6103 4724 6137
rect 4724 6103 4752 6137
rect 4818 6103 4852 6137
rect 4918 6103 4952 6137
rect 5018 6103 5052 6137
rect 5118 6103 5152 6137
rect 5218 6103 5252 6137
rect 5318 6103 5352 6137
rect 5418 6103 5452 6137
rect 5518 6103 5552 6137
rect 5618 6103 5652 6137
rect 5718 6103 5752 6137
rect 5818 6103 5852 6137
rect 5918 6103 5952 6137
rect 6018 6103 6046 6137
rect 6046 6103 6052 6137
rect 6118 6103 6124 6137
rect 6124 6103 6152 6137
rect 6218 6103 6246 6137
rect 6246 6103 6252 6137
rect 6318 6103 6324 6137
rect 6324 6103 6352 6137
rect 6418 6103 6446 6137
rect 6446 6103 6452 6137
rect 6516 6118 6524 6152
rect 6524 6118 6550 6152
rect 6720 6088 6746 6122
rect 6746 6088 6754 6122
rect 18 5963 52 5997
rect 118 5963 152 5997
rect 218 5963 252 5997
rect 318 5963 352 5997
rect 418 5963 446 5997
rect 446 5963 452 5997
rect 518 5963 524 5997
rect 524 5963 552 5997
rect 618 5963 652 5997
rect 718 5963 752 5997
rect 818 5963 852 5997
rect 918 5963 952 5997
rect 1018 5963 1052 5997
rect 1118 5963 1152 5997
rect 1218 5963 1252 5997
rect 1318 5963 1346 5997
rect 1346 5963 1352 5997
rect 1418 5963 1424 5997
rect 1424 5963 1452 5997
rect 1518 5963 1552 5997
rect 1618 5963 1652 5997
rect 1718 5963 1752 5997
rect 1818 5963 1852 5997
rect 1918 5963 1952 5997
rect 2018 5963 2052 5997
rect 2118 5963 2152 5997
rect 2218 5963 2252 5997
rect 2318 5963 2352 5997
rect 2418 5963 2452 5997
rect 2518 5963 2552 5997
rect 2618 5963 2652 5997
rect 2718 5963 2752 5997
rect 2818 5963 2852 5997
rect 2918 5963 2952 5997
rect 3018 5963 3052 5997
rect 3118 5963 3152 5997
rect 3218 5963 3252 5997
rect 3318 5963 3346 5997
rect 3346 5963 3352 5997
rect 3418 5963 3424 5997
rect 3424 5963 3452 5997
rect 3518 5963 3552 5997
rect 3618 5963 3652 5997
rect 3718 5963 3752 5997
rect 3818 5963 3852 5997
rect 3918 5963 3952 5997
rect 4018 5963 4052 5997
rect 4118 5963 4152 5997
rect 4218 5963 4252 5997
rect 4318 5963 4352 5997
rect 4418 5963 4452 5997
rect 4518 5963 4552 5997
rect 4618 5963 4652 5997
rect 4718 5963 4752 5997
rect 4818 5963 4852 5997
rect 4918 5963 4952 5997
rect 5018 5963 5052 5997
rect 5118 5963 5152 5997
rect 5218 5963 5246 5997
rect 5246 5963 5252 5997
rect 5318 5963 5324 5997
rect 5324 5963 5352 5997
rect 5418 5963 5452 5997
rect 5518 5963 5552 5997
rect 5618 5963 5652 5997
rect 5718 5963 5752 5997
rect 5818 5963 5846 5997
rect 5846 5963 5852 5997
rect 5918 5963 5924 5997
rect 5924 5963 5952 5997
rect 6018 5963 6052 5997
rect 6118 5963 6152 5997
rect 6218 5963 6252 5997
rect 6318 5963 6352 5997
rect 6418 5963 6446 5997
rect 6446 5963 6452 5997
rect 6516 5978 6524 6012
rect 6524 5978 6550 6012
rect 6720 5948 6746 5982
rect 6746 5948 6754 5982
rect 18 5823 24 5857
rect 24 5823 52 5857
rect 118 5823 152 5857
rect 218 5823 252 5857
rect 318 5823 352 5857
rect 418 5823 452 5857
rect 518 5823 552 5857
rect 618 5823 652 5857
rect 718 5823 752 5857
rect 818 5823 852 5857
rect 918 5823 952 5857
rect 1018 5823 1052 5857
rect 1118 5823 1152 5857
rect 1218 5823 1252 5857
rect 1318 5823 1352 5857
rect 1418 5823 1452 5857
rect 1518 5823 1552 5857
rect 1618 5823 1652 5857
rect 1718 5823 1752 5857
rect 1818 5823 1852 5857
rect 1918 5823 1952 5857
rect 2018 5823 2046 5857
rect 2046 5823 2052 5857
rect 2118 5823 2124 5857
rect 2124 5823 2152 5857
rect 2218 5823 2252 5857
rect 2318 5823 2352 5857
rect 2418 5823 2452 5857
rect 2518 5823 2552 5857
rect 2618 5823 2652 5857
rect 2718 5823 2752 5857
rect 2818 5823 2852 5857
rect 2918 5823 2952 5857
rect 3018 5823 3052 5857
rect 3118 5823 3152 5857
rect 3218 5823 3252 5857
rect 3318 5823 3352 5857
rect 3418 5823 3446 5857
rect 3446 5823 3452 5857
rect 3518 5823 3524 5857
rect 3524 5823 3552 5857
rect 3618 5823 3652 5857
rect 3718 5823 3752 5857
rect 3818 5823 3852 5857
rect 3918 5823 3952 5857
rect 4018 5823 4052 5857
rect 4118 5823 4146 5857
rect 4146 5823 4152 5857
rect 4218 5823 4224 5857
rect 4224 5823 4252 5857
rect 4318 5823 4352 5857
rect 4418 5823 4452 5857
rect 4518 5823 4552 5857
rect 4618 5823 4652 5857
rect 4718 5823 4752 5857
rect 4818 5823 4852 5857
rect 4918 5823 4952 5857
rect 5018 5823 5052 5857
rect 5118 5823 5152 5857
rect 5218 5823 5252 5857
rect 5318 5823 5352 5857
rect 5418 5823 5452 5857
rect 5518 5823 5552 5857
rect 5618 5823 5652 5857
rect 5718 5823 5746 5857
rect 5746 5823 5752 5857
rect 5818 5823 5824 5857
rect 5824 5823 5852 5857
rect 5918 5823 5946 5857
rect 5946 5823 5952 5857
rect 6018 5823 6024 5857
rect 6024 5823 6052 5857
rect 6118 5823 6152 5857
rect 6218 5823 6252 5857
rect 6318 5823 6352 5857
rect 6418 5823 6452 5857
rect 6516 5838 6524 5872
rect 6524 5838 6550 5872
rect 6720 5808 6746 5842
rect 6746 5808 6754 5842
rect 18 5683 52 5717
rect 118 5683 152 5717
rect 218 5683 252 5717
rect 318 5683 346 5717
rect 346 5683 352 5717
rect 418 5683 424 5717
rect 424 5683 452 5717
rect 518 5683 552 5717
rect 618 5683 652 5717
rect 718 5683 752 5717
rect 818 5683 852 5717
rect 918 5683 952 5717
rect 1018 5683 1046 5717
rect 1046 5683 1052 5717
rect 1118 5683 1124 5717
rect 1124 5683 1152 5717
rect 1218 5683 1252 5717
rect 1318 5683 1352 5717
rect 1418 5683 1452 5717
rect 1518 5683 1552 5717
rect 1618 5683 1652 5717
rect 1718 5683 1752 5717
rect 1818 5683 1852 5717
rect 1918 5683 1952 5717
rect 2018 5683 2052 5717
rect 2118 5683 2152 5717
rect 2218 5683 2252 5717
rect 2318 5683 2352 5717
rect 2418 5683 2452 5717
rect 2518 5683 2552 5717
rect 2618 5683 2652 5717
rect 2718 5683 2752 5717
rect 2818 5683 2846 5717
rect 2846 5683 2852 5717
rect 2918 5683 2924 5717
rect 2924 5683 2952 5717
rect 3018 5683 3046 5717
rect 3046 5683 3052 5717
rect 3118 5683 3124 5717
rect 3124 5683 3152 5717
rect 3218 5683 3246 5717
rect 3246 5683 3252 5717
rect 3318 5683 3324 5717
rect 3324 5683 3352 5717
rect 3418 5683 3446 5717
rect 3446 5683 3452 5717
rect 3518 5683 3524 5717
rect 3524 5683 3552 5717
rect 3618 5683 3646 5717
rect 3646 5683 3652 5717
rect 3718 5683 3724 5717
rect 3724 5683 3752 5717
rect 3818 5683 3852 5717
rect 3918 5683 3952 5717
rect 4018 5683 4052 5717
rect 4118 5683 4146 5717
rect 4146 5683 4152 5717
rect 4218 5683 4224 5717
rect 4224 5683 4252 5717
rect 4318 5683 4346 5717
rect 4346 5683 4352 5717
rect 4418 5683 4424 5717
rect 4424 5683 4452 5717
rect 4518 5683 4546 5717
rect 4546 5683 4552 5717
rect 4618 5683 4624 5717
rect 4624 5683 4652 5717
rect 4718 5683 4752 5717
rect 4818 5683 4852 5717
rect 4918 5683 4952 5717
rect 5018 5683 5052 5717
rect 5118 5683 5152 5717
rect 5218 5683 5252 5717
rect 5318 5683 5352 5717
rect 5418 5683 5452 5717
rect 5518 5683 5546 5717
rect 5546 5683 5552 5717
rect 5618 5683 5624 5717
rect 5624 5683 5652 5717
rect 5718 5683 5752 5717
rect 5818 5683 5852 5717
rect 5918 5683 5952 5717
rect 6018 5683 6052 5717
rect 6118 5683 6152 5717
rect 6218 5683 6252 5717
rect 6318 5683 6352 5717
rect 6418 5683 6452 5717
rect 6516 5698 6524 5732
rect 6524 5698 6550 5732
rect 6720 5668 6746 5702
rect 6746 5668 6754 5702
rect 18 5543 52 5577
rect 118 5543 152 5577
rect 218 5543 252 5577
rect 318 5543 352 5577
rect 418 5543 452 5577
rect 518 5543 552 5577
rect 618 5543 652 5577
rect 718 5543 752 5577
rect 818 5543 852 5577
rect 918 5543 952 5577
rect 1018 5543 1052 5577
rect 1118 5543 1146 5577
rect 1146 5543 1152 5577
rect 1218 5543 1224 5577
rect 1224 5543 1252 5577
rect 1318 5543 1346 5577
rect 1346 5543 1352 5577
rect 1418 5543 1424 5577
rect 1424 5543 1452 5577
rect 1518 5543 1552 5577
rect 1618 5543 1652 5577
rect 1718 5543 1752 5577
rect 1818 5543 1852 5577
rect 1918 5543 1946 5577
rect 1946 5543 1952 5577
rect 2018 5543 2024 5577
rect 2024 5543 2052 5577
rect 2118 5543 2152 5577
rect 2218 5543 2246 5577
rect 2246 5543 2252 5577
rect 2318 5543 2324 5577
rect 2324 5543 2352 5577
rect 2418 5543 2452 5577
rect 2518 5543 2552 5577
rect 2618 5543 2652 5577
rect 2718 5543 2752 5577
rect 2818 5543 2852 5577
rect 2918 5543 2952 5577
rect 3018 5543 3052 5577
rect 3118 5543 3152 5577
rect 3218 5543 3252 5577
rect 3318 5543 3352 5577
rect 3418 5543 3452 5577
rect 3518 5543 3552 5577
rect 3618 5543 3652 5577
rect 3718 5543 3752 5577
rect 3818 5543 3852 5577
rect 3918 5543 3952 5577
rect 4018 5543 4046 5577
rect 4046 5543 4052 5577
rect 4118 5543 4124 5577
rect 4124 5543 4152 5577
rect 4218 5543 4252 5577
rect 4318 5543 4352 5577
rect 4418 5543 4452 5577
rect 4518 5543 4552 5577
rect 4618 5543 4652 5577
rect 4718 5543 4752 5577
rect 4818 5543 4852 5577
rect 4918 5543 4952 5577
rect 5018 5543 5052 5577
rect 5118 5543 5152 5577
rect 5218 5543 5252 5577
rect 5318 5543 5352 5577
rect 5418 5543 5452 5577
rect 5518 5543 5552 5577
rect 5618 5543 5652 5577
rect 5718 5543 5752 5577
rect 5818 5543 5852 5577
rect 5918 5543 5952 5577
rect 6018 5543 6052 5577
rect 6118 5543 6152 5577
rect 6218 5543 6252 5577
rect 6318 5543 6352 5577
rect 6418 5543 6452 5577
rect 6516 5558 6524 5592
rect 6524 5558 6550 5592
rect 6720 5528 6746 5562
rect 6746 5528 6754 5562
rect 18 5403 24 5437
rect 24 5403 52 5437
rect 118 5403 152 5437
rect 218 5403 252 5437
rect 318 5403 352 5437
rect 418 5403 446 5437
rect 446 5403 452 5437
rect 518 5403 524 5437
rect 524 5403 552 5437
rect 618 5403 652 5437
rect 718 5403 752 5437
rect 818 5403 852 5437
rect 918 5403 952 5437
rect 1018 5403 1052 5437
rect 1118 5403 1152 5437
rect 1218 5403 1252 5437
rect 1318 5403 1352 5437
rect 1418 5403 1446 5437
rect 1446 5403 1452 5437
rect 1518 5403 1524 5437
rect 1524 5403 1552 5437
rect 1618 5403 1652 5437
rect 1718 5403 1746 5437
rect 1746 5403 1752 5437
rect 1818 5403 1824 5437
rect 1824 5403 1852 5437
rect 1918 5403 1952 5437
rect 2018 5403 2052 5437
rect 2118 5403 2152 5437
rect 2218 5403 2246 5437
rect 2246 5403 2252 5437
rect 2318 5403 2324 5437
rect 2324 5403 2352 5437
rect 2418 5403 2452 5437
rect 2518 5403 2552 5437
rect 2618 5403 2652 5437
rect 2718 5403 2752 5437
rect 2818 5403 2852 5437
rect 2918 5403 2952 5437
rect 3018 5403 3052 5437
rect 3118 5403 3152 5437
rect 3218 5403 3252 5437
rect 3318 5403 3352 5437
rect 3418 5403 3452 5437
rect 3518 5403 3552 5437
rect 3618 5403 3652 5437
rect 3718 5403 3746 5437
rect 3746 5403 3752 5437
rect 3818 5403 3824 5437
rect 3824 5403 3852 5437
rect 3918 5403 3952 5437
rect 4018 5403 4052 5437
rect 4118 5403 4152 5437
rect 4218 5403 4252 5437
rect 4318 5403 4352 5437
rect 4418 5403 4452 5437
rect 4518 5403 4552 5437
rect 4618 5403 4652 5437
rect 4718 5403 4752 5437
rect 4818 5403 4852 5437
rect 4918 5403 4952 5437
rect 5018 5403 5052 5437
rect 5118 5403 5146 5437
rect 5146 5403 5152 5437
rect 5218 5403 5224 5437
rect 5224 5403 5252 5437
rect 5318 5403 5346 5437
rect 5346 5403 5352 5437
rect 5418 5403 5424 5437
rect 5424 5403 5452 5437
rect 5518 5403 5546 5437
rect 5546 5403 5552 5437
rect 5618 5403 5624 5437
rect 5624 5403 5652 5437
rect 5718 5403 5746 5437
rect 5746 5403 5752 5437
rect 5818 5403 5824 5437
rect 5824 5403 5852 5437
rect 5918 5403 5952 5437
rect 6018 5403 6052 5437
rect 6118 5403 6152 5437
rect 6218 5403 6252 5437
rect 6318 5403 6352 5437
rect 6418 5403 6452 5437
rect 6516 5418 6524 5452
rect 6524 5418 6550 5452
rect 6720 5388 6746 5422
rect 6746 5388 6754 5422
rect 18 5263 52 5297
rect 118 5263 152 5297
rect 218 5263 252 5297
rect 318 5263 352 5297
rect 418 5263 452 5297
rect 518 5263 552 5297
rect 618 5263 652 5297
rect 718 5263 752 5297
rect 818 5263 852 5297
rect 918 5263 952 5297
rect 1018 5263 1052 5297
rect 1118 5263 1152 5297
rect 1218 5263 1252 5297
rect 1318 5263 1352 5297
rect 1418 5263 1452 5297
rect 1518 5263 1552 5297
rect 1618 5263 1652 5297
rect 1718 5263 1752 5297
rect 1818 5263 1852 5297
rect 1918 5263 1952 5297
rect 2018 5263 2052 5297
rect 2118 5263 2146 5297
rect 2146 5263 2152 5297
rect 2218 5263 2224 5297
rect 2224 5263 2252 5297
rect 2318 5263 2346 5297
rect 2346 5263 2352 5297
rect 2418 5263 2424 5297
rect 2424 5263 2452 5297
rect 2518 5263 2552 5297
rect 2618 5263 2646 5297
rect 2646 5263 2652 5297
rect 2718 5263 2724 5297
rect 2724 5263 2752 5297
rect 2818 5263 2852 5297
rect 2918 5263 2946 5297
rect 2946 5263 2952 5297
rect 3018 5263 3024 5297
rect 3024 5263 3052 5297
rect 3118 5263 3146 5297
rect 3146 5263 3152 5297
rect 3218 5263 3224 5297
rect 3224 5263 3252 5297
rect 3318 5263 3352 5297
rect 3418 5263 3452 5297
rect 3518 5263 3552 5297
rect 3618 5263 3652 5297
rect 3718 5263 3752 5297
rect 3818 5263 3852 5297
rect 3918 5263 3952 5297
rect 4018 5263 4052 5297
rect 4118 5263 4152 5297
rect 4218 5263 4252 5297
rect 4318 5263 4352 5297
rect 4418 5263 4452 5297
rect 4518 5263 4552 5297
rect 4618 5263 4652 5297
rect 4718 5263 4752 5297
rect 4818 5263 4852 5297
rect 4918 5263 4952 5297
rect 5018 5263 5052 5297
rect 5118 5263 5152 5297
rect 5218 5263 5246 5297
rect 5246 5263 5252 5297
rect 5318 5263 5324 5297
rect 5324 5263 5352 5297
rect 5418 5263 5446 5297
rect 5446 5263 5452 5297
rect 5518 5263 5524 5297
rect 5524 5263 5552 5297
rect 5618 5263 5652 5297
rect 5718 5263 5752 5297
rect 5818 5263 5852 5297
rect 5918 5263 5952 5297
rect 6018 5263 6052 5297
rect 6118 5263 6152 5297
rect 6218 5263 6252 5297
rect 6318 5263 6352 5297
rect 6418 5263 6446 5297
rect 6446 5263 6452 5297
rect 6516 5278 6524 5312
rect 6524 5278 6550 5312
rect 6720 5248 6746 5282
rect 6746 5248 6754 5282
rect 18 5123 52 5157
rect 118 5123 152 5157
rect 218 5123 252 5157
rect 318 5123 352 5157
rect 418 5123 452 5157
rect 518 5123 552 5157
rect 618 5123 652 5157
rect 718 5123 752 5157
rect 818 5123 852 5157
rect 918 5123 952 5157
rect 1018 5123 1052 5157
rect 1118 5123 1152 5157
rect 1218 5123 1252 5157
rect 1318 5123 1346 5157
rect 1346 5123 1352 5157
rect 1418 5123 1424 5157
rect 1424 5123 1452 5157
rect 1518 5123 1552 5157
rect 1618 5123 1652 5157
rect 1718 5123 1752 5157
rect 1818 5123 1852 5157
rect 1918 5123 1952 5157
rect 2018 5123 2052 5157
rect 2118 5123 2146 5157
rect 2146 5123 2152 5157
rect 2218 5123 2224 5157
rect 2224 5123 2252 5157
rect 2318 5123 2352 5157
rect 2418 5123 2452 5157
rect 2518 5123 2552 5157
rect 2618 5123 2652 5157
rect 2718 5123 2752 5157
rect 2818 5123 2852 5157
rect 2918 5123 2952 5157
rect 3018 5123 3052 5157
rect 3118 5123 3152 5157
rect 3218 5123 3252 5157
rect 3318 5123 3352 5157
rect 3418 5123 3452 5157
rect 3518 5123 3552 5157
rect 3618 5123 3652 5157
rect 3718 5123 3752 5157
rect 3818 5123 3852 5157
rect 3918 5123 3952 5157
rect 4018 5123 4052 5157
rect 4118 5123 4152 5157
rect 4218 5123 4252 5157
rect 4318 5123 4346 5157
rect 4346 5123 4352 5157
rect 4418 5123 4424 5157
rect 4424 5123 4452 5157
rect 4518 5123 4552 5157
rect 4618 5123 4652 5157
rect 4718 5123 4746 5157
rect 4746 5123 4752 5157
rect 4818 5123 4824 5157
rect 4824 5123 4852 5157
rect 4918 5123 4952 5157
rect 5018 5123 5052 5157
rect 5118 5123 5152 5157
rect 5218 5123 5252 5157
rect 5318 5123 5352 5157
rect 5418 5123 5452 5157
rect 5518 5123 5552 5157
rect 5618 5123 5652 5157
rect 5718 5123 5746 5157
rect 5746 5123 5752 5157
rect 5818 5123 5824 5157
rect 5824 5123 5852 5157
rect 5918 5123 5952 5157
rect 6018 5123 6052 5157
rect 6118 5123 6152 5157
rect 6218 5123 6252 5157
rect 6318 5123 6352 5157
rect 6418 5123 6452 5157
rect 6516 5138 6524 5172
rect 6524 5138 6550 5172
rect 6720 5108 6746 5142
rect 6746 5108 6754 5142
rect 118 4983 152 5017
rect 318 4983 352 5017
rect 518 4983 552 5017
rect 718 4983 752 5017
rect 918 4983 952 5017
rect 1118 4983 1152 5017
rect 1318 4983 1352 5017
rect 1518 4983 1552 5017
rect 1718 4983 1752 5017
rect 1918 4983 1952 5017
rect 2118 4983 2152 5017
rect 2318 4983 2352 5017
rect 2518 4983 2552 5017
rect 2718 4983 2752 5017
rect 2918 4983 2952 5017
rect 3118 4983 3152 5017
rect 3318 4983 3352 5017
rect 3518 4983 3552 5017
rect 3718 4983 3752 5017
rect 3918 4983 3952 5017
rect 4118 4983 4152 5017
rect 4318 4983 4352 5017
rect 4518 4983 4552 5017
rect 4718 4983 4752 5017
rect 4918 4983 4952 5017
rect 5118 4983 5152 5017
rect 5318 4983 5352 5017
rect 5518 4983 5552 5017
rect 5718 4983 5752 5017
rect 5918 4983 5952 5017
rect 6118 4983 6152 5017
rect 6318 4983 6352 5017
rect 18 4860 52 4894
rect 218 4876 252 4910
rect 418 4860 452 4894
rect 618 4876 652 4910
rect 818 4860 852 4894
rect 1018 4876 1052 4910
rect 1218 4860 1252 4894
rect 1418 4876 1452 4910
rect 1618 4860 1652 4894
rect 1818 4876 1852 4910
rect 2018 4860 2052 4894
rect 2218 4876 2252 4910
rect 2418 4860 2452 4894
rect 2618 4876 2652 4910
rect 2818 4860 2852 4894
rect 3018 4876 3052 4910
rect 3218 4860 3252 4894
rect 3418 4876 3452 4910
rect 3618 4860 3652 4894
rect 3818 4876 3852 4910
rect 4018 4860 4052 4894
rect 4218 4876 4252 4910
rect 4418 4860 4452 4894
rect 4618 4876 4652 4910
rect 4818 4860 4852 4894
rect 5018 4876 5052 4910
rect 5218 4860 5252 4894
rect 5418 4876 5452 4910
rect 5618 4860 5652 4894
rect 5818 4876 5852 4910
rect 6018 4860 6052 4894
rect 6218 4876 6252 4910
rect 6516 4857 6550 4891
rect 6720 4879 6754 4913
rect 6878 4874 6912 4908
rect 6978 4874 7012 4908
rect 7078 4874 7112 4908
rect 7178 4874 7212 4908
rect 7278 4874 7312 4908
rect 7378 4874 7412 4908
rect 18 4753 24 4787
rect 24 4753 52 4787
rect 118 4753 152 4787
rect 218 4753 246 4787
rect 246 4753 252 4787
rect 318 4753 324 4787
rect 324 4753 352 4787
rect 418 4753 452 4787
rect 518 4753 552 4787
rect 618 4753 652 4787
rect 718 4753 752 4787
rect 818 4753 852 4787
rect 918 4753 952 4787
rect 1018 4753 1052 4787
rect 1118 4753 1146 4787
rect 1146 4753 1152 4787
rect 1218 4753 1224 4787
rect 1224 4753 1252 4787
rect 1318 4753 1352 4787
rect 1418 4753 1452 4787
rect 1518 4753 1552 4787
rect 1618 4753 1652 4787
rect 1718 4753 1752 4787
rect 1818 4753 1852 4787
rect 1918 4753 1952 4787
rect 2018 4753 2052 4787
rect 2118 4753 2152 4787
rect 2218 4753 2252 4787
rect 2318 4753 2352 4787
rect 2418 4753 2452 4787
rect 2518 4753 2552 4787
rect 2618 4753 2652 4787
rect 2718 4753 2752 4787
rect 2818 4753 2846 4787
rect 2846 4753 2852 4787
rect 2918 4753 2924 4787
rect 2924 4753 2952 4787
rect 3018 4753 3052 4787
rect 3118 4753 3152 4787
rect 3218 4753 3252 4787
rect 3318 4753 3352 4787
rect 3418 4753 3452 4787
rect 3518 4753 3552 4787
rect 3618 4753 3652 4787
rect 3718 4753 3752 4787
rect 3818 4753 3852 4787
rect 3918 4753 3952 4787
rect 4018 4753 4052 4787
rect 4118 4753 4152 4787
rect 4218 4753 4252 4787
rect 4318 4753 4352 4787
rect 4418 4753 4452 4787
rect 4518 4753 4552 4787
rect 4618 4753 4646 4787
rect 4646 4753 4652 4787
rect 4718 4753 4724 4787
rect 4724 4753 4752 4787
rect 4818 4753 4852 4787
rect 4918 4753 4952 4787
rect 5018 4753 5052 4787
rect 5118 4753 5152 4787
rect 5218 4753 5252 4787
rect 5318 4753 5352 4787
rect 5418 4753 5446 4787
rect 5446 4753 5452 4787
rect 5518 4753 5524 4787
rect 5524 4753 5552 4787
rect 5618 4753 5652 4787
rect 5718 4753 5752 4787
rect 5818 4753 5852 4787
rect 5918 4753 5946 4787
rect 5946 4753 5952 4787
rect 6018 4753 6024 4787
rect 6024 4753 6052 4787
rect 6118 4753 6146 4787
rect 6146 4753 6152 4787
rect 6218 4753 6224 4787
rect 6224 4753 6252 4787
rect 6318 4753 6352 4787
rect 6418 4753 6452 4787
rect 6516 4768 6524 4802
rect 6524 4768 6550 4802
rect 6720 4738 6746 4772
rect 6746 4738 6754 4772
rect 18 4613 24 4647
rect 24 4613 52 4647
rect 118 4613 152 4647
rect 218 4613 252 4647
rect 318 4613 352 4647
rect 418 4613 452 4647
rect 518 4613 552 4647
rect 618 4613 652 4647
rect 718 4613 752 4647
rect 818 4613 852 4647
rect 918 4613 952 4647
rect 1018 4613 1052 4647
rect 1118 4613 1152 4647
rect 1218 4613 1252 4647
rect 1318 4613 1352 4647
rect 1418 4613 1452 4647
rect 1518 4613 1552 4647
rect 1618 4613 1652 4647
rect 1718 4613 1752 4647
rect 1818 4613 1846 4647
rect 1846 4613 1852 4647
rect 1918 4613 1924 4647
rect 1924 4613 1952 4647
rect 2018 4613 2046 4647
rect 2046 4613 2052 4647
rect 2118 4613 2124 4647
rect 2124 4613 2152 4647
rect 2218 4613 2252 4647
rect 2318 4613 2352 4647
rect 2418 4613 2452 4647
rect 2518 4613 2552 4647
rect 2618 4613 2652 4647
rect 2718 4613 2752 4647
rect 2818 4613 2852 4647
rect 2918 4613 2952 4647
rect 3018 4613 3052 4647
rect 3118 4613 3152 4647
rect 3218 4613 3246 4647
rect 3246 4613 3252 4647
rect 3318 4613 3324 4647
rect 3324 4613 3352 4647
rect 3418 4613 3452 4647
rect 3518 4613 3552 4647
rect 3618 4613 3652 4647
rect 3718 4613 3752 4647
rect 3818 4613 3852 4647
rect 3918 4613 3952 4647
rect 4018 4613 4052 4647
rect 4118 4613 4152 4647
rect 4218 4613 4252 4647
rect 4318 4613 4352 4647
rect 4418 4613 4452 4647
rect 4518 4613 4546 4647
rect 4546 4613 4552 4647
rect 4618 4613 4624 4647
rect 4624 4613 4652 4647
rect 4718 4613 4752 4647
rect 4818 4613 4852 4647
rect 4918 4613 4952 4647
rect 5018 4613 5052 4647
rect 5118 4613 5152 4647
rect 5218 4613 5252 4647
rect 5318 4613 5352 4647
rect 5418 4613 5452 4647
rect 5518 4613 5552 4647
rect 5618 4613 5652 4647
rect 5718 4613 5752 4647
rect 5818 4613 5852 4647
rect 5918 4613 5952 4647
rect 6018 4613 6046 4647
rect 6046 4613 6052 4647
rect 6118 4613 6124 4647
rect 6124 4613 6152 4647
rect 6218 4613 6246 4647
rect 6246 4613 6252 4647
rect 6318 4613 6324 4647
rect 6324 4613 6352 4647
rect 6418 4613 6446 4647
rect 6446 4613 6452 4647
rect 6516 4628 6524 4662
rect 6524 4628 6550 4662
rect 6720 4598 6746 4632
rect 6746 4598 6754 4632
rect 18 4473 24 4507
rect 24 4473 52 4507
rect 118 4473 146 4507
rect 146 4473 152 4507
rect 218 4473 224 4507
rect 224 4473 252 4507
rect 318 4473 352 4507
rect 418 4473 452 4507
rect 518 4473 552 4507
rect 618 4473 652 4507
rect 718 4473 752 4507
rect 818 4473 852 4507
rect 918 4473 952 4507
rect 1018 4473 1052 4507
rect 1118 4473 1152 4507
rect 1218 4473 1252 4507
rect 1318 4473 1352 4507
rect 1418 4473 1452 4507
rect 1518 4473 1552 4507
rect 1618 4473 1646 4507
rect 1646 4473 1652 4507
rect 1718 4473 1724 4507
rect 1724 4473 1752 4507
rect 1818 4473 1852 4507
rect 1918 4473 1952 4507
rect 2018 4473 2052 4507
rect 2118 4473 2152 4507
rect 2218 4473 2252 4507
rect 2318 4473 2352 4507
rect 2418 4473 2446 4507
rect 2446 4473 2452 4507
rect 2518 4473 2524 4507
rect 2524 4473 2552 4507
rect 2618 4473 2652 4507
rect 2718 4473 2752 4507
rect 2818 4473 2852 4507
rect 2918 4473 2952 4507
rect 3018 4473 3052 4507
rect 3118 4473 3152 4507
rect 3218 4473 3252 4507
rect 3318 4473 3346 4507
rect 3346 4473 3352 4507
rect 3418 4473 3424 4507
rect 3424 4473 3452 4507
rect 3518 4473 3552 4507
rect 3618 4473 3652 4507
rect 3718 4473 3752 4507
rect 3818 4473 3852 4507
rect 3918 4473 3952 4507
rect 4018 4473 4052 4507
rect 4118 4473 4152 4507
rect 4218 4473 4252 4507
rect 4318 4473 4346 4507
rect 4346 4473 4352 4507
rect 4418 4473 4424 4507
rect 4424 4473 4452 4507
rect 4518 4473 4552 4507
rect 4618 4473 4652 4507
rect 4718 4473 4752 4507
rect 4818 4473 4852 4507
rect 4918 4473 4952 4507
rect 5018 4473 5052 4507
rect 5118 4473 5152 4507
rect 5218 4473 5246 4507
rect 5246 4473 5252 4507
rect 5318 4473 5324 4507
rect 5324 4473 5352 4507
rect 5418 4473 5452 4507
rect 5518 4473 5552 4507
rect 5618 4473 5652 4507
rect 5718 4473 5746 4507
rect 5746 4473 5752 4507
rect 5818 4473 5824 4507
rect 5824 4473 5852 4507
rect 5918 4473 5952 4507
rect 6018 4473 6052 4507
rect 6118 4473 6152 4507
rect 6218 4473 6246 4507
rect 6246 4473 6252 4507
rect 6318 4473 6324 4507
rect 6324 4473 6352 4507
rect 6418 4473 6446 4507
rect 6446 4473 6452 4507
rect 6516 4488 6524 4522
rect 6524 4488 6550 4522
rect 6720 4458 6746 4492
rect 6746 4458 6754 4492
rect 18 4333 24 4367
rect 24 4333 52 4367
rect 118 4333 152 4367
rect 218 4333 252 4367
rect 318 4333 352 4367
rect 418 4333 446 4367
rect 446 4333 452 4367
rect 518 4333 524 4367
rect 524 4333 552 4367
rect 618 4333 652 4367
rect 718 4333 746 4367
rect 746 4333 752 4367
rect 818 4333 824 4367
rect 824 4333 852 4367
rect 918 4333 952 4367
rect 1018 4333 1052 4367
rect 1118 4333 1152 4367
rect 1218 4333 1252 4367
rect 1318 4333 1352 4367
rect 1418 4333 1452 4367
rect 1518 4333 1552 4367
rect 1618 4333 1652 4367
rect 1718 4333 1752 4367
rect 1818 4333 1852 4367
rect 1918 4333 1952 4367
rect 2018 4333 2052 4367
rect 2118 4333 2152 4367
rect 2218 4333 2252 4367
rect 2318 4333 2352 4367
rect 2418 4333 2446 4367
rect 2446 4333 2452 4367
rect 2518 4333 2524 4367
rect 2524 4333 2552 4367
rect 2618 4333 2652 4367
rect 2718 4333 2752 4367
rect 2818 4333 2846 4367
rect 2846 4333 2852 4367
rect 2918 4333 2924 4367
rect 2924 4333 2952 4367
rect 3018 4333 3052 4367
rect 3118 4333 3152 4367
rect 3218 4333 3246 4367
rect 3246 4333 3252 4367
rect 3318 4333 3324 4367
rect 3324 4333 3352 4367
rect 3418 4333 3452 4367
rect 3518 4333 3552 4367
rect 3618 4333 3652 4367
rect 3718 4333 3752 4367
rect 3818 4333 3852 4367
rect 3918 4333 3952 4367
rect 4018 4333 4052 4367
rect 4118 4333 4152 4367
rect 4218 4333 4252 4367
rect 4318 4333 4352 4367
rect 4418 4333 4452 4367
rect 4518 4333 4552 4367
rect 4618 4333 4652 4367
rect 4718 4333 4752 4367
rect 4818 4333 4852 4367
rect 4918 4333 4952 4367
rect 5018 4333 5046 4367
rect 5046 4333 5052 4367
rect 5118 4333 5124 4367
rect 5124 4333 5152 4367
rect 5218 4333 5252 4367
rect 5318 4333 5352 4367
rect 5418 4333 5446 4367
rect 5446 4333 5452 4367
rect 5518 4333 5524 4367
rect 5524 4333 5552 4367
rect 5618 4333 5652 4367
rect 5718 4333 5752 4367
rect 5818 4333 5852 4367
rect 5918 4333 5952 4367
rect 6018 4333 6046 4367
rect 6046 4333 6052 4367
rect 6118 4333 6124 4367
rect 6124 4333 6152 4367
rect 6218 4333 6246 4367
rect 6246 4333 6252 4367
rect 6318 4333 6324 4367
rect 6324 4333 6352 4367
rect 6418 4333 6446 4367
rect 6446 4333 6452 4367
rect 6516 4348 6524 4382
rect 6524 4348 6550 4382
rect 6720 4318 6746 4352
rect 6746 4318 6754 4352
rect 18 4193 24 4227
rect 24 4193 52 4227
rect 118 4193 146 4227
rect 146 4193 152 4227
rect 218 4193 224 4227
rect 224 4193 252 4227
rect 318 4193 346 4227
rect 346 4193 352 4227
rect 418 4193 424 4227
rect 424 4193 452 4227
rect 518 4193 552 4227
rect 618 4193 652 4227
rect 718 4193 752 4227
rect 818 4193 852 4227
rect 918 4193 952 4227
rect 1018 4193 1052 4227
rect 1118 4193 1152 4227
rect 1218 4193 1252 4227
rect 1318 4193 1352 4227
rect 1418 4193 1446 4227
rect 1446 4193 1452 4227
rect 1518 4193 1524 4227
rect 1524 4193 1552 4227
rect 1618 4193 1652 4227
rect 1718 4193 1752 4227
rect 1818 4193 1852 4227
rect 1918 4193 1952 4227
rect 2018 4193 2052 4227
rect 2118 4193 2152 4227
rect 2218 4193 2252 4227
rect 2318 4193 2352 4227
rect 2418 4193 2452 4227
rect 2518 4193 2552 4227
rect 2618 4193 2652 4227
rect 2718 4193 2752 4227
rect 2818 4193 2852 4227
rect 2918 4193 2952 4227
rect 3018 4193 3052 4227
rect 3118 4193 3152 4227
rect 3218 4193 3252 4227
rect 3318 4193 3352 4227
rect 3418 4193 3446 4227
rect 3446 4193 3452 4227
rect 3518 4193 3524 4227
rect 3524 4193 3552 4227
rect 3618 4193 3646 4227
rect 3646 4193 3652 4227
rect 3718 4193 3724 4227
rect 3724 4193 3752 4227
rect 3818 4193 3852 4227
rect 3918 4193 3952 4227
rect 4018 4193 4052 4227
rect 4118 4193 4152 4227
rect 4218 4193 4252 4227
rect 4318 4193 4352 4227
rect 4418 4193 4446 4227
rect 4446 4193 4452 4227
rect 4518 4193 4524 4227
rect 4524 4193 4552 4227
rect 4618 4193 4652 4227
rect 4718 4193 4752 4227
rect 4818 4193 4852 4227
rect 4918 4193 4952 4227
rect 5018 4193 5046 4227
rect 5046 4193 5052 4227
rect 5118 4193 5124 4227
rect 5124 4193 5152 4227
rect 5218 4193 5252 4227
rect 5318 4193 5352 4227
rect 5418 4193 5446 4227
rect 5446 4193 5452 4227
rect 5518 4193 5524 4227
rect 5524 4193 5552 4227
rect 5618 4193 5652 4227
rect 5718 4193 5752 4227
rect 5818 4193 5846 4227
rect 5846 4193 5852 4227
rect 5918 4193 5924 4227
rect 5924 4193 5952 4227
rect 6018 4193 6052 4227
rect 6118 4193 6152 4227
rect 6218 4193 6252 4227
rect 6318 4193 6352 4227
rect 6418 4193 6446 4227
rect 6446 4193 6452 4227
rect 6516 4208 6524 4242
rect 6524 4208 6550 4242
rect 6720 4178 6746 4212
rect 6746 4178 6754 4212
rect 18 4053 24 4087
rect 24 4053 52 4087
rect 118 4053 152 4087
rect 218 4053 252 4087
rect 318 4053 352 4087
rect 418 4053 446 4087
rect 446 4053 452 4087
rect 518 4053 524 4087
rect 524 4053 552 4087
rect 618 4053 646 4087
rect 646 4053 652 4087
rect 718 4053 724 4087
rect 724 4053 752 4087
rect 818 4053 852 4087
rect 918 4053 952 4087
rect 1018 4053 1052 4087
rect 1118 4053 1152 4087
rect 1218 4053 1252 4087
rect 1318 4053 1352 4087
rect 1418 4053 1452 4087
rect 1518 4053 1546 4087
rect 1546 4053 1552 4087
rect 1618 4053 1624 4087
rect 1624 4053 1652 4087
rect 1718 4053 1746 4087
rect 1746 4053 1752 4087
rect 1818 4053 1824 4087
rect 1824 4053 1852 4087
rect 1918 4053 1946 4087
rect 1946 4053 1952 4087
rect 2018 4053 2024 4087
rect 2024 4053 2052 4087
rect 2118 4053 2152 4087
rect 2218 4053 2246 4087
rect 2246 4053 2252 4087
rect 2318 4053 2324 4087
rect 2324 4053 2352 4087
rect 2418 4053 2446 4087
rect 2446 4053 2452 4087
rect 2518 4053 2524 4087
rect 2524 4053 2552 4087
rect 2618 4053 2652 4087
rect 2718 4053 2752 4087
rect 2818 4053 2852 4087
rect 2918 4053 2952 4087
rect 3018 4053 3052 4087
rect 3118 4053 3152 4087
rect 3218 4053 3246 4087
rect 3246 4053 3252 4087
rect 3318 4053 3324 4087
rect 3324 4053 3352 4087
rect 3418 4053 3446 4087
rect 3446 4053 3452 4087
rect 3518 4053 3524 4087
rect 3524 4053 3552 4087
rect 3618 4053 3652 4087
rect 3718 4053 3752 4087
rect 3818 4053 3852 4087
rect 3918 4053 3952 4087
rect 4018 4053 4052 4087
rect 4118 4053 4152 4087
rect 4218 4053 4252 4087
rect 4318 4053 4352 4087
rect 4418 4053 4452 4087
rect 4518 4053 4552 4087
rect 4618 4053 4652 4087
rect 4718 4053 4746 4087
rect 4746 4053 4752 4087
rect 4818 4053 4824 4087
rect 4824 4053 4852 4087
rect 4918 4053 4952 4087
rect 5018 4053 5052 4087
rect 5118 4053 5152 4087
rect 5218 4053 5252 4087
rect 5318 4053 5352 4087
rect 5418 4053 5452 4087
rect 5518 4053 5552 4087
rect 5618 4053 5646 4087
rect 5646 4053 5652 4087
rect 5718 4053 5724 4087
rect 5724 4053 5752 4087
rect 5818 4053 5852 4087
rect 5918 4053 5952 4087
rect 6018 4053 6052 4087
rect 6118 4053 6152 4087
rect 6218 4053 6252 4087
rect 6318 4053 6352 4087
rect 6418 4053 6446 4087
rect 6446 4053 6452 4087
rect 6516 4068 6524 4102
rect 6524 4068 6550 4102
rect 6720 4038 6746 4072
rect 6746 4038 6754 4072
rect 18 3913 52 3947
rect 118 3913 152 3947
rect 218 3913 252 3947
rect 318 3913 352 3947
rect 418 3913 452 3947
rect 518 3913 546 3947
rect 546 3913 552 3947
rect 618 3913 624 3947
rect 624 3913 652 3947
rect 718 3913 752 3947
rect 818 3913 852 3947
rect 918 3913 952 3947
rect 1018 3913 1052 3947
rect 1118 3913 1152 3947
rect 1218 3913 1252 3947
rect 1318 3913 1352 3947
rect 1418 3913 1452 3947
rect 1518 3913 1552 3947
rect 1618 3913 1652 3947
rect 1718 3913 1752 3947
rect 1818 3913 1852 3947
rect 1918 3913 1952 3947
rect 2018 3913 2052 3947
rect 2118 3913 2146 3947
rect 2146 3913 2152 3947
rect 2218 3913 2224 3947
rect 2224 3913 2252 3947
rect 2318 3913 2352 3947
rect 2418 3913 2452 3947
rect 2518 3913 2552 3947
rect 2618 3913 2652 3947
rect 2718 3913 2752 3947
rect 2818 3913 2852 3947
rect 2918 3913 2952 3947
rect 3018 3913 3052 3947
rect 3118 3913 3152 3947
rect 3218 3913 3246 3947
rect 3246 3913 3252 3947
rect 3318 3913 3324 3947
rect 3324 3913 3352 3947
rect 3418 3913 3452 3947
rect 3518 3913 3552 3947
rect 3618 3913 3652 3947
rect 3718 3913 3752 3947
rect 3818 3913 3852 3947
rect 3918 3913 3952 3947
rect 4018 3913 4052 3947
rect 4118 3913 4146 3947
rect 4146 3913 4152 3947
rect 4218 3913 4224 3947
rect 4224 3913 4252 3947
rect 4318 3913 4352 3947
rect 4418 3913 4452 3947
rect 4518 3913 4546 3947
rect 4546 3913 4552 3947
rect 4618 3913 4624 3947
rect 4624 3913 4652 3947
rect 4718 3913 4752 3947
rect 4818 3913 4852 3947
rect 4918 3913 4952 3947
rect 5018 3913 5052 3947
rect 5118 3913 5152 3947
rect 5218 3913 5252 3947
rect 5318 3913 5352 3947
rect 5418 3913 5452 3947
rect 5518 3913 5552 3947
rect 5618 3913 5652 3947
rect 5718 3913 5752 3947
rect 5818 3913 5852 3947
rect 5918 3913 5952 3947
rect 6018 3913 6046 3947
rect 6046 3913 6052 3947
rect 6118 3913 6124 3947
rect 6124 3913 6152 3947
rect 6218 3913 6252 3947
rect 6318 3913 6352 3947
rect 6418 3913 6452 3947
rect 6516 3928 6524 3962
rect 6524 3928 6550 3962
rect 6720 3898 6746 3932
rect 6746 3898 6754 3932
rect 18 3773 52 3807
rect 118 3773 152 3807
rect 218 3773 252 3807
rect 318 3773 352 3807
rect 418 3773 452 3807
rect 518 3773 552 3807
rect 618 3773 652 3807
rect 718 3773 752 3807
rect 818 3773 852 3807
rect 918 3773 952 3807
rect 1018 3773 1052 3807
rect 1118 3773 1152 3807
rect 1218 3773 1246 3807
rect 1246 3773 1252 3807
rect 1318 3773 1324 3807
rect 1324 3773 1352 3807
rect 1418 3773 1446 3807
rect 1446 3773 1452 3807
rect 1518 3773 1524 3807
rect 1524 3773 1552 3807
rect 1618 3773 1652 3807
rect 1718 3773 1746 3807
rect 1746 3773 1752 3807
rect 1818 3773 1824 3807
rect 1824 3773 1852 3807
rect 1918 3773 1952 3807
rect 2018 3773 2052 3807
rect 2118 3773 2152 3807
rect 2218 3773 2252 3807
rect 2318 3773 2352 3807
rect 2418 3773 2452 3807
rect 2518 3773 2552 3807
rect 2618 3773 2652 3807
rect 2718 3773 2752 3807
rect 2818 3773 2852 3807
rect 2918 3773 2952 3807
rect 3018 3773 3052 3807
rect 3118 3773 3152 3807
rect 3218 3773 3252 3807
rect 3318 3773 3352 3807
rect 3418 3773 3446 3807
rect 3446 3773 3452 3807
rect 3518 3773 3524 3807
rect 3524 3773 3552 3807
rect 3618 3773 3652 3807
rect 3718 3773 3752 3807
rect 3818 3773 3852 3807
rect 3918 3773 3952 3807
rect 4018 3773 4052 3807
rect 4118 3773 4152 3807
rect 4218 3773 4252 3807
rect 4318 3773 4352 3807
rect 4418 3773 4452 3807
rect 4518 3773 4552 3807
rect 4618 3773 4652 3807
rect 4718 3773 4746 3807
rect 4746 3773 4752 3807
rect 4818 3773 4824 3807
rect 4824 3773 4852 3807
rect 4918 3773 4952 3807
rect 5018 3773 5052 3807
rect 5118 3773 5152 3807
rect 5218 3773 5252 3807
rect 5318 3773 5352 3807
rect 5418 3773 5452 3807
rect 5518 3773 5552 3807
rect 5618 3773 5646 3807
rect 5646 3773 5652 3807
rect 5718 3773 5724 3807
rect 5724 3773 5752 3807
rect 5818 3773 5852 3807
rect 5918 3773 5952 3807
rect 6018 3773 6052 3807
rect 6118 3773 6152 3807
rect 6218 3773 6252 3807
rect 6318 3773 6352 3807
rect 6418 3773 6452 3807
rect 6516 3788 6524 3822
rect 6524 3788 6550 3822
rect 6720 3758 6746 3792
rect 6746 3758 6754 3792
rect 18 3650 52 3684
rect 218 3666 252 3700
rect 418 3650 452 3684
rect 618 3666 652 3700
rect 818 3650 852 3684
rect 1018 3666 1052 3700
rect 1218 3650 1252 3684
rect 1418 3666 1452 3700
rect 1618 3650 1652 3684
rect 1818 3666 1852 3700
rect 2018 3650 2052 3684
rect 2218 3666 2252 3700
rect 2418 3650 2452 3684
rect 2618 3666 2652 3700
rect 2818 3650 2852 3684
rect 3018 3666 3052 3700
rect 3218 3650 3252 3684
rect 3418 3666 3452 3700
rect 3618 3650 3652 3684
rect 3818 3666 3852 3700
rect 4018 3650 4052 3684
rect 4218 3666 4252 3700
rect 4418 3650 4452 3684
rect 4618 3666 4652 3700
rect 4818 3650 4852 3684
rect 5018 3666 5052 3700
rect 5218 3650 5252 3684
rect 5418 3666 5452 3700
rect 5618 3650 5652 3684
rect 5818 3666 5852 3700
rect 6018 3650 6052 3684
rect 6218 3666 6252 3700
rect 6516 3647 6550 3681
rect 6720 3669 6754 3703
rect 6878 3664 6912 3698
rect 6978 3664 7012 3698
rect 7078 3664 7112 3698
rect 7178 3664 7212 3698
rect 7278 3664 7312 3698
rect 7378 3664 7412 3698
rect 18 3543 52 3577
rect 118 3543 152 3577
rect 218 3543 246 3577
rect 246 3543 252 3577
rect 318 3543 324 3577
rect 324 3543 352 3577
rect 418 3543 452 3577
rect 518 3543 552 3577
rect 618 3543 652 3577
rect 718 3543 752 3577
rect 818 3543 852 3577
rect 918 3543 952 3577
rect 1018 3543 1052 3577
rect 1118 3543 1152 3577
rect 1218 3543 1252 3577
rect 1318 3543 1346 3577
rect 1346 3543 1352 3577
rect 1418 3543 1424 3577
rect 1424 3543 1452 3577
rect 1518 3543 1546 3577
rect 1546 3543 1552 3577
rect 1618 3543 1624 3577
rect 1624 3543 1652 3577
rect 1718 3543 1752 3577
rect 1818 3543 1852 3577
rect 1918 3543 1952 3577
rect 2018 3543 2052 3577
rect 2118 3543 2152 3577
rect 2218 3543 2246 3577
rect 2246 3543 2252 3577
rect 2318 3543 2324 3577
rect 2324 3543 2352 3577
rect 2418 3543 2452 3577
rect 2518 3543 2552 3577
rect 2618 3543 2652 3577
rect 2718 3543 2752 3577
rect 2818 3543 2852 3577
rect 2918 3543 2952 3577
rect 3018 3543 3052 3577
rect 3118 3543 3152 3577
rect 3218 3543 3252 3577
rect 3318 3543 3352 3577
rect 3418 3543 3452 3577
rect 3518 3543 3546 3577
rect 3546 3543 3552 3577
rect 3618 3543 3624 3577
rect 3624 3543 3652 3577
rect 3718 3543 3746 3577
rect 3746 3543 3752 3577
rect 3818 3543 3824 3577
rect 3824 3543 3852 3577
rect 3918 3543 3952 3577
rect 4018 3543 4052 3577
rect 4118 3543 4152 3577
rect 4218 3543 4246 3577
rect 4246 3543 4252 3577
rect 4318 3543 4324 3577
rect 4324 3543 4352 3577
rect 4418 3543 4452 3577
rect 4518 3543 4552 3577
rect 4618 3543 4652 3577
rect 4718 3543 4746 3577
rect 4746 3543 4752 3577
rect 4818 3543 4824 3577
rect 4824 3543 4852 3577
rect 4918 3543 4952 3577
rect 5018 3543 5052 3577
rect 5118 3543 5152 3577
rect 5218 3543 5246 3577
rect 5246 3543 5252 3577
rect 5318 3543 5324 3577
rect 5324 3543 5352 3577
rect 5418 3543 5452 3577
rect 5518 3543 5552 3577
rect 5618 3543 5652 3577
rect 5718 3543 5752 3577
rect 5818 3543 5852 3577
rect 5918 3543 5952 3577
rect 6018 3543 6052 3577
rect 6118 3543 6152 3577
rect 6218 3543 6252 3577
rect 6318 3543 6352 3577
rect 6418 3543 6446 3577
rect 6446 3543 6452 3577
rect 6516 3558 6524 3592
rect 6524 3558 6550 3592
rect 6720 3528 6746 3562
rect 6746 3528 6754 3562
rect 18 3403 52 3437
rect 118 3403 152 3437
rect 218 3403 252 3437
rect 318 3403 352 3437
rect 418 3403 452 3437
rect 518 3403 546 3437
rect 546 3403 552 3437
rect 618 3403 624 3437
rect 624 3403 652 3437
rect 718 3403 746 3437
rect 746 3403 752 3437
rect 818 3403 824 3437
rect 824 3403 852 3437
rect 918 3403 952 3437
rect 1018 3403 1052 3437
rect 1118 3403 1152 3437
rect 1218 3403 1252 3437
rect 1318 3403 1352 3437
rect 1418 3403 1452 3437
rect 1518 3403 1552 3437
rect 1618 3403 1652 3437
rect 1718 3403 1752 3437
rect 1818 3403 1852 3437
rect 1918 3403 1946 3437
rect 1946 3403 1952 3437
rect 2018 3403 2024 3437
rect 2024 3403 2052 3437
rect 2118 3403 2152 3437
rect 2218 3403 2252 3437
rect 2318 3403 2352 3437
rect 2418 3403 2452 3437
rect 2518 3403 2552 3437
rect 2618 3403 2652 3437
rect 2718 3403 2752 3437
rect 2818 3403 2846 3437
rect 2846 3403 2852 3437
rect 2918 3403 2924 3437
rect 2924 3403 2952 3437
rect 3018 3403 3052 3437
rect 3118 3403 3152 3437
rect 3218 3403 3252 3437
rect 3318 3403 3352 3437
rect 3418 3403 3452 3437
rect 3518 3403 3552 3437
rect 3618 3403 3652 3437
rect 3718 3403 3752 3437
rect 3818 3403 3852 3437
rect 3918 3403 3952 3437
rect 4018 3403 4052 3437
rect 4118 3403 4152 3437
rect 4218 3403 4252 3437
rect 4318 3403 4352 3437
rect 4418 3403 4452 3437
rect 4518 3403 4552 3437
rect 4618 3403 4652 3437
rect 4718 3403 4752 3437
rect 4818 3403 4852 3437
rect 4918 3403 4952 3437
rect 5018 3403 5052 3437
rect 5118 3403 5152 3437
rect 5218 3403 5252 3437
rect 5318 3403 5352 3437
rect 5418 3403 5452 3437
rect 5518 3403 5552 3437
rect 5618 3403 5652 3437
rect 5718 3403 5752 3437
rect 5818 3403 5852 3437
rect 5918 3403 5946 3437
rect 5946 3403 5952 3437
rect 6018 3403 6024 3437
rect 6024 3403 6052 3437
rect 6118 3403 6152 3437
rect 6218 3403 6252 3437
rect 6318 3403 6352 3437
rect 6418 3403 6452 3437
rect 6516 3418 6524 3452
rect 6524 3418 6550 3452
rect 6720 3388 6746 3422
rect 6746 3388 6754 3422
rect 18 3263 24 3297
rect 24 3263 52 3297
rect 118 3263 152 3297
rect 218 3263 252 3297
rect 318 3263 352 3297
rect 418 3263 452 3297
rect 518 3263 552 3297
rect 618 3263 652 3297
rect 718 3263 752 3297
rect 818 3263 852 3297
rect 918 3263 952 3297
rect 1018 3263 1052 3297
rect 1118 3263 1152 3297
rect 1218 3263 1246 3297
rect 1246 3263 1252 3297
rect 1318 3263 1324 3297
rect 1324 3263 1352 3297
rect 1418 3263 1452 3297
rect 1518 3263 1552 3297
rect 1618 3263 1652 3297
rect 1718 3263 1752 3297
rect 1818 3263 1852 3297
rect 1918 3263 1952 3297
rect 2018 3263 2052 3297
rect 2118 3263 2152 3297
rect 2218 3263 2252 3297
rect 2318 3263 2352 3297
rect 2418 3263 2452 3297
rect 2518 3263 2552 3297
rect 2618 3263 2652 3297
rect 2718 3263 2746 3297
rect 2746 3263 2752 3297
rect 2818 3263 2824 3297
rect 2824 3263 2852 3297
rect 2918 3263 2946 3297
rect 2946 3263 2952 3297
rect 3018 3263 3024 3297
rect 3024 3263 3052 3297
rect 3118 3263 3152 3297
rect 3218 3263 3252 3297
rect 3318 3263 3352 3297
rect 3418 3263 3452 3297
rect 3518 3263 3552 3297
rect 3618 3263 3652 3297
rect 3718 3263 3752 3297
rect 3818 3263 3852 3297
rect 3918 3263 3952 3297
rect 4018 3263 4052 3297
rect 4118 3263 4152 3297
rect 4218 3263 4252 3297
rect 4318 3263 4346 3297
rect 4346 3263 4352 3297
rect 4418 3263 4424 3297
rect 4424 3263 4452 3297
rect 4518 3263 4552 3297
rect 4618 3263 4652 3297
rect 4718 3263 4752 3297
rect 4818 3263 4846 3297
rect 4846 3263 4852 3297
rect 4918 3263 4924 3297
rect 4924 3263 4952 3297
rect 5018 3263 5052 3297
rect 5118 3263 5152 3297
rect 5218 3263 5252 3297
rect 5318 3263 5352 3297
rect 5418 3263 5452 3297
rect 5518 3263 5546 3297
rect 5546 3263 5552 3297
rect 5618 3263 5624 3297
rect 5624 3263 5652 3297
rect 5718 3263 5752 3297
rect 5818 3263 5852 3297
rect 5918 3263 5952 3297
rect 6018 3263 6052 3297
rect 6118 3263 6152 3297
rect 6218 3263 6252 3297
rect 6318 3263 6352 3297
rect 6418 3263 6452 3297
rect 6516 3278 6524 3312
rect 6524 3278 6550 3312
rect 6720 3248 6746 3282
rect 6746 3248 6754 3282
rect 18 3123 52 3157
rect 118 3123 152 3157
rect 218 3123 252 3157
rect 318 3123 352 3157
rect 418 3123 446 3157
rect 446 3123 452 3157
rect 518 3123 524 3157
rect 524 3123 552 3157
rect 618 3123 652 3157
rect 718 3123 752 3157
rect 818 3123 852 3157
rect 918 3123 952 3157
rect 1018 3123 1052 3157
rect 1118 3123 1146 3157
rect 1146 3123 1152 3157
rect 1218 3123 1224 3157
rect 1224 3123 1252 3157
rect 1318 3123 1352 3157
rect 1418 3123 1452 3157
rect 1518 3123 1552 3157
rect 1618 3123 1652 3157
rect 1718 3123 1752 3157
rect 1818 3123 1852 3157
rect 1918 3123 1952 3157
rect 2018 3123 2052 3157
rect 2118 3123 2152 3157
rect 2218 3123 2252 3157
rect 2318 3123 2352 3157
rect 2418 3123 2446 3157
rect 2446 3123 2452 3157
rect 2518 3123 2524 3157
rect 2524 3123 2552 3157
rect 2618 3123 2652 3157
rect 2718 3123 2752 3157
rect 2818 3123 2852 3157
rect 2918 3123 2952 3157
rect 3018 3123 3052 3157
rect 3118 3123 3152 3157
rect 3218 3123 3246 3157
rect 3246 3123 3252 3157
rect 3318 3123 3324 3157
rect 3324 3123 3352 3157
rect 3418 3123 3452 3157
rect 3518 3123 3552 3157
rect 3618 3123 3646 3157
rect 3646 3123 3652 3157
rect 3718 3123 3724 3157
rect 3724 3123 3752 3157
rect 3818 3123 3852 3157
rect 3918 3123 3952 3157
rect 4018 3123 4052 3157
rect 4118 3123 4152 3157
rect 4218 3123 4246 3157
rect 4246 3123 4252 3157
rect 4318 3123 4324 3157
rect 4324 3123 4352 3157
rect 4418 3123 4452 3157
rect 4518 3123 4546 3157
rect 4546 3123 4552 3157
rect 4618 3123 4624 3157
rect 4624 3123 4652 3157
rect 4718 3123 4746 3157
rect 4746 3123 4752 3157
rect 4818 3123 4824 3157
rect 4824 3123 4852 3157
rect 4918 3123 4952 3157
rect 5018 3123 5046 3157
rect 5046 3123 5052 3157
rect 5118 3123 5124 3157
rect 5124 3123 5152 3157
rect 5218 3123 5252 3157
rect 5318 3123 5352 3157
rect 5418 3123 5452 3157
rect 5518 3123 5546 3157
rect 5546 3123 5552 3157
rect 5618 3123 5624 3157
rect 5624 3123 5652 3157
rect 5718 3123 5746 3157
rect 5746 3123 5752 3157
rect 5818 3123 5824 3157
rect 5824 3123 5852 3157
rect 5918 3123 5952 3157
rect 6018 3123 6052 3157
rect 6118 3123 6152 3157
rect 6218 3123 6252 3157
rect 6318 3123 6352 3157
rect 6418 3123 6452 3157
rect 6516 3138 6524 3172
rect 6524 3138 6550 3172
rect 6720 3108 6746 3142
rect 6746 3108 6754 3142
rect 18 2983 52 3017
rect 118 2983 152 3017
rect 218 2983 252 3017
rect 318 2983 352 3017
rect 418 2983 452 3017
rect 518 2983 552 3017
rect 618 2983 652 3017
rect 718 2983 752 3017
rect 818 2983 852 3017
rect 918 2983 952 3017
rect 1018 2983 1052 3017
rect 1118 2983 1152 3017
rect 1218 2983 1252 3017
rect 1318 2983 1352 3017
rect 1418 2983 1452 3017
rect 1518 2983 1552 3017
rect 1618 2983 1652 3017
rect 1718 2983 1752 3017
rect 1818 2983 1852 3017
rect 1918 2983 1952 3017
rect 2018 2983 2052 3017
rect 2118 2983 2152 3017
rect 2218 2983 2252 3017
rect 2318 2983 2352 3017
rect 2418 2983 2452 3017
rect 2518 2983 2552 3017
rect 2618 2983 2652 3017
rect 2718 2983 2752 3017
rect 2818 2983 2852 3017
rect 2918 2983 2952 3017
rect 3018 2983 3052 3017
rect 3118 2983 3152 3017
rect 3218 2983 3252 3017
rect 3318 2983 3346 3017
rect 3346 2983 3352 3017
rect 3418 2983 3424 3017
rect 3424 2983 3452 3017
rect 3518 2983 3552 3017
rect 3618 2983 3652 3017
rect 3718 2983 3752 3017
rect 3818 2983 3846 3017
rect 3846 2983 3852 3017
rect 3918 2983 3924 3017
rect 3924 2983 3952 3017
rect 4018 2983 4046 3017
rect 4046 2983 4052 3017
rect 4118 2983 4124 3017
rect 4124 2983 4152 3017
rect 4218 2983 4252 3017
rect 4318 2983 4352 3017
rect 4418 2983 4452 3017
rect 4518 2983 4546 3017
rect 4546 2983 4552 3017
rect 4618 2983 4624 3017
rect 4624 2983 4652 3017
rect 4718 2983 4752 3017
rect 4818 2983 4852 3017
rect 4918 2983 4952 3017
rect 5018 2983 5052 3017
rect 5118 2983 5152 3017
rect 5218 2983 5252 3017
rect 5318 2983 5352 3017
rect 5418 2983 5452 3017
rect 5518 2983 5552 3017
rect 5618 2983 5652 3017
rect 5718 2983 5752 3017
rect 5818 2983 5852 3017
rect 5918 2983 5946 3017
rect 5946 2983 5952 3017
rect 6018 2983 6024 3017
rect 6024 2983 6052 3017
rect 6118 2983 6152 3017
rect 6218 2983 6252 3017
rect 6318 2983 6352 3017
rect 6418 2983 6452 3017
rect 6516 2998 6524 3032
rect 6524 2998 6550 3032
rect 6720 2968 6746 3002
rect 6746 2968 6754 3002
rect 18 2843 52 2877
rect 118 2843 152 2877
rect 218 2843 252 2877
rect 318 2843 346 2877
rect 346 2843 352 2877
rect 418 2843 424 2877
rect 424 2843 452 2877
rect 518 2843 552 2877
rect 618 2843 652 2877
rect 718 2843 746 2877
rect 746 2843 752 2877
rect 818 2843 824 2877
rect 824 2843 852 2877
rect 918 2843 952 2877
rect 1018 2843 1052 2877
rect 1118 2843 1152 2877
rect 1218 2843 1252 2877
rect 1318 2843 1352 2877
rect 1418 2843 1446 2877
rect 1446 2843 1452 2877
rect 1518 2843 1524 2877
rect 1524 2843 1552 2877
rect 1618 2843 1652 2877
rect 1718 2843 1752 2877
rect 1818 2843 1852 2877
rect 1918 2843 1952 2877
rect 2018 2843 2052 2877
rect 2118 2843 2146 2877
rect 2146 2843 2152 2877
rect 2218 2843 2224 2877
rect 2224 2843 2252 2877
rect 2318 2843 2346 2877
rect 2346 2843 2352 2877
rect 2418 2843 2424 2877
rect 2424 2843 2452 2877
rect 2518 2843 2546 2877
rect 2546 2843 2552 2877
rect 2618 2843 2624 2877
rect 2624 2843 2652 2877
rect 2718 2843 2752 2877
rect 2818 2843 2852 2877
rect 2918 2843 2952 2877
rect 3018 2843 3046 2877
rect 3046 2843 3052 2877
rect 3118 2843 3124 2877
rect 3124 2843 3152 2877
rect 3218 2843 3252 2877
rect 3318 2843 3352 2877
rect 3418 2843 3452 2877
rect 3518 2843 3552 2877
rect 3618 2843 3652 2877
rect 3718 2843 3752 2877
rect 3818 2843 3852 2877
rect 3918 2843 3952 2877
rect 4018 2843 4052 2877
rect 4118 2843 4152 2877
rect 4218 2843 4252 2877
rect 4318 2843 4352 2877
rect 4418 2843 4452 2877
rect 4518 2843 4552 2877
rect 4618 2843 4652 2877
rect 4718 2843 4752 2877
rect 4818 2843 4852 2877
rect 4918 2843 4952 2877
rect 5018 2843 5052 2877
rect 5118 2843 5152 2877
rect 5218 2843 5252 2877
rect 5318 2843 5352 2877
rect 5418 2843 5452 2877
rect 5518 2843 5552 2877
rect 5618 2843 5652 2877
rect 5718 2843 5752 2877
rect 5818 2843 5852 2877
rect 5918 2843 5952 2877
rect 6018 2843 6046 2877
rect 6046 2843 6052 2877
rect 6118 2843 6124 2877
rect 6124 2843 6152 2877
rect 6218 2843 6252 2877
rect 6318 2843 6352 2877
rect 6418 2843 6446 2877
rect 6446 2843 6452 2877
rect 6516 2858 6524 2892
rect 6524 2858 6550 2892
rect 6720 2828 6746 2862
rect 6746 2828 6754 2862
rect 18 2703 52 2737
rect 118 2703 152 2737
rect 218 2703 252 2737
rect 318 2703 352 2737
rect 418 2703 452 2737
rect 518 2703 552 2737
rect 618 2703 652 2737
rect 718 2703 752 2737
rect 818 2703 852 2737
rect 918 2703 952 2737
rect 1018 2703 1052 2737
rect 1118 2703 1152 2737
rect 1218 2703 1252 2737
rect 1318 2703 1346 2737
rect 1346 2703 1352 2737
rect 1418 2703 1424 2737
rect 1424 2703 1452 2737
rect 1518 2703 1546 2737
rect 1546 2703 1552 2737
rect 1618 2703 1624 2737
rect 1624 2703 1652 2737
rect 1718 2703 1752 2737
rect 1818 2703 1852 2737
rect 1918 2703 1952 2737
rect 2018 2703 2046 2737
rect 2046 2703 2052 2737
rect 2118 2703 2124 2737
rect 2124 2703 2152 2737
rect 2218 2703 2252 2737
rect 2318 2703 2352 2737
rect 2418 2703 2452 2737
rect 2518 2703 2552 2737
rect 2618 2703 2652 2737
rect 2718 2703 2752 2737
rect 2818 2703 2846 2737
rect 2846 2703 2852 2737
rect 2918 2703 2924 2737
rect 2924 2703 2952 2737
rect 3018 2703 3052 2737
rect 3118 2703 3146 2737
rect 3146 2703 3152 2737
rect 3218 2703 3224 2737
rect 3224 2703 3252 2737
rect 3318 2703 3352 2737
rect 3418 2703 3452 2737
rect 3518 2703 3552 2737
rect 3618 2703 3652 2737
rect 3718 2703 3752 2737
rect 3818 2703 3852 2737
rect 3918 2703 3952 2737
rect 4018 2703 4052 2737
rect 4118 2703 4152 2737
rect 4218 2703 4252 2737
rect 4318 2703 4352 2737
rect 4418 2703 4446 2737
rect 4446 2703 4452 2737
rect 4518 2703 4524 2737
rect 4524 2703 4552 2737
rect 4618 2703 4646 2737
rect 4646 2703 4652 2737
rect 4718 2703 4724 2737
rect 4724 2703 4752 2737
rect 4818 2703 4852 2737
rect 4918 2703 4952 2737
rect 5018 2703 5052 2737
rect 5118 2703 5152 2737
rect 5218 2703 5252 2737
rect 5318 2703 5352 2737
rect 5418 2703 5446 2737
rect 5446 2703 5452 2737
rect 5518 2703 5524 2737
rect 5524 2703 5552 2737
rect 5618 2703 5652 2737
rect 5718 2703 5752 2737
rect 5818 2703 5852 2737
rect 5918 2703 5952 2737
rect 6018 2703 6052 2737
rect 6118 2703 6152 2737
rect 6218 2703 6252 2737
rect 6318 2703 6352 2737
rect 6418 2703 6452 2737
rect 6516 2718 6524 2752
rect 6524 2718 6550 2752
rect 6720 2688 6746 2722
rect 6746 2688 6754 2722
rect 18 2563 52 2597
rect 118 2563 152 2597
rect 218 2563 252 2597
rect 318 2563 352 2597
rect 418 2563 452 2597
rect 518 2563 552 2597
rect 618 2563 652 2597
rect 718 2563 752 2597
rect 818 2563 852 2597
rect 918 2563 952 2597
rect 1018 2563 1052 2597
rect 1118 2563 1152 2597
rect 1218 2563 1252 2597
rect 1318 2563 1352 2597
rect 1418 2563 1452 2597
rect 1518 2563 1546 2597
rect 1546 2563 1552 2597
rect 1618 2563 1624 2597
rect 1624 2563 1652 2597
rect 1718 2563 1752 2597
rect 1818 2563 1852 2597
rect 1918 2563 1952 2597
rect 2018 2563 2052 2597
rect 2118 2563 2146 2597
rect 2146 2563 2152 2597
rect 2218 2563 2224 2597
rect 2224 2563 2252 2597
rect 2318 2563 2352 2597
rect 2418 2563 2446 2597
rect 2446 2563 2452 2597
rect 2518 2563 2524 2597
rect 2524 2563 2552 2597
rect 2618 2563 2646 2597
rect 2646 2563 2652 2597
rect 2718 2563 2724 2597
rect 2724 2563 2752 2597
rect 2818 2563 2852 2597
rect 2918 2563 2952 2597
rect 3018 2563 3052 2597
rect 3118 2563 3152 2597
rect 3218 2563 3246 2597
rect 3246 2563 3252 2597
rect 3318 2563 3324 2597
rect 3324 2563 3352 2597
rect 3418 2563 3446 2597
rect 3446 2563 3452 2597
rect 3518 2563 3524 2597
rect 3524 2563 3552 2597
rect 3618 2563 3652 2597
rect 3718 2563 3752 2597
rect 3818 2563 3852 2597
rect 3918 2563 3952 2597
rect 4018 2563 4052 2597
rect 4118 2563 4152 2597
rect 4218 2563 4252 2597
rect 4318 2563 4352 2597
rect 4418 2563 4452 2597
rect 4518 2563 4552 2597
rect 4618 2563 4652 2597
rect 4718 2563 4752 2597
rect 4818 2563 4852 2597
rect 4918 2563 4952 2597
rect 5018 2563 5052 2597
rect 5118 2563 5152 2597
rect 5218 2563 5252 2597
rect 5318 2563 5352 2597
rect 5418 2563 5452 2597
rect 5518 2563 5546 2597
rect 5546 2563 5552 2597
rect 5618 2563 5624 2597
rect 5624 2563 5652 2597
rect 5718 2563 5752 2597
rect 5818 2563 5852 2597
rect 5918 2563 5952 2597
rect 6018 2563 6052 2597
rect 6118 2563 6152 2597
rect 6218 2563 6252 2597
rect 6318 2563 6352 2597
rect 6418 2563 6452 2597
rect 6516 2578 6524 2612
rect 6524 2578 6550 2612
rect 6720 2548 6746 2582
rect 6746 2548 6754 2582
rect 18 2440 52 2474
rect 218 2456 252 2490
rect 418 2440 452 2474
rect 618 2456 652 2490
rect 818 2440 852 2474
rect 1018 2456 1052 2490
rect 1218 2440 1252 2474
rect 1418 2456 1452 2490
rect 1618 2440 1652 2474
rect 1818 2456 1852 2490
rect 2018 2440 2052 2474
rect 2218 2456 2252 2490
rect 2418 2440 2452 2474
rect 2618 2456 2652 2490
rect 2818 2440 2852 2474
rect 3018 2456 3052 2490
rect 3218 2440 3252 2474
rect 3418 2456 3452 2490
rect 3618 2440 3652 2474
rect 3818 2456 3852 2490
rect 4018 2440 4052 2474
rect 4218 2456 4252 2490
rect 4418 2440 4452 2474
rect 4618 2456 4652 2490
rect 4818 2440 4852 2474
rect 5018 2456 5052 2490
rect 5218 2440 5252 2474
rect 5418 2456 5452 2490
rect 5618 2440 5652 2474
rect 5818 2456 5852 2490
rect 6018 2440 6052 2474
rect 6218 2456 6252 2490
rect 6516 2437 6550 2471
rect 6720 2459 6754 2493
rect 6878 2454 6912 2488
rect 6978 2454 7012 2488
rect 7078 2454 7112 2488
rect 7178 2454 7212 2488
rect 7278 2454 7312 2488
rect 7378 2454 7412 2488
rect 18 2333 52 2367
rect 118 2333 152 2367
rect 218 2333 252 2367
rect 318 2333 352 2367
rect 418 2333 452 2367
rect 518 2333 552 2367
rect 618 2333 652 2367
rect 718 2333 752 2367
rect 818 2333 852 2367
rect 918 2333 952 2367
rect 1018 2333 1052 2367
rect 1118 2333 1152 2367
rect 1218 2333 1252 2367
rect 1318 2333 1352 2367
rect 1418 2333 1452 2367
rect 1518 2333 1552 2367
rect 1618 2333 1652 2367
rect 1718 2333 1752 2367
rect 1818 2333 1852 2367
rect 1918 2333 1952 2367
rect 2018 2333 2052 2367
rect 2118 2333 2152 2367
rect 2218 2333 2252 2367
rect 2318 2333 2352 2367
rect 2418 2333 2452 2367
rect 2518 2333 2552 2367
rect 2618 2333 2652 2367
rect 2718 2333 2752 2367
rect 2818 2333 2852 2367
rect 2918 2333 2952 2367
rect 3018 2333 3052 2367
rect 3118 2333 3152 2367
rect 3218 2333 3252 2367
rect 3318 2333 3352 2367
rect 3418 2333 3452 2367
rect 3518 2333 3552 2367
rect 3618 2333 3652 2367
rect 3718 2333 3752 2367
rect 3818 2333 3852 2367
rect 3918 2333 3952 2367
rect 4018 2333 4052 2367
rect 4118 2333 4152 2367
rect 4218 2333 4252 2367
rect 4318 2333 4352 2367
rect 4418 2333 4452 2367
rect 4518 2333 4552 2367
rect 4618 2333 4652 2367
rect 4718 2333 4752 2367
rect 4818 2333 4852 2367
rect 4918 2333 4952 2367
rect 5018 2333 5052 2367
rect 5118 2333 5152 2367
rect 5218 2333 5252 2367
rect 5318 2333 5352 2367
rect 5418 2333 5446 2367
rect 5446 2333 5452 2367
rect 5518 2333 5524 2367
rect 5524 2333 5552 2367
rect 5618 2333 5652 2367
rect 5718 2333 5752 2367
rect 5818 2333 5852 2367
rect 5918 2333 5952 2367
rect 6018 2333 6052 2367
rect 6118 2333 6152 2367
rect 6218 2333 6252 2367
rect 6318 2333 6352 2367
rect 6418 2333 6446 2367
rect 6446 2333 6452 2367
rect 6516 2348 6524 2382
rect 6524 2348 6550 2382
rect 6720 2318 6746 2352
rect 6746 2318 6754 2352
rect 18 2193 24 2227
rect 24 2193 52 2227
rect 118 2193 152 2227
rect 218 2193 246 2227
rect 246 2193 252 2227
rect 318 2193 324 2227
rect 324 2193 352 2227
rect 418 2193 452 2227
rect 518 2193 552 2227
rect 618 2193 652 2227
rect 718 2193 752 2227
rect 818 2193 852 2227
rect 918 2193 952 2227
rect 1018 2193 1052 2227
rect 1118 2193 1152 2227
rect 1218 2193 1252 2227
rect 1318 2193 1346 2227
rect 1346 2193 1352 2227
rect 1418 2193 1424 2227
rect 1424 2193 1452 2227
rect 1518 2193 1546 2227
rect 1546 2193 1552 2227
rect 1618 2193 1624 2227
rect 1624 2193 1652 2227
rect 1718 2193 1752 2227
rect 1818 2193 1846 2227
rect 1846 2193 1852 2227
rect 1918 2193 1924 2227
rect 1924 2193 1952 2227
rect 2018 2193 2052 2227
rect 2118 2193 2152 2227
rect 2218 2193 2246 2227
rect 2246 2193 2252 2227
rect 2318 2193 2324 2227
rect 2324 2193 2352 2227
rect 2418 2193 2452 2227
rect 2518 2193 2552 2227
rect 2618 2193 2652 2227
rect 2718 2193 2752 2227
rect 2818 2193 2846 2227
rect 2846 2193 2852 2227
rect 2918 2193 2924 2227
rect 2924 2193 2952 2227
rect 3018 2193 3052 2227
rect 3118 2193 3152 2227
rect 3218 2193 3252 2227
rect 3318 2193 3352 2227
rect 3418 2193 3452 2227
rect 3518 2193 3546 2227
rect 3546 2193 3552 2227
rect 3618 2193 3624 2227
rect 3624 2193 3652 2227
rect 3718 2193 3752 2227
rect 3818 2193 3852 2227
rect 3918 2193 3952 2227
rect 4018 2193 4052 2227
rect 4118 2193 4152 2227
rect 4218 2193 4246 2227
rect 4246 2193 4252 2227
rect 4318 2193 4324 2227
rect 4324 2193 4352 2227
rect 4418 2193 4446 2227
rect 4446 2193 4452 2227
rect 4518 2193 4524 2227
rect 4524 2193 4552 2227
rect 4618 2193 4652 2227
rect 4718 2193 4752 2227
rect 4818 2193 4852 2227
rect 4918 2193 4952 2227
rect 5018 2193 5052 2227
rect 5118 2193 5152 2227
rect 5218 2193 5252 2227
rect 5318 2193 5352 2227
rect 5418 2193 5452 2227
rect 5518 2193 5552 2227
rect 5618 2193 5652 2227
rect 5718 2193 5752 2227
rect 5818 2193 5852 2227
rect 5918 2193 5952 2227
rect 6018 2193 6052 2227
rect 6118 2193 6152 2227
rect 6218 2193 6252 2227
rect 6318 2193 6352 2227
rect 6418 2193 6446 2227
rect 6446 2193 6452 2227
rect 6516 2208 6524 2242
rect 6524 2208 6550 2242
rect 6720 2178 6746 2212
rect 6746 2178 6754 2212
rect 18 2053 24 2087
rect 24 2053 52 2087
rect 118 2053 152 2087
rect 218 2053 252 2087
rect 318 2053 346 2087
rect 346 2053 352 2087
rect 418 2053 424 2087
rect 424 2053 452 2087
rect 518 2053 552 2087
rect 618 2053 652 2087
rect 718 2053 752 2087
rect 818 2053 852 2087
rect 918 2053 952 2087
rect 1018 2053 1052 2087
rect 1118 2053 1152 2087
rect 1218 2053 1252 2087
rect 1318 2053 1346 2087
rect 1346 2053 1352 2087
rect 1418 2053 1424 2087
rect 1424 2053 1452 2087
rect 1518 2053 1546 2087
rect 1546 2053 1552 2087
rect 1618 2053 1624 2087
rect 1624 2053 1652 2087
rect 1718 2053 1752 2087
rect 1818 2053 1846 2087
rect 1846 2053 1852 2087
rect 1918 2053 1924 2087
rect 1924 2053 1952 2087
rect 2018 2053 2052 2087
rect 2118 2053 2152 2087
rect 2218 2053 2246 2087
rect 2246 2053 2252 2087
rect 2318 2053 2324 2087
rect 2324 2053 2352 2087
rect 2418 2053 2446 2087
rect 2446 2053 2452 2087
rect 2518 2053 2524 2087
rect 2524 2053 2552 2087
rect 2618 2053 2652 2087
rect 2718 2053 2752 2087
rect 2818 2053 2852 2087
rect 2918 2053 2952 2087
rect 3018 2053 3052 2087
rect 3118 2053 3152 2087
rect 3218 2053 3252 2087
rect 3318 2053 3346 2087
rect 3346 2053 3352 2087
rect 3418 2053 3424 2087
rect 3424 2053 3452 2087
rect 3518 2053 3552 2087
rect 3618 2053 3646 2087
rect 3646 2053 3652 2087
rect 3718 2053 3724 2087
rect 3724 2053 3752 2087
rect 3818 2053 3852 2087
rect 3918 2053 3946 2087
rect 3946 2053 3952 2087
rect 4018 2053 4024 2087
rect 4024 2053 4052 2087
rect 4118 2053 4152 2087
rect 4218 2053 4252 2087
rect 4318 2053 4352 2087
rect 4418 2053 4446 2087
rect 4446 2053 4452 2087
rect 4518 2053 4524 2087
rect 4524 2053 4552 2087
rect 4618 2053 4652 2087
rect 4718 2053 4752 2087
rect 4818 2053 4852 2087
rect 4918 2053 4952 2087
rect 5018 2053 5052 2087
rect 5118 2053 5152 2087
rect 5218 2053 5252 2087
rect 5318 2053 5352 2087
rect 5418 2053 5452 2087
rect 5518 2053 5552 2087
rect 5618 2053 5652 2087
rect 5718 2053 5752 2087
rect 5818 2053 5852 2087
rect 5918 2053 5952 2087
rect 6018 2053 6052 2087
rect 6118 2053 6152 2087
rect 6218 2053 6252 2087
rect 6318 2053 6352 2087
rect 6418 2053 6452 2087
rect 6516 2068 6524 2102
rect 6524 2068 6550 2102
rect 6720 2038 6746 2072
rect 6746 2038 6754 2072
rect 18 1913 52 1947
rect 118 1913 152 1947
rect 218 1913 252 1947
rect 318 1913 346 1947
rect 346 1913 352 1947
rect 418 1913 424 1947
rect 424 1913 452 1947
rect 518 1913 552 1947
rect 618 1913 652 1947
rect 718 1913 752 1947
rect 818 1913 852 1947
rect 918 1913 952 1947
rect 1018 1913 1052 1947
rect 1118 1913 1152 1947
rect 1218 1913 1252 1947
rect 1318 1913 1352 1947
rect 1418 1913 1446 1947
rect 1446 1913 1452 1947
rect 1518 1913 1524 1947
rect 1524 1913 1552 1947
rect 1618 1913 1652 1947
rect 1718 1913 1752 1947
rect 1818 1913 1852 1947
rect 1918 1913 1952 1947
rect 2018 1913 2052 1947
rect 2118 1913 2152 1947
rect 2218 1913 2252 1947
rect 2318 1913 2352 1947
rect 2418 1913 2446 1947
rect 2446 1913 2452 1947
rect 2518 1913 2524 1947
rect 2524 1913 2552 1947
rect 2618 1913 2652 1947
rect 2718 1913 2752 1947
rect 2818 1913 2852 1947
rect 2918 1913 2952 1947
rect 3018 1913 3046 1947
rect 3046 1913 3052 1947
rect 3118 1913 3124 1947
rect 3124 1913 3152 1947
rect 3218 1913 3252 1947
rect 3318 1913 3352 1947
rect 3418 1913 3452 1947
rect 3518 1913 3552 1947
rect 3618 1913 3652 1947
rect 3718 1913 3752 1947
rect 3818 1913 3846 1947
rect 3846 1913 3852 1947
rect 3918 1913 3924 1947
rect 3924 1913 3952 1947
rect 4018 1913 4052 1947
rect 4118 1913 4152 1947
rect 4218 1913 4252 1947
rect 4318 1913 4352 1947
rect 4418 1913 4446 1947
rect 4446 1913 4452 1947
rect 4518 1913 4524 1947
rect 4524 1913 4552 1947
rect 4618 1913 4652 1947
rect 4718 1913 4752 1947
rect 4818 1913 4852 1947
rect 4918 1913 4946 1947
rect 4946 1913 4952 1947
rect 5018 1913 5024 1947
rect 5024 1913 5052 1947
rect 5118 1913 5146 1947
rect 5146 1913 5152 1947
rect 5218 1913 5224 1947
rect 5224 1913 5252 1947
rect 5318 1913 5346 1947
rect 5346 1913 5352 1947
rect 5418 1913 5424 1947
rect 5424 1913 5452 1947
rect 5518 1913 5552 1947
rect 5618 1913 5652 1947
rect 5718 1913 5746 1947
rect 5746 1913 5752 1947
rect 5818 1913 5824 1947
rect 5824 1913 5852 1947
rect 5918 1913 5952 1947
rect 6018 1913 6046 1947
rect 6046 1913 6052 1947
rect 6118 1913 6124 1947
rect 6124 1913 6152 1947
rect 6218 1913 6252 1947
rect 6318 1913 6352 1947
rect 6418 1913 6452 1947
rect 6516 1928 6524 1962
rect 6524 1928 6550 1962
rect 6720 1898 6746 1932
rect 6746 1898 6754 1932
rect 18 1773 52 1807
rect 118 1773 152 1807
rect 218 1773 252 1807
rect 318 1773 352 1807
rect 418 1773 452 1807
rect 518 1773 552 1807
rect 618 1773 652 1807
rect 718 1773 752 1807
rect 818 1773 852 1807
rect 918 1773 946 1807
rect 946 1773 952 1807
rect 1018 1773 1024 1807
rect 1024 1773 1052 1807
rect 1118 1773 1152 1807
rect 1218 1773 1252 1807
rect 1318 1773 1352 1807
rect 1418 1773 1452 1807
rect 1518 1773 1552 1807
rect 1618 1773 1652 1807
rect 1718 1773 1752 1807
rect 1818 1773 1846 1807
rect 1846 1773 1852 1807
rect 1918 1773 1924 1807
rect 1924 1773 1952 1807
rect 2018 1773 2052 1807
rect 2118 1773 2152 1807
rect 2218 1773 2252 1807
rect 2318 1773 2352 1807
rect 2418 1773 2452 1807
rect 2518 1773 2552 1807
rect 2618 1773 2652 1807
rect 2718 1773 2752 1807
rect 2818 1773 2852 1807
rect 2918 1773 2952 1807
rect 3018 1773 3052 1807
rect 3118 1773 3152 1807
rect 3218 1773 3252 1807
rect 3318 1773 3352 1807
rect 3418 1773 3446 1807
rect 3446 1773 3452 1807
rect 3518 1773 3524 1807
rect 3524 1773 3552 1807
rect 3618 1773 3646 1807
rect 3646 1773 3652 1807
rect 3718 1773 3724 1807
rect 3724 1773 3752 1807
rect 3818 1773 3852 1807
rect 3918 1773 3946 1807
rect 3946 1773 3952 1807
rect 4018 1773 4024 1807
rect 4024 1773 4052 1807
rect 4118 1773 4152 1807
rect 4218 1773 4252 1807
rect 4318 1773 4352 1807
rect 4418 1773 4452 1807
rect 4518 1773 4552 1807
rect 4618 1773 4652 1807
rect 4718 1773 4752 1807
rect 4818 1773 4846 1807
rect 4846 1773 4852 1807
rect 4918 1773 4924 1807
rect 4924 1773 4952 1807
rect 5018 1773 5052 1807
rect 5118 1773 5152 1807
rect 5218 1773 5252 1807
rect 5318 1773 5352 1807
rect 5418 1773 5452 1807
rect 5518 1773 5552 1807
rect 5618 1773 5652 1807
rect 5718 1773 5752 1807
rect 5818 1773 5852 1807
rect 5918 1773 5952 1807
rect 6018 1773 6052 1807
rect 6118 1773 6152 1807
rect 6218 1773 6252 1807
rect 6318 1773 6352 1807
rect 6418 1773 6452 1807
rect 6516 1788 6524 1822
rect 6524 1788 6550 1822
rect 6720 1758 6746 1792
rect 6746 1758 6754 1792
rect 18 1633 24 1667
rect 24 1633 52 1667
rect 118 1633 146 1667
rect 146 1633 152 1667
rect 218 1633 224 1667
rect 224 1633 252 1667
rect 318 1633 352 1667
rect 418 1633 452 1667
rect 518 1633 552 1667
rect 618 1633 652 1667
rect 718 1633 746 1667
rect 746 1633 752 1667
rect 818 1633 824 1667
rect 824 1633 852 1667
rect 918 1633 946 1667
rect 946 1633 952 1667
rect 1018 1633 1024 1667
rect 1024 1633 1052 1667
rect 1118 1633 1152 1667
rect 1218 1633 1252 1667
rect 1318 1633 1352 1667
rect 1418 1633 1452 1667
rect 1518 1633 1546 1667
rect 1546 1633 1552 1667
rect 1618 1633 1624 1667
rect 1624 1633 1652 1667
rect 1718 1633 1746 1667
rect 1746 1633 1752 1667
rect 1818 1633 1824 1667
rect 1824 1633 1852 1667
rect 1918 1633 1946 1667
rect 1946 1633 1952 1667
rect 2018 1633 2024 1667
rect 2024 1633 2052 1667
rect 2118 1633 2152 1667
rect 2218 1633 2252 1667
rect 2318 1633 2352 1667
rect 2418 1633 2452 1667
rect 2518 1633 2552 1667
rect 2618 1633 2646 1667
rect 2646 1633 2652 1667
rect 2718 1633 2724 1667
rect 2724 1633 2752 1667
rect 2818 1633 2852 1667
rect 2918 1633 2952 1667
rect 3018 1633 3052 1667
rect 3118 1633 3152 1667
rect 3218 1633 3252 1667
rect 3318 1633 3352 1667
rect 3418 1633 3446 1667
rect 3446 1633 3452 1667
rect 3518 1633 3524 1667
rect 3524 1633 3552 1667
rect 3618 1633 3652 1667
rect 3718 1633 3746 1667
rect 3746 1633 3752 1667
rect 3818 1633 3824 1667
rect 3824 1633 3852 1667
rect 3918 1633 3952 1667
rect 4018 1633 4052 1667
rect 4118 1633 4152 1667
rect 4218 1633 4252 1667
rect 4318 1633 4352 1667
rect 4418 1633 4446 1667
rect 4446 1633 4452 1667
rect 4518 1633 4524 1667
rect 4524 1633 4552 1667
rect 4618 1633 4652 1667
rect 4718 1633 4752 1667
rect 4818 1633 4852 1667
rect 4918 1633 4952 1667
rect 5018 1633 5052 1667
rect 5118 1633 5152 1667
rect 5218 1633 5252 1667
rect 5318 1633 5346 1667
rect 5346 1633 5352 1667
rect 5418 1633 5424 1667
rect 5424 1633 5452 1667
rect 5518 1633 5552 1667
rect 5618 1633 5652 1667
rect 5718 1633 5746 1667
rect 5746 1633 5752 1667
rect 5818 1633 5824 1667
rect 5824 1633 5852 1667
rect 5918 1633 5946 1667
rect 5946 1633 5952 1667
rect 6018 1633 6024 1667
rect 6024 1633 6052 1667
rect 6118 1633 6152 1667
rect 6218 1633 6252 1667
rect 6318 1633 6352 1667
rect 6418 1633 6452 1667
rect 6516 1648 6524 1682
rect 6524 1648 6550 1682
rect 6720 1618 6746 1652
rect 6746 1618 6754 1652
rect 18 1493 24 1527
rect 24 1493 52 1527
rect 118 1493 146 1527
rect 146 1493 152 1527
rect 218 1493 224 1527
rect 224 1493 252 1527
rect 318 1493 352 1527
rect 418 1493 446 1527
rect 446 1493 452 1527
rect 518 1493 524 1527
rect 524 1493 552 1527
rect 618 1493 652 1527
rect 718 1493 752 1527
rect 818 1493 852 1527
rect 918 1493 952 1527
rect 1018 1493 1052 1527
rect 1118 1493 1152 1527
rect 1218 1493 1252 1527
rect 1318 1493 1352 1527
rect 1418 1493 1452 1527
rect 1518 1493 1552 1527
rect 1618 1493 1646 1527
rect 1646 1493 1652 1527
rect 1718 1493 1724 1527
rect 1724 1493 1752 1527
rect 1818 1493 1852 1527
rect 1918 1493 1952 1527
rect 2018 1493 2052 1527
rect 2118 1493 2152 1527
rect 2218 1493 2252 1527
rect 2318 1493 2352 1527
rect 2418 1493 2452 1527
rect 2518 1493 2552 1527
rect 2618 1493 2652 1527
rect 2718 1493 2752 1527
rect 2818 1493 2852 1527
rect 2918 1493 2952 1527
rect 3018 1493 3052 1527
rect 3118 1493 3152 1527
rect 3218 1493 3252 1527
rect 3318 1493 3352 1527
rect 3418 1493 3452 1527
rect 3518 1493 3552 1527
rect 3618 1493 3652 1527
rect 3718 1493 3752 1527
rect 3818 1493 3852 1527
rect 3918 1493 3952 1527
rect 4018 1493 4052 1527
rect 4118 1493 4146 1527
rect 4146 1493 4152 1527
rect 4218 1493 4224 1527
rect 4224 1493 4252 1527
rect 4318 1493 4352 1527
rect 4418 1493 4446 1527
rect 4446 1493 4452 1527
rect 4518 1493 4524 1527
rect 4524 1493 4552 1527
rect 4618 1493 4652 1527
rect 4718 1493 4752 1527
rect 4818 1493 4852 1527
rect 4918 1493 4952 1527
rect 5018 1493 5046 1527
rect 5046 1493 5052 1527
rect 5118 1493 5124 1527
rect 5124 1493 5152 1527
rect 5218 1493 5246 1527
rect 5246 1493 5252 1527
rect 5318 1493 5324 1527
rect 5324 1493 5352 1527
rect 5418 1493 5446 1527
rect 5446 1493 5452 1527
rect 5518 1493 5524 1527
rect 5524 1493 5552 1527
rect 5618 1493 5652 1527
rect 5718 1493 5746 1527
rect 5746 1493 5752 1527
rect 5818 1493 5824 1527
rect 5824 1493 5852 1527
rect 5918 1493 5946 1527
rect 5946 1493 5952 1527
rect 6018 1493 6024 1527
rect 6024 1493 6052 1527
rect 6118 1493 6152 1527
rect 6218 1493 6246 1527
rect 6246 1493 6252 1527
rect 6318 1493 6324 1527
rect 6324 1493 6352 1527
rect 6418 1493 6446 1527
rect 6446 1493 6452 1527
rect 6516 1508 6524 1542
rect 6524 1508 6550 1542
rect 6720 1478 6746 1512
rect 6746 1478 6754 1512
rect 18 1353 52 1387
rect 118 1353 152 1387
rect 218 1353 246 1387
rect 246 1353 252 1387
rect 318 1353 324 1387
rect 324 1353 352 1387
rect 418 1353 452 1387
rect 518 1353 546 1387
rect 546 1353 552 1387
rect 618 1353 624 1387
rect 624 1353 652 1387
rect 718 1353 752 1387
rect 818 1353 852 1387
rect 918 1353 952 1387
rect 1018 1353 1052 1387
rect 1118 1353 1152 1387
rect 1218 1353 1252 1387
rect 1318 1353 1352 1387
rect 1418 1353 1452 1387
rect 1518 1353 1546 1387
rect 1546 1353 1552 1387
rect 1618 1353 1624 1387
rect 1624 1353 1652 1387
rect 1718 1353 1746 1387
rect 1746 1353 1752 1387
rect 1818 1353 1824 1387
rect 1824 1353 1852 1387
rect 1918 1353 1952 1387
rect 2018 1353 2052 1387
rect 2118 1353 2152 1387
rect 2218 1353 2252 1387
rect 2318 1353 2352 1387
rect 2418 1353 2452 1387
rect 2518 1353 2552 1387
rect 2618 1353 2652 1387
rect 2718 1353 2752 1387
rect 2818 1353 2852 1387
rect 2918 1353 2946 1387
rect 2946 1353 2952 1387
rect 3018 1353 3024 1387
rect 3024 1353 3052 1387
rect 3118 1353 3152 1387
rect 3218 1353 3252 1387
rect 3318 1353 3352 1387
rect 3418 1353 3452 1387
rect 3518 1353 3546 1387
rect 3546 1353 3552 1387
rect 3618 1353 3624 1387
rect 3624 1353 3652 1387
rect 3718 1353 3752 1387
rect 3818 1353 3846 1387
rect 3846 1353 3852 1387
rect 3918 1353 3924 1387
rect 3924 1353 3952 1387
rect 4018 1353 4052 1387
rect 4118 1353 4152 1387
rect 4218 1353 4252 1387
rect 4318 1353 4352 1387
rect 4418 1353 4452 1387
rect 4518 1353 4552 1387
rect 4618 1353 4652 1387
rect 4718 1353 4752 1387
rect 4818 1353 4846 1387
rect 4846 1353 4852 1387
rect 4918 1353 4924 1387
rect 4924 1353 4952 1387
rect 5018 1353 5046 1387
rect 5046 1353 5052 1387
rect 5118 1353 5124 1387
rect 5124 1353 5152 1387
rect 5218 1353 5252 1387
rect 5318 1353 5352 1387
rect 5418 1353 5452 1387
rect 5518 1353 5552 1387
rect 5618 1353 5652 1387
rect 5718 1353 5752 1387
rect 5818 1353 5852 1387
rect 5918 1353 5952 1387
rect 6018 1353 6052 1387
rect 6118 1353 6146 1387
rect 6146 1353 6152 1387
rect 6218 1353 6224 1387
rect 6224 1353 6252 1387
rect 6318 1353 6352 1387
rect 6418 1353 6452 1387
rect 6516 1368 6524 1402
rect 6524 1368 6550 1402
rect 6720 1338 6746 1372
rect 6746 1338 6754 1372
rect 18 1230 52 1264
rect 218 1246 252 1280
rect 418 1230 452 1264
rect 618 1246 652 1280
rect 818 1230 852 1264
rect 1018 1246 1052 1280
rect 1218 1230 1252 1264
rect 1418 1246 1452 1280
rect 1618 1230 1652 1264
rect 1818 1246 1852 1280
rect 2018 1230 2052 1264
rect 2218 1246 2252 1280
rect 2418 1230 2452 1264
rect 2618 1246 2652 1280
rect 2818 1230 2852 1264
rect 3018 1246 3052 1280
rect 3218 1230 3252 1264
rect 3418 1246 3452 1280
rect 3618 1230 3652 1264
rect 3818 1246 3852 1280
rect 4018 1230 4052 1264
rect 4218 1246 4252 1280
rect 4418 1230 4452 1264
rect 4618 1246 4652 1280
rect 4818 1230 4852 1264
rect 5018 1246 5052 1280
rect 5218 1230 5252 1264
rect 5418 1246 5452 1280
rect 5618 1230 5652 1264
rect 5818 1246 5852 1280
rect 6018 1230 6052 1264
rect 6218 1246 6252 1280
rect 6516 1227 6550 1261
rect 6720 1249 6754 1283
rect 6878 1244 6912 1278
rect 6978 1244 7012 1278
rect 7078 1244 7112 1278
rect 7178 1244 7212 1278
rect 7278 1244 7312 1278
rect 7378 1244 7412 1278
rect 18 1123 52 1157
rect 118 1123 152 1157
rect 218 1123 252 1157
rect 318 1123 346 1157
rect 346 1123 352 1157
rect 418 1123 424 1157
rect 424 1123 452 1157
rect 518 1123 546 1157
rect 546 1123 552 1157
rect 618 1123 624 1157
rect 624 1123 652 1157
rect 718 1123 746 1157
rect 746 1123 752 1157
rect 818 1123 824 1157
rect 824 1123 852 1157
rect 918 1123 952 1157
rect 1018 1123 1052 1157
rect 1118 1123 1152 1157
rect 1218 1123 1246 1157
rect 1246 1123 1252 1157
rect 1318 1123 1324 1157
rect 1324 1123 1352 1157
rect 1418 1123 1452 1157
rect 1518 1123 1552 1157
rect 1618 1123 1652 1157
rect 1718 1123 1752 1157
rect 1818 1123 1852 1157
rect 1918 1123 1952 1157
rect 2018 1123 2052 1157
rect 2118 1123 2152 1157
rect 2218 1123 2252 1157
rect 2318 1123 2352 1157
rect 2418 1123 2452 1157
rect 2518 1123 2546 1157
rect 2546 1123 2552 1157
rect 2618 1123 2624 1157
rect 2624 1123 2652 1157
rect 2718 1123 2746 1157
rect 2746 1123 2752 1157
rect 2818 1123 2824 1157
rect 2824 1123 2852 1157
rect 2918 1123 2952 1157
rect 3018 1123 3052 1157
rect 3118 1123 3152 1157
rect 3218 1123 3252 1157
rect 3318 1123 3352 1157
rect 3418 1123 3452 1157
rect 3518 1123 3552 1157
rect 3618 1123 3652 1157
rect 3718 1123 3752 1157
rect 3818 1123 3852 1157
rect 3918 1123 3952 1157
rect 4018 1123 4052 1157
rect 4118 1123 4152 1157
rect 4218 1123 4246 1157
rect 4246 1123 4252 1157
rect 4318 1123 4324 1157
rect 4324 1123 4352 1157
rect 4418 1123 4452 1157
rect 4518 1123 4552 1157
rect 4618 1123 4652 1157
rect 4718 1123 4752 1157
rect 4818 1123 4852 1157
rect 4918 1123 4952 1157
rect 5018 1123 5052 1157
rect 5118 1123 5152 1157
rect 5218 1123 5252 1157
rect 5318 1123 5352 1157
rect 5418 1123 5446 1157
rect 5446 1123 5452 1157
rect 5518 1123 5524 1157
rect 5524 1123 5552 1157
rect 5618 1123 5652 1157
rect 5718 1123 5752 1157
rect 5818 1123 5852 1157
rect 5918 1123 5946 1157
rect 5946 1123 5952 1157
rect 6018 1123 6024 1157
rect 6024 1123 6052 1157
rect 6118 1123 6152 1157
rect 6218 1123 6252 1157
rect 6318 1123 6352 1157
rect 6418 1123 6446 1157
rect 6446 1123 6452 1157
rect 6516 1138 6524 1172
rect 6524 1138 6550 1172
rect 6720 1108 6746 1142
rect 6746 1108 6754 1142
rect 18 983 52 1017
rect 118 983 152 1017
rect 218 983 252 1017
rect 318 983 352 1017
rect 418 983 452 1017
rect 518 983 552 1017
rect 618 983 652 1017
rect 718 983 752 1017
rect 818 983 852 1017
rect 918 983 946 1017
rect 946 983 952 1017
rect 1018 983 1024 1017
rect 1024 983 1052 1017
rect 1118 983 1146 1017
rect 1146 983 1152 1017
rect 1218 983 1224 1017
rect 1224 983 1252 1017
rect 1318 983 1352 1017
rect 1418 983 1452 1017
rect 1518 983 1552 1017
rect 1618 983 1652 1017
rect 1718 983 1752 1017
rect 1818 983 1852 1017
rect 1918 983 1952 1017
rect 2018 983 2052 1017
rect 2118 983 2146 1017
rect 2146 983 2152 1017
rect 2218 983 2224 1017
rect 2224 983 2252 1017
rect 2318 983 2352 1017
rect 2418 983 2446 1017
rect 2446 983 2452 1017
rect 2518 983 2524 1017
rect 2524 983 2552 1017
rect 2618 983 2652 1017
rect 2718 983 2752 1017
rect 2818 983 2852 1017
rect 2918 983 2952 1017
rect 3018 983 3052 1017
rect 3118 983 3152 1017
rect 3218 983 3252 1017
rect 3318 983 3352 1017
rect 3418 983 3452 1017
rect 3518 983 3552 1017
rect 3618 983 3652 1017
rect 3718 983 3752 1017
rect 3818 983 3852 1017
rect 3918 983 3952 1017
rect 4018 983 4052 1017
rect 4118 983 4152 1017
rect 4218 983 4246 1017
rect 4246 983 4252 1017
rect 4318 983 4324 1017
rect 4324 983 4352 1017
rect 4418 983 4452 1017
rect 4518 983 4552 1017
rect 4618 983 4652 1017
rect 4718 983 4752 1017
rect 4818 983 4846 1017
rect 4846 983 4852 1017
rect 4918 983 4924 1017
rect 4924 983 4952 1017
rect 5018 983 5046 1017
rect 5046 983 5052 1017
rect 5118 983 5124 1017
rect 5124 983 5152 1017
rect 5218 983 5252 1017
rect 5318 983 5352 1017
rect 5418 983 5452 1017
rect 5518 983 5552 1017
rect 5618 983 5652 1017
rect 5718 983 5752 1017
rect 5818 983 5852 1017
rect 5918 983 5952 1017
rect 6018 983 6052 1017
rect 6118 983 6152 1017
rect 6218 983 6246 1017
rect 6246 983 6252 1017
rect 6318 983 6324 1017
rect 6324 983 6352 1017
rect 6418 983 6446 1017
rect 6446 983 6452 1017
rect 6516 998 6524 1032
rect 6524 998 6550 1032
rect 6720 968 6746 1002
rect 6746 968 6754 1002
rect 18 843 52 877
rect 118 843 152 877
rect 218 843 252 877
rect 318 843 352 877
rect 418 843 452 877
rect 518 843 552 877
rect 618 843 652 877
rect 718 843 752 877
rect 818 843 852 877
rect 918 843 952 877
rect 1018 843 1046 877
rect 1046 843 1052 877
rect 1118 843 1124 877
rect 1124 843 1152 877
rect 1218 843 1252 877
rect 1318 843 1352 877
rect 1418 843 1452 877
rect 1518 843 1552 877
rect 1618 843 1652 877
rect 1718 843 1746 877
rect 1746 843 1752 877
rect 1818 843 1824 877
rect 1824 843 1852 877
rect 1918 843 1952 877
rect 2018 843 2052 877
rect 2118 843 2152 877
rect 2218 843 2252 877
rect 2318 843 2352 877
rect 2418 843 2452 877
rect 2518 843 2552 877
rect 2618 843 2652 877
rect 2718 843 2752 877
rect 2818 843 2852 877
rect 2918 843 2952 877
rect 3018 843 3052 877
rect 3118 843 3152 877
rect 3218 843 3252 877
rect 3318 843 3352 877
rect 3418 843 3452 877
rect 3518 843 3552 877
rect 3618 843 3652 877
rect 3718 843 3752 877
rect 3818 843 3852 877
rect 3918 843 3952 877
rect 4018 843 4052 877
rect 4118 843 4152 877
rect 4218 843 4252 877
rect 4318 843 4346 877
rect 4346 843 4352 877
rect 4418 843 4424 877
rect 4424 843 4452 877
rect 4518 843 4546 877
rect 4546 843 4552 877
rect 4618 843 4624 877
rect 4624 843 4652 877
rect 4718 843 4752 877
rect 4818 843 4852 877
rect 4918 843 4952 877
rect 5018 843 5052 877
rect 5118 843 5152 877
rect 5218 843 5252 877
rect 5318 843 5352 877
rect 5418 843 5452 877
rect 5518 843 5552 877
rect 5618 843 5652 877
rect 5718 843 5752 877
rect 5818 843 5852 877
rect 5918 843 5952 877
rect 6018 843 6052 877
rect 6118 843 6152 877
rect 6218 843 6252 877
rect 6318 843 6352 877
rect 6418 843 6452 877
rect 6516 858 6524 892
rect 6524 858 6550 892
rect 6720 828 6746 862
rect 6746 828 6754 862
rect 18 703 24 737
rect 24 703 52 737
rect 118 703 152 737
rect 218 703 252 737
rect 318 703 352 737
rect 418 703 452 737
rect 518 703 552 737
rect 618 703 652 737
rect 718 703 752 737
rect 818 703 852 737
rect 918 703 946 737
rect 946 703 952 737
rect 1018 703 1024 737
rect 1024 703 1052 737
rect 1118 703 1152 737
rect 1218 703 1252 737
rect 1318 703 1352 737
rect 1418 703 1452 737
rect 1518 703 1552 737
rect 1618 703 1652 737
rect 1718 703 1752 737
rect 1818 703 1852 737
rect 1918 703 1952 737
rect 2018 703 2046 737
rect 2046 703 2052 737
rect 2118 703 2124 737
rect 2124 703 2152 737
rect 2218 703 2246 737
rect 2246 703 2252 737
rect 2318 703 2324 737
rect 2324 703 2352 737
rect 2418 703 2452 737
rect 2518 703 2552 737
rect 2618 703 2652 737
rect 2718 703 2752 737
rect 2818 703 2852 737
rect 2918 703 2952 737
rect 3018 703 3052 737
rect 3118 703 3152 737
rect 3218 703 3252 737
rect 3318 703 3352 737
rect 3418 703 3452 737
rect 3518 703 3552 737
rect 3618 703 3652 737
rect 3718 703 3752 737
rect 3818 703 3852 737
rect 3918 703 3952 737
rect 4018 703 4052 737
rect 4118 703 4152 737
rect 4218 703 4252 737
rect 4318 703 4352 737
rect 4418 703 4446 737
rect 4446 703 4452 737
rect 4518 703 4524 737
rect 4524 703 4552 737
rect 4618 703 4652 737
rect 4718 703 4752 737
rect 4818 703 4852 737
rect 4918 703 4952 737
rect 5018 703 5052 737
rect 5118 703 5152 737
rect 5218 703 5252 737
rect 5318 703 5352 737
rect 5418 703 5452 737
rect 5518 703 5546 737
rect 5546 703 5552 737
rect 5618 703 5624 737
rect 5624 703 5652 737
rect 5718 703 5746 737
rect 5746 703 5752 737
rect 5818 703 5824 737
rect 5824 703 5852 737
rect 5918 703 5952 737
rect 6018 703 6052 737
rect 6118 703 6152 737
rect 6218 703 6252 737
rect 6318 703 6352 737
rect 6418 703 6452 737
rect 6516 718 6524 752
rect 6524 718 6550 752
rect 6720 688 6746 722
rect 6746 688 6754 722
rect 18 563 52 597
rect 118 563 152 597
rect 218 563 252 597
rect 318 563 352 597
rect 418 563 452 597
rect 518 563 546 597
rect 546 563 552 597
rect 618 563 624 597
rect 624 563 652 597
rect 718 563 752 597
rect 818 563 852 597
rect 918 563 952 597
rect 1018 563 1046 597
rect 1046 563 1052 597
rect 1118 563 1124 597
rect 1124 563 1152 597
rect 1218 563 1252 597
rect 1318 563 1352 597
rect 1418 563 1452 597
rect 1518 563 1552 597
rect 1618 563 1652 597
rect 1718 563 1752 597
rect 1818 563 1852 597
rect 1918 563 1952 597
rect 2018 563 2052 597
rect 2118 563 2152 597
rect 2218 563 2252 597
rect 2318 563 2352 597
rect 2418 563 2452 597
rect 2518 563 2552 597
rect 2618 563 2652 597
rect 2718 563 2752 597
rect 2818 563 2852 597
rect 2918 563 2952 597
rect 3018 563 3052 597
rect 3118 563 3152 597
rect 3218 563 3252 597
rect 3318 563 3352 597
rect 3418 563 3452 597
rect 3518 563 3552 597
rect 3618 563 3652 597
rect 3718 563 3746 597
rect 3746 563 3752 597
rect 3818 563 3824 597
rect 3824 563 3852 597
rect 3918 563 3952 597
rect 4018 563 4046 597
rect 4046 563 4052 597
rect 4118 563 4124 597
rect 4124 563 4152 597
rect 4218 563 4246 597
rect 4246 563 4252 597
rect 4318 563 4324 597
rect 4324 563 4352 597
rect 4418 563 4452 597
rect 4518 563 4552 597
rect 4618 563 4646 597
rect 4646 563 4652 597
rect 4718 563 4724 597
rect 4724 563 4752 597
rect 4818 563 4852 597
rect 4918 563 4952 597
rect 5018 563 5052 597
rect 5118 563 5152 597
rect 5218 563 5246 597
rect 5246 563 5252 597
rect 5318 563 5324 597
rect 5324 563 5352 597
rect 5418 563 5452 597
rect 5518 563 5552 597
rect 5618 563 5652 597
rect 5718 563 5752 597
rect 5818 563 5852 597
rect 5918 563 5952 597
rect 6018 563 6046 597
rect 6046 563 6052 597
rect 6118 563 6124 597
rect 6124 563 6152 597
rect 6218 563 6252 597
rect 6318 563 6352 597
rect 6418 563 6446 597
rect 6446 563 6452 597
rect 6516 578 6524 612
rect 6524 578 6550 612
rect 6720 548 6746 582
rect 6746 548 6754 582
rect 18 423 52 457
rect 118 423 152 457
rect 218 423 246 457
rect 246 423 252 457
rect 318 423 324 457
rect 324 423 352 457
rect 418 423 446 457
rect 446 423 452 457
rect 518 423 524 457
rect 524 423 552 457
rect 618 423 652 457
rect 718 423 752 457
rect 818 423 852 457
rect 918 423 952 457
rect 1018 423 1052 457
rect 1118 423 1152 457
rect 1218 423 1252 457
rect 1318 423 1352 457
rect 1418 423 1446 457
rect 1446 423 1452 457
rect 1518 423 1524 457
rect 1524 423 1552 457
rect 1618 423 1652 457
rect 1718 423 1752 457
rect 1818 423 1852 457
rect 1918 423 1952 457
rect 2018 423 2052 457
rect 2118 423 2152 457
rect 2218 423 2252 457
rect 2318 423 2352 457
rect 2418 423 2452 457
rect 2518 423 2552 457
rect 2618 423 2652 457
rect 2718 423 2752 457
rect 2818 423 2852 457
rect 2918 423 2952 457
rect 3018 423 3046 457
rect 3046 423 3052 457
rect 3118 423 3124 457
rect 3124 423 3152 457
rect 3218 423 3246 457
rect 3246 423 3252 457
rect 3318 423 3324 457
rect 3324 423 3352 457
rect 3418 423 3452 457
rect 3518 423 3546 457
rect 3546 423 3552 457
rect 3618 423 3624 457
rect 3624 423 3652 457
rect 3718 423 3746 457
rect 3746 423 3752 457
rect 3818 423 3824 457
rect 3824 423 3852 457
rect 3918 423 3952 457
rect 4018 423 4052 457
rect 4118 423 4152 457
rect 4218 423 4252 457
rect 4318 423 4352 457
rect 4418 423 4452 457
rect 4518 423 4552 457
rect 4618 423 4652 457
rect 4718 423 4752 457
rect 4818 423 4852 457
rect 4918 423 4952 457
rect 5018 423 5052 457
rect 5118 423 5152 457
rect 5218 423 5252 457
rect 5318 423 5352 457
rect 5418 423 5452 457
rect 5518 423 5546 457
rect 5546 423 5552 457
rect 5618 423 5624 457
rect 5624 423 5652 457
rect 5718 423 5752 457
rect 5818 423 5852 457
rect 5918 423 5952 457
rect 6018 423 6052 457
rect 6118 423 6152 457
rect 6218 423 6246 457
rect 6246 423 6252 457
rect 6318 423 6324 457
rect 6324 423 6352 457
rect 6418 423 6446 457
rect 6446 423 6452 457
rect 6516 438 6524 472
rect 6524 438 6550 472
rect 6720 408 6746 442
rect 6746 408 6754 442
rect 18 283 52 317
rect 118 283 152 317
rect 218 283 252 317
rect 318 283 352 317
rect 418 283 452 317
rect 518 283 552 317
rect 618 283 646 317
rect 646 283 652 317
rect 718 283 724 317
rect 724 283 752 317
rect 818 283 852 317
rect 918 283 952 317
rect 1018 283 1052 317
rect 1118 283 1152 317
rect 1218 283 1252 317
rect 1318 283 1352 317
rect 1418 283 1452 317
rect 1518 283 1546 317
rect 1546 283 1552 317
rect 1618 283 1624 317
rect 1624 283 1652 317
rect 1718 283 1752 317
rect 1818 283 1852 317
rect 1918 283 1952 317
rect 2018 283 2052 317
rect 2118 283 2152 317
rect 2218 283 2246 317
rect 2246 283 2252 317
rect 2318 283 2324 317
rect 2324 283 2352 317
rect 2418 283 2446 317
rect 2446 283 2452 317
rect 2518 283 2524 317
rect 2524 283 2552 317
rect 2618 283 2646 317
rect 2646 283 2652 317
rect 2718 283 2724 317
rect 2724 283 2752 317
rect 2818 283 2846 317
rect 2846 283 2852 317
rect 2918 283 2924 317
rect 2924 283 2952 317
rect 3018 283 3052 317
rect 3118 283 3152 317
rect 3218 283 3252 317
rect 3318 283 3352 317
rect 3418 283 3452 317
rect 3518 283 3546 317
rect 3546 283 3552 317
rect 3618 283 3624 317
rect 3624 283 3652 317
rect 3718 283 3752 317
rect 3818 283 3852 317
rect 3918 283 3952 317
rect 4018 283 4052 317
rect 4118 283 4152 317
rect 4218 283 4252 317
rect 4318 283 4352 317
rect 4418 283 4452 317
rect 4518 283 4552 317
rect 4618 283 4652 317
rect 4718 283 4752 317
rect 4818 283 4852 317
rect 4918 283 4952 317
rect 5018 283 5052 317
rect 5118 283 5152 317
rect 5218 283 5252 317
rect 5318 283 5352 317
rect 5418 283 5452 317
rect 5518 283 5552 317
rect 5618 283 5646 317
rect 5646 283 5652 317
rect 5718 283 5724 317
rect 5724 283 5752 317
rect 5818 283 5852 317
rect 5918 283 5952 317
rect 6018 283 6052 317
rect 6118 283 6152 317
rect 6218 283 6252 317
rect 6318 283 6352 317
rect 6418 283 6446 317
rect 6446 283 6452 317
rect 6516 298 6524 332
rect 6524 298 6550 332
rect 6720 268 6746 302
rect 6746 268 6754 302
rect 18 143 24 177
rect 24 143 52 177
rect 118 143 152 177
rect 218 143 252 177
rect 318 143 352 177
rect 418 143 452 177
rect 518 143 552 177
rect 618 143 652 177
rect 718 143 752 177
rect 818 143 846 177
rect 846 143 852 177
rect 918 143 924 177
rect 924 143 952 177
rect 1018 143 1052 177
rect 1118 143 1152 177
rect 1218 143 1252 177
rect 1318 143 1352 177
rect 1418 143 1452 177
rect 1518 143 1552 177
rect 1618 143 1652 177
rect 1718 143 1752 177
rect 1818 143 1852 177
rect 1918 143 1946 177
rect 1946 143 1952 177
rect 2018 143 2024 177
rect 2024 143 2052 177
rect 2118 143 2152 177
rect 2218 143 2252 177
rect 2318 143 2352 177
rect 2418 143 2452 177
rect 2518 143 2552 177
rect 2618 143 2652 177
rect 2718 143 2752 177
rect 2818 143 2852 177
rect 2918 143 2952 177
rect 3018 143 3052 177
rect 3118 143 3152 177
rect 3218 143 3252 177
rect 3318 143 3352 177
rect 3418 143 3452 177
rect 3518 143 3546 177
rect 3546 143 3552 177
rect 3618 143 3624 177
rect 3624 143 3652 177
rect 3718 143 3752 177
rect 3818 143 3852 177
rect 3918 143 3952 177
rect 4018 143 4052 177
rect 4118 143 4152 177
rect 4218 143 4252 177
rect 4318 143 4352 177
rect 4418 143 4452 177
rect 4518 143 4552 177
rect 4618 143 4652 177
rect 4718 143 4746 177
rect 4746 143 4752 177
rect 4818 143 4824 177
rect 4824 143 4852 177
rect 4918 143 4952 177
rect 5018 143 5052 177
rect 5118 143 5152 177
rect 5218 143 5252 177
rect 5318 143 5352 177
rect 5418 143 5452 177
rect 5518 143 5552 177
rect 5618 143 5652 177
rect 5718 143 5752 177
rect 5818 143 5852 177
rect 5918 143 5952 177
rect 6018 143 6052 177
rect 6118 143 6146 177
rect 6146 143 6152 177
rect 6218 143 6224 177
rect 6224 143 6252 177
rect 6318 143 6352 177
rect 6418 143 6446 177
rect 6446 143 6452 177
rect 6516 158 6524 192
rect 6524 158 6550 192
rect 6720 128 6746 162
rect 6746 128 6754 162
rect 18 20 52 54
rect 218 36 252 70
rect 418 20 452 54
rect 618 36 652 70
rect 818 20 852 54
rect 1018 36 1052 70
rect 1218 20 1252 54
rect 1418 36 1452 70
rect 1618 20 1652 54
rect 1818 36 1852 70
rect 2018 20 2052 54
rect 2218 36 2252 70
rect 2418 20 2452 54
rect 2618 36 2652 70
rect 2818 20 2852 54
rect 3018 36 3052 70
rect 3218 20 3252 54
rect 3418 36 3452 70
rect 3618 20 3652 54
rect 3818 36 3852 70
rect 4018 20 4052 54
rect 4218 36 4252 70
rect 4418 20 4452 54
rect 4618 36 4652 70
rect 4818 20 4852 54
rect 5018 36 5052 70
rect 5218 20 5252 54
rect 5418 36 5452 70
rect 5618 20 5652 54
rect 5818 36 5852 70
rect 6018 20 6052 54
rect 6218 36 6252 70
rect 6516 17 6550 51
rect 6720 39 6754 73
rect 6878 34 6912 68
rect 6978 34 7012 68
rect 7078 34 7112 68
rect 7178 34 7212 68
rect 7278 34 7312 68
rect 7378 34 7412 68
rect -82 -94 -48 -60
rect 118 -94 152 -60
rect -82 -149 -48 -132
rect -82 -166 -48 -149
rect 18 -149 52 -133
rect 18 -167 52 -149
rect 318 -94 352 -60
rect 118 -149 152 -132
rect 118 -166 152 -149
rect 218 -149 252 -133
rect 218 -167 252 -149
rect 518 -94 552 -60
rect 318 -149 352 -132
rect 318 -166 352 -149
rect 418 -149 452 -133
rect 418 -167 452 -149
rect 718 -94 752 -60
rect 518 -149 552 -132
rect 518 -166 552 -149
rect 618 -149 652 -133
rect 618 -167 652 -149
rect 918 -94 952 -60
rect 718 -149 752 -132
rect 718 -166 752 -149
rect 818 -149 852 -133
rect 818 -167 852 -149
rect 1118 -94 1152 -60
rect 918 -149 952 -132
rect 918 -166 952 -149
rect 1018 -149 1052 -133
rect 1018 -167 1052 -149
rect 1318 -94 1352 -60
rect 1118 -149 1152 -132
rect 1118 -166 1152 -149
rect 1218 -149 1252 -133
rect 1218 -167 1252 -149
rect 1518 -94 1552 -60
rect 1318 -149 1352 -132
rect 1318 -166 1352 -149
rect 1418 -149 1452 -133
rect 1418 -167 1452 -149
rect 1718 -94 1752 -60
rect 1518 -149 1552 -132
rect 1518 -166 1552 -149
rect 1618 -149 1652 -133
rect 1618 -167 1652 -149
rect 1918 -94 1952 -60
rect 1718 -149 1752 -132
rect 1718 -166 1752 -149
rect 1818 -149 1852 -133
rect 1818 -167 1852 -149
rect 2118 -94 2152 -60
rect 1918 -149 1952 -132
rect 1918 -166 1952 -149
rect 2018 -149 2052 -133
rect 2018 -167 2052 -149
rect 2318 -94 2352 -60
rect 2118 -149 2152 -132
rect 2118 -166 2152 -149
rect 2218 -149 2252 -133
rect 2218 -167 2252 -149
rect 2518 -94 2552 -60
rect 2318 -149 2352 -132
rect 2318 -166 2352 -149
rect 2418 -149 2452 -133
rect 2418 -167 2452 -149
rect 2718 -94 2752 -60
rect 2518 -149 2552 -132
rect 2518 -166 2552 -149
rect 2618 -149 2652 -133
rect 2618 -167 2652 -149
rect 2918 -94 2952 -60
rect 2718 -149 2752 -132
rect 2718 -166 2752 -149
rect 2818 -149 2852 -133
rect 2818 -167 2852 -149
rect 3118 -94 3152 -60
rect 2918 -149 2952 -132
rect 2918 -166 2952 -149
rect 3018 -149 3052 -133
rect 3018 -167 3052 -149
rect 3318 -94 3352 -60
rect 3118 -149 3152 -132
rect 3118 -166 3152 -149
rect 3218 -149 3252 -133
rect 3218 -167 3252 -149
rect 3518 -94 3552 -60
rect 3318 -149 3352 -132
rect 3318 -166 3352 -149
rect 3418 -149 3452 -133
rect 3418 -167 3452 -149
rect 3718 -94 3752 -60
rect 3518 -149 3552 -132
rect 3518 -166 3552 -149
rect 3618 -149 3652 -133
rect 3618 -167 3652 -149
rect 3918 -94 3952 -60
rect 3718 -149 3752 -132
rect 3718 -166 3752 -149
rect 3818 -149 3852 -133
rect 3818 -167 3852 -149
rect 4118 -94 4152 -60
rect 3918 -149 3952 -132
rect 3918 -166 3952 -149
rect 4018 -149 4052 -133
rect 4018 -167 4052 -149
rect 4318 -94 4352 -60
rect 4118 -149 4152 -132
rect 4118 -166 4152 -149
rect 4218 -149 4252 -133
rect 4218 -167 4252 -149
rect 4518 -94 4552 -60
rect 4318 -149 4352 -132
rect 4318 -166 4352 -149
rect 4418 -149 4452 -133
rect 4418 -167 4452 -149
rect 4718 -94 4752 -60
rect 4518 -149 4552 -132
rect 4518 -166 4552 -149
rect 4618 -149 4652 -133
rect 4618 -167 4652 -149
rect 4918 -94 4952 -60
rect 4718 -149 4752 -132
rect 4718 -166 4752 -149
rect 4818 -149 4852 -133
rect 4818 -167 4852 -149
rect 5118 -94 5152 -60
rect 4918 -149 4952 -132
rect 4918 -166 4952 -149
rect 5018 -149 5052 -133
rect 5018 -167 5052 -149
rect 5318 -94 5352 -60
rect 5118 -149 5152 -132
rect 5118 -166 5152 -149
rect 5218 -149 5252 -133
rect 5218 -167 5252 -149
rect 5518 -94 5552 -60
rect 5318 -149 5352 -132
rect 5318 -166 5352 -149
rect 5418 -149 5452 -133
rect 5418 -167 5452 -149
rect 5718 -94 5752 -60
rect 5518 -149 5552 -132
rect 5518 -166 5552 -149
rect 5618 -149 5652 -133
rect 5618 -167 5652 -149
rect 5918 -94 5952 -60
rect 5718 -149 5752 -132
rect 5718 -166 5752 -149
rect 5818 -149 5852 -133
rect 5818 -167 5852 -149
rect 6118 -94 6152 -60
rect 5918 -149 5952 -132
rect 5918 -166 5952 -149
rect 6018 -149 6052 -133
rect 6018 -167 6052 -149
rect 6318 -94 6352 -60
rect 8158 -42 8162 -8
rect 8162 -42 8192 -8
rect 8230 -42 8264 -8
rect 8442 -42 8447 -8
rect 8447 -42 8476 -8
rect 8514 -42 8515 -8
rect 8515 -42 8548 -8
rect 8586 -42 8617 -8
rect 8617 -42 8620 -8
rect 8658 -42 8685 -8
rect 8685 -42 8692 -8
rect 8849 -42 8857 -8
rect 8857 -42 8883 -8
rect 8921 -42 8925 -8
rect 8925 -42 8955 -8
rect 8993 -42 9027 -8
rect 9065 -42 9095 -8
rect 9095 -42 9099 -8
rect 9277 -42 9278 -8
rect 9278 -42 9311 -8
rect 9349 -42 9380 -8
rect 9380 -42 9383 -8
rect 6118 -149 6152 -132
rect 6118 -166 6152 -149
rect 6218 -149 6252 -133
rect 6218 -167 6252 -149
rect 6318 -149 6352 -132
rect 8160 -142 8162 -108
rect 8162 -142 8194 -108
rect 8232 -142 8264 -108
rect 8264 -142 8266 -108
rect 6318 -166 6352 -149
rect 8441 -142 8447 -108
rect 8447 -142 8475 -108
rect 8513 -142 8515 -108
rect 8515 -142 8547 -108
rect 8585 -142 8617 -108
rect 8617 -142 8619 -108
rect 8657 -142 8685 -108
rect 8685 -142 8691 -108
rect 8851 -142 8857 -108
rect 8857 -142 8885 -108
rect 8923 -142 8925 -108
rect 8925 -142 8957 -108
rect 8995 -142 9027 -108
rect 9027 -142 9029 -108
rect 9067 -142 9095 -108
rect 9095 -142 9101 -108
rect 9276 -142 9278 -108
rect 9278 -142 9310 -108
rect 9348 -142 9380 -108
rect 9380 -142 9382 -108
rect 8158 -242 8162 -208
rect 8162 -242 8192 -208
rect 8230 -242 8264 -208
rect 8334 -242 8368 -208
rect 8442 -242 8447 -208
rect 8447 -242 8476 -208
rect 8514 -242 8515 -208
rect 8515 -242 8548 -208
rect 8586 -242 8617 -208
rect 8617 -242 8620 -208
rect 8658 -242 8685 -208
rect 8685 -242 8692 -208
rect 8849 -242 8857 -208
rect 8857 -242 8883 -208
rect 8921 -242 8925 -208
rect 8925 -242 8955 -208
rect 8993 -242 9027 -208
rect 9065 -242 9095 -208
rect 9095 -242 9099 -208
rect 9174 -242 9208 -208
rect 9277 -242 9278 -208
rect 9278 -242 9311 -208
rect 9349 -242 9380 -208
rect 9380 -242 9383 -208
rect -66 -282 -32 -248
rect 134 -282 168 -248
rect 334 -282 368 -248
rect 534 -282 568 -248
rect 734 -282 768 -248
rect 934 -282 968 -248
rect 1134 -282 1168 -248
rect 1334 -282 1368 -248
rect 1534 -282 1568 -248
rect 1734 -282 1768 -248
rect 1934 -282 1968 -248
rect 2134 -282 2168 -248
rect 2334 -282 2368 -248
rect 2534 -282 2568 -248
rect 2734 -282 2768 -248
rect 2934 -282 2968 -248
rect 3134 -282 3168 -248
rect 3334 -282 3368 -248
rect 3534 -282 3568 -248
rect 3734 -282 3768 -248
rect 3934 -282 3968 -248
rect 4134 -282 4168 -248
rect 4334 -282 4368 -248
rect 4534 -282 4568 -248
rect 4734 -282 4768 -248
rect 4934 -282 4968 -248
rect 5134 -282 5168 -248
rect 5334 -282 5368 -248
rect 5534 -282 5568 -248
rect 5734 -282 5768 -248
rect 5934 -282 5968 -248
rect 6134 -282 6168 -248
rect -82 -397 -48 -363
rect -82 -465 -48 -435
rect -82 -469 -48 -465
rect 18 -397 52 -363
rect 18 -465 52 -435
rect 18 -469 52 -465
rect 118 -397 152 -363
rect 118 -465 152 -435
rect 118 -469 152 -465
rect -118 -595 -84 -561
rect -46 -595 -12 -561
rect 44 -664 78 -630
rect 218 -397 252 -363
rect 218 -465 252 -435
rect 218 -469 252 -465
rect 318 -397 352 -363
rect 318 -465 352 -435
rect 318 -469 352 -465
rect 418 -397 452 -363
rect 418 -465 452 -435
rect 418 -469 452 -465
rect 518 -397 552 -363
rect 518 -465 552 -435
rect 518 -469 552 -465
rect 282 -595 316 -561
rect 354 -595 388 -561
rect 192 -664 226 -630
rect 444 -664 478 -630
rect 618 -397 652 -363
rect 618 -465 652 -435
rect 618 -469 652 -465
rect 718 -397 752 -363
rect 718 -465 752 -435
rect 718 -469 752 -465
rect 818 -397 852 -363
rect 818 -465 852 -435
rect 818 -469 852 -465
rect 918 -397 952 -363
rect 918 -465 952 -435
rect 918 -469 952 -465
rect 682 -595 716 -561
rect 754 -595 788 -561
rect 592 -664 626 -630
rect 844 -664 878 -630
rect 1018 -397 1052 -363
rect 1018 -465 1052 -435
rect 1018 -469 1052 -465
rect 1118 -397 1152 -363
rect 1118 -465 1152 -435
rect 1118 -469 1152 -465
rect 1218 -397 1252 -363
rect 1218 -465 1252 -435
rect 1218 -469 1252 -465
rect 1318 -397 1352 -363
rect 1318 -465 1352 -435
rect 1318 -469 1352 -465
rect 1082 -595 1116 -561
rect 1154 -595 1188 -561
rect 992 -664 1026 -630
rect 1244 -664 1278 -630
rect 1418 -397 1452 -363
rect 1418 -465 1452 -435
rect 1418 -469 1452 -465
rect 1518 -397 1552 -363
rect 1518 -465 1552 -435
rect 1518 -469 1552 -465
rect 1618 -397 1652 -363
rect 1618 -465 1652 -435
rect 1618 -469 1652 -465
rect 1718 -397 1752 -363
rect 1718 -465 1752 -435
rect 1718 -469 1752 -465
rect 1482 -595 1516 -561
rect 1554 -595 1588 -561
rect 1392 -664 1426 -630
rect 1644 -664 1678 -630
rect 1818 -397 1852 -363
rect 1818 -465 1852 -435
rect 1818 -469 1852 -465
rect 1918 -397 1952 -363
rect 1918 -465 1952 -435
rect 1918 -469 1952 -465
rect 2018 -397 2052 -363
rect 2018 -465 2052 -435
rect 2018 -469 2052 -465
rect 2118 -397 2152 -363
rect 2118 -465 2152 -435
rect 2118 -469 2152 -465
rect 1882 -595 1916 -561
rect 1954 -595 1988 -561
rect 1792 -664 1826 -630
rect 2044 -664 2078 -630
rect 2218 -397 2252 -363
rect 2218 -465 2252 -435
rect 2218 -469 2252 -465
rect 2318 -397 2352 -363
rect 2318 -465 2352 -435
rect 2318 -469 2352 -465
rect 2418 -397 2452 -363
rect 2418 -465 2452 -435
rect 2418 -469 2452 -465
rect 2518 -397 2552 -363
rect 2518 -465 2552 -435
rect 2518 -469 2552 -465
rect 2282 -595 2316 -561
rect 2354 -595 2388 -561
rect 2192 -664 2226 -630
rect 2444 -664 2478 -630
rect 2618 -397 2652 -363
rect 2618 -465 2652 -435
rect 2618 -469 2652 -465
rect 2718 -397 2752 -363
rect 2718 -465 2752 -435
rect 2718 -469 2752 -465
rect 2818 -397 2852 -363
rect 2818 -465 2852 -435
rect 2818 -469 2852 -465
rect 2918 -397 2952 -363
rect 2918 -465 2952 -435
rect 2918 -469 2952 -465
rect 2682 -595 2716 -561
rect 2754 -595 2788 -561
rect 2592 -664 2626 -630
rect 2844 -664 2878 -630
rect 3018 -397 3052 -363
rect 3018 -465 3052 -435
rect 3018 -469 3052 -465
rect 3118 -397 3152 -363
rect 3118 -465 3152 -435
rect 3118 -469 3152 -465
rect 3218 -397 3252 -363
rect 3218 -465 3252 -435
rect 3218 -469 3252 -465
rect 3318 -397 3352 -363
rect 3318 -465 3352 -435
rect 3318 -469 3352 -465
rect 3082 -595 3116 -561
rect 3154 -595 3188 -561
rect 2992 -664 3026 -630
rect 3244 -664 3278 -630
rect 3418 -397 3452 -363
rect 3418 -465 3452 -435
rect 3418 -469 3452 -465
rect 3518 -397 3552 -363
rect 3518 -465 3552 -435
rect 3518 -469 3552 -465
rect 3618 -397 3652 -363
rect 3618 -465 3652 -435
rect 3618 -469 3652 -465
rect 3718 -397 3752 -363
rect 3718 -465 3752 -435
rect 3718 -469 3752 -465
rect 3482 -595 3516 -561
rect 3554 -595 3588 -561
rect 3392 -664 3426 -630
rect 3644 -664 3678 -630
rect 3818 -397 3852 -363
rect 3818 -465 3852 -435
rect 3818 -469 3852 -465
rect 3918 -397 3952 -363
rect 3918 -465 3952 -435
rect 3918 -469 3952 -465
rect 4018 -397 4052 -363
rect 4018 -465 4052 -435
rect 4018 -469 4052 -465
rect 4118 -397 4152 -363
rect 4118 -465 4152 -435
rect 4118 -469 4152 -465
rect 3882 -595 3916 -561
rect 3954 -595 3988 -561
rect 3792 -664 3826 -630
rect 4044 -664 4078 -630
rect 4218 -397 4252 -363
rect 4218 -465 4252 -435
rect 4218 -469 4252 -465
rect 4318 -397 4352 -363
rect 4318 -465 4352 -435
rect 4318 -469 4352 -465
rect 4418 -397 4452 -363
rect 4418 -465 4452 -435
rect 4418 -469 4452 -465
rect 4518 -397 4552 -363
rect 4518 -465 4552 -435
rect 4518 -469 4552 -465
rect 4282 -595 4316 -561
rect 4354 -595 4388 -561
rect 4192 -664 4226 -630
rect 4444 -664 4478 -630
rect 4618 -397 4652 -363
rect 4618 -465 4652 -435
rect 4618 -469 4652 -465
rect 4718 -397 4752 -363
rect 4718 -465 4752 -435
rect 4718 -469 4752 -465
rect 4818 -397 4852 -363
rect 4818 -465 4852 -435
rect 4818 -469 4852 -465
rect 4918 -397 4952 -363
rect 4918 -465 4952 -435
rect 4918 -469 4952 -465
rect 4682 -595 4716 -561
rect 4754 -595 4788 -561
rect 4592 -664 4626 -630
rect 4844 -664 4878 -630
rect 5018 -397 5052 -363
rect 5018 -465 5052 -435
rect 5018 -469 5052 -465
rect 5118 -397 5152 -363
rect 5118 -465 5152 -435
rect 5118 -469 5152 -465
rect 5218 -397 5252 -363
rect 5218 -465 5252 -435
rect 5218 -469 5252 -465
rect 5318 -397 5352 -363
rect 5318 -465 5352 -435
rect 5318 -469 5352 -465
rect 5082 -595 5116 -561
rect 5154 -595 5188 -561
rect 4992 -664 5026 -630
rect 5244 -664 5278 -630
rect 5418 -397 5452 -363
rect 5418 -465 5452 -435
rect 5418 -469 5452 -465
rect 5518 -397 5552 -363
rect 5518 -465 5552 -435
rect 5518 -469 5552 -465
rect 5618 -397 5652 -363
rect 5618 -465 5652 -435
rect 5618 -469 5652 -465
rect 5718 -397 5752 -363
rect 5718 -465 5752 -435
rect 5718 -469 5752 -465
rect 5482 -595 5516 -561
rect 5554 -595 5588 -561
rect 5392 -664 5426 -630
rect 5644 -664 5678 -630
rect 5818 -397 5852 -363
rect 5818 -465 5852 -435
rect 5818 -469 5852 -465
rect 5918 -397 5952 -363
rect 5918 -465 5952 -435
rect 5918 -469 5952 -465
rect 6018 -397 6052 -363
rect 6018 -465 6052 -435
rect 6018 -469 6052 -465
rect 6118 -397 6152 -363
rect 6118 -465 6152 -435
rect 6118 -469 6152 -465
rect 5882 -595 5916 -561
rect 5954 -595 5988 -561
rect 5792 -664 5826 -630
rect 6044 -664 6078 -630
rect 6218 -397 6252 -363
rect 6218 -465 6252 -435
rect 6218 -469 6252 -465
rect 8160 -342 8162 -308
rect 8162 -342 8194 -308
rect 8232 -342 8264 -308
rect 8264 -342 8266 -308
rect 6318 -397 6352 -363
rect 8441 -342 8447 -308
rect 8447 -342 8475 -308
rect 8513 -342 8515 -308
rect 8515 -342 8547 -308
rect 8585 -342 8617 -308
rect 8617 -342 8619 -308
rect 8657 -342 8685 -308
rect 8685 -342 8691 -308
rect 8851 -342 8857 -308
rect 8857 -342 8885 -308
rect 8923 -342 8925 -308
rect 8925 -342 8957 -308
rect 8995 -342 9027 -308
rect 9027 -342 9029 -308
rect 9067 -342 9095 -308
rect 9095 -342 9101 -308
rect 9276 -342 9278 -308
rect 9278 -342 9310 -308
rect 9348 -342 9380 -308
rect 9380 -342 9382 -308
rect 6318 -465 6352 -435
rect 8158 -442 8162 -408
rect 8162 -442 8192 -408
rect 8230 -442 8264 -408
rect 8334 -442 8368 -408
rect 8442 -442 8447 -408
rect 8447 -442 8476 -408
rect 8514 -442 8515 -408
rect 8515 -442 8548 -408
rect 8586 -442 8617 -408
rect 8617 -442 8620 -408
rect 8658 -442 8685 -408
rect 8685 -442 8692 -408
rect 8849 -442 8857 -408
rect 8857 -442 8883 -408
rect 8921 -442 8925 -408
rect 8925 -442 8955 -408
rect 8993 -442 9027 -408
rect 9065 -442 9095 -408
rect 9095 -442 9099 -408
rect 9174 -442 9208 -408
rect 9277 -442 9278 -408
rect 9278 -442 9311 -408
rect 9349 -442 9380 -408
rect 9380 -442 9383 -408
rect 6318 -469 6352 -465
rect 8160 -542 8162 -508
rect 8162 -542 8194 -508
rect 8232 -542 8264 -508
rect 8264 -542 8266 -508
rect 8441 -542 8447 -508
rect 8447 -542 8475 -508
rect 8513 -542 8515 -508
rect 8515 -542 8547 -508
rect 8585 -542 8617 -508
rect 8617 -542 8619 -508
rect 8657 -542 8685 -508
rect 8685 -542 8691 -508
rect 8851 -542 8857 -508
rect 8857 -542 8885 -508
rect 8923 -542 8925 -508
rect 8925 -542 8957 -508
rect 8995 -542 9027 -508
rect 9027 -542 9029 -508
rect 9067 -542 9095 -508
rect 9095 -542 9101 -508
rect 6282 -595 6316 -561
rect 6354 -595 6388 -561
rect 9276 -542 9278 -508
rect 9278 -542 9310 -508
rect 9348 -542 9380 -508
rect 9380 -542 9382 -508
rect 6192 -664 6226 -630
rect 8158 -642 8162 -608
rect 8162 -642 8192 -608
rect 8230 -642 8264 -608
rect 8334 -642 8368 -608
rect 8442 -642 8447 -608
rect 8447 -642 8476 -608
rect 8514 -642 8515 -608
rect 8515 -642 8548 -608
rect 8586 -642 8617 -608
rect 8617 -642 8620 -608
rect 8658 -642 8685 -608
rect 8685 -642 8692 -608
rect 8849 -642 8857 -608
rect 8857 -642 8883 -608
rect 8921 -642 8925 -608
rect 8925 -642 8955 -608
rect 8993 -642 9027 -608
rect 9065 -642 9095 -608
rect 9095 -642 9099 -608
rect 9174 -642 9208 -608
rect 9277 -642 9278 -608
rect 9278 -642 9311 -608
rect 9349 -642 9380 -608
rect 9380 -642 9383 -608
rect 8160 -742 8162 -708
rect 8162 -742 8194 -708
rect 8232 -742 8264 -708
rect 8264 -742 8266 -708
rect 8441 -742 8447 -708
rect 8447 -742 8475 -708
rect 8513 -742 8515 -708
rect 8515 -742 8547 -708
rect 8585 -742 8617 -708
rect 8617 -742 8619 -708
rect 8657 -742 8685 -708
rect 8685 -742 8691 -708
rect 8851 -742 8857 -708
rect 8857 -742 8885 -708
rect 8923 -742 8925 -708
rect 8925 -742 8957 -708
rect 8995 -742 9027 -708
rect 9027 -742 9029 -708
rect 9067 -742 9095 -708
rect 9095 -742 9101 -708
rect 9276 -742 9278 -708
rect 9278 -742 9310 -708
rect 9348 -742 9380 -708
rect 9380 -742 9382 -708
rect -4 -858 30 -837
rect 68 -858 102 -837
rect -4 -871 -2 -858
rect -2 -871 30 -858
rect 68 -871 100 -858
rect 100 -871 102 -858
rect -82 -942 -48 -908
rect 168 -858 202 -837
rect 240 -858 274 -837
rect 168 -871 170 -858
rect 170 -871 202 -858
rect 240 -871 272 -858
rect 272 -871 274 -858
rect 396 -858 430 -837
rect 468 -858 502 -837
rect 396 -871 398 -858
rect 398 -871 430 -858
rect 468 -871 500 -858
rect 500 -871 502 -858
rect -82 -1042 -48 -1008
rect -82 -1142 -48 -1108
rect 568 -858 602 -837
rect 640 -858 674 -837
rect 568 -871 570 -858
rect 570 -871 602 -858
rect 640 -871 672 -858
rect 672 -871 674 -858
rect 796 -858 830 -837
rect 868 -858 902 -837
rect 796 -871 798 -858
rect 798 -871 830 -858
rect 868 -871 900 -858
rect 900 -871 902 -858
rect 718 -942 752 -908
rect 968 -858 1002 -837
rect 1040 -858 1074 -837
rect 968 -871 970 -858
rect 970 -871 1002 -858
rect 1040 -871 1072 -858
rect 1072 -871 1074 -858
rect 1196 -858 1230 -837
rect 1268 -858 1302 -837
rect 1196 -871 1198 -858
rect 1198 -871 1230 -858
rect 1268 -871 1300 -858
rect 1300 -871 1302 -858
rect 718 -1042 752 -1008
rect 718 -1142 752 -1108
rect -82 -1242 -48 -1208
rect -82 -1342 -48 -1308
rect 1368 -858 1402 -837
rect 1440 -858 1474 -837
rect 1368 -871 1370 -858
rect 1370 -871 1402 -858
rect 1440 -871 1472 -858
rect 1472 -871 1474 -858
rect 1596 -858 1630 -837
rect 1668 -858 1702 -837
rect 1596 -871 1598 -858
rect 1598 -871 1630 -858
rect 1668 -871 1700 -858
rect 1700 -871 1702 -858
rect 1518 -942 1552 -908
rect 1768 -858 1802 -837
rect 1840 -858 1874 -837
rect 1768 -871 1770 -858
rect 1770 -871 1802 -858
rect 1840 -871 1872 -858
rect 1872 -871 1874 -858
rect 1996 -858 2030 -837
rect 2068 -858 2102 -837
rect 1996 -871 1998 -858
rect 1998 -871 2030 -858
rect 2068 -871 2100 -858
rect 2100 -871 2102 -858
rect 1518 -1042 1552 -1008
rect 1518 -1142 1552 -1108
rect 718 -1242 752 -1208
rect 2168 -858 2202 -837
rect 2240 -858 2274 -837
rect 2168 -871 2170 -858
rect 2170 -871 2202 -858
rect 2240 -871 2272 -858
rect 2272 -871 2274 -858
rect 2396 -858 2430 -837
rect 2468 -858 2502 -837
rect 2396 -871 2398 -858
rect 2398 -871 2430 -858
rect 2468 -871 2500 -858
rect 2500 -871 2502 -858
rect 2318 -942 2352 -908
rect 2568 -858 2602 -837
rect 2640 -858 2674 -837
rect 2568 -871 2570 -858
rect 2570 -871 2602 -858
rect 2640 -871 2672 -858
rect 2672 -871 2674 -858
rect 2796 -858 2830 -837
rect 2868 -858 2902 -837
rect 2796 -871 2798 -858
rect 2798 -871 2830 -858
rect 2868 -871 2900 -858
rect 2900 -871 2902 -858
rect 2318 -1042 2352 -1008
rect 2318 -1142 2352 -1108
rect 1518 -1242 1552 -1208
rect 718 -1342 752 -1308
rect 1518 -1342 1552 -1308
rect -82 -1442 -48 -1408
rect 718 -1442 752 -1408
rect -82 -1542 -48 -1508
rect 718 -1542 752 -1508
rect 2968 -858 3002 -837
rect 3040 -858 3074 -837
rect 2968 -871 2970 -858
rect 2970 -871 3002 -858
rect 3040 -871 3072 -858
rect 3072 -871 3074 -858
rect 3196 -858 3230 -837
rect 3268 -858 3302 -837
rect 3196 -871 3198 -858
rect 3198 -871 3230 -858
rect 3268 -871 3300 -858
rect 3300 -871 3302 -858
rect 3118 -942 3152 -908
rect 3368 -858 3402 -837
rect 3440 -858 3474 -837
rect 3368 -871 3370 -858
rect 3370 -871 3402 -858
rect 3440 -871 3472 -858
rect 3472 -871 3474 -858
rect 3596 -858 3630 -837
rect 3668 -858 3702 -837
rect 3596 -871 3598 -858
rect 3598 -871 3630 -858
rect 3668 -871 3700 -858
rect 3700 -871 3702 -858
rect 3118 -1042 3152 -1008
rect 3118 -1142 3152 -1108
rect 2318 -1242 2352 -1208
rect 3768 -858 3802 -837
rect 3840 -858 3874 -837
rect 3768 -871 3770 -858
rect 3770 -871 3802 -858
rect 3840 -871 3872 -858
rect 3872 -871 3874 -858
rect 3996 -858 4030 -837
rect 4068 -858 4102 -837
rect 3996 -871 3998 -858
rect 3998 -871 4030 -858
rect 4068 -871 4100 -858
rect 4100 -871 4102 -858
rect 3918 -942 3952 -908
rect 4168 -858 4202 -837
rect 4240 -858 4274 -837
rect 4168 -871 4170 -858
rect 4170 -871 4202 -858
rect 4240 -871 4272 -858
rect 4272 -871 4274 -858
rect 4396 -858 4430 -837
rect 4468 -858 4502 -837
rect 4396 -871 4398 -858
rect 4398 -871 4430 -858
rect 4468 -871 4500 -858
rect 4500 -871 4502 -858
rect 3918 -1042 3952 -1008
rect 3918 -1142 3952 -1108
rect 3118 -1242 3152 -1208
rect 2318 -1342 2352 -1308
rect 3118 -1342 3152 -1308
rect 1518 -1442 1552 -1408
rect 2318 -1442 2352 -1408
rect 4568 -858 4602 -837
rect 4640 -858 4674 -837
rect 4568 -871 4570 -858
rect 4570 -871 4602 -858
rect 4640 -871 4672 -858
rect 4672 -871 4674 -858
rect 4796 -858 4830 -837
rect 4868 -858 4902 -837
rect 4796 -871 4798 -858
rect 4798 -871 4830 -858
rect 4868 -871 4900 -858
rect 4900 -871 4902 -858
rect 4718 -942 4752 -908
rect 4968 -858 5002 -837
rect 5040 -858 5074 -837
rect 4968 -871 4970 -858
rect 4970 -871 5002 -858
rect 5040 -871 5072 -858
rect 5072 -871 5074 -858
rect 5196 -858 5230 -837
rect 5268 -858 5302 -837
rect 5196 -871 5198 -858
rect 5198 -871 5230 -858
rect 5268 -871 5300 -858
rect 5300 -871 5302 -858
rect 4718 -1042 4752 -1008
rect 4718 -1142 4752 -1108
rect 3918 -1242 3952 -1208
rect 5368 -858 5402 -837
rect 5440 -858 5474 -837
rect 5368 -871 5370 -858
rect 5370 -871 5402 -858
rect 5440 -871 5472 -858
rect 5472 -871 5474 -858
rect 5596 -858 5630 -837
rect 5668 -858 5702 -837
rect 5596 -871 5598 -858
rect 5598 -871 5630 -858
rect 5668 -871 5700 -858
rect 5700 -871 5702 -858
rect 5518 -942 5552 -908
rect 5768 -858 5802 -837
rect 5840 -858 5874 -837
rect 5768 -871 5770 -858
rect 5770 -871 5802 -858
rect 5840 -871 5872 -858
rect 5872 -871 5874 -858
rect 5996 -858 6030 -837
rect 6068 -858 6102 -837
rect 5996 -871 5998 -858
rect 5998 -871 6030 -858
rect 6068 -871 6100 -858
rect 6100 -871 6102 -858
rect 5518 -1042 5552 -1008
rect 5518 -1142 5552 -1108
rect 4718 -1242 4752 -1208
rect 3918 -1342 3952 -1308
rect 4718 -1342 4752 -1308
rect 3118 -1442 3152 -1408
rect 3918 -1442 3952 -1408
rect 1518 -1542 1552 -1508
rect 2318 -1542 2352 -1508
rect 3118 -1542 3152 -1508
rect -82 -1642 -48 -1608
rect 718 -1642 752 -1608
rect 1518 -1642 1552 -1608
rect -82 -1742 -48 -1708
rect 718 -1742 752 -1708
rect 1518 -1742 1552 -1708
rect 2318 -1642 2352 -1608
rect 2318 -1742 2352 -1708
rect 3918 -1542 3952 -1508
rect 6168 -858 6202 -837
rect 6240 -858 6274 -837
rect 6168 -871 6170 -858
rect 6170 -871 6202 -858
rect 6240 -871 6272 -858
rect 6272 -871 6274 -858
rect 8158 -842 8162 -808
rect 8162 -842 8192 -808
rect 8230 -842 8264 -808
rect 8334 -842 8368 -808
rect 8442 -842 8447 -808
rect 8447 -842 8476 -808
rect 8514 -842 8515 -808
rect 8515 -842 8548 -808
rect 8586 -842 8617 -808
rect 8617 -842 8620 -808
rect 8658 -842 8685 -808
rect 8685 -842 8692 -808
rect 8849 -842 8857 -808
rect 8857 -842 8883 -808
rect 8921 -842 8925 -808
rect 8925 -842 8955 -808
rect 8993 -842 9027 -808
rect 9065 -842 9095 -808
rect 9095 -842 9099 -808
rect 9174 -842 9208 -808
rect 9277 -842 9278 -808
rect 9278 -842 9311 -808
rect 9349 -842 9380 -808
rect 9380 -842 9383 -808
rect 6318 -942 6352 -908
rect 8160 -942 8162 -908
rect 8162 -942 8194 -908
rect 8232 -942 8264 -908
rect 8264 -942 8266 -908
rect 8441 -942 8447 -908
rect 8447 -942 8475 -908
rect 8513 -942 8515 -908
rect 8515 -942 8547 -908
rect 8585 -942 8617 -908
rect 8617 -942 8619 -908
rect 8657 -942 8685 -908
rect 8685 -942 8691 -908
rect 8851 -942 8857 -908
rect 8857 -942 8885 -908
rect 8923 -942 8925 -908
rect 8925 -942 8957 -908
rect 8995 -942 9027 -908
rect 9027 -942 9029 -908
rect 9067 -942 9095 -908
rect 9095 -942 9101 -908
rect 9276 -942 9278 -908
rect 9278 -942 9310 -908
rect 9348 -942 9380 -908
rect 9380 -942 9382 -908
rect 6318 -1042 6352 -1008
rect 8158 -1042 8162 -1008
rect 8162 -1042 8192 -1008
rect 8230 -1042 8264 -1008
rect 8334 -1042 8368 -1008
rect 8442 -1042 8447 -1008
rect 8447 -1042 8476 -1008
rect 8514 -1042 8515 -1008
rect 8515 -1042 8548 -1008
rect 8586 -1042 8617 -1008
rect 8617 -1042 8620 -1008
rect 8658 -1042 8685 -1008
rect 8685 -1042 8692 -1008
rect 8849 -1042 8857 -1008
rect 8857 -1042 8883 -1008
rect 8921 -1042 8925 -1008
rect 8925 -1042 8955 -1008
rect 8993 -1042 9027 -1008
rect 9065 -1042 9095 -1008
rect 9095 -1042 9099 -1008
rect 9174 -1042 9208 -1008
rect 9277 -1042 9278 -1008
rect 9278 -1042 9311 -1008
rect 9349 -1042 9380 -1008
rect 9380 -1042 9383 -1008
rect 6318 -1142 6352 -1108
rect 8160 -1142 8162 -1108
rect 8162 -1142 8194 -1108
rect 8232 -1142 8264 -1108
rect 8264 -1142 8266 -1108
rect 5518 -1242 5552 -1208
rect 8441 -1142 8447 -1108
rect 8447 -1142 8475 -1108
rect 8513 -1142 8515 -1108
rect 8515 -1142 8547 -1108
rect 8585 -1142 8617 -1108
rect 8617 -1142 8619 -1108
rect 8657 -1142 8685 -1108
rect 8685 -1142 8691 -1108
rect 8851 -1142 8857 -1108
rect 8857 -1142 8885 -1108
rect 8923 -1142 8925 -1108
rect 8925 -1142 8957 -1108
rect 8995 -1142 9027 -1108
rect 9027 -1142 9029 -1108
rect 9067 -1142 9095 -1108
rect 9095 -1142 9101 -1108
rect 9276 -1142 9278 -1108
rect 9278 -1142 9310 -1108
rect 9348 -1142 9380 -1108
rect 9380 -1142 9382 -1108
rect 6318 -1242 6352 -1208
rect 8158 -1242 8162 -1208
rect 8162 -1242 8192 -1208
rect 8230 -1242 8264 -1208
rect 8334 -1242 8368 -1208
rect 8442 -1242 8447 -1208
rect 8447 -1242 8476 -1208
rect 8514 -1242 8515 -1208
rect 8515 -1242 8548 -1208
rect 8586 -1242 8617 -1208
rect 8617 -1242 8620 -1208
rect 8658 -1242 8685 -1208
rect 8685 -1242 8692 -1208
rect 8849 -1242 8857 -1208
rect 8857 -1242 8883 -1208
rect 8921 -1242 8925 -1208
rect 8925 -1242 8955 -1208
rect 8993 -1242 9027 -1208
rect 9065 -1242 9095 -1208
rect 9095 -1242 9099 -1208
rect 9174 -1242 9208 -1208
rect 9277 -1242 9278 -1208
rect 9278 -1242 9311 -1208
rect 9349 -1242 9380 -1208
rect 9380 -1242 9383 -1208
rect 5518 -1342 5552 -1308
rect 6318 -1342 6352 -1308
rect 8160 -1342 8162 -1308
rect 8162 -1342 8194 -1308
rect 8232 -1342 8264 -1308
rect 8264 -1342 8266 -1308
rect 4718 -1442 4752 -1408
rect 5518 -1442 5552 -1408
rect 8441 -1342 8447 -1308
rect 8447 -1342 8475 -1308
rect 8513 -1342 8515 -1308
rect 8515 -1342 8547 -1308
rect 8585 -1342 8617 -1308
rect 8617 -1342 8619 -1308
rect 8657 -1342 8685 -1308
rect 8685 -1342 8691 -1308
rect 8851 -1342 8857 -1308
rect 8857 -1342 8885 -1308
rect 8923 -1342 8925 -1308
rect 8925 -1342 8957 -1308
rect 8995 -1342 9027 -1308
rect 9027 -1342 9029 -1308
rect 9067 -1342 9095 -1308
rect 9095 -1342 9101 -1308
rect 9276 -1342 9278 -1308
rect 9278 -1342 9310 -1308
rect 9348 -1342 9380 -1308
rect 9380 -1342 9382 -1308
rect 6318 -1442 6352 -1408
rect 8158 -1442 8162 -1408
rect 8162 -1442 8192 -1408
rect 8230 -1442 8264 -1408
rect 8334 -1442 8368 -1408
rect 8442 -1442 8447 -1408
rect 8447 -1442 8476 -1408
rect 8514 -1442 8515 -1408
rect 8515 -1442 8548 -1408
rect 8586 -1442 8617 -1408
rect 8617 -1442 8620 -1408
rect 8658 -1442 8685 -1408
rect 8685 -1442 8692 -1408
rect 8849 -1442 8857 -1408
rect 8857 -1442 8883 -1408
rect 8921 -1442 8925 -1408
rect 8925 -1442 8955 -1408
rect 8993 -1442 9027 -1408
rect 9065 -1442 9095 -1408
rect 9095 -1442 9099 -1408
rect 9174 -1442 9208 -1408
rect 9277 -1442 9278 -1408
rect 9278 -1442 9311 -1408
rect 9349 -1442 9380 -1408
rect 9380 -1442 9383 -1408
rect 4718 -1542 4752 -1508
rect 5518 -1542 5552 -1508
rect 6318 -1542 6352 -1508
rect 8160 -1542 8162 -1508
rect 8162 -1542 8194 -1508
rect 8232 -1542 8264 -1508
rect 8264 -1542 8266 -1508
rect 3118 -1642 3152 -1608
rect 3918 -1642 3952 -1608
rect 4718 -1642 4752 -1608
rect 5518 -1642 5552 -1608
rect 8441 -1542 8447 -1508
rect 8447 -1542 8475 -1508
rect 8513 -1542 8515 -1508
rect 8515 -1542 8547 -1508
rect 8585 -1542 8617 -1508
rect 8617 -1542 8619 -1508
rect 8657 -1542 8685 -1508
rect 8685 -1542 8691 -1508
rect 8851 -1542 8857 -1508
rect 8857 -1542 8885 -1508
rect 8923 -1542 8925 -1508
rect 8925 -1542 8957 -1508
rect 8995 -1542 9027 -1508
rect 9027 -1542 9029 -1508
rect 9067 -1542 9095 -1508
rect 9095 -1542 9101 -1508
rect 9276 -1542 9278 -1508
rect 9278 -1542 9310 -1508
rect 9348 -1542 9380 -1508
rect 9380 -1542 9382 -1508
rect 6318 -1642 6352 -1608
rect 8158 -1642 8162 -1608
rect 8162 -1642 8192 -1608
rect 8230 -1642 8264 -1608
rect 8334 -1642 8368 -1608
rect 8442 -1642 8447 -1608
rect 8447 -1642 8476 -1608
rect 8514 -1642 8515 -1608
rect 8515 -1642 8548 -1608
rect 8586 -1642 8617 -1608
rect 8617 -1642 8620 -1608
rect 8658 -1642 8685 -1608
rect 8685 -1642 8692 -1608
rect 8849 -1642 8857 -1608
rect 8857 -1642 8883 -1608
rect 8921 -1642 8925 -1608
rect 8925 -1642 8955 -1608
rect 8993 -1642 9027 -1608
rect 9065 -1642 9095 -1608
rect 9095 -1642 9099 -1608
rect 9174 -1642 9208 -1608
rect 9277 -1642 9278 -1608
rect 9278 -1642 9311 -1608
rect 9349 -1642 9380 -1608
rect 9380 -1642 9383 -1608
rect 3118 -1742 3152 -1708
rect 3918 -1742 3952 -1708
rect 4718 -1742 4752 -1708
rect 5518 -1742 5552 -1708
rect 6318 -1742 6352 -1708
rect 8160 -1742 8162 -1708
rect 8162 -1742 8194 -1708
rect 8232 -1742 8264 -1708
rect 8264 -1742 8266 -1708
rect -82 -1842 -48 -1808
rect 718 -1842 752 -1808
rect 1518 -1842 1552 -1808
rect 2318 -1842 2352 -1808
rect 3118 -1842 3152 -1808
rect 3918 -1842 3952 -1808
rect 4718 -1842 4752 -1808
rect 5518 -1842 5552 -1808
rect 8441 -1742 8447 -1708
rect 8447 -1742 8475 -1708
rect 8513 -1742 8515 -1708
rect 8515 -1742 8547 -1708
rect 8585 -1742 8617 -1708
rect 8617 -1742 8619 -1708
rect 8657 -1742 8685 -1708
rect 8685 -1742 8691 -1708
rect 8851 -1742 8857 -1708
rect 8857 -1742 8885 -1708
rect 8923 -1742 8925 -1708
rect 8925 -1742 8957 -1708
rect 8995 -1742 9027 -1708
rect 9027 -1742 9029 -1708
rect 9067 -1742 9095 -1708
rect 9095 -1742 9101 -1708
rect 9276 -1742 9278 -1708
rect 9278 -1742 9310 -1708
rect 9348 -1742 9380 -1708
rect 9380 -1742 9382 -1708
rect 6318 -1842 6352 -1808
rect 8158 -1842 8162 -1808
rect 8162 -1842 8192 -1808
rect 8230 -1842 8264 -1808
rect 8334 -1842 8368 -1808
rect 8442 -1842 8447 -1808
rect 8447 -1842 8476 -1808
rect 8514 -1842 8515 -1808
rect 8515 -1842 8548 -1808
rect 8586 -1842 8617 -1808
rect 8617 -1842 8620 -1808
rect 8658 -1842 8685 -1808
rect 8685 -1842 8692 -1808
rect 8849 -1842 8857 -1808
rect 8857 -1842 8883 -1808
rect 8921 -1842 8925 -1808
rect 8925 -1842 8955 -1808
rect 8993 -1842 9027 -1808
rect 9065 -1842 9095 -1808
rect 9095 -1842 9099 -1808
rect 9174 -1842 9208 -1808
rect 9277 -1842 9278 -1808
rect 9278 -1842 9311 -1808
rect 9349 -1842 9380 -1808
rect 9380 -1842 9383 -1808
rect -4 -1969 30 -1935
rect 68 -1969 102 -1935
rect 168 -1969 202 -1935
rect 240 -1969 274 -1935
rect 396 -1969 430 -1935
rect 468 -1969 502 -1935
rect 568 -1969 602 -1935
rect 640 -1969 674 -1935
rect 796 -1969 830 -1935
rect 868 -1969 902 -1935
rect 968 -1969 1002 -1935
rect 1040 -1969 1074 -1935
rect 1196 -1969 1230 -1935
rect 1268 -1969 1302 -1935
rect 1368 -1969 1402 -1935
rect 1440 -1969 1474 -1935
rect 1596 -1969 1630 -1935
rect 1668 -1969 1702 -1935
rect 1768 -1969 1802 -1935
rect 1840 -1969 1874 -1935
rect 1996 -1969 2030 -1935
rect 2068 -1969 2102 -1935
rect 2168 -1969 2202 -1935
rect 2240 -1969 2274 -1935
rect 2396 -1969 2430 -1935
rect 2468 -1969 2502 -1935
rect 2568 -1969 2602 -1935
rect 2640 -1969 2674 -1935
rect 2796 -1969 2830 -1935
rect 2868 -1969 2902 -1935
rect 2968 -1969 3002 -1935
rect 3040 -1969 3074 -1935
rect 3196 -1969 3230 -1935
rect 3268 -1969 3302 -1935
rect 3368 -1969 3402 -1935
rect 3440 -1969 3474 -1935
rect 3596 -1969 3630 -1935
rect 3668 -1969 3702 -1935
rect 3768 -1969 3802 -1935
rect 3840 -1969 3874 -1935
rect 3996 -1969 4030 -1935
rect 4068 -1969 4102 -1935
rect 4168 -1969 4202 -1935
rect 4240 -1969 4274 -1935
rect 4396 -1969 4430 -1935
rect 4468 -1969 4502 -1935
rect 4568 -1969 4602 -1935
rect 4640 -1969 4674 -1935
rect 4796 -1969 4830 -1935
rect 4868 -1969 4902 -1935
rect 4968 -1969 5002 -1935
rect 5040 -1969 5074 -1935
rect 5196 -1969 5230 -1935
rect 5268 -1969 5302 -1935
rect 5368 -1969 5402 -1935
rect 5440 -1969 5474 -1935
rect 5596 -1969 5630 -1935
rect 5668 -1969 5702 -1935
rect 5768 -1969 5802 -1935
rect 5840 -1969 5874 -1935
rect 5996 -1969 6030 -1935
rect 6068 -1969 6102 -1935
rect 6168 -1969 6202 -1935
rect 6240 -1969 6274 -1935
<< metal1 >>
rect 108 10020 162 10050
rect 308 10020 362 10050
rect 508 10020 562 10050
rect 708 10020 762 10050
rect 908 10020 962 10050
rect 1108 10020 1162 10050
rect 1308 10020 1362 10050
rect 1508 10020 1562 10050
rect 1708 10020 1762 10050
rect 1908 10020 1962 10050
rect 2108 10020 2162 10050
rect 2308 10020 2362 10050
rect 2508 10020 2562 10050
rect 2708 10020 2762 10050
rect 2908 10020 2962 10050
rect 3108 10020 3162 10050
rect 3308 10020 3362 10050
rect 3508 10020 3562 10050
rect 3708 10020 3762 10050
rect 3908 10020 3962 10050
rect 4108 10020 4162 10050
rect 4308 10020 4362 10050
rect 4508 10020 4562 10050
rect 4708 10020 4762 10050
rect 4908 10020 4962 10050
rect 5108 10020 5162 10050
rect 5308 10020 5362 10050
rect 5508 10020 5562 10050
rect 5708 10020 5762 10050
rect 5908 10020 5962 10050
rect 6108 10020 6162 10050
rect 6308 10020 6362 10050
rect 35 9997 6435 10020
rect 35 9963 118 9997
rect 152 9963 318 9997
rect 352 9963 518 9997
rect 552 9963 718 9997
rect 752 9963 918 9997
rect 952 9963 1118 9997
rect 1152 9963 1318 9997
rect 1352 9963 1518 9997
rect 1552 9963 1718 9997
rect 1752 9963 1918 9997
rect 1952 9963 2118 9997
rect 2152 9963 2318 9997
rect 2352 9963 2518 9997
rect 2552 9963 2718 9997
rect 2752 9963 2918 9997
rect 2952 9963 3118 9997
rect 3152 9963 3318 9997
rect 3352 9963 3518 9997
rect 3552 9963 3718 9997
rect 3752 9963 3918 9997
rect 3952 9963 4118 9997
rect 4152 9963 4318 9997
rect 4352 9963 4518 9997
rect 4552 9963 4718 9997
rect 4752 9963 4918 9997
rect 4952 9963 5118 9997
rect 5152 9963 5318 9997
rect 5352 9963 5518 9997
rect 5552 9963 5718 9997
rect 5752 9963 5918 9997
rect 5952 9963 6118 9997
rect 6152 9963 6318 9997
rect 6352 9963 6435 9997
rect 35 9940 6435 9963
rect 2 9883 68 9884
rect 2 9831 9 9883
rect 61 9831 68 9883
rect 2 9830 68 9831
rect 8 9767 62 9779
rect 8 9741 18 9767
rect 52 9741 62 9767
rect 8 9689 9 9741
rect 61 9689 62 9741
rect 8 9682 62 9689
rect 108 9767 162 9940
rect 202 9899 268 9900
rect 202 9847 209 9899
rect 261 9847 268 9899
rect 202 9846 268 9847
rect 108 9733 118 9767
rect 152 9733 162 9767
rect 8 9627 62 9639
rect 8 9601 18 9627
rect 52 9601 62 9627
rect 8 9549 9 9601
rect 61 9549 62 9601
rect 8 9542 62 9549
rect 108 9627 162 9733
rect 208 9811 262 9818
rect 208 9759 209 9811
rect 261 9759 262 9811
rect 208 9733 218 9759
rect 252 9733 262 9759
rect 208 9721 262 9733
rect 308 9767 362 9940
rect 402 9883 468 9884
rect 402 9831 409 9883
rect 461 9831 468 9883
rect 402 9830 468 9831
rect 308 9733 318 9767
rect 352 9733 362 9767
rect 108 9593 118 9627
rect 152 9593 162 9627
rect 8 9487 62 9499
rect 8 9461 18 9487
rect 52 9461 62 9487
rect 8 9409 9 9461
rect 61 9409 62 9461
rect 8 9402 62 9409
rect 108 9487 162 9593
rect 208 9671 262 9678
rect 208 9619 209 9671
rect 261 9619 262 9671
rect 208 9593 218 9619
rect 252 9593 262 9619
rect 208 9581 262 9593
rect 308 9627 362 9733
rect 408 9767 462 9779
rect 408 9741 418 9767
rect 452 9741 462 9767
rect 408 9689 409 9741
rect 461 9689 462 9741
rect 408 9682 462 9689
rect 508 9767 562 9940
rect 602 9899 668 9900
rect 602 9847 609 9899
rect 661 9847 668 9899
rect 602 9846 668 9847
rect 508 9733 518 9767
rect 552 9733 562 9767
rect 308 9593 318 9627
rect 352 9593 362 9627
rect 108 9453 118 9487
rect 152 9453 162 9487
rect 8 9347 62 9359
rect 8 9321 18 9347
rect 52 9321 62 9347
rect 8 9269 9 9321
rect 61 9269 62 9321
rect 8 9262 62 9269
rect 108 9347 162 9453
rect 208 9531 262 9538
rect 208 9479 209 9531
rect 261 9479 262 9531
rect 208 9453 218 9479
rect 252 9453 262 9479
rect 208 9441 262 9453
rect 308 9487 362 9593
rect 408 9627 462 9639
rect 408 9601 418 9627
rect 452 9601 462 9627
rect 408 9549 409 9601
rect 461 9549 462 9601
rect 408 9542 462 9549
rect 508 9627 562 9733
rect 608 9811 662 9818
rect 608 9759 609 9811
rect 661 9759 662 9811
rect 608 9733 618 9759
rect 652 9733 662 9759
rect 608 9721 662 9733
rect 708 9767 762 9940
rect 802 9883 868 9884
rect 802 9831 809 9883
rect 861 9831 868 9883
rect 802 9830 868 9831
rect 708 9733 718 9767
rect 752 9733 762 9767
rect 508 9593 518 9627
rect 552 9593 562 9627
rect 308 9453 318 9487
rect 352 9453 362 9487
rect 108 9313 118 9347
rect 152 9313 162 9347
rect 8 9207 62 9219
rect 8 9181 18 9207
rect 52 9181 62 9207
rect 8 9129 9 9181
rect 61 9129 62 9181
rect 8 9122 62 9129
rect 108 9207 162 9313
rect 208 9391 262 9398
rect 208 9339 209 9391
rect 261 9339 262 9391
rect 208 9313 218 9339
rect 252 9313 262 9339
rect 208 9301 262 9313
rect 308 9347 362 9453
rect 408 9487 462 9499
rect 408 9461 418 9487
rect 452 9461 462 9487
rect 408 9409 409 9461
rect 461 9409 462 9461
rect 408 9402 462 9409
rect 508 9487 562 9593
rect 608 9671 662 9678
rect 608 9619 609 9671
rect 661 9619 662 9671
rect 608 9593 618 9619
rect 652 9593 662 9619
rect 608 9581 662 9593
rect 708 9627 762 9733
rect 808 9767 862 9779
rect 808 9741 818 9767
rect 852 9741 862 9767
rect 808 9689 809 9741
rect 861 9689 862 9741
rect 808 9682 862 9689
rect 908 9767 962 9940
rect 1002 9899 1068 9900
rect 1002 9847 1009 9899
rect 1061 9847 1068 9899
rect 1002 9846 1068 9847
rect 908 9733 918 9767
rect 952 9733 962 9767
rect 708 9593 718 9627
rect 752 9593 762 9627
rect 508 9453 518 9487
rect 552 9453 562 9487
rect 308 9313 318 9347
rect 352 9313 362 9347
rect 108 9173 118 9207
rect 152 9173 162 9207
rect 8 9067 62 9079
rect 8 9041 18 9067
rect 52 9041 62 9067
rect 8 8989 9 9041
rect 61 8989 62 9041
rect 8 8982 62 8989
rect 108 9067 162 9173
rect 208 9251 262 9258
rect 208 9199 209 9251
rect 261 9199 262 9251
rect 208 9173 218 9199
rect 252 9173 262 9199
rect 208 9161 262 9173
rect 308 9207 362 9313
rect 408 9347 462 9359
rect 408 9321 418 9347
rect 452 9321 462 9347
rect 408 9269 409 9321
rect 461 9269 462 9321
rect 408 9262 462 9269
rect 508 9347 562 9453
rect 608 9531 662 9538
rect 608 9479 609 9531
rect 661 9479 662 9531
rect 608 9453 618 9479
rect 652 9453 662 9479
rect 608 9441 662 9453
rect 708 9487 762 9593
rect 808 9627 862 9639
rect 808 9601 818 9627
rect 852 9601 862 9627
rect 808 9549 809 9601
rect 861 9549 862 9601
rect 808 9542 862 9549
rect 908 9627 962 9733
rect 1008 9811 1062 9818
rect 1008 9759 1009 9811
rect 1061 9759 1062 9811
rect 1008 9733 1018 9759
rect 1052 9733 1062 9759
rect 1008 9721 1062 9733
rect 1108 9767 1162 9940
rect 1202 9883 1268 9884
rect 1202 9831 1209 9883
rect 1261 9831 1268 9883
rect 1202 9830 1268 9831
rect 1108 9733 1118 9767
rect 1152 9733 1162 9767
rect 908 9593 918 9627
rect 952 9593 962 9627
rect 708 9453 718 9487
rect 752 9453 762 9487
rect 508 9313 518 9347
rect 552 9313 562 9347
rect 308 9173 318 9207
rect 352 9173 362 9207
rect 108 9033 118 9067
rect 152 9033 162 9067
rect 8 8927 62 8939
rect 8 8901 18 8927
rect 52 8901 62 8927
rect 8 8849 9 8901
rect 61 8849 62 8901
rect 8 8842 62 8849
rect 108 8927 162 9033
rect 208 9111 262 9118
rect 208 9059 209 9111
rect 261 9059 262 9111
rect 208 9033 218 9059
rect 252 9033 262 9059
rect 208 9021 262 9033
rect 308 9067 362 9173
rect 408 9207 462 9219
rect 408 9181 418 9207
rect 452 9181 462 9207
rect 408 9129 409 9181
rect 461 9129 462 9181
rect 408 9122 462 9129
rect 508 9207 562 9313
rect 608 9391 662 9398
rect 608 9339 609 9391
rect 661 9339 662 9391
rect 608 9313 618 9339
rect 652 9313 662 9339
rect 608 9301 662 9313
rect 708 9347 762 9453
rect 808 9487 862 9499
rect 808 9461 818 9487
rect 852 9461 862 9487
rect 808 9409 809 9461
rect 861 9409 862 9461
rect 808 9402 862 9409
rect 908 9487 962 9593
rect 1008 9671 1062 9678
rect 1008 9619 1009 9671
rect 1061 9619 1062 9671
rect 1008 9593 1018 9619
rect 1052 9593 1062 9619
rect 1008 9581 1062 9593
rect 1108 9627 1162 9733
rect 1208 9767 1262 9779
rect 1208 9741 1218 9767
rect 1252 9741 1262 9767
rect 1208 9689 1209 9741
rect 1261 9689 1262 9741
rect 1208 9682 1262 9689
rect 1308 9767 1362 9940
rect 1402 9899 1468 9900
rect 1402 9847 1409 9899
rect 1461 9847 1468 9899
rect 1402 9846 1468 9847
rect 1308 9733 1318 9767
rect 1352 9733 1362 9767
rect 1108 9593 1118 9627
rect 1152 9593 1162 9627
rect 908 9453 918 9487
rect 952 9453 962 9487
rect 708 9313 718 9347
rect 752 9313 762 9347
rect 508 9173 518 9207
rect 552 9173 562 9207
rect 308 9033 318 9067
rect 352 9033 362 9067
rect 108 8893 118 8927
rect 152 8893 162 8927
rect 8 8787 62 8799
rect 8 8761 18 8787
rect 52 8761 62 8787
rect 8 8709 9 8761
rect 61 8709 62 8761
rect 8 8702 62 8709
rect 108 8787 162 8893
rect 208 8971 262 8978
rect 208 8919 209 8971
rect 261 8919 262 8971
rect 208 8893 218 8919
rect 252 8893 262 8919
rect 208 8881 262 8893
rect 308 8927 362 9033
rect 408 9067 462 9079
rect 408 9041 418 9067
rect 452 9041 462 9067
rect 408 8989 409 9041
rect 461 8989 462 9041
rect 408 8982 462 8989
rect 508 9067 562 9173
rect 608 9251 662 9258
rect 608 9199 609 9251
rect 661 9199 662 9251
rect 608 9173 618 9199
rect 652 9173 662 9199
rect 608 9161 662 9173
rect 708 9207 762 9313
rect 808 9347 862 9359
rect 808 9321 818 9347
rect 852 9321 862 9347
rect 808 9269 809 9321
rect 861 9269 862 9321
rect 808 9262 862 9269
rect 908 9347 962 9453
rect 1008 9531 1062 9538
rect 1008 9479 1009 9531
rect 1061 9479 1062 9531
rect 1008 9453 1018 9479
rect 1052 9453 1062 9479
rect 1008 9441 1062 9453
rect 1108 9487 1162 9593
rect 1208 9627 1262 9639
rect 1208 9601 1218 9627
rect 1252 9601 1262 9627
rect 1208 9549 1209 9601
rect 1261 9549 1262 9601
rect 1208 9542 1262 9549
rect 1308 9627 1362 9733
rect 1408 9811 1462 9818
rect 1408 9759 1409 9811
rect 1461 9759 1462 9811
rect 1408 9733 1418 9759
rect 1452 9733 1462 9759
rect 1408 9721 1462 9733
rect 1508 9767 1562 9940
rect 1602 9883 1668 9884
rect 1602 9831 1609 9883
rect 1661 9831 1668 9883
rect 1602 9830 1668 9831
rect 1508 9733 1518 9767
rect 1552 9733 1562 9767
rect 1308 9593 1318 9627
rect 1352 9593 1362 9627
rect 1108 9453 1118 9487
rect 1152 9453 1162 9487
rect 908 9313 918 9347
rect 952 9313 962 9347
rect 708 9173 718 9207
rect 752 9173 762 9207
rect 508 9033 518 9067
rect 552 9033 562 9067
rect 308 8893 318 8927
rect 352 8893 362 8927
rect 108 8753 118 8787
rect 152 8753 162 8787
rect 2 8673 68 8674
rect 2 8621 9 8673
rect 61 8621 68 8673
rect 2 8620 68 8621
rect 8 8557 62 8569
rect 8 8531 18 8557
rect 52 8531 62 8557
rect 8 8479 9 8531
rect 61 8479 62 8531
rect 8 8472 62 8479
rect 108 8557 162 8753
rect 208 8831 262 8838
rect 208 8779 209 8831
rect 261 8779 262 8831
rect 208 8753 218 8779
rect 252 8753 262 8779
rect 208 8741 262 8753
rect 308 8787 362 8893
rect 408 8927 462 8939
rect 408 8901 418 8927
rect 452 8901 462 8927
rect 408 8849 409 8901
rect 461 8849 462 8901
rect 408 8842 462 8849
rect 508 8927 562 9033
rect 608 9111 662 9118
rect 608 9059 609 9111
rect 661 9059 662 9111
rect 608 9033 618 9059
rect 652 9033 662 9059
rect 608 9021 662 9033
rect 708 9067 762 9173
rect 808 9207 862 9219
rect 808 9181 818 9207
rect 852 9181 862 9207
rect 808 9129 809 9181
rect 861 9129 862 9181
rect 808 9122 862 9129
rect 908 9207 962 9313
rect 1008 9391 1062 9398
rect 1008 9339 1009 9391
rect 1061 9339 1062 9391
rect 1008 9313 1018 9339
rect 1052 9313 1062 9339
rect 1008 9301 1062 9313
rect 1108 9347 1162 9453
rect 1208 9487 1262 9499
rect 1208 9461 1218 9487
rect 1252 9461 1262 9487
rect 1208 9409 1209 9461
rect 1261 9409 1262 9461
rect 1208 9402 1262 9409
rect 1308 9487 1362 9593
rect 1408 9671 1462 9678
rect 1408 9619 1409 9671
rect 1461 9619 1462 9671
rect 1408 9593 1418 9619
rect 1452 9593 1462 9619
rect 1408 9581 1462 9593
rect 1508 9627 1562 9733
rect 1608 9767 1662 9779
rect 1608 9741 1618 9767
rect 1652 9741 1662 9767
rect 1608 9689 1609 9741
rect 1661 9689 1662 9741
rect 1608 9682 1662 9689
rect 1708 9767 1762 9940
rect 1802 9899 1868 9900
rect 1802 9847 1809 9899
rect 1861 9847 1868 9899
rect 1802 9846 1868 9847
rect 1708 9733 1718 9767
rect 1752 9733 1762 9767
rect 1508 9593 1518 9627
rect 1552 9593 1562 9627
rect 1308 9453 1318 9487
rect 1352 9453 1362 9487
rect 1108 9313 1118 9347
rect 1152 9313 1162 9347
rect 908 9173 918 9207
rect 952 9173 962 9207
rect 708 9033 718 9067
rect 752 9033 762 9067
rect 508 8893 518 8927
rect 552 8893 562 8927
rect 308 8753 318 8787
rect 352 8753 362 8787
rect 202 8689 268 8690
rect 202 8637 209 8689
rect 261 8637 268 8689
rect 202 8636 268 8637
rect 108 8523 118 8557
rect 152 8523 162 8557
rect 8 8417 62 8429
rect 8 8391 18 8417
rect 52 8391 62 8417
rect 8 8339 9 8391
rect 61 8339 62 8391
rect 8 8332 62 8339
rect 108 8417 162 8523
rect 208 8601 262 8608
rect 208 8549 209 8601
rect 261 8549 262 8601
rect 208 8523 218 8549
rect 252 8523 262 8549
rect 208 8511 262 8523
rect 308 8557 362 8753
rect 408 8787 462 8799
rect 408 8761 418 8787
rect 452 8761 462 8787
rect 408 8709 409 8761
rect 461 8709 462 8761
rect 408 8702 462 8709
rect 508 8787 562 8893
rect 608 8971 662 8978
rect 608 8919 609 8971
rect 661 8919 662 8971
rect 608 8893 618 8919
rect 652 8893 662 8919
rect 608 8881 662 8893
rect 708 8927 762 9033
rect 808 9067 862 9079
rect 808 9041 818 9067
rect 852 9041 862 9067
rect 808 8989 809 9041
rect 861 8989 862 9041
rect 808 8982 862 8989
rect 908 9067 962 9173
rect 1008 9251 1062 9258
rect 1008 9199 1009 9251
rect 1061 9199 1062 9251
rect 1008 9173 1018 9199
rect 1052 9173 1062 9199
rect 1008 9161 1062 9173
rect 1108 9207 1162 9313
rect 1208 9347 1262 9359
rect 1208 9321 1218 9347
rect 1252 9321 1262 9347
rect 1208 9269 1209 9321
rect 1261 9269 1262 9321
rect 1208 9262 1262 9269
rect 1308 9347 1362 9453
rect 1408 9531 1462 9538
rect 1408 9479 1409 9531
rect 1461 9479 1462 9531
rect 1408 9453 1418 9479
rect 1452 9453 1462 9479
rect 1408 9441 1462 9453
rect 1508 9487 1562 9593
rect 1608 9627 1662 9639
rect 1608 9601 1618 9627
rect 1652 9601 1662 9627
rect 1608 9549 1609 9601
rect 1661 9549 1662 9601
rect 1608 9542 1662 9549
rect 1708 9627 1762 9733
rect 1808 9811 1862 9818
rect 1808 9759 1809 9811
rect 1861 9759 1862 9811
rect 1808 9733 1818 9759
rect 1852 9733 1862 9759
rect 1808 9721 1862 9733
rect 1908 9767 1962 9940
rect 2002 9883 2068 9884
rect 2002 9831 2009 9883
rect 2061 9831 2068 9883
rect 2002 9830 2068 9831
rect 1908 9733 1918 9767
rect 1952 9733 1962 9767
rect 1708 9593 1718 9627
rect 1752 9593 1762 9627
rect 1508 9453 1518 9487
rect 1552 9453 1562 9487
rect 1308 9313 1318 9347
rect 1352 9313 1362 9347
rect 1108 9173 1118 9207
rect 1152 9173 1162 9207
rect 908 9033 918 9067
rect 952 9033 962 9067
rect 708 8893 718 8927
rect 752 8893 762 8927
rect 508 8753 518 8787
rect 552 8753 562 8787
rect 402 8673 468 8674
rect 402 8621 409 8673
rect 461 8621 468 8673
rect 402 8620 468 8621
rect 308 8523 318 8557
rect 352 8523 362 8557
rect 108 8383 118 8417
rect 152 8383 162 8417
rect 8 8277 62 8289
rect 8 8251 18 8277
rect 52 8251 62 8277
rect 8 8199 9 8251
rect 61 8199 62 8251
rect 8 8192 62 8199
rect 108 8277 162 8383
rect 208 8461 262 8468
rect 208 8409 209 8461
rect 261 8409 262 8461
rect 208 8383 218 8409
rect 252 8383 262 8409
rect 208 8371 262 8383
rect 308 8417 362 8523
rect 408 8557 462 8569
rect 408 8531 418 8557
rect 452 8531 462 8557
rect 408 8479 409 8531
rect 461 8479 462 8531
rect 408 8472 462 8479
rect 508 8557 562 8753
rect 608 8831 662 8838
rect 608 8779 609 8831
rect 661 8779 662 8831
rect 608 8753 618 8779
rect 652 8753 662 8779
rect 608 8741 662 8753
rect 708 8787 762 8893
rect 808 8927 862 8939
rect 808 8901 818 8927
rect 852 8901 862 8927
rect 808 8849 809 8901
rect 861 8849 862 8901
rect 808 8842 862 8849
rect 908 8927 962 9033
rect 1008 9111 1062 9118
rect 1008 9059 1009 9111
rect 1061 9059 1062 9111
rect 1008 9033 1018 9059
rect 1052 9033 1062 9059
rect 1008 9021 1062 9033
rect 1108 9067 1162 9173
rect 1208 9207 1262 9219
rect 1208 9181 1218 9207
rect 1252 9181 1262 9207
rect 1208 9129 1209 9181
rect 1261 9129 1262 9181
rect 1208 9122 1262 9129
rect 1308 9207 1362 9313
rect 1408 9391 1462 9398
rect 1408 9339 1409 9391
rect 1461 9339 1462 9391
rect 1408 9313 1418 9339
rect 1452 9313 1462 9339
rect 1408 9301 1462 9313
rect 1508 9347 1562 9453
rect 1608 9487 1662 9499
rect 1608 9461 1618 9487
rect 1652 9461 1662 9487
rect 1608 9409 1609 9461
rect 1661 9409 1662 9461
rect 1608 9402 1662 9409
rect 1708 9487 1762 9593
rect 1808 9671 1862 9678
rect 1808 9619 1809 9671
rect 1861 9619 1862 9671
rect 1808 9593 1818 9619
rect 1852 9593 1862 9619
rect 1808 9581 1862 9593
rect 1908 9627 1962 9733
rect 2008 9767 2062 9779
rect 2008 9741 2018 9767
rect 2052 9741 2062 9767
rect 2008 9689 2009 9741
rect 2061 9689 2062 9741
rect 2008 9682 2062 9689
rect 2108 9767 2162 9940
rect 2202 9899 2268 9900
rect 2202 9847 2209 9899
rect 2261 9847 2268 9899
rect 2202 9846 2268 9847
rect 2108 9733 2118 9767
rect 2152 9733 2162 9767
rect 1908 9593 1918 9627
rect 1952 9593 1962 9627
rect 1708 9453 1718 9487
rect 1752 9453 1762 9487
rect 1508 9313 1518 9347
rect 1552 9313 1562 9347
rect 1308 9173 1318 9207
rect 1352 9173 1362 9207
rect 1108 9033 1118 9067
rect 1152 9033 1162 9067
rect 908 8893 918 8927
rect 952 8893 962 8927
rect 708 8753 718 8787
rect 752 8753 762 8787
rect 602 8689 668 8690
rect 602 8637 609 8689
rect 661 8637 668 8689
rect 602 8636 668 8637
rect 508 8523 518 8557
rect 552 8523 562 8557
rect 308 8383 318 8417
rect 352 8383 362 8417
rect 108 8243 118 8277
rect 152 8243 162 8277
rect 8 8137 62 8149
rect 8 8111 18 8137
rect 52 8111 62 8137
rect 8 8059 9 8111
rect 61 8059 62 8111
rect 8 8052 62 8059
rect 108 8137 162 8243
rect 208 8321 262 8328
rect 208 8269 209 8321
rect 261 8269 262 8321
rect 208 8243 218 8269
rect 252 8243 262 8269
rect 208 8231 262 8243
rect 308 8277 362 8383
rect 408 8417 462 8429
rect 408 8391 418 8417
rect 452 8391 462 8417
rect 408 8339 409 8391
rect 461 8339 462 8391
rect 408 8332 462 8339
rect 508 8417 562 8523
rect 608 8601 662 8608
rect 608 8549 609 8601
rect 661 8549 662 8601
rect 608 8523 618 8549
rect 652 8523 662 8549
rect 608 8511 662 8523
rect 708 8557 762 8753
rect 808 8787 862 8799
rect 808 8761 818 8787
rect 852 8761 862 8787
rect 808 8709 809 8761
rect 861 8709 862 8761
rect 808 8702 862 8709
rect 908 8787 962 8893
rect 1008 8971 1062 8978
rect 1008 8919 1009 8971
rect 1061 8919 1062 8971
rect 1008 8893 1018 8919
rect 1052 8893 1062 8919
rect 1008 8881 1062 8893
rect 1108 8927 1162 9033
rect 1208 9067 1262 9079
rect 1208 9041 1218 9067
rect 1252 9041 1262 9067
rect 1208 8989 1209 9041
rect 1261 8989 1262 9041
rect 1208 8982 1262 8989
rect 1308 9067 1362 9173
rect 1408 9251 1462 9258
rect 1408 9199 1409 9251
rect 1461 9199 1462 9251
rect 1408 9173 1418 9199
rect 1452 9173 1462 9199
rect 1408 9161 1462 9173
rect 1508 9207 1562 9313
rect 1608 9347 1662 9359
rect 1608 9321 1618 9347
rect 1652 9321 1662 9347
rect 1608 9269 1609 9321
rect 1661 9269 1662 9321
rect 1608 9262 1662 9269
rect 1708 9347 1762 9453
rect 1808 9531 1862 9538
rect 1808 9479 1809 9531
rect 1861 9479 1862 9531
rect 1808 9453 1818 9479
rect 1852 9453 1862 9479
rect 1808 9441 1862 9453
rect 1908 9487 1962 9593
rect 2008 9627 2062 9639
rect 2008 9601 2018 9627
rect 2052 9601 2062 9627
rect 2008 9549 2009 9601
rect 2061 9549 2062 9601
rect 2008 9542 2062 9549
rect 2108 9627 2162 9733
rect 2208 9811 2262 9818
rect 2208 9759 2209 9811
rect 2261 9759 2262 9811
rect 2208 9733 2218 9759
rect 2252 9733 2262 9759
rect 2208 9721 2262 9733
rect 2308 9767 2362 9940
rect 2402 9883 2468 9884
rect 2402 9831 2409 9883
rect 2461 9831 2468 9883
rect 2402 9830 2468 9831
rect 2308 9733 2318 9767
rect 2352 9733 2362 9767
rect 2108 9593 2118 9627
rect 2152 9593 2162 9627
rect 1908 9453 1918 9487
rect 1952 9453 1962 9487
rect 1708 9313 1718 9347
rect 1752 9313 1762 9347
rect 1508 9173 1518 9207
rect 1552 9173 1562 9207
rect 1308 9033 1318 9067
rect 1352 9033 1362 9067
rect 1108 8893 1118 8927
rect 1152 8893 1162 8927
rect 908 8753 918 8787
rect 952 8753 962 8787
rect 802 8673 868 8674
rect 802 8621 809 8673
rect 861 8621 868 8673
rect 802 8620 868 8621
rect 708 8523 718 8557
rect 752 8523 762 8557
rect 508 8383 518 8417
rect 552 8383 562 8417
rect 308 8243 318 8277
rect 352 8243 362 8277
rect 108 8103 118 8137
rect 152 8103 162 8137
rect 8 7997 62 8009
rect 8 7971 18 7997
rect 52 7971 62 7997
rect 8 7919 9 7971
rect 61 7919 62 7971
rect 8 7912 62 7919
rect 108 7997 162 8103
rect 208 8181 262 8188
rect 208 8129 209 8181
rect 261 8129 262 8181
rect 208 8103 218 8129
rect 252 8103 262 8129
rect 208 8091 262 8103
rect 308 8137 362 8243
rect 408 8277 462 8289
rect 408 8251 418 8277
rect 452 8251 462 8277
rect 408 8199 409 8251
rect 461 8199 462 8251
rect 408 8192 462 8199
rect 508 8277 562 8383
rect 608 8461 662 8468
rect 608 8409 609 8461
rect 661 8409 662 8461
rect 608 8383 618 8409
rect 652 8383 662 8409
rect 608 8371 662 8383
rect 708 8417 762 8523
rect 808 8557 862 8569
rect 808 8531 818 8557
rect 852 8531 862 8557
rect 808 8479 809 8531
rect 861 8479 862 8531
rect 808 8472 862 8479
rect 908 8557 962 8753
rect 1008 8831 1062 8838
rect 1008 8779 1009 8831
rect 1061 8779 1062 8831
rect 1008 8753 1018 8779
rect 1052 8753 1062 8779
rect 1008 8741 1062 8753
rect 1108 8787 1162 8893
rect 1208 8927 1262 8939
rect 1208 8901 1218 8927
rect 1252 8901 1262 8927
rect 1208 8849 1209 8901
rect 1261 8849 1262 8901
rect 1208 8842 1262 8849
rect 1308 8927 1362 9033
rect 1408 9111 1462 9118
rect 1408 9059 1409 9111
rect 1461 9059 1462 9111
rect 1408 9033 1418 9059
rect 1452 9033 1462 9059
rect 1408 9021 1462 9033
rect 1508 9067 1562 9173
rect 1608 9207 1662 9219
rect 1608 9181 1618 9207
rect 1652 9181 1662 9207
rect 1608 9129 1609 9181
rect 1661 9129 1662 9181
rect 1608 9122 1662 9129
rect 1708 9207 1762 9313
rect 1808 9391 1862 9398
rect 1808 9339 1809 9391
rect 1861 9339 1862 9391
rect 1808 9313 1818 9339
rect 1852 9313 1862 9339
rect 1808 9301 1862 9313
rect 1908 9347 1962 9453
rect 2008 9487 2062 9499
rect 2008 9461 2018 9487
rect 2052 9461 2062 9487
rect 2008 9409 2009 9461
rect 2061 9409 2062 9461
rect 2008 9402 2062 9409
rect 2108 9487 2162 9593
rect 2208 9671 2262 9678
rect 2208 9619 2209 9671
rect 2261 9619 2262 9671
rect 2208 9593 2218 9619
rect 2252 9593 2262 9619
rect 2208 9581 2262 9593
rect 2308 9627 2362 9733
rect 2408 9767 2462 9779
rect 2408 9741 2418 9767
rect 2452 9741 2462 9767
rect 2408 9689 2409 9741
rect 2461 9689 2462 9741
rect 2408 9682 2462 9689
rect 2508 9767 2562 9940
rect 2602 9899 2668 9900
rect 2602 9847 2609 9899
rect 2661 9847 2668 9899
rect 2602 9846 2668 9847
rect 2508 9733 2518 9767
rect 2552 9733 2562 9767
rect 2308 9593 2318 9627
rect 2352 9593 2362 9627
rect 2108 9453 2118 9487
rect 2152 9453 2162 9487
rect 1908 9313 1918 9347
rect 1952 9313 1962 9347
rect 1708 9173 1718 9207
rect 1752 9173 1762 9207
rect 1508 9033 1518 9067
rect 1552 9033 1562 9067
rect 1308 8893 1318 8927
rect 1352 8893 1362 8927
rect 1108 8753 1118 8787
rect 1152 8753 1162 8787
rect 1002 8689 1068 8690
rect 1002 8637 1009 8689
rect 1061 8637 1068 8689
rect 1002 8636 1068 8637
rect 908 8523 918 8557
rect 952 8523 962 8557
rect 708 8383 718 8417
rect 752 8383 762 8417
rect 508 8243 518 8277
rect 552 8243 562 8277
rect 308 8103 318 8137
rect 352 8103 362 8137
rect 108 7963 118 7997
rect 152 7963 162 7997
rect 8 7857 62 7869
rect 8 7831 18 7857
rect 52 7831 62 7857
rect 8 7779 9 7831
rect 61 7779 62 7831
rect 8 7772 62 7779
rect 108 7857 162 7963
rect 208 8041 262 8048
rect 208 7989 209 8041
rect 261 7989 262 8041
rect 208 7963 218 7989
rect 252 7963 262 7989
rect 208 7951 262 7963
rect 308 7997 362 8103
rect 408 8137 462 8149
rect 408 8111 418 8137
rect 452 8111 462 8137
rect 408 8059 409 8111
rect 461 8059 462 8111
rect 408 8052 462 8059
rect 508 8137 562 8243
rect 608 8321 662 8328
rect 608 8269 609 8321
rect 661 8269 662 8321
rect 608 8243 618 8269
rect 652 8243 662 8269
rect 608 8231 662 8243
rect 708 8277 762 8383
rect 808 8417 862 8429
rect 808 8391 818 8417
rect 852 8391 862 8417
rect 808 8339 809 8391
rect 861 8339 862 8391
rect 808 8332 862 8339
rect 908 8417 962 8523
rect 1008 8601 1062 8608
rect 1008 8549 1009 8601
rect 1061 8549 1062 8601
rect 1008 8523 1018 8549
rect 1052 8523 1062 8549
rect 1008 8511 1062 8523
rect 1108 8557 1162 8753
rect 1208 8787 1262 8799
rect 1208 8761 1218 8787
rect 1252 8761 1262 8787
rect 1208 8709 1209 8761
rect 1261 8709 1262 8761
rect 1208 8702 1262 8709
rect 1308 8787 1362 8893
rect 1408 8971 1462 8978
rect 1408 8919 1409 8971
rect 1461 8919 1462 8971
rect 1408 8893 1418 8919
rect 1452 8893 1462 8919
rect 1408 8881 1462 8893
rect 1508 8927 1562 9033
rect 1608 9067 1662 9079
rect 1608 9041 1618 9067
rect 1652 9041 1662 9067
rect 1608 8989 1609 9041
rect 1661 8989 1662 9041
rect 1608 8982 1662 8989
rect 1708 9067 1762 9173
rect 1808 9251 1862 9258
rect 1808 9199 1809 9251
rect 1861 9199 1862 9251
rect 1808 9173 1818 9199
rect 1852 9173 1862 9199
rect 1808 9161 1862 9173
rect 1908 9207 1962 9313
rect 2008 9347 2062 9359
rect 2008 9321 2018 9347
rect 2052 9321 2062 9347
rect 2008 9269 2009 9321
rect 2061 9269 2062 9321
rect 2008 9262 2062 9269
rect 2108 9347 2162 9453
rect 2208 9531 2262 9538
rect 2208 9479 2209 9531
rect 2261 9479 2262 9531
rect 2208 9453 2218 9479
rect 2252 9453 2262 9479
rect 2208 9441 2262 9453
rect 2308 9487 2362 9593
rect 2408 9627 2462 9639
rect 2408 9601 2418 9627
rect 2452 9601 2462 9627
rect 2408 9549 2409 9601
rect 2461 9549 2462 9601
rect 2408 9542 2462 9549
rect 2508 9627 2562 9733
rect 2608 9811 2662 9818
rect 2608 9759 2609 9811
rect 2661 9759 2662 9811
rect 2608 9733 2618 9759
rect 2652 9733 2662 9759
rect 2608 9721 2662 9733
rect 2708 9767 2762 9940
rect 2802 9883 2868 9884
rect 2802 9831 2809 9883
rect 2861 9831 2868 9883
rect 2802 9830 2868 9831
rect 2708 9733 2718 9767
rect 2752 9733 2762 9767
rect 2508 9593 2518 9627
rect 2552 9593 2562 9627
rect 2308 9453 2318 9487
rect 2352 9453 2362 9487
rect 2108 9313 2118 9347
rect 2152 9313 2162 9347
rect 1908 9173 1918 9207
rect 1952 9173 1962 9207
rect 1708 9033 1718 9067
rect 1752 9033 1762 9067
rect 1508 8893 1518 8927
rect 1552 8893 1562 8927
rect 1308 8753 1318 8787
rect 1352 8753 1362 8787
rect 1202 8673 1268 8674
rect 1202 8621 1209 8673
rect 1261 8621 1268 8673
rect 1202 8620 1268 8621
rect 1108 8523 1118 8557
rect 1152 8523 1162 8557
rect 908 8383 918 8417
rect 952 8383 962 8417
rect 708 8243 718 8277
rect 752 8243 762 8277
rect 508 8103 518 8137
rect 552 8103 562 8137
rect 308 7963 318 7997
rect 352 7963 362 7997
rect 108 7823 118 7857
rect 152 7823 162 7857
rect 8 7717 62 7729
rect 8 7691 18 7717
rect 52 7691 62 7717
rect 8 7639 9 7691
rect 61 7639 62 7691
rect 8 7632 62 7639
rect 108 7717 162 7823
rect 208 7901 262 7908
rect 208 7849 209 7901
rect 261 7849 262 7901
rect 208 7823 218 7849
rect 252 7823 262 7849
rect 208 7811 262 7823
rect 308 7857 362 7963
rect 408 7997 462 8009
rect 408 7971 418 7997
rect 452 7971 462 7997
rect 408 7919 409 7971
rect 461 7919 462 7971
rect 408 7912 462 7919
rect 508 7997 562 8103
rect 608 8181 662 8188
rect 608 8129 609 8181
rect 661 8129 662 8181
rect 608 8103 618 8129
rect 652 8103 662 8129
rect 608 8091 662 8103
rect 708 8137 762 8243
rect 808 8277 862 8289
rect 808 8251 818 8277
rect 852 8251 862 8277
rect 808 8199 809 8251
rect 861 8199 862 8251
rect 808 8192 862 8199
rect 908 8277 962 8383
rect 1008 8461 1062 8468
rect 1008 8409 1009 8461
rect 1061 8409 1062 8461
rect 1008 8383 1018 8409
rect 1052 8383 1062 8409
rect 1008 8371 1062 8383
rect 1108 8417 1162 8523
rect 1208 8557 1262 8569
rect 1208 8531 1218 8557
rect 1252 8531 1262 8557
rect 1208 8479 1209 8531
rect 1261 8479 1262 8531
rect 1208 8472 1262 8479
rect 1308 8557 1362 8753
rect 1408 8831 1462 8838
rect 1408 8779 1409 8831
rect 1461 8779 1462 8831
rect 1408 8753 1418 8779
rect 1452 8753 1462 8779
rect 1408 8741 1462 8753
rect 1508 8787 1562 8893
rect 1608 8927 1662 8939
rect 1608 8901 1618 8927
rect 1652 8901 1662 8927
rect 1608 8849 1609 8901
rect 1661 8849 1662 8901
rect 1608 8842 1662 8849
rect 1708 8927 1762 9033
rect 1808 9111 1862 9118
rect 1808 9059 1809 9111
rect 1861 9059 1862 9111
rect 1808 9033 1818 9059
rect 1852 9033 1862 9059
rect 1808 9021 1862 9033
rect 1908 9067 1962 9173
rect 2008 9207 2062 9219
rect 2008 9181 2018 9207
rect 2052 9181 2062 9207
rect 2008 9129 2009 9181
rect 2061 9129 2062 9181
rect 2008 9122 2062 9129
rect 2108 9207 2162 9313
rect 2208 9391 2262 9398
rect 2208 9339 2209 9391
rect 2261 9339 2262 9391
rect 2208 9313 2218 9339
rect 2252 9313 2262 9339
rect 2208 9301 2262 9313
rect 2308 9347 2362 9453
rect 2408 9487 2462 9499
rect 2408 9461 2418 9487
rect 2452 9461 2462 9487
rect 2408 9409 2409 9461
rect 2461 9409 2462 9461
rect 2408 9402 2462 9409
rect 2508 9487 2562 9593
rect 2608 9671 2662 9678
rect 2608 9619 2609 9671
rect 2661 9619 2662 9671
rect 2608 9593 2618 9619
rect 2652 9593 2662 9619
rect 2608 9581 2662 9593
rect 2708 9627 2762 9733
rect 2808 9767 2862 9779
rect 2808 9741 2818 9767
rect 2852 9741 2862 9767
rect 2808 9689 2809 9741
rect 2861 9689 2862 9741
rect 2808 9682 2862 9689
rect 2908 9767 2962 9940
rect 3002 9899 3068 9900
rect 3002 9847 3009 9899
rect 3061 9847 3068 9899
rect 3002 9846 3068 9847
rect 2908 9733 2918 9767
rect 2952 9733 2962 9767
rect 2708 9593 2718 9627
rect 2752 9593 2762 9627
rect 2508 9453 2518 9487
rect 2552 9453 2562 9487
rect 2308 9313 2318 9347
rect 2352 9313 2362 9347
rect 2108 9173 2118 9207
rect 2152 9173 2162 9207
rect 1908 9033 1918 9067
rect 1952 9033 1962 9067
rect 1708 8893 1718 8927
rect 1752 8893 1762 8927
rect 1508 8753 1518 8787
rect 1552 8753 1562 8787
rect 1402 8689 1468 8690
rect 1402 8637 1409 8689
rect 1461 8637 1468 8689
rect 1402 8636 1468 8637
rect 1308 8523 1318 8557
rect 1352 8523 1362 8557
rect 1108 8383 1118 8417
rect 1152 8383 1162 8417
rect 908 8243 918 8277
rect 952 8243 962 8277
rect 708 8103 718 8137
rect 752 8103 762 8137
rect 508 7963 518 7997
rect 552 7963 562 7997
rect 308 7823 318 7857
rect 352 7823 362 7857
rect 108 7683 118 7717
rect 152 7683 162 7717
rect 8 7577 62 7589
rect 8 7551 18 7577
rect 52 7551 62 7577
rect 8 7499 9 7551
rect 61 7499 62 7551
rect 8 7492 62 7499
rect 108 7577 162 7683
rect 208 7761 262 7768
rect 208 7709 209 7761
rect 261 7709 262 7761
rect 208 7683 218 7709
rect 252 7683 262 7709
rect 208 7671 262 7683
rect 308 7717 362 7823
rect 408 7857 462 7869
rect 408 7831 418 7857
rect 452 7831 462 7857
rect 408 7779 409 7831
rect 461 7779 462 7831
rect 408 7772 462 7779
rect 508 7857 562 7963
rect 608 8041 662 8048
rect 608 7989 609 8041
rect 661 7989 662 8041
rect 608 7963 618 7989
rect 652 7963 662 7989
rect 608 7951 662 7963
rect 708 7997 762 8103
rect 808 8137 862 8149
rect 808 8111 818 8137
rect 852 8111 862 8137
rect 808 8059 809 8111
rect 861 8059 862 8111
rect 808 8052 862 8059
rect 908 8137 962 8243
rect 1008 8321 1062 8328
rect 1008 8269 1009 8321
rect 1061 8269 1062 8321
rect 1008 8243 1018 8269
rect 1052 8243 1062 8269
rect 1008 8231 1062 8243
rect 1108 8277 1162 8383
rect 1208 8417 1262 8429
rect 1208 8391 1218 8417
rect 1252 8391 1262 8417
rect 1208 8339 1209 8391
rect 1261 8339 1262 8391
rect 1208 8332 1262 8339
rect 1308 8417 1362 8523
rect 1408 8601 1462 8608
rect 1408 8549 1409 8601
rect 1461 8549 1462 8601
rect 1408 8523 1418 8549
rect 1452 8523 1462 8549
rect 1408 8511 1462 8523
rect 1508 8557 1562 8753
rect 1608 8787 1662 8799
rect 1608 8761 1618 8787
rect 1652 8761 1662 8787
rect 1608 8709 1609 8761
rect 1661 8709 1662 8761
rect 1608 8702 1662 8709
rect 1708 8787 1762 8893
rect 1808 8971 1862 8978
rect 1808 8919 1809 8971
rect 1861 8919 1862 8971
rect 1808 8893 1818 8919
rect 1852 8893 1862 8919
rect 1808 8881 1862 8893
rect 1908 8927 1962 9033
rect 2008 9067 2062 9079
rect 2008 9041 2018 9067
rect 2052 9041 2062 9067
rect 2008 8989 2009 9041
rect 2061 8989 2062 9041
rect 2008 8982 2062 8989
rect 2108 9067 2162 9173
rect 2208 9251 2262 9258
rect 2208 9199 2209 9251
rect 2261 9199 2262 9251
rect 2208 9173 2218 9199
rect 2252 9173 2262 9199
rect 2208 9161 2262 9173
rect 2308 9207 2362 9313
rect 2408 9347 2462 9359
rect 2408 9321 2418 9347
rect 2452 9321 2462 9347
rect 2408 9269 2409 9321
rect 2461 9269 2462 9321
rect 2408 9262 2462 9269
rect 2508 9347 2562 9453
rect 2608 9531 2662 9538
rect 2608 9479 2609 9531
rect 2661 9479 2662 9531
rect 2608 9453 2618 9479
rect 2652 9453 2662 9479
rect 2608 9441 2662 9453
rect 2708 9487 2762 9593
rect 2808 9627 2862 9639
rect 2808 9601 2818 9627
rect 2852 9601 2862 9627
rect 2808 9549 2809 9601
rect 2861 9549 2862 9601
rect 2808 9542 2862 9549
rect 2908 9627 2962 9733
rect 3008 9811 3062 9818
rect 3008 9759 3009 9811
rect 3061 9759 3062 9811
rect 3008 9733 3018 9759
rect 3052 9733 3062 9759
rect 3008 9721 3062 9733
rect 3108 9767 3162 9940
rect 3202 9883 3268 9884
rect 3202 9831 3209 9883
rect 3261 9831 3268 9883
rect 3202 9830 3268 9831
rect 3108 9733 3118 9767
rect 3152 9733 3162 9767
rect 2908 9593 2918 9627
rect 2952 9593 2962 9627
rect 2708 9453 2718 9487
rect 2752 9453 2762 9487
rect 2508 9313 2518 9347
rect 2552 9313 2562 9347
rect 2308 9173 2318 9207
rect 2352 9173 2362 9207
rect 2108 9033 2118 9067
rect 2152 9033 2162 9067
rect 1908 8893 1918 8927
rect 1952 8893 1962 8927
rect 1708 8753 1718 8787
rect 1752 8753 1762 8787
rect 1602 8673 1668 8674
rect 1602 8621 1609 8673
rect 1661 8621 1668 8673
rect 1602 8620 1668 8621
rect 1508 8523 1518 8557
rect 1552 8523 1562 8557
rect 1308 8383 1318 8417
rect 1352 8383 1362 8417
rect 1108 8243 1118 8277
rect 1152 8243 1162 8277
rect 908 8103 918 8137
rect 952 8103 962 8137
rect 708 7963 718 7997
rect 752 7963 762 7997
rect 508 7823 518 7857
rect 552 7823 562 7857
rect 308 7683 318 7717
rect 352 7683 362 7717
rect 108 7543 118 7577
rect 152 7543 162 7577
rect 2 7463 68 7464
rect 2 7411 9 7463
rect 61 7411 68 7463
rect 2 7410 68 7411
rect 8 7347 62 7359
rect 8 7321 18 7347
rect 52 7321 62 7347
rect 8 7269 9 7321
rect 61 7269 62 7321
rect 8 7262 62 7269
rect 108 7347 162 7543
rect 208 7621 262 7628
rect 208 7569 209 7621
rect 261 7569 262 7621
rect 208 7543 218 7569
rect 252 7543 262 7569
rect 208 7531 262 7543
rect 308 7577 362 7683
rect 408 7717 462 7729
rect 408 7691 418 7717
rect 452 7691 462 7717
rect 408 7639 409 7691
rect 461 7639 462 7691
rect 408 7632 462 7639
rect 508 7717 562 7823
rect 608 7901 662 7908
rect 608 7849 609 7901
rect 661 7849 662 7901
rect 608 7823 618 7849
rect 652 7823 662 7849
rect 608 7811 662 7823
rect 708 7857 762 7963
rect 808 7997 862 8009
rect 808 7971 818 7997
rect 852 7971 862 7997
rect 808 7919 809 7971
rect 861 7919 862 7971
rect 808 7912 862 7919
rect 908 7997 962 8103
rect 1008 8181 1062 8188
rect 1008 8129 1009 8181
rect 1061 8129 1062 8181
rect 1008 8103 1018 8129
rect 1052 8103 1062 8129
rect 1008 8091 1062 8103
rect 1108 8137 1162 8243
rect 1208 8277 1262 8289
rect 1208 8251 1218 8277
rect 1252 8251 1262 8277
rect 1208 8199 1209 8251
rect 1261 8199 1262 8251
rect 1208 8192 1262 8199
rect 1308 8277 1362 8383
rect 1408 8461 1462 8468
rect 1408 8409 1409 8461
rect 1461 8409 1462 8461
rect 1408 8383 1418 8409
rect 1452 8383 1462 8409
rect 1408 8371 1462 8383
rect 1508 8417 1562 8523
rect 1608 8557 1662 8569
rect 1608 8531 1618 8557
rect 1652 8531 1662 8557
rect 1608 8479 1609 8531
rect 1661 8479 1662 8531
rect 1608 8472 1662 8479
rect 1708 8557 1762 8753
rect 1808 8831 1862 8838
rect 1808 8779 1809 8831
rect 1861 8779 1862 8831
rect 1808 8753 1818 8779
rect 1852 8753 1862 8779
rect 1808 8741 1862 8753
rect 1908 8787 1962 8893
rect 2008 8927 2062 8939
rect 2008 8901 2018 8927
rect 2052 8901 2062 8927
rect 2008 8849 2009 8901
rect 2061 8849 2062 8901
rect 2008 8842 2062 8849
rect 2108 8927 2162 9033
rect 2208 9111 2262 9118
rect 2208 9059 2209 9111
rect 2261 9059 2262 9111
rect 2208 9033 2218 9059
rect 2252 9033 2262 9059
rect 2208 9021 2262 9033
rect 2308 9067 2362 9173
rect 2408 9207 2462 9219
rect 2408 9181 2418 9207
rect 2452 9181 2462 9207
rect 2408 9129 2409 9181
rect 2461 9129 2462 9181
rect 2408 9122 2462 9129
rect 2508 9207 2562 9313
rect 2608 9391 2662 9398
rect 2608 9339 2609 9391
rect 2661 9339 2662 9391
rect 2608 9313 2618 9339
rect 2652 9313 2662 9339
rect 2608 9301 2662 9313
rect 2708 9347 2762 9453
rect 2808 9487 2862 9499
rect 2808 9461 2818 9487
rect 2852 9461 2862 9487
rect 2808 9409 2809 9461
rect 2861 9409 2862 9461
rect 2808 9402 2862 9409
rect 2908 9487 2962 9593
rect 3008 9671 3062 9678
rect 3008 9619 3009 9671
rect 3061 9619 3062 9671
rect 3008 9593 3018 9619
rect 3052 9593 3062 9619
rect 3008 9581 3062 9593
rect 3108 9627 3162 9733
rect 3208 9767 3262 9779
rect 3208 9741 3218 9767
rect 3252 9741 3262 9767
rect 3208 9689 3209 9741
rect 3261 9689 3262 9741
rect 3208 9682 3262 9689
rect 3308 9767 3362 9940
rect 3402 9899 3468 9900
rect 3402 9847 3409 9899
rect 3461 9847 3468 9899
rect 3402 9846 3468 9847
rect 3308 9733 3318 9767
rect 3352 9733 3362 9767
rect 3108 9593 3118 9627
rect 3152 9593 3162 9627
rect 2908 9453 2918 9487
rect 2952 9453 2962 9487
rect 2708 9313 2718 9347
rect 2752 9313 2762 9347
rect 2508 9173 2518 9207
rect 2552 9173 2562 9207
rect 2308 9033 2318 9067
rect 2352 9033 2362 9067
rect 2108 8893 2118 8927
rect 2152 8893 2162 8927
rect 1908 8753 1918 8787
rect 1952 8753 1962 8787
rect 1802 8689 1868 8690
rect 1802 8637 1809 8689
rect 1861 8637 1868 8689
rect 1802 8636 1868 8637
rect 1708 8523 1718 8557
rect 1752 8523 1762 8557
rect 1508 8383 1518 8417
rect 1552 8383 1562 8417
rect 1308 8243 1318 8277
rect 1352 8243 1362 8277
rect 1108 8103 1118 8137
rect 1152 8103 1162 8137
rect 908 7963 918 7997
rect 952 7963 962 7997
rect 708 7823 718 7857
rect 752 7823 762 7857
rect 508 7683 518 7717
rect 552 7683 562 7717
rect 308 7543 318 7577
rect 352 7543 362 7577
rect 202 7479 268 7480
rect 202 7427 209 7479
rect 261 7427 268 7479
rect 202 7426 268 7427
rect 108 7313 118 7347
rect 152 7313 162 7347
rect 8 7207 62 7219
rect 8 7181 18 7207
rect 52 7181 62 7207
rect 8 7129 9 7181
rect 61 7129 62 7181
rect 8 7122 62 7129
rect 108 7207 162 7313
rect 208 7391 262 7398
rect 208 7339 209 7391
rect 261 7339 262 7391
rect 208 7313 218 7339
rect 252 7313 262 7339
rect 208 7301 262 7313
rect 308 7347 362 7543
rect 408 7577 462 7589
rect 408 7551 418 7577
rect 452 7551 462 7577
rect 408 7499 409 7551
rect 461 7499 462 7551
rect 408 7492 462 7499
rect 508 7577 562 7683
rect 608 7761 662 7768
rect 608 7709 609 7761
rect 661 7709 662 7761
rect 608 7683 618 7709
rect 652 7683 662 7709
rect 608 7671 662 7683
rect 708 7717 762 7823
rect 808 7857 862 7869
rect 808 7831 818 7857
rect 852 7831 862 7857
rect 808 7779 809 7831
rect 861 7779 862 7831
rect 808 7772 862 7779
rect 908 7857 962 7963
rect 1008 8041 1062 8048
rect 1008 7989 1009 8041
rect 1061 7989 1062 8041
rect 1008 7963 1018 7989
rect 1052 7963 1062 7989
rect 1008 7951 1062 7963
rect 1108 7997 1162 8103
rect 1208 8137 1262 8149
rect 1208 8111 1218 8137
rect 1252 8111 1262 8137
rect 1208 8059 1209 8111
rect 1261 8059 1262 8111
rect 1208 8052 1262 8059
rect 1308 8137 1362 8243
rect 1408 8321 1462 8328
rect 1408 8269 1409 8321
rect 1461 8269 1462 8321
rect 1408 8243 1418 8269
rect 1452 8243 1462 8269
rect 1408 8231 1462 8243
rect 1508 8277 1562 8383
rect 1608 8417 1662 8429
rect 1608 8391 1618 8417
rect 1652 8391 1662 8417
rect 1608 8339 1609 8391
rect 1661 8339 1662 8391
rect 1608 8332 1662 8339
rect 1708 8417 1762 8523
rect 1808 8601 1862 8608
rect 1808 8549 1809 8601
rect 1861 8549 1862 8601
rect 1808 8523 1818 8549
rect 1852 8523 1862 8549
rect 1808 8511 1862 8523
rect 1908 8557 1962 8753
rect 2008 8787 2062 8799
rect 2008 8761 2018 8787
rect 2052 8761 2062 8787
rect 2008 8709 2009 8761
rect 2061 8709 2062 8761
rect 2008 8702 2062 8709
rect 2108 8787 2162 8893
rect 2208 8971 2262 8978
rect 2208 8919 2209 8971
rect 2261 8919 2262 8971
rect 2208 8893 2218 8919
rect 2252 8893 2262 8919
rect 2208 8881 2262 8893
rect 2308 8927 2362 9033
rect 2408 9067 2462 9079
rect 2408 9041 2418 9067
rect 2452 9041 2462 9067
rect 2408 8989 2409 9041
rect 2461 8989 2462 9041
rect 2408 8982 2462 8989
rect 2508 9067 2562 9173
rect 2608 9251 2662 9258
rect 2608 9199 2609 9251
rect 2661 9199 2662 9251
rect 2608 9173 2618 9199
rect 2652 9173 2662 9199
rect 2608 9161 2662 9173
rect 2708 9207 2762 9313
rect 2808 9347 2862 9359
rect 2808 9321 2818 9347
rect 2852 9321 2862 9347
rect 2808 9269 2809 9321
rect 2861 9269 2862 9321
rect 2808 9262 2862 9269
rect 2908 9347 2962 9453
rect 3008 9531 3062 9538
rect 3008 9479 3009 9531
rect 3061 9479 3062 9531
rect 3008 9453 3018 9479
rect 3052 9453 3062 9479
rect 3008 9441 3062 9453
rect 3108 9487 3162 9593
rect 3208 9627 3262 9639
rect 3208 9601 3218 9627
rect 3252 9601 3262 9627
rect 3208 9549 3209 9601
rect 3261 9549 3262 9601
rect 3208 9542 3262 9549
rect 3308 9627 3362 9733
rect 3408 9811 3462 9818
rect 3408 9759 3409 9811
rect 3461 9759 3462 9811
rect 3408 9733 3418 9759
rect 3452 9733 3462 9759
rect 3408 9721 3462 9733
rect 3508 9767 3562 9940
rect 3602 9883 3668 9884
rect 3602 9831 3609 9883
rect 3661 9831 3668 9883
rect 3602 9830 3668 9831
rect 3508 9733 3518 9767
rect 3552 9733 3562 9767
rect 3308 9593 3318 9627
rect 3352 9593 3362 9627
rect 3108 9453 3118 9487
rect 3152 9453 3162 9487
rect 2908 9313 2918 9347
rect 2952 9313 2962 9347
rect 2708 9173 2718 9207
rect 2752 9173 2762 9207
rect 2508 9033 2518 9067
rect 2552 9033 2562 9067
rect 2308 8893 2318 8927
rect 2352 8893 2362 8927
rect 2108 8753 2118 8787
rect 2152 8753 2162 8787
rect 2002 8673 2068 8674
rect 2002 8621 2009 8673
rect 2061 8621 2068 8673
rect 2002 8620 2068 8621
rect 1908 8523 1918 8557
rect 1952 8523 1962 8557
rect 1708 8383 1718 8417
rect 1752 8383 1762 8417
rect 1508 8243 1518 8277
rect 1552 8243 1562 8277
rect 1308 8103 1318 8137
rect 1352 8103 1362 8137
rect 1108 7963 1118 7997
rect 1152 7963 1162 7997
rect 908 7823 918 7857
rect 952 7823 962 7857
rect 708 7683 718 7717
rect 752 7683 762 7717
rect 508 7543 518 7577
rect 552 7543 562 7577
rect 402 7463 468 7464
rect 402 7411 409 7463
rect 461 7411 468 7463
rect 402 7410 468 7411
rect 308 7313 318 7347
rect 352 7313 362 7347
rect 108 7173 118 7207
rect 152 7173 162 7207
rect 8 7067 62 7079
rect 8 7041 18 7067
rect 52 7041 62 7067
rect 8 6989 9 7041
rect 61 6989 62 7041
rect 8 6982 62 6989
rect 108 7067 162 7173
rect 208 7251 262 7258
rect 208 7199 209 7251
rect 261 7199 262 7251
rect 208 7173 218 7199
rect 252 7173 262 7199
rect 208 7161 262 7173
rect 308 7207 362 7313
rect 408 7347 462 7359
rect 408 7321 418 7347
rect 452 7321 462 7347
rect 408 7269 409 7321
rect 461 7269 462 7321
rect 408 7262 462 7269
rect 508 7347 562 7543
rect 608 7621 662 7628
rect 608 7569 609 7621
rect 661 7569 662 7621
rect 608 7543 618 7569
rect 652 7543 662 7569
rect 608 7531 662 7543
rect 708 7577 762 7683
rect 808 7717 862 7729
rect 808 7691 818 7717
rect 852 7691 862 7717
rect 808 7639 809 7691
rect 861 7639 862 7691
rect 808 7632 862 7639
rect 908 7717 962 7823
rect 1008 7901 1062 7908
rect 1008 7849 1009 7901
rect 1061 7849 1062 7901
rect 1008 7823 1018 7849
rect 1052 7823 1062 7849
rect 1008 7811 1062 7823
rect 1108 7857 1162 7963
rect 1208 7997 1262 8009
rect 1208 7971 1218 7997
rect 1252 7971 1262 7997
rect 1208 7919 1209 7971
rect 1261 7919 1262 7971
rect 1208 7912 1262 7919
rect 1308 7997 1362 8103
rect 1408 8181 1462 8188
rect 1408 8129 1409 8181
rect 1461 8129 1462 8181
rect 1408 8103 1418 8129
rect 1452 8103 1462 8129
rect 1408 8091 1462 8103
rect 1508 8137 1562 8243
rect 1608 8277 1662 8289
rect 1608 8251 1618 8277
rect 1652 8251 1662 8277
rect 1608 8199 1609 8251
rect 1661 8199 1662 8251
rect 1608 8192 1662 8199
rect 1708 8277 1762 8383
rect 1808 8461 1862 8468
rect 1808 8409 1809 8461
rect 1861 8409 1862 8461
rect 1808 8383 1818 8409
rect 1852 8383 1862 8409
rect 1808 8371 1862 8383
rect 1908 8417 1962 8523
rect 2008 8557 2062 8569
rect 2008 8531 2018 8557
rect 2052 8531 2062 8557
rect 2008 8479 2009 8531
rect 2061 8479 2062 8531
rect 2008 8472 2062 8479
rect 2108 8557 2162 8753
rect 2208 8831 2262 8838
rect 2208 8779 2209 8831
rect 2261 8779 2262 8831
rect 2208 8753 2218 8779
rect 2252 8753 2262 8779
rect 2208 8741 2262 8753
rect 2308 8787 2362 8893
rect 2408 8927 2462 8939
rect 2408 8901 2418 8927
rect 2452 8901 2462 8927
rect 2408 8849 2409 8901
rect 2461 8849 2462 8901
rect 2408 8842 2462 8849
rect 2508 8927 2562 9033
rect 2608 9111 2662 9118
rect 2608 9059 2609 9111
rect 2661 9059 2662 9111
rect 2608 9033 2618 9059
rect 2652 9033 2662 9059
rect 2608 9021 2662 9033
rect 2708 9067 2762 9173
rect 2808 9207 2862 9219
rect 2808 9181 2818 9207
rect 2852 9181 2862 9207
rect 2808 9129 2809 9181
rect 2861 9129 2862 9181
rect 2808 9122 2862 9129
rect 2908 9207 2962 9313
rect 3008 9391 3062 9398
rect 3008 9339 3009 9391
rect 3061 9339 3062 9391
rect 3008 9313 3018 9339
rect 3052 9313 3062 9339
rect 3008 9301 3062 9313
rect 3108 9347 3162 9453
rect 3208 9487 3262 9499
rect 3208 9461 3218 9487
rect 3252 9461 3262 9487
rect 3208 9409 3209 9461
rect 3261 9409 3262 9461
rect 3208 9402 3262 9409
rect 3308 9487 3362 9593
rect 3408 9671 3462 9678
rect 3408 9619 3409 9671
rect 3461 9619 3462 9671
rect 3408 9593 3418 9619
rect 3452 9593 3462 9619
rect 3408 9581 3462 9593
rect 3508 9627 3562 9733
rect 3608 9767 3662 9779
rect 3608 9741 3618 9767
rect 3652 9741 3662 9767
rect 3608 9689 3609 9741
rect 3661 9689 3662 9741
rect 3608 9682 3662 9689
rect 3708 9767 3762 9940
rect 3802 9899 3868 9900
rect 3802 9847 3809 9899
rect 3861 9847 3868 9899
rect 3802 9846 3868 9847
rect 3708 9733 3718 9767
rect 3752 9733 3762 9767
rect 3508 9593 3518 9627
rect 3552 9593 3562 9627
rect 3308 9453 3318 9487
rect 3352 9453 3362 9487
rect 3108 9313 3118 9347
rect 3152 9313 3162 9347
rect 2908 9173 2918 9207
rect 2952 9173 2962 9207
rect 2708 9033 2718 9067
rect 2752 9033 2762 9067
rect 2508 8893 2518 8927
rect 2552 8893 2562 8927
rect 2308 8753 2318 8787
rect 2352 8753 2362 8787
rect 2202 8689 2268 8690
rect 2202 8637 2209 8689
rect 2261 8637 2268 8689
rect 2202 8636 2268 8637
rect 2108 8523 2118 8557
rect 2152 8523 2162 8557
rect 1908 8383 1918 8417
rect 1952 8383 1962 8417
rect 1708 8243 1718 8277
rect 1752 8243 1762 8277
rect 1508 8103 1518 8137
rect 1552 8103 1562 8137
rect 1308 7963 1318 7997
rect 1352 7963 1362 7997
rect 1108 7823 1118 7857
rect 1152 7823 1162 7857
rect 908 7683 918 7717
rect 952 7683 962 7717
rect 708 7543 718 7577
rect 752 7543 762 7577
rect 602 7479 668 7480
rect 602 7427 609 7479
rect 661 7427 668 7479
rect 602 7426 668 7427
rect 508 7313 518 7347
rect 552 7313 562 7347
rect 308 7173 318 7207
rect 352 7173 362 7207
rect 108 7033 118 7067
rect 152 7033 162 7067
rect 8 6927 62 6939
rect 8 6901 18 6927
rect 52 6901 62 6927
rect 8 6849 9 6901
rect 61 6849 62 6901
rect 8 6842 62 6849
rect 108 6927 162 7033
rect 208 7111 262 7118
rect 208 7059 209 7111
rect 261 7059 262 7111
rect 208 7033 218 7059
rect 252 7033 262 7059
rect 208 7021 262 7033
rect 308 7067 362 7173
rect 408 7207 462 7219
rect 408 7181 418 7207
rect 452 7181 462 7207
rect 408 7129 409 7181
rect 461 7129 462 7181
rect 408 7122 462 7129
rect 508 7207 562 7313
rect 608 7391 662 7398
rect 608 7339 609 7391
rect 661 7339 662 7391
rect 608 7313 618 7339
rect 652 7313 662 7339
rect 608 7301 662 7313
rect 708 7347 762 7543
rect 808 7577 862 7589
rect 808 7551 818 7577
rect 852 7551 862 7577
rect 808 7499 809 7551
rect 861 7499 862 7551
rect 808 7492 862 7499
rect 908 7577 962 7683
rect 1008 7761 1062 7768
rect 1008 7709 1009 7761
rect 1061 7709 1062 7761
rect 1008 7683 1018 7709
rect 1052 7683 1062 7709
rect 1008 7671 1062 7683
rect 1108 7717 1162 7823
rect 1208 7857 1262 7869
rect 1208 7831 1218 7857
rect 1252 7831 1262 7857
rect 1208 7779 1209 7831
rect 1261 7779 1262 7831
rect 1208 7772 1262 7779
rect 1308 7857 1362 7963
rect 1408 8041 1462 8048
rect 1408 7989 1409 8041
rect 1461 7989 1462 8041
rect 1408 7963 1418 7989
rect 1452 7963 1462 7989
rect 1408 7951 1462 7963
rect 1508 7997 1562 8103
rect 1608 8137 1662 8149
rect 1608 8111 1618 8137
rect 1652 8111 1662 8137
rect 1608 8059 1609 8111
rect 1661 8059 1662 8111
rect 1608 8052 1662 8059
rect 1708 8137 1762 8243
rect 1808 8321 1862 8328
rect 1808 8269 1809 8321
rect 1861 8269 1862 8321
rect 1808 8243 1818 8269
rect 1852 8243 1862 8269
rect 1808 8231 1862 8243
rect 1908 8277 1962 8383
rect 2008 8417 2062 8429
rect 2008 8391 2018 8417
rect 2052 8391 2062 8417
rect 2008 8339 2009 8391
rect 2061 8339 2062 8391
rect 2008 8332 2062 8339
rect 2108 8417 2162 8523
rect 2208 8601 2262 8608
rect 2208 8549 2209 8601
rect 2261 8549 2262 8601
rect 2208 8523 2218 8549
rect 2252 8523 2262 8549
rect 2208 8511 2262 8523
rect 2308 8557 2362 8753
rect 2408 8787 2462 8799
rect 2408 8761 2418 8787
rect 2452 8761 2462 8787
rect 2408 8709 2409 8761
rect 2461 8709 2462 8761
rect 2408 8702 2462 8709
rect 2508 8787 2562 8893
rect 2608 8971 2662 8978
rect 2608 8919 2609 8971
rect 2661 8919 2662 8971
rect 2608 8893 2618 8919
rect 2652 8893 2662 8919
rect 2608 8881 2662 8893
rect 2708 8927 2762 9033
rect 2808 9067 2862 9079
rect 2808 9041 2818 9067
rect 2852 9041 2862 9067
rect 2808 8989 2809 9041
rect 2861 8989 2862 9041
rect 2808 8982 2862 8989
rect 2908 9067 2962 9173
rect 3008 9251 3062 9258
rect 3008 9199 3009 9251
rect 3061 9199 3062 9251
rect 3008 9173 3018 9199
rect 3052 9173 3062 9199
rect 3008 9161 3062 9173
rect 3108 9207 3162 9313
rect 3208 9347 3262 9359
rect 3208 9321 3218 9347
rect 3252 9321 3262 9347
rect 3208 9269 3209 9321
rect 3261 9269 3262 9321
rect 3208 9262 3262 9269
rect 3308 9347 3362 9453
rect 3408 9531 3462 9538
rect 3408 9479 3409 9531
rect 3461 9479 3462 9531
rect 3408 9453 3418 9479
rect 3452 9453 3462 9479
rect 3408 9441 3462 9453
rect 3508 9487 3562 9593
rect 3608 9627 3662 9639
rect 3608 9601 3618 9627
rect 3652 9601 3662 9627
rect 3608 9549 3609 9601
rect 3661 9549 3662 9601
rect 3608 9542 3662 9549
rect 3708 9627 3762 9733
rect 3808 9811 3862 9818
rect 3808 9759 3809 9811
rect 3861 9759 3862 9811
rect 3808 9733 3818 9759
rect 3852 9733 3862 9759
rect 3808 9721 3862 9733
rect 3908 9767 3962 9940
rect 4002 9883 4068 9884
rect 4002 9831 4009 9883
rect 4061 9831 4068 9883
rect 4002 9830 4068 9831
rect 3908 9733 3918 9767
rect 3952 9733 3962 9767
rect 3708 9593 3718 9627
rect 3752 9593 3762 9627
rect 3508 9453 3518 9487
rect 3552 9453 3562 9487
rect 3308 9313 3318 9347
rect 3352 9313 3362 9347
rect 3108 9173 3118 9207
rect 3152 9173 3162 9207
rect 2908 9033 2918 9067
rect 2952 9033 2962 9067
rect 2708 8893 2718 8927
rect 2752 8893 2762 8927
rect 2508 8753 2518 8787
rect 2552 8753 2562 8787
rect 2402 8673 2468 8674
rect 2402 8621 2409 8673
rect 2461 8621 2468 8673
rect 2402 8620 2468 8621
rect 2308 8523 2318 8557
rect 2352 8523 2362 8557
rect 2108 8383 2118 8417
rect 2152 8383 2162 8417
rect 1908 8243 1918 8277
rect 1952 8243 1962 8277
rect 1708 8103 1718 8137
rect 1752 8103 1762 8137
rect 1508 7963 1518 7997
rect 1552 7963 1562 7997
rect 1308 7823 1318 7857
rect 1352 7823 1362 7857
rect 1108 7683 1118 7717
rect 1152 7683 1162 7717
rect 908 7543 918 7577
rect 952 7543 962 7577
rect 802 7463 868 7464
rect 802 7411 809 7463
rect 861 7411 868 7463
rect 802 7410 868 7411
rect 708 7313 718 7347
rect 752 7313 762 7347
rect 508 7173 518 7207
rect 552 7173 562 7207
rect 308 7033 318 7067
rect 352 7033 362 7067
rect 108 6893 118 6927
rect 152 6893 162 6927
rect 8 6787 62 6799
rect 8 6761 18 6787
rect 52 6761 62 6787
rect 8 6709 9 6761
rect 61 6709 62 6761
rect 8 6702 62 6709
rect 108 6787 162 6893
rect 208 6971 262 6978
rect 208 6919 209 6971
rect 261 6919 262 6971
rect 208 6893 218 6919
rect 252 6893 262 6919
rect 208 6881 262 6893
rect 308 6927 362 7033
rect 408 7067 462 7079
rect 408 7041 418 7067
rect 452 7041 462 7067
rect 408 6989 409 7041
rect 461 6989 462 7041
rect 408 6982 462 6989
rect 508 7067 562 7173
rect 608 7251 662 7258
rect 608 7199 609 7251
rect 661 7199 662 7251
rect 608 7173 618 7199
rect 652 7173 662 7199
rect 608 7161 662 7173
rect 708 7207 762 7313
rect 808 7347 862 7359
rect 808 7321 818 7347
rect 852 7321 862 7347
rect 808 7269 809 7321
rect 861 7269 862 7321
rect 808 7262 862 7269
rect 908 7347 962 7543
rect 1008 7621 1062 7628
rect 1008 7569 1009 7621
rect 1061 7569 1062 7621
rect 1008 7543 1018 7569
rect 1052 7543 1062 7569
rect 1008 7531 1062 7543
rect 1108 7577 1162 7683
rect 1208 7717 1262 7729
rect 1208 7691 1218 7717
rect 1252 7691 1262 7717
rect 1208 7639 1209 7691
rect 1261 7639 1262 7691
rect 1208 7632 1262 7639
rect 1308 7717 1362 7823
rect 1408 7901 1462 7908
rect 1408 7849 1409 7901
rect 1461 7849 1462 7901
rect 1408 7823 1418 7849
rect 1452 7823 1462 7849
rect 1408 7811 1462 7823
rect 1508 7857 1562 7963
rect 1608 7997 1662 8009
rect 1608 7971 1618 7997
rect 1652 7971 1662 7997
rect 1608 7919 1609 7971
rect 1661 7919 1662 7971
rect 1608 7912 1662 7919
rect 1708 7997 1762 8103
rect 1808 8181 1862 8188
rect 1808 8129 1809 8181
rect 1861 8129 1862 8181
rect 1808 8103 1818 8129
rect 1852 8103 1862 8129
rect 1808 8091 1862 8103
rect 1908 8137 1962 8243
rect 2008 8277 2062 8289
rect 2008 8251 2018 8277
rect 2052 8251 2062 8277
rect 2008 8199 2009 8251
rect 2061 8199 2062 8251
rect 2008 8192 2062 8199
rect 2108 8277 2162 8383
rect 2208 8461 2262 8468
rect 2208 8409 2209 8461
rect 2261 8409 2262 8461
rect 2208 8383 2218 8409
rect 2252 8383 2262 8409
rect 2208 8371 2262 8383
rect 2308 8417 2362 8523
rect 2408 8557 2462 8569
rect 2408 8531 2418 8557
rect 2452 8531 2462 8557
rect 2408 8479 2409 8531
rect 2461 8479 2462 8531
rect 2408 8472 2462 8479
rect 2508 8557 2562 8753
rect 2608 8831 2662 8838
rect 2608 8779 2609 8831
rect 2661 8779 2662 8831
rect 2608 8753 2618 8779
rect 2652 8753 2662 8779
rect 2608 8741 2662 8753
rect 2708 8787 2762 8893
rect 2808 8927 2862 8939
rect 2808 8901 2818 8927
rect 2852 8901 2862 8927
rect 2808 8849 2809 8901
rect 2861 8849 2862 8901
rect 2808 8842 2862 8849
rect 2908 8927 2962 9033
rect 3008 9111 3062 9118
rect 3008 9059 3009 9111
rect 3061 9059 3062 9111
rect 3008 9033 3018 9059
rect 3052 9033 3062 9059
rect 3008 9021 3062 9033
rect 3108 9067 3162 9173
rect 3208 9207 3262 9219
rect 3208 9181 3218 9207
rect 3252 9181 3262 9207
rect 3208 9129 3209 9181
rect 3261 9129 3262 9181
rect 3208 9122 3262 9129
rect 3308 9207 3362 9313
rect 3408 9391 3462 9398
rect 3408 9339 3409 9391
rect 3461 9339 3462 9391
rect 3408 9313 3418 9339
rect 3452 9313 3462 9339
rect 3408 9301 3462 9313
rect 3508 9347 3562 9453
rect 3608 9487 3662 9499
rect 3608 9461 3618 9487
rect 3652 9461 3662 9487
rect 3608 9409 3609 9461
rect 3661 9409 3662 9461
rect 3608 9402 3662 9409
rect 3708 9487 3762 9593
rect 3808 9671 3862 9678
rect 3808 9619 3809 9671
rect 3861 9619 3862 9671
rect 3808 9593 3818 9619
rect 3852 9593 3862 9619
rect 3808 9581 3862 9593
rect 3908 9627 3962 9733
rect 4008 9767 4062 9779
rect 4008 9741 4018 9767
rect 4052 9741 4062 9767
rect 4008 9689 4009 9741
rect 4061 9689 4062 9741
rect 4008 9682 4062 9689
rect 4108 9767 4162 9940
rect 4202 9899 4268 9900
rect 4202 9847 4209 9899
rect 4261 9847 4268 9899
rect 4202 9846 4268 9847
rect 4108 9733 4118 9767
rect 4152 9733 4162 9767
rect 3908 9593 3918 9627
rect 3952 9593 3962 9627
rect 3708 9453 3718 9487
rect 3752 9453 3762 9487
rect 3508 9313 3518 9347
rect 3552 9313 3562 9347
rect 3308 9173 3318 9207
rect 3352 9173 3362 9207
rect 3108 9033 3118 9067
rect 3152 9033 3162 9067
rect 2908 8893 2918 8927
rect 2952 8893 2962 8927
rect 2708 8753 2718 8787
rect 2752 8753 2762 8787
rect 2602 8689 2668 8690
rect 2602 8637 2609 8689
rect 2661 8637 2668 8689
rect 2602 8636 2668 8637
rect 2508 8523 2518 8557
rect 2552 8523 2562 8557
rect 2308 8383 2318 8417
rect 2352 8383 2362 8417
rect 2108 8243 2118 8277
rect 2152 8243 2162 8277
rect 1908 8103 1918 8137
rect 1952 8103 1962 8137
rect 1708 7963 1718 7997
rect 1752 7963 1762 7997
rect 1508 7823 1518 7857
rect 1552 7823 1562 7857
rect 1308 7683 1318 7717
rect 1352 7683 1362 7717
rect 1108 7543 1118 7577
rect 1152 7543 1162 7577
rect 1002 7479 1068 7480
rect 1002 7427 1009 7479
rect 1061 7427 1068 7479
rect 1002 7426 1068 7427
rect 908 7313 918 7347
rect 952 7313 962 7347
rect 708 7173 718 7207
rect 752 7173 762 7207
rect 508 7033 518 7067
rect 552 7033 562 7067
rect 308 6893 318 6927
rect 352 6893 362 6927
rect 108 6753 118 6787
rect 152 6753 162 6787
rect 8 6647 62 6659
rect 8 6621 18 6647
rect 52 6621 62 6647
rect 8 6569 9 6621
rect 61 6569 62 6621
rect 8 6562 62 6569
rect 108 6647 162 6753
rect 208 6831 262 6838
rect 208 6779 209 6831
rect 261 6779 262 6831
rect 208 6753 218 6779
rect 252 6753 262 6779
rect 208 6741 262 6753
rect 308 6787 362 6893
rect 408 6927 462 6939
rect 408 6901 418 6927
rect 452 6901 462 6927
rect 408 6849 409 6901
rect 461 6849 462 6901
rect 408 6842 462 6849
rect 508 6927 562 7033
rect 608 7111 662 7118
rect 608 7059 609 7111
rect 661 7059 662 7111
rect 608 7033 618 7059
rect 652 7033 662 7059
rect 608 7021 662 7033
rect 708 7067 762 7173
rect 808 7207 862 7219
rect 808 7181 818 7207
rect 852 7181 862 7207
rect 808 7129 809 7181
rect 861 7129 862 7181
rect 808 7122 862 7129
rect 908 7207 962 7313
rect 1008 7391 1062 7398
rect 1008 7339 1009 7391
rect 1061 7339 1062 7391
rect 1008 7313 1018 7339
rect 1052 7313 1062 7339
rect 1008 7301 1062 7313
rect 1108 7347 1162 7543
rect 1208 7577 1262 7589
rect 1208 7551 1218 7577
rect 1252 7551 1262 7577
rect 1208 7499 1209 7551
rect 1261 7499 1262 7551
rect 1208 7492 1262 7499
rect 1308 7577 1362 7683
rect 1408 7761 1462 7768
rect 1408 7709 1409 7761
rect 1461 7709 1462 7761
rect 1408 7683 1418 7709
rect 1452 7683 1462 7709
rect 1408 7671 1462 7683
rect 1508 7717 1562 7823
rect 1608 7857 1662 7869
rect 1608 7831 1618 7857
rect 1652 7831 1662 7857
rect 1608 7779 1609 7831
rect 1661 7779 1662 7831
rect 1608 7772 1662 7779
rect 1708 7857 1762 7963
rect 1808 8041 1862 8048
rect 1808 7989 1809 8041
rect 1861 7989 1862 8041
rect 1808 7963 1818 7989
rect 1852 7963 1862 7989
rect 1808 7951 1862 7963
rect 1908 7997 1962 8103
rect 2008 8137 2062 8149
rect 2008 8111 2018 8137
rect 2052 8111 2062 8137
rect 2008 8059 2009 8111
rect 2061 8059 2062 8111
rect 2008 8052 2062 8059
rect 2108 8137 2162 8243
rect 2208 8321 2262 8328
rect 2208 8269 2209 8321
rect 2261 8269 2262 8321
rect 2208 8243 2218 8269
rect 2252 8243 2262 8269
rect 2208 8231 2262 8243
rect 2308 8277 2362 8383
rect 2408 8417 2462 8429
rect 2408 8391 2418 8417
rect 2452 8391 2462 8417
rect 2408 8339 2409 8391
rect 2461 8339 2462 8391
rect 2408 8332 2462 8339
rect 2508 8417 2562 8523
rect 2608 8601 2662 8608
rect 2608 8549 2609 8601
rect 2661 8549 2662 8601
rect 2608 8523 2618 8549
rect 2652 8523 2662 8549
rect 2608 8511 2662 8523
rect 2708 8557 2762 8753
rect 2808 8787 2862 8799
rect 2808 8761 2818 8787
rect 2852 8761 2862 8787
rect 2808 8709 2809 8761
rect 2861 8709 2862 8761
rect 2808 8702 2862 8709
rect 2908 8787 2962 8893
rect 3008 8971 3062 8978
rect 3008 8919 3009 8971
rect 3061 8919 3062 8971
rect 3008 8893 3018 8919
rect 3052 8893 3062 8919
rect 3008 8881 3062 8893
rect 3108 8927 3162 9033
rect 3208 9067 3262 9079
rect 3208 9041 3218 9067
rect 3252 9041 3262 9067
rect 3208 8989 3209 9041
rect 3261 8989 3262 9041
rect 3208 8982 3262 8989
rect 3308 9067 3362 9173
rect 3408 9251 3462 9258
rect 3408 9199 3409 9251
rect 3461 9199 3462 9251
rect 3408 9173 3418 9199
rect 3452 9173 3462 9199
rect 3408 9161 3462 9173
rect 3508 9207 3562 9313
rect 3608 9347 3662 9359
rect 3608 9321 3618 9347
rect 3652 9321 3662 9347
rect 3608 9269 3609 9321
rect 3661 9269 3662 9321
rect 3608 9262 3662 9269
rect 3708 9347 3762 9453
rect 3808 9531 3862 9538
rect 3808 9479 3809 9531
rect 3861 9479 3862 9531
rect 3808 9453 3818 9479
rect 3852 9453 3862 9479
rect 3808 9441 3862 9453
rect 3908 9487 3962 9593
rect 4008 9627 4062 9639
rect 4008 9601 4018 9627
rect 4052 9601 4062 9627
rect 4008 9549 4009 9601
rect 4061 9549 4062 9601
rect 4008 9542 4062 9549
rect 4108 9627 4162 9733
rect 4208 9811 4262 9818
rect 4208 9759 4209 9811
rect 4261 9759 4262 9811
rect 4208 9733 4218 9759
rect 4252 9733 4262 9759
rect 4208 9721 4262 9733
rect 4308 9767 4362 9940
rect 4402 9883 4468 9884
rect 4402 9831 4409 9883
rect 4461 9831 4468 9883
rect 4402 9830 4468 9831
rect 4308 9733 4318 9767
rect 4352 9733 4362 9767
rect 4108 9593 4118 9627
rect 4152 9593 4162 9627
rect 3908 9453 3918 9487
rect 3952 9453 3962 9487
rect 3708 9313 3718 9347
rect 3752 9313 3762 9347
rect 3508 9173 3518 9207
rect 3552 9173 3562 9207
rect 3308 9033 3318 9067
rect 3352 9033 3362 9067
rect 3108 8893 3118 8927
rect 3152 8893 3162 8927
rect 2908 8753 2918 8787
rect 2952 8753 2962 8787
rect 2802 8673 2868 8674
rect 2802 8621 2809 8673
rect 2861 8621 2868 8673
rect 2802 8620 2868 8621
rect 2708 8523 2718 8557
rect 2752 8523 2762 8557
rect 2508 8383 2518 8417
rect 2552 8383 2562 8417
rect 2308 8243 2318 8277
rect 2352 8243 2362 8277
rect 2108 8103 2118 8137
rect 2152 8103 2162 8137
rect 1908 7963 1918 7997
rect 1952 7963 1962 7997
rect 1708 7823 1718 7857
rect 1752 7823 1762 7857
rect 1508 7683 1518 7717
rect 1552 7683 1562 7717
rect 1308 7543 1318 7577
rect 1352 7543 1362 7577
rect 1202 7463 1268 7464
rect 1202 7411 1209 7463
rect 1261 7411 1268 7463
rect 1202 7410 1268 7411
rect 1108 7313 1118 7347
rect 1152 7313 1162 7347
rect 908 7173 918 7207
rect 952 7173 962 7207
rect 708 7033 718 7067
rect 752 7033 762 7067
rect 508 6893 518 6927
rect 552 6893 562 6927
rect 308 6753 318 6787
rect 352 6753 362 6787
rect 108 6613 118 6647
rect 152 6613 162 6647
rect 8 6507 62 6519
rect 8 6481 18 6507
rect 52 6481 62 6507
rect 8 6429 9 6481
rect 61 6429 62 6481
rect 8 6422 62 6429
rect 108 6507 162 6613
rect 208 6691 262 6698
rect 208 6639 209 6691
rect 261 6639 262 6691
rect 208 6613 218 6639
rect 252 6613 262 6639
rect 208 6601 262 6613
rect 308 6647 362 6753
rect 408 6787 462 6799
rect 408 6761 418 6787
rect 452 6761 462 6787
rect 408 6709 409 6761
rect 461 6709 462 6761
rect 408 6702 462 6709
rect 508 6787 562 6893
rect 608 6971 662 6978
rect 608 6919 609 6971
rect 661 6919 662 6971
rect 608 6893 618 6919
rect 652 6893 662 6919
rect 608 6881 662 6893
rect 708 6927 762 7033
rect 808 7067 862 7079
rect 808 7041 818 7067
rect 852 7041 862 7067
rect 808 6989 809 7041
rect 861 6989 862 7041
rect 808 6982 862 6989
rect 908 7067 962 7173
rect 1008 7251 1062 7258
rect 1008 7199 1009 7251
rect 1061 7199 1062 7251
rect 1008 7173 1018 7199
rect 1052 7173 1062 7199
rect 1008 7161 1062 7173
rect 1108 7207 1162 7313
rect 1208 7347 1262 7359
rect 1208 7321 1218 7347
rect 1252 7321 1262 7347
rect 1208 7269 1209 7321
rect 1261 7269 1262 7321
rect 1208 7262 1262 7269
rect 1308 7347 1362 7543
rect 1408 7621 1462 7628
rect 1408 7569 1409 7621
rect 1461 7569 1462 7621
rect 1408 7543 1418 7569
rect 1452 7543 1462 7569
rect 1408 7531 1462 7543
rect 1508 7577 1562 7683
rect 1608 7717 1662 7729
rect 1608 7691 1618 7717
rect 1652 7691 1662 7717
rect 1608 7639 1609 7691
rect 1661 7639 1662 7691
rect 1608 7632 1662 7639
rect 1708 7717 1762 7823
rect 1808 7901 1862 7908
rect 1808 7849 1809 7901
rect 1861 7849 1862 7901
rect 1808 7823 1818 7849
rect 1852 7823 1862 7849
rect 1808 7811 1862 7823
rect 1908 7857 1962 7963
rect 2008 7997 2062 8009
rect 2008 7971 2018 7997
rect 2052 7971 2062 7997
rect 2008 7919 2009 7971
rect 2061 7919 2062 7971
rect 2008 7912 2062 7919
rect 2108 7997 2162 8103
rect 2208 8181 2262 8188
rect 2208 8129 2209 8181
rect 2261 8129 2262 8181
rect 2208 8103 2218 8129
rect 2252 8103 2262 8129
rect 2208 8091 2262 8103
rect 2308 8137 2362 8243
rect 2408 8277 2462 8289
rect 2408 8251 2418 8277
rect 2452 8251 2462 8277
rect 2408 8199 2409 8251
rect 2461 8199 2462 8251
rect 2408 8192 2462 8199
rect 2508 8277 2562 8383
rect 2608 8461 2662 8468
rect 2608 8409 2609 8461
rect 2661 8409 2662 8461
rect 2608 8383 2618 8409
rect 2652 8383 2662 8409
rect 2608 8371 2662 8383
rect 2708 8417 2762 8523
rect 2808 8557 2862 8569
rect 2808 8531 2818 8557
rect 2852 8531 2862 8557
rect 2808 8479 2809 8531
rect 2861 8479 2862 8531
rect 2808 8472 2862 8479
rect 2908 8557 2962 8753
rect 3008 8831 3062 8838
rect 3008 8779 3009 8831
rect 3061 8779 3062 8831
rect 3008 8753 3018 8779
rect 3052 8753 3062 8779
rect 3008 8741 3062 8753
rect 3108 8787 3162 8893
rect 3208 8927 3262 8939
rect 3208 8901 3218 8927
rect 3252 8901 3262 8927
rect 3208 8849 3209 8901
rect 3261 8849 3262 8901
rect 3208 8842 3262 8849
rect 3308 8927 3362 9033
rect 3408 9111 3462 9118
rect 3408 9059 3409 9111
rect 3461 9059 3462 9111
rect 3408 9033 3418 9059
rect 3452 9033 3462 9059
rect 3408 9021 3462 9033
rect 3508 9067 3562 9173
rect 3608 9207 3662 9219
rect 3608 9181 3618 9207
rect 3652 9181 3662 9207
rect 3608 9129 3609 9181
rect 3661 9129 3662 9181
rect 3608 9122 3662 9129
rect 3708 9207 3762 9313
rect 3808 9391 3862 9398
rect 3808 9339 3809 9391
rect 3861 9339 3862 9391
rect 3808 9313 3818 9339
rect 3852 9313 3862 9339
rect 3808 9301 3862 9313
rect 3908 9347 3962 9453
rect 4008 9487 4062 9499
rect 4008 9461 4018 9487
rect 4052 9461 4062 9487
rect 4008 9409 4009 9461
rect 4061 9409 4062 9461
rect 4008 9402 4062 9409
rect 4108 9487 4162 9593
rect 4208 9671 4262 9678
rect 4208 9619 4209 9671
rect 4261 9619 4262 9671
rect 4208 9593 4218 9619
rect 4252 9593 4262 9619
rect 4208 9581 4262 9593
rect 4308 9627 4362 9733
rect 4408 9767 4462 9779
rect 4408 9741 4418 9767
rect 4452 9741 4462 9767
rect 4408 9689 4409 9741
rect 4461 9689 4462 9741
rect 4408 9682 4462 9689
rect 4508 9767 4562 9940
rect 4602 9899 4668 9900
rect 4602 9847 4609 9899
rect 4661 9847 4668 9899
rect 4602 9846 4668 9847
rect 4508 9733 4518 9767
rect 4552 9733 4562 9767
rect 4308 9593 4318 9627
rect 4352 9593 4362 9627
rect 4108 9453 4118 9487
rect 4152 9453 4162 9487
rect 3908 9313 3918 9347
rect 3952 9313 3962 9347
rect 3708 9173 3718 9207
rect 3752 9173 3762 9207
rect 3508 9033 3518 9067
rect 3552 9033 3562 9067
rect 3308 8893 3318 8927
rect 3352 8893 3362 8927
rect 3108 8753 3118 8787
rect 3152 8753 3162 8787
rect 3002 8689 3068 8690
rect 3002 8637 3009 8689
rect 3061 8637 3068 8689
rect 3002 8636 3068 8637
rect 2908 8523 2918 8557
rect 2952 8523 2962 8557
rect 2708 8383 2718 8417
rect 2752 8383 2762 8417
rect 2508 8243 2518 8277
rect 2552 8243 2562 8277
rect 2308 8103 2318 8137
rect 2352 8103 2362 8137
rect 2108 7963 2118 7997
rect 2152 7963 2162 7997
rect 1908 7823 1918 7857
rect 1952 7823 1962 7857
rect 1708 7683 1718 7717
rect 1752 7683 1762 7717
rect 1508 7543 1518 7577
rect 1552 7543 1562 7577
rect 1402 7479 1468 7480
rect 1402 7427 1409 7479
rect 1461 7427 1468 7479
rect 1402 7426 1468 7427
rect 1308 7313 1318 7347
rect 1352 7313 1362 7347
rect 1108 7173 1118 7207
rect 1152 7173 1162 7207
rect 908 7033 918 7067
rect 952 7033 962 7067
rect 708 6893 718 6927
rect 752 6893 762 6927
rect 508 6753 518 6787
rect 552 6753 562 6787
rect 308 6613 318 6647
rect 352 6613 362 6647
rect 108 6473 118 6507
rect 152 6473 162 6507
rect 8 6367 62 6379
rect 8 6341 18 6367
rect 52 6341 62 6367
rect 8 6289 9 6341
rect 61 6289 62 6341
rect 8 6282 62 6289
rect 108 6367 162 6473
rect 208 6551 262 6558
rect 208 6499 209 6551
rect 261 6499 262 6551
rect 208 6473 218 6499
rect 252 6473 262 6499
rect 208 6461 262 6473
rect 308 6507 362 6613
rect 408 6647 462 6659
rect 408 6621 418 6647
rect 452 6621 462 6647
rect 408 6569 409 6621
rect 461 6569 462 6621
rect 408 6562 462 6569
rect 508 6647 562 6753
rect 608 6831 662 6838
rect 608 6779 609 6831
rect 661 6779 662 6831
rect 608 6753 618 6779
rect 652 6753 662 6779
rect 608 6741 662 6753
rect 708 6787 762 6893
rect 808 6927 862 6939
rect 808 6901 818 6927
rect 852 6901 862 6927
rect 808 6849 809 6901
rect 861 6849 862 6901
rect 808 6842 862 6849
rect 908 6927 962 7033
rect 1008 7111 1062 7118
rect 1008 7059 1009 7111
rect 1061 7059 1062 7111
rect 1008 7033 1018 7059
rect 1052 7033 1062 7059
rect 1008 7021 1062 7033
rect 1108 7067 1162 7173
rect 1208 7207 1262 7219
rect 1208 7181 1218 7207
rect 1252 7181 1262 7207
rect 1208 7129 1209 7181
rect 1261 7129 1262 7181
rect 1208 7122 1262 7129
rect 1308 7207 1362 7313
rect 1408 7391 1462 7398
rect 1408 7339 1409 7391
rect 1461 7339 1462 7391
rect 1408 7313 1418 7339
rect 1452 7313 1462 7339
rect 1408 7301 1462 7313
rect 1508 7347 1562 7543
rect 1608 7577 1662 7589
rect 1608 7551 1618 7577
rect 1652 7551 1662 7577
rect 1608 7499 1609 7551
rect 1661 7499 1662 7551
rect 1608 7492 1662 7499
rect 1708 7577 1762 7683
rect 1808 7761 1862 7768
rect 1808 7709 1809 7761
rect 1861 7709 1862 7761
rect 1808 7683 1818 7709
rect 1852 7683 1862 7709
rect 1808 7671 1862 7683
rect 1908 7717 1962 7823
rect 2008 7857 2062 7869
rect 2008 7831 2018 7857
rect 2052 7831 2062 7857
rect 2008 7779 2009 7831
rect 2061 7779 2062 7831
rect 2008 7772 2062 7779
rect 2108 7857 2162 7963
rect 2208 8041 2262 8048
rect 2208 7989 2209 8041
rect 2261 7989 2262 8041
rect 2208 7963 2218 7989
rect 2252 7963 2262 7989
rect 2208 7951 2262 7963
rect 2308 7997 2362 8103
rect 2408 8137 2462 8149
rect 2408 8111 2418 8137
rect 2452 8111 2462 8137
rect 2408 8059 2409 8111
rect 2461 8059 2462 8111
rect 2408 8052 2462 8059
rect 2508 8137 2562 8243
rect 2608 8321 2662 8328
rect 2608 8269 2609 8321
rect 2661 8269 2662 8321
rect 2608 8243 2618 8269
rect 2652 8243 2662 8269
rect 2608 8231 2662 8243
rect 2708 8277 2762 8383
rect 2808 8417 2862 8429
rect 2808 8391 2818 8417
rect 2852 8391 2862 8417
rect 2808 8339 2809 8391
rect 2861 8339 2862 8391
rect 2808 8332 2862 8339
rect 2908 8417 2962 8523
rect 3008 8601 3062 8608
rect 3008 8549 3009 8601
rect 3061 8549 3062 8601
rect 3008 8523 3018 8549
rect 3052 8523 3062 8549
rect 3008 8511 3062 8523
rect 3108 8557 3162 8753
rect 3208 8787 3262 8799
rect 3208 8761 3218 8787
rect 3252 8761 3262 8787
rect 3208 8709 3209 8761
rect 3261 8709 3262 8761
rect 3208 8702 3262 8709
rect 3308 8787 3362 8893
rect 3408 8971 3462 8978
rect 3408 8919 3409 8971
rect 3461 8919 3462 8971
rect 3408 8893 3418 8919
rect 3452 8893 3462 8919
rect 3408 8881 3462 8893
rect 3508 8927 3562 9033
rect 3608 9067 3662 9079
rect 3608 9041 3618 9067
rect 3652 9041 3662 9067
rect 3608 8989 3609 9041
rect 3661 8989 3662 9041
rect 3608 8982 3662 8989
rect 3708 9067 3762 9173
rect 3808 9251 3862 9258
rect 3808 9199 3809 9251
rect 3861 9199 3862 9251
rect 3808 9173 3818 9199
rect 3852 9173 3862 9199
rect 3808 9161 3862 9173
rect 3908 9207 3962 9313
rect 4008 9347 4062 9359
rect 4008 9321 4018 9347
rect 4052 9321 4062 9347
rect 4008 9269 4009 9321
rect 4061 9269 4062 9321
rect 4008 9262 4062 9269
rect 4108 9347 4162 9453
rect 4208 9531 4262 9538
rect 4208 9479 4209 9531
rect 4261 9479 4262 9531
rect 4208 9453 4218 9479
rect 4252 9453 4262 9479
rect 4208 9441 4262 9453
rect 4308 9487 4362 9593
rect 4408 9627 4462 9639
rect 4408 9601 4418 9627
rect 4452 9601 4462 9627
rect 4408 9549 4409 9601
rect 4461 9549 4462 9601
rect 4408 9542 4462 9549
rect 4508 9627 4562 9733
rect 4608 9811 4662 9818
rect 4608 9759 4609 9811
rect 4661 9759 4662 9811
rect 4608 9733 4618 9759
rect 4652 9733 4662 9759
rect 4608 9721 4662 9733
rect 4708 9767 4762 9940
rect 4802 9883 4868 9884
rect 4802 9831 4809 9883
rect 4861 9831 4868 9883
rect 4802 9830 4868 9831
rect 4708 9733 4718 9767
rect 4752 9733 4762 9767
rect 4508 9593 4518 9627
rect 4552 9593 4562 9627
rect 4308 9453 4318 9487
rect 4352 9453 4362 9487
rect 4108 9313 4118 9347
rect 4152 9313 4162 9347
rect 3908 9173 3918 9207
rect 3952 9173 3962 9207
rect 3708 9033 3718 9067
rect 3752 9033 3762 9067
rect 3508 8893 3518 8927
rect 3552 8893 3562 8927
rect 3308 8753 3318 8787
rect 3352 8753 3362 8787
rect 3202 8673 3268 8674
rect 3202 8621 3209 8673
rect 3261 8621 3268 8673
rect 3202 8620 3268 8621
rect 3108 8523 3118 8557
rect 3152 8523 3162 8557
rect 2908 8383 2918 8417
rect 2952 8383 2962 8417
rect 2708 8243 2718 8277
rect 2752 8243 2762 8277
rect 2508 8103 2518 8137
rect 2552 8103 2562 8137
rect 2308 7963 2318 7997
rect 2352 7963 2362 7997
rect 2108 7823 2118 7857
rect 2152 7823 2162 7857
rect 1908 7683 1918 7717
rect 1952 7683 1962 7717
rect 1708 7543 1718 7577
rect 1752 7543 1762 7577
rect 1602 7463 1668 7464
rect 1602 7411 1609 7463
rect 1661 7411 1668 7463
rect 1602 7410 1668 7411
rect 1508 7313 1518 7347
rect 1552 7313 1562 7347
rect 1308 7173 1318 7207
rect 1352 7173 1362 7207
rect 1108 7033 1118 7067
rect 1152 7033 1162 7067
rect 908 6893 918 6927
rect 952 6893 962 6927
rect 708 6753 718 6787
rect 752 6753 762 6787
rect 508 6613 518 6647
rect 552 6613 562 6647
rect 308 6473 318 6507
rect 352 6473 362 6507
rect 108 6333 118 6367
rect 152 6333 162 6367
rect 2 6253 68 6254
rect 2 6201 9 6253
rect 61 6201 68 6253
rect 2 6200 68 6201
rect 8 6137 62 6149
rect 8 6111 18 6137
rect 52 6111 62 6137
rect 8 6059 9 6111
rect 61 6059 62 6111
rect 8 6052 62 6059
rect 108 6137 162 6333
rect 208 6411 262 6418
rect 208 6359 209 6411
rect 261 6359 262 6411
rect 208 6333 218 6359
rect 252 6333 262 6359
rect 208 6321 262 6333
rect 308 6367 362 6473
rect 408 6507 462 6519
rect 408 6481 418 6507
rect 452 6481 462 6507
rect 408 6429 409 6481
rect 461 6429 462 6481
rect 408 6422 462 6429
rect 508 6507 562 6613
rect 608 6691 662 6698
rect 608 6639 609 6691
rect 661 6639 662 6691
rect 608 6613 618 6639
rect 652 6613 662 6639
rect 608 6601 662 6613
rect 708 6647 762 6753
rect 808 6787 862 6799
rect 808 6761 818 6787
rect 852 6761 862 6787
rect 808 6709 809 6761
rect 861 6709 862 6761
rect 808 6702 862 6709
rect 908 6787 962 6893
rect 1008 6971 1062 6978
rect 1008 6919 1009 6971
rect 1061 6919 1062 6971
rect 1008 6893 1018 6919
rect 1052 6893 1062 6919
rect 1008 6881 1062 6893
rect 1108 6927 1162 7033
rect 1208 7067 1262 7079
rect 1208 7041 1218 7067
rect 1252 7041 1262 7067
rect 1208 6989 1209 7041
rect 1261 6989 1262 7041
rect 1208 6982 1262 6989
rect 1308 7067 1362 7173
rect 1408 7251 1462 7258
rect 1408 7199 1409 7251
rect 1461 7199 1462 7251
rect 1408 7173 1418 7199
rect 1452 7173 1462 7199
rect 1408 7161 1462 7173
rect 1508 7207 1562 7313
rect 1608 7347 1662 7359
rect 1608 7321 1618 7347
rect 1652 7321 1662 7347
rect 1608 7269 1609 7321
rect 1661 7269 1662 7321
rect 1608 7262 1662 7269
rect 1708 7347 1762 7543
rect 1808 7621 1862 7628
rect 1808 7569 1809 7621
rect 1861 7569 1862 7621
rect 1808 7543 1818 7569
rect 1852 7543 1862 7569
rect 1808 7531 1862 7543
rect 1908 7577 1962 7683
rect 2008 7717 2062 7729
rect 2008 7691 2018 7717
rect 2052 7691 2062 7717
rect 2008 7639 2009 7691
rect 2061 7639 2062 7691
rect 2008 7632 2062 7639
rect 2108 7717 2162 7823
rect 2208 7901 2262 7908
rect 2208 7849 2209 7901
rect 2261 7849 2262 7901
rect 2208 7823 2218 7849
rect 2252 7823 2262 7849
rect 2208 7811 2262 7823
rect 2308 7857 2362 7963
rect 2408 7997 2462 8009
rect 2408 7971 2418 7997
rect 2452 7971 2462 7997
rect 2408 7919 2409 7971
rect 2461 7919 2462 7971
rect 2408 7912 2462 7919
rect 2508 7997 2562 8103
rect 2608 8181 2662 8188
rect 2608 8129 2609 8181
rect 2661 8129 2662 8181
rect 2608 8103 2618 8129
rect 2652 8103 2662 8129
rect 2608 8091 2662 8103
rect 2708 8137 2762 8243
rect 2808 8277 2862 8289
rect 2808 8251 2818 8277
rect 2852 8251 2862 8277
rect 2808 8199 2809 8251
rect 2861 8199 2862 8251
rect 2808 8192 2862 8199
rect 2908 8277 2962 8383
rect 3008 8461 3062 8468
rect 3008 8409 3009 8461
rect 3061 8409 3062 8461
rect 3008 8383 3018 8409
rect 3052 8383 3062 8409
rect 3008 8371 3062 8383
rect 3108 8417 3162 8523
rect 3208 8557 3262 8569
rect 3208 8531 3218 8557
rect 3252 8531 3262 8557
rect 3208 8479 3209 8531
rect 3261 8479 3262 8531
rect 3208 8472 3262 8479
rect 3308 8557 3362 8753
rect 3408 8831 3462 8838
rect 3408 8779 3409 8831
rect 3461 8779 3462 8831
rect 3408 8753 3418 8779
rect 3452 8753 3462 8779
rect 3408 8741 3462 8753
rect 3508 8787 3562 8893
rect 3608 8927 3662 8939
rect 3608 8901 3618 8927
rect 3652 8901 3662 8927
rect 3608 8849 3609 8901
rect 3661 8849 3662 8901
rect 3608 8842 3662 8849
rect 3708 8927 3762 9033
rect 3808 9111 3862 9118
rect 3808 9059 3809 9111
rect 3861 9059 3862 9111
rect 3808 9033 3818 9059
rect 3852 9033 3862 9059
rect 3808 9021 3862 9033
rect 3908 9067 3962 9173
rect 4008 9207 4062 9219
rect 4008 9181 4018 9207
rect 4052 9181 4062 9207
rect 4008 9129 4009 9181
rect 4061 9129 4062 9181
rect 4008 9122 4062 9129
rect 4108 9207 4162 9313
rect 4208 9391 4262 9398
rect 4208 9339 4209 9391
rect 4261 9339 4262 9391
rect 4208 9313 4218 9339
rect 4252 9313 4262 9339
rect 4208 9301 4262 9313
rect 4308 9347 4362 9453
rect 4408 9487 4462 9499
rect 4408 9461 4418 9487
rect 4452 9461 4462 9487
rect 4408 9409 4409 9461
rect 4461 9409 4462 9461
rect 4408 9402 4462 9409
rect 4508 9487 4562 9593
rect 4608 9671 4662 9678
rect 4608 9619 4609 9671
rect 4661 9619 4662 9671
rect 4608 9593 4618 9619
rect 4652 9593 4662 9619
rect 4608 9581 4662 9593
rect 4708 9627 4762 9733
rect 4808 9767 4862 9779
rect 4808 9741 4818 9767
rect 4852 9741 4862 9767
rect 4808 9689 4809 9741
rect 4861 9689 4862 9741
rect 4808 9682 4862 9689
rect 4908 9767 4962 9940
rect 5002 9899 5068 9900
rect 5002 9847 5009 9899
rect 5061 9847 5068 9899
rect 5002 9846 5068 9847
rect 4908 9733 4918 9767
rect 4952 9733 4962 9767
rect 4708 9593 4718 9627
rect 4752 9593 4762 9627
rect 4508 9453 4518 9487
rect 4552 9453 4562 9487
rect 4308 9313 4318 9347
rect 4352 9313 4362 9347
rect 4108 9173 4118 9207
rect 4152 9173 4162 9207
rect 3908 9033 3918 9067
rect 3952 9033 3962 9067
rect 3708 8893 3718 8927
rect 3752 8893 3762 8927
rect 3508 8753 3518 8787
rect 3552 8753 3562 8787
rect 3402 8689 3468 8690
rect 3402 8637 3409 8689
rect 3461 8637 3468 8689
rect 3402 8636 3468 8637
rect 3308 8523 3318 8557
rect 3352 8523 3362 8557
rect 3108 8383 3118 8417
rect 3152 8383 3162 8417
rect 2908 8243 2918 8277
rect 2952 8243 2962 8277
rect 2708 8103 2718 8137
rect 2752 8103 2762 8137
rect 2508 7963 2518 7997
rect 2552 7963 2562 7997
rect 2308 7823 2318 7857
rect 2352 7823 2362 7857
rect 2108 7683 2118 7717
rect 2152 7683 2162 7717
rect 1908 7543 1918 7577
rect 1952 7543 1962 7577
rect 1802 7479 1868 7480
rect 1802 7427 1809 7479
rect 1861 7427 1868 7479
rect 1802 7426 1868 7427
rect 1708 7313 1718 7347
rect 1752 7313 1762 7347
rect 1508 7173 1518 7207
rect 1552 7173 1562 7207
rect 1308 7033 1318 7067
rect 1352 7033 1362 7067
rect 1108 6893 1118 6927
rect 1152 6893 1162 6927
rect 908 6753 918 6787
rect 952 6753 962 6787
rect 708 6613 718 6647
rect 752 6613 762 6647
rect 508 6473 518 6507
rect 552 6473 562 6507
rect 308 6333 318 6367
rect 352 6333 362 6367
rect 202 6269 268 6270
rect 202 6217 209 6269
rect 261 6217 268 6269
rect 202 6216 268 6217
rect 108 6103 118 6137
rect 152 6103 162 6137
rect 8 5997 62 6009
rect 8 5971 18 5997
rect 52 5971 62 5997
rect 8 5919 9 5971
rect 61 5919 62 5971
rect 8 5912 62 5919
rect 108 5997 162 6103
rect 208 6181 262 6188
rect 208 6129 209 6181
rect 261 6129 262 6181
rect 208 6103 218 6129
rect 252 6103 262 6129
rect 208 6091 262 6103
rect 308 6137 362 6333
rect 408 6367 462 6379
rect 408 6341 418 6367
rect 452 6341 462 6367
rect 408 6289 409 6341
rect 461 6289 462 6341
rect 408 6282 462 6289
rect 508 6367 562 6473
rect 608 6551 662 6558
rect 608 6499 609 6551
rect 661 6499 662 6551
rect 608 6473 618 6499
rect 652 6473 662 6499
rect 608 6461 662 6473
rect 708 6507 762 6613
rect 808 6647 862 6659
rect 808 6621 818 6647
rect 852 6621 862 6647
rect 808 6569 809 6621
rect 861 6569 862 6621
rect 808 6562 862 6569
rect 908 6647 962 6753
rect 1008 6831 1062 6838
rect 1008 6779 1009 6831
rect 1061 6779 1062 6831
rect 1008 6753 1018 6779
rect 1052 6753 1062 6779
rect 1008 6741 1062 6753
rect 1108 6787 1162 6893
rect 1208 6927 1262 6939
rect 1208 6901 1218 6927
rect 1252 6901 1262 6927
rect 1208 6849 1209 6901
rect 1261 6849 1262 6901
rect 1208 6842 1262 6849
rect 1308 6927 1362 7033
rect 1408 7111 1462 7118
rect 1408 7059 1409 7111
rect 1461 7059 1462 7111
rect 1408 7033 1418 7059
rect 1452 7033 1462 7059
rect 1408 7021 1462 7033
rect 1508 7067 1562 7173
rect 1608 7207 1662 7219
rect 1608 7181 1618 7207
rect 1652 7181 1662 7207
rect 1608 7129 1609 7181
rect 1661 7129 1662 7181
rect 1608 7122 1662 7129
rect 1708 7207 1762 7313
rect 1808 7391 1862 7398
rect 1808 7339 1809 7391
rect 1861 7339 1862 7391
rect 1808 7313 1818 7339
rect 1852 7313 1862 7339
rect 1808 7301 1862 7313
rect 1908 7347 1962 7543
rect 2008 7577 2062 7589
rect 2008 7551 2018 7577
rect 2052 7551 2062 7577
rect 2008 7499 2009 7551
rect 2061 7499 2062 7551
rect 2008 7492 2062 7499
rect 2108 7577 2162 7683
rect 2208 7761 2262 7768
rect 2208 7709 2209 7761
rect 2261 7709 2262 7761
rect 2208 7683 2218 7709
rect 2252 7683 2262 7709
rect 2208 7671 2262 7683
rect 2308 7717 2362 7823
rect 2408 7857 2462 7869
rect 2408 7831 2418 7857
rect 2452 7831 2462 7857
rect 2408 7779 2409 7831
rect 2461 7779 2462 7831
rect 2408 7772 2462 7779
rect 2508 7857 2562 7963
rect 2608 8041 2662 8048
rect 2608 7989 2609 8041
rect 2661 7989 2662 8041
rect 2608 7963 2618 7989
rect 2652 7963 2662 7989
rect 2608 7951 2662 7963
rect 2708 7997 2762 8103
rect 2808 8137 2862 8149
rect 2808 8111 2818 8137
rect 2852 8111 2862 8137
rect 2808 8059 2809 8111
rect 2861 8059 2862 8111
rect 2808 8052 2862 8059
rect 2908 8137 2962 8243
rect 3008 8321 3062 8328
rect 3008 8269 3009 8321
rect 3061 8269 3062 8321
rect 3008 8243 3018 8269
rect 3052 8243 3062 8269
rect 3008 8231 3062 8243
rect 3108 8277 3162 8383
rect 3208 8417 3262 8429
rect 3208 8391 3218 8417
rect 3252 8391 3262 8417
rect 3208 8339 3209 8391
rect 3261 8339 3262 8391
rect 3208 8332 3262 8339
rect 3308 8417 3362 8523
rect 3408 8601 3462 8608
rect 3408 8549 3409 8601
rect 3461 8549 3462 8601
rect 3408 8523 3418 8549
rect 3452 8523 3462 8549
rect 3408 8511 3462 8523
rect 3508 8557 3562 8753
rect 3608 8787 3662 8799
rect 3608 8761 3618 8787
rect 3652 8761 3662 8787
rect 3608 8709 3609 8761
rect 3661 8709 3662 8761
rect 3608 8702 3662 8709
rect 3708 8787 3762 8893
rect 3808 8971 3862 8978
rect 3808 8919 3809 8971
rect 3861 8919 3862 8971
rect 3808 8893 3818 8919
rect 3852 8893 3862 8919
rect 3808 8881 3862 8893
rect 3908 8927 3962 9033
rect 4008 9067 4062 9079
rect 4008 9041 4018 9067
rect 4052 9041 4062 9067
rect 4008 8989 4009 9041
rect 4061 8989 4062 9041
rect 4008 8982 4062 8989
rect 4108 9067 4162 9173
rect 4208 9251 4262 9258
rect 4208 9199 4209 9251
rect 4261 9199 4262 9251
rect 4208 9173 4218 9199
rect 4252 9173 4262 9199
rect 4208 9161 4262 9173
rect 4308 9207 4362 9313
rect 4408 9347 4462 9359
rect 4408 9321 4418 9347
rect 4452 9321 4462 9347
rect 4408 9269 4409 9321
rect 4461 9269 4462 9321
rect 4408 9262 4462 9269
rect 4508 9347 4562 9453
rect 4608 9531 4662 9538
rect 4608 9479 4609 9531
rect 4661 9479 4662 9531
rect 4608 9453 4618 9479
rect 4652 9453 4662 9479
rect 4608 9441 4662 9453
rect 4708 9487 4762 9593
rect 4808 9627 4862 9639
rect 4808 9601 4818 9627
rect 4852 9601 4862 9627
rect 4808 9549 4809 9601
rect 4861 9549 4862 9601
rect 4808 9542 4862 9549
rect 4908 9627 4962 9733
rect 5008 9811 5062 9818
rect 5008 9759 5009 9811
rect 5061 9759 5062 9811
rect 5008 9733 5018 9759
rect 5052 9733 5062 9759
rect 5008 9721 5062 9733
rect 5108 9767 5162 9940
rect 5202 9883 5268 9884
rect 5202 9831 5209 9883
rect 5261 9831 5268 9883
rect 5202 9830 5268 9831
rect 5108 9733 5118 9767
rect 5152 9733 5162 9767
rect 4908 9593 4918 9627
rect 4952 9593 4962 9627
rect 4708 9453 4718 9487
rect 4752 9453 4762 9487
rect 4508 9313 4518 9347
rect 4552 9313 4562 9347
rect 4308 9173 4318 9207
rect 4352 9173 4362 9207
rect 4108 9033 4118 9067
rect 4152 9033 4162 9067
rect 3908 8893 3918 8927
rect 3952 8893 3962 8927
rect 3708 8753 3718 8787
rect 3752 8753 3762 8787
rect 3602 8673 3668 8674
rect 3602 8621 3609 8673
rect 3661 8621 3668 8673
rect 3602 8620 3668 8621
rect 3508 8523 3518 8557
rect 3552 8523 3562 8557
rect 3308 8383 3318 8417
rect 3352 8383 3362 8417
rect 3108 8243 3118 8277
rect 3152 8243 3162 8277
rect 2908 8103 2918 8137
rect 2952 8103 2962 8137
rect 2708 7963 2718 7997
rect 2752 7963 2762 7997
rect 2508 7823 2518 7857
rect 2552 7823 2562 7857
rect 2308 7683 2318 7717
rect 2352 7683 2362 7717
rect 2108 7543 2118 7577
rect 2152 7543 2162 7577
rect 2002 7463 2068 7464
rect 2002 7411 2009 7463
rect 2061 7411 2068 7463
rect 2002 7410 2068 7411
rect 1908 7313 1918 7347
rect 1952 7313 1962 7347
rect 1708 7173 1718 7207
rect 1752 7173 1762 7207
rect 1508 7033 1518 7067
rect 1552 7033 1562 7067
rect 1308 6893 1318 6927
rect 1352 6893 1362 6927
rect 1108 6753 1118 6787
rect 1152 6753 1162 6787
rect 908 6613 918 6647
rect 952 6613 962 6647
rect 708 6473 718 6507
rect 752 6473 762 6507
rect 508 6333 518 6367
rect 552 6333 562 6367
rect 402 6253 468 6254
rect 402 6201 409 6253
rect 461 6201 468 6253
rect 402 6200 468 6201
rect 308 6103 318 6137
rect 352 6103 362 6137
rect 108 5963 118 5997
rect 152 5963 162 5997
rect 8 5857 62 5869
rect 8 5831 18 5857
rect 52 5831 62 5857
rect 8 5779 9 5831
rect 61 5779 62 5831
rect 8 5772 62 5779
rect 108 5857 162 5963
rect 208 6041 262 6048
rect 208 5989 209 6041
rect 261 5989 262 6041
rect 208 5963 218 5989
rect 252 5963 262 5989
rect 208 5951 262 5963
rect 308 5997 362 6103
rect 408 6137 462 6149
rect 408 6111 418 6137
rect 452 6111 462 6137
rect 408 6059 409 6111
rect 461 6059 462 6111
rect 408 6052 462 6059
rect 508 6137 562 6333
rect 608 6411 662 6418
rect 608 6359 609 6411
rect 661 6359 662 6411
rect 608 6333 618 6359
rect 652 6333 662 6359
rect 608 6321 662 6333
rect 708 6367 762 6473
rect 808 6507 862 6519
rect 808 6481 818 6507
rect 852 6481 862 6507
rect 808 6429 809 6481
rect 861 6429 862 6481
rect 808 6422 862 6429
rect 908 6507 962 6613
rect 1008 6691 1062 6698
rect 1008 6639 1009 6691
rect 1061 6639 1062 6691
rect 1008 6613 1018 6639
rect 1052 6613 1062 6639
rect 1008 6601 1062 6613
rect 1108 6647 1162 6753
rect 1208 6787 1262 6799
rect 1208 6761 1218 6787
rect 1252 6761 1262 6787
rect 1208 6709 1209 6761
rect 1261 6709 1262 6761
rect 1208 6702 1262 6709
rect 1308 6787 1362 6893
rect 1408 6971 1462 6978
rect 1408 6919 1409 6971
rect 1461 6919 1462 6971
rect 1408 6893 1418 6919
rect 1452 6893 1462 6919
rect 1408 6881 1462 6893
rect 1508 6927 1562 7033
rect 1608 7067 1662 7079
rect 1608 7041 1618 7067
rect 1652 7041 1662 7067
rect 1608 6989 1609 7041
rect 1661 6989 1662 7041
rect 1608 6982 1662 6989
rect 1708 7067 1762 7173
rect 1808 7251 1862 7258
rect 1808 7199 1809 7251
rect 1861 7199 1862 7251
rect 1808 7173 1818 7199
rect 1852 7173 1862 7199
rect 1808 7161 1862 7173
rect 1908 7207 1962 7313
rect 2008 7347 2062 7359
rect 2008 7321 2018 7347
rect 2052 7321 2062 7347
rect 2008 7269 2009 7321
rect 2061 7269 2062 7321
rect 2008 7262 2062 7269
rect 2108 7347 2162 7543
rect 2208 7621 2262 7628
rect 2208 7569 2209 7621
rect 2261 7569 2262 7621
rect 2208 7543 2218 7569
rect 2252 7543 2262 7569
rect 2208 7531 2262 7543
rect 2308 7577 2362 7683
rect 2408 7717 2462 7729
rect 2408 7691 2418 7717
rect 2452 7691 2462 7717
rect 2408 7639 2409 7691
rect 2461 7639 2462 7691
rect 2408 7632 2462 7639
rect 2508 7717 2562 7823
rect 2608 7901 2662 7908
rect 2608 7849 2609 7901
rect 2661 7849 2662 7901
rect 2608 7823 2618 7849
rect 2652 7823 2662 7849
rect 2608 7811 2662 7823
rect 2708 7857 2762 7963
rect 2808 7997 2862 8009
rect 2808 7971 2818 7997
rect 2852 7971 2862 7997
rect 2808 7919 2809 7971
rect 2861 7919 2862 7971
rect 2808 7912 2862 7919
rect 2908 7997 2962 8103
rect 3008 8181 3062 8188
rect 3008 8129 3009 8181
rect 3061 8129 3062 8181
rect 3008 8103 3018 8129
rect 3052 8103 3062 8129
rect 3008 8091 3062 8103
rect 3108 8137 3162 8243
rect 3208 8277 3262 8289
rect 3208 8251 3218 8277
rect 3252 8251 3262 8277
rect 3208 8199 3209 8251
rect 3261 8199 3262 8251
rect 3208 8192 3262 8199
rect 3308 8277 3362 8383
rect 3408 8461 3462 8468
rect 3408 8409 3409 8461
rect 3461 8409 3462 8461
rect 3408 8383 3418 8409
rect 3452 8383 3462 8409
rect 3408 8371 3462 8383
rect 3508 8417 3562 8523
rect 3608 8557 3662 8569
rect 3608 8531 3618 8557
rect 3652 8531 3662 8557
rect 3608 8479 3609 8531
rect 3661 8479 3662 8531
rect 3608 8472 3662 8479
rect 3708 8557 3762 8753
rect 3808 8831 3862 8838
rect 3808 8779 3809 8831
rect 3861 8779 3862 8831
rect 3808 8753 3818 8779
rect 3852 8753 3862 8779
rect 3808 8741 3862 8753
rect 3908 8787 3962 8893
rect 4008 8927 4062 8939
rect 4008 8901 4018 8927
rect 4052 8901 4062 8927
rect 4008 8849 4009 8901
rect 4061 8849 4062 8901
rect 4008 8842 4062 8849
rect 4108 8927 4162 9033
rect 4208 9111 4262 9118
rect 4208 9059 4209 9111
rect 4261 9059 4262 9111
rect 4208 9033 4218 9059
rect 4252 9033 4262 9059
rect 4208 9021 4262 9033
rect 4308 9067 4362 9173
rect 4408 9207 4462 9219
rect 4408 9181 4418 9207
rect 4452 9181 4462 9207
rect 4408 9129 4409 9181
rect 4461 9129 4462 9181
rect 4408 9122 4462 9129
rect 4508 9207 4562 9313
rect 4608 9391 4662 9398
rect 4608 9339 4609 9391
rect 4661 9339 4662 9391
rect 4608 9313 4618 9339
rect 4652 9313 4662 9339
rect 4608 9301 4662 9313
rect 4708 9347 4762 9453
rect 4808 9487 4862 9499
rect 4808 9461 4818 9487
rect 4852 9461 4862 9487
rect 4808 9409 4809 9461
rect 4861 9409 4862 9461
rect 4808 9402 4862 9409
rect 4908 9487 4962 9593
rect 5008 9671 5062 9678
rect 5008 9619 5009 9671
rect 5061 9619 5062 9671
rect 5008 9593 5018 9619
rect 5052 9593 5062 9619
rect 5008 9581 5062 9593
rect 5108 9627 5162 9733
rect 5208 9767 5262 9779
rect 5208 9741 5218 9767
rect 5252 9741 5262 9767
rect 5208 9689 5209 9741
rect 5261 9689 5262 9741
rect 5208 9682 5262 9689
rect 5308 9767 5362 9940
rect 5402 9899 5468 9900
rect 5402 9847 5409 9899
rect 5461 9847 5468 9899
rect 5402 9846 5468 9847
rect 5308 9733 5318 9767
rect 5352 9733 5362 9767
rect 5108 9593 5118 9627
rect 5152 9593 5162 9627
rect 4908 9453 4918 9487
rect 4952 9453 4962 9487
rect 4708 9313 4718 9347
rect 4752 9313 4762 9347
rect 4508 9173 4518 9207
rect 4552 9173 4562 9207
rect 4308 9033 4318 9067
rect 4352 9033 4362 9067
rect 4108 8893 4118 8927
rect 4152 8893 4162 8927
rect 3908 8753 3918 8787
rect 3952 8753 3962 8787
rect 3802 8689 3868 8690
rect 3802 8637 3809 8689
rect 3861 8637 3868 8689
rect 3802 8636 3868 8637
rect 3708 8523 3718 8557
rect 3752 8523 3762 8557
rect 3508 8383 3518 8417
rect 3552 8383 3562 8417
rect 3308 8243 3318 8277
rect 3352 8243 3362 8277
rect 3108 8103 3118 8137
rect 3152 8103 3162 8137
rect 2908 7963 2918 7997
rect 2952 7963 2962 7997
rect 2708 7823 2718 7857
rect 2752 7823 2762 7857
rect 2508 7683 2518 7717
rect 2552 7683 2562 7717
rect 2308 7543 2318 7577
rect 2352 7543 2362 7577
rect 2202 7479 2268 7480
rect 2202 7427 2209 7479
rect 2261 7427 2268 7479
rect 2202 7426 2268 7427
rect 2108 7313 2118 7347
rect 2152 7313 2162 7347
rect 1908 7173 1918 7207
rect 1952 7173 1962 7207
rect 1708 7033 1718 7067
rect 1752 7033 1762 7067
rect 1508 6893 1518 6927
rect 1552 6893 1562 6927
rect 1308 6753 1318 6787
rect 1352 6753 1362 6787
rect 1108 6613 1118 6647
rect 1152 6613 1162 6647
rect 908 6473 918 6507
rect 952 6473 962 6507
rect 708 6333 718 6367
rect 752 6333 762 6367
rect 602 6269 668 6270
rect 602 6217 609 6269
rect 661 6217 668 6269
rect 602 6216 668 6217
rect 508 6103 518 6137
rect 552 6103 562 6137
rect 308 5963 318 5997
rect 352 5963 362 5997
rect 108 5823 118 5857
rect 152 5823 162 5857
rect 8 5717 62 5729
rect 8 5691 18 5717
rect 52 5691 62 5717
rect 8 5639 9 5691
rect 61 5639 62 5691
rect 8 5632 62 5639
rect 108 5717 162 5823
rect 208 5901 262 5908
rect 208 5849 209 5901
rect 261 5849 262 5901
rect 208 5823 218 5849
rect 252 5823 262 5849
rect 208 5811 262 5823
rect 308 5857 362 5963
rect 408 5997 462 6009
rect 408 5971 418 5997
rect 452 5971 462 5997
rect 408 5919 409 5971
rect 461 5919 462 5971
rect 408 5912 462 5919
rect 508 5997 562 6103
rect 608 6181 662 6188
rect 608 6129 609 6181
rect 661 6129 662 6181
rect 608 6103 618 6129
rect 652 6103 662 6129
rect 608 6091 662 6103
rect 708 6137 762 6333
rect 808 6367 862 6379
rect 808 6341 818 6367
rect 852 6341 862 6367
rect 808 6289 809 6341
rect 861 6289 862 6341
rect 808 6282 862 6289
rect 908 6367 962 6473
rect 1008 6551 1062 6558
rect 1008 6499 1009 6551
rect 1061 6499 1062 6551
rect 1008 6473 1018 6499
rect 1052 6473 1062 6499
rect 1008 6461 1062 6473
rect 1108 6507 1162 6613
rect 1208 6647 1262 6659
rect 1208 6621 1218 6647
rect 1252 6621 1262 6647
rect 1208 6569 1209 6621
rect 1261 6569 1262 6621
rect 1208 6562 1262 6569
rect 1308 6647 1362 6753
rect 1408 6831 1462 6838
rect 1408 6779 1409 6831
rect 1461 6779 1462 6831
rect 1408 6753 1418 6779
rect 1452 6753 1462 6779
rect 1408 6741 1462 6753
rect 1508 6787 1562 6893
rect 1608 6927 1662 6939
rect 1608 6901 1618 6927
rect 1652 6901 1662 6927
rect 1608 6849 1609 6901
rect 1661 6849 1662 6901
rect 1608 6842 1662 6849
rect 1708 6927 1762 7033
rect 1808 7111 1862 7118
rect 1808 7059 1809 7111
rect 1861 7059 1862 7111
rect 1808 7033 1818 7059
rect 1852 7033 1862 7059
rect 1808 7021 1862 7033
rect 1908 7067 1962 7173
rect 2008 7207 2062 7219
rect 2008 7181 2018 7207
rect 2052 7181 2062 7207
rect 2008 7129 2009 7181
rect 2061 7129 2062 7181
rect 2008 7122 2062 7129
rect 2108 7207 2162 7313
rect 2208 7391 2262 7398
rect 2208 7339 2209 7391
rect 2261 7339 2262 7391
rect 2208 7313 2218 7339
rect 2252 7313 2262 7339
rect 2208 7301 2262 7313
rect 2308 7347 2362 7543
rect 2408 7577 2462 7589
rect 2408 7551 2418 7577
rect 2452 7551 2462 7577
rect 2408 7499 2409 7551
rect 2461 7499 2462 7551
rect 2408 7492 2462 7499
rect 2508 7577 2562 7683
rect 2608 7761 2662 7768
rect 2608 7709 2609 7761
rect 2661 7709 2662 7761
rect 2608 7683 2618 7709
rect 2652 7683 2662 7709
rect 2608 7671 2662 7683
rect 2708 7717 2762 7823
rect 2808 7857 2862 7869
rect 2808 7831 2818 7857
rect 2852 7831 2862 7857
rect 2808 7779 2809 7831
rect 2861 7779 2862 7831
rect 2808 7772 2862 7779
rect 2908 7857 2962 7963
rect 3008 8041 3062 8048
rect 3008 7989 3009 8041
rect 3061 7989 3062 8041
rect 3008 7963 3018 7989
rect 3052 7963 3062 7989
rect 3008 7951 3062 7963
rect 3108 7997 3162 8103
rect 3208 8137 3262 8149
rect 3208 8111 3218 8137
rect 3252 8111 3262 8137
rect 3208 8059 3209 8111
rect 3261 8059 3262 8111
rect 3208 8052 3262 8059
rect 3308 8137 3362 8243
rect 3408 8321 3462 8328
rect 3408 8269 3409 8321
rect 3461 8269 3462 8321
rect 3408 8243 3418 8269
rect 3452 8243 3462 8269
rect 3408 8231 3462 8243
rect 3508 8277 3562 8383
rect 3608 8417 3662 8429
rect 3608 8391 3618 8417
rect 3652 8391 3662 8417
rect 3608 8339 3609 8391
rect 3661 8339 3662 8391
rect 3608 8332 3662 8339
rect 3708 8417 3762 8523
rect 3808 8601 3862 8608
rect 3808 8549 3809 8601
rect 3861 8549 3862 8601
rect 3808 8523 3818 8549
rect 3852 8523 3862 8549
rect 3808 8511 3862 8523
rect 3908 8557 3962 8753
rect 4008 8787 4062 8799
rect 4008 8761 4018 8787
rect 4052 8761 4062 8787
rect 4008 8709 4009 8761
rect 4061 8709 4062 8761
rect 4008 8702 4062 8709
rect 4108 8787 4162 8893
rect 4208 8971 4262 8978
rect 4208 8919 4209 8971
rect 4261 8919 4262 8971
rect 4208 8893 4218 8919
rect 4252 8893 4262 8919
rect 4208 8881 4262 8893
rect 4308 8927 4362 9033
rect 4408 9067 4462 9079
rect 4408 9041 4418 9067
rect 4452 9041 4462 9067
rect 4408 8989 4409 9041
rect 4461 8989 4462 9041
rect 4408 8982 4462 8989
rect 4508 9067 4562 9173
rect 4608 9251 4662 9258
rect 4608 9199 4609 9251
rect 4661 9199 4662 9251
rect 4608 9173 4618 9199
rect 4652 9173 4662 9199
rect 4608 9161 4662 9173
rect 4708 9207 4762 9313
rect 4808 9347 4862 9359
rect 4808 9321 4818 9347
rect 4852 9321 4862 9347
rect 4808 9269 4809 9321
rect 4861 9269 4862 9321
rect 4808 9262 4862 9269
rect 4908 9347 4962 9453
rect 5008 9531 5062 9538
rect 5008 9479 5009 9531
rect 5061 9479 5062 9531
rect 5008 9453 5018 9479
rect 5052 9453 5062 9479
rect 5008 9441 5062 9453
rect 5108 9487 5162 9593
rect 5208 9627 5262 9639
rect 5208 9601 5218 9627
rect 5252 9601 5262 9627
rect 5208 9549 5209 9601
rect 5261 9549 5262 9601
rect 5208 9542 5262 9549
rect 5308 9627 5362 9733
rect 5408 9811 5462 9818
rect 5408 9759 5409 9811
rect 5461 9759 5462 9811
rect 5408 9733 5418 9759
rect 5452 9733 5462 9759
rect 5408 9721 5462 9733
rect 5508 9767 5562 9940
rect 5602 9883 5668 9884
rect 5602 9831 5609 9883
rect 5661 9831 5668 9883
rect 5602 9830 5668 9831
rect 5508 9733 5518 9767
rect 5552 9733 5562 9767
rect 5308 9593 5318 9627
rect 5352 9593 5362 9627
rect 5108 9453 5118 9487
rect 5152 9453 5162 9487
rect 4908 9313 4918 9347
rect 4952 9313 4962 9347
rect 4708 9173 4718 9207
rect 4752 9173 4762 9207
rect 4508 9033 4518 9067
rect 4552 9033 4562 9067
rect 4308 8893 4318 8927
rect 4352 8893 4362 8927
rect 4108 8753 4118 8787
rect 4152 8753 4162 8787
rect 4002 8673 4068 8674
rect 4002 8621 4009 8673
rect 4061 8621 4068 8673
rect 4002 8620 4068 8621
rect 3908 8523 3918 8557
rect 3952 8523 3962 8557
rect 3708 8383 3718 8417
rect 3752 8383 3762 8417
rect 3508 8243 3518 8277
rect 3552 8243 3562 8277
rect 3308 8103 3318 8137
rect 3352 8103 3362 8137
rect 3108 7963 3118 7997
rect 3152 7963 3162 7997
rect 2908 7823 2918 7857
rect 2952 7823 2962 7857
rect 2708 7683 2718 7717
rect 2752 7683 2762 7717
rect 2508 7543 2518 7577
rect 2552 7543 2562 7577
rect 2402 7463 2468 7464
rect 2402 7411 2409 7463
rect 2461 7411 2468 7463
rect 2402 7410 2468 7411
rect 2308 7313 2318 7347
rect 2352 7313 2362 7347
rect 2108 7173 2118 7207
rect 2152 7173 2162 7207
rect 1908 7033 1918 7067
rect 1952 7033 1962 7067
rect 1708 6893 1718 6927
rect 1752 6893 1762 6927
rect 1508 6753 1518 6787
rect 1552 6753 1562 6787
rect 1308 6613 1318 6647
rect 1352 6613 1362 6647
rect 1108 6473 1118 6507
rect 1152 6473 1162 6507
rect 908 6333 918 6367
rect 952 6333 962 6367
rect 802 6253 868 6254
rect 802 6201 809 6253
rect 861 6201 868 6253
rect 802 6200 868 6201
rect 708 6103 718 6137
rect 752 6103 762 6137
rect 508 5963 518 5997
rect 552 5963 562 5997
rect 308 5823 318 5857
rect 352 5823 362 5857
rect 108 5683 118 5717
rect 152 5683 162 5717
rect 8 5577 62 5589
rect 8 5551 18 5577
rect 52 5551 62 5577
rect 8 5499 9 5551
rect 61 5499 62 5551
rect 8 5492 62 5499
rect 108 5577 162 5683
rect 208 5761 262 5768
rect 208 5709 209 5761
rect 261 5709 262 5761
rect 208 5683 218 5709
rect 252 5683 262 5709
rect 208 5671 262 5683
rect 308 5717 362 5823
rect 408 5857 462 5869
rect 408 5831 418 5857
rect 452 5831 462 5857
rect 408 5779 409 5831
rect 461 5779 462 5831
rect 408 5772 462 5779
rect 508 5857 562 5963
rect 608 6041 662 6048
rect 608 5989 609 6041
rect 661 5989 662 6041
rect 608 5963 618 5989
rect 652 5963 662 5989
rect 608 5951 662 5963
rect 708 5997 762 6103
rect 808 6137 862 6149
rect 808 6111 818 6137
rect 852 6111 862 6137
rect 808 6059 809 6111
rect 861 6059 862 6111
rect 808 6052 862 6059
rect 908 6137 962 6333
rect 1008 6411 1062 6418
rect 1008 6359 1009 6411
rect 1061 6359 1062 6411
rect 1008 6333 1018 6359
rect 1052 6333 1062 6359
rect 1008 6321 1062 6333
rect 1108 6367 1162 6473
rect 1208 6507 1262 6519
rect 1208 6481 1218 6507
rect 1252 6481 1262 6507
rect 1208 6429 1209 6481
rect 1261 6429 1262 6481
rect 1208 6422 1262 6429
rect 1308 6507 1362 6613
rect 1408 6691 1462 6698
rect 1408 6639 1409 6691
rect 1461 6639 1462 6691
rect 1408 6613 1418 6639
rect 1452 6613 1462 6639
rect 1408 6601 1462 6613
rect 1508 6647 1562 6753
rect 1608 6787 1662 6799
rect 1608 6761 1618 6787
rect 1652 6761 1662 6787
rect 1608 6709 1609 6761
rect 1661 6709 1662 6761
rect 1608 6702 1662 6709
rect 1708 6787 1762 6893
rect 1808 6971 1862 6978
rect 1808 6919 1809 6971
rect 1861 6919 1862 6971
rect 1808 6893 1818 6919
rect 1852 6893 1862 6919
rect 1808 6881 1862 6893
rect 1908 6927 1962 7033
rect 2008 7067 2062 7079
rect 2008 7041 2018 7067
rect 2052 7041 2062 7067
rect 2008 6989 2009 7041
rect 2061 6989 2062 7041
rect 2008 6982 2062 6989
rect 2108 7067 2162 7173
rect 2208 7251 2262 7258
rect 2208 7199 2209 7251
rect 2261 7199 2262 7251
rect 2208 7173 2218 7199
rect 2252 7173 2262 7199
rect 2208 7161 2262 7173
rect 2308 7207 2362 7313
rect 2408 7347 2462 7359
rect 2408 7321 2418 7347
rect 2452 7321 2462 7347
rect 2408 7269 2409 7321
rect 2461 7269 2462 7321
rect 2408 7262 2462 7269
rect 2508 7347 2562 7543
rect 2608 7621 2662 7628
rect 2608 7569 2609 7621
rect 2661 7569 2662 7621
rect 2608 7543 2618 7569
rect 2652 7543 2662 7569
rect 2608 7531 2662 7543
rect 2708 7577 2762 7683
rect 2808 7717 2862 7729
rect 2808 7691 2818 7717
rect 2852 7691 2862 7717
rect 2808 7639 2809 7691
rect 2861 7639 2862 7691
rect 2808 7632 2862 7639
rect 2908 7717 2962 7823
rect 3008 7901 3062 7908
rect 3008 7849 3009 7901
rect 3061 7849 3062 7901
rect 3008 7823 3018 7849
rect 3052 7823 3062 7849
rect 3008 7811 3062 7823
rect 3108 7857 3162 7963
rect 3208 7997 3262 8009
rect 3208 7971 3218 7997
rect 3252 7971 3262 7997
rect 3208 7919 3209 7971
rect 3261 7919 3262 7971
rect 3208 7912 3262 7919
rect 3308 7997 3362 8103
rect 3408 8181 3462 8188
rect 3408 8129 3409 8181
rect 3461 8129 3462 8181
rect 3408 8103 3418 8129
rect 3452 8103 3462 8129
rect 3408 8091 3462 8103
rect 3508 8137 3562 8243
rect 3608 8277 3662 8289
rect 3608 8251 3618 8277
rect 3652 8251 3662 8277
rect 3608 8199 3609 8251
rect 3661 8199 3662 8251
rect 3608 8192 3662 8199
rect 3708 8277 3762 8383
rect 3808 8461 3862 8468
rect 3808 8409 3809 8461
rect 3861 8409 3862 8461
rect 3808 8383 3818 8409
rect 3852 8383 3862 8409
rect 3808 8371 3862 8383
rect 3908 8417 3962 8523
rect 4008 8557 4062 8569
rect 4008 8531 4018 8557
rect 4052 8531 4062 8557
rect 4008 8479 4009 8531
rect 4061 8479 4062 8531
rect 4008 8472 4062 8479
rect 4108 8557 4162 8753
rect 4208 8831 4262 8838
rect 4208 8779 4209 8831
rect 4261 8779 4262 8831
rect 4208 8753 4218 8779
rect 4252 8753 4262 8779
rect 4208 8741 4262 8753
rect 4308 8787 4362 8893
rect 4408 8927 4462 8939
rect 4408 8901 4418 8927
rect 4452 8901 4462 8927
rect 4408 8849 4409 8901
rect 4461 8849 4462 8901
rect 4408 8842 4462 8849
rect 4508 8927 4562 9033
rect 4608 9111 4662 9118
rect 4608 9059 4609 9111
rect 4661 9059 4662 9111
rect 4608 9033 4618 9059
rect 4652 9033 4662 9059
rect 4608 9021 4662 9033
rect 4708 9067 4762 9173
rect 4808 9207 4862 9219
rect 4808 9181 4818 9207
rect 4852 9181 4862 9207
rect 4808 9129 4809 9181
rect 4861 9129 4862 9181
rect 4808 9122 4862 9129
rect 4908 9207 4962 9313
rect 5008 9391 5062 9398
rect 5008 9339 5009 9391
rect 5061 9339 5062 9391
rect 5008 9313 5018 9339
rect 5052 9313 5062 9339
rect 5008 9301 5062 9313
rect 5108 9347 5162 9453
rect 5208 9487 5262 9499
rect 5208 9461 5218 9487
rect 5252 9461 5262 9487
rect 5208 9409 5209 9461
rect 5261 9409 5262 9461
rect 5208 9402 5262 9409
rect 5308 9487 5362 9593
rect 5408 9671 5462 9678
rect 5408 9619 5409 9671
rect 5461 9619 5462 9671
rect 5408 9593 5418 9619
rect 5452 9593 5462 9619
rect 5408 9581 5462 9593
rect 5508 9627 5562 9733
rect 5608 9767 5662 9779
rect 5608 9741 5618 9767
rect 5652 9741 5662 9767
rect 5608 9689 5609 9741
rect 5661 9689 5662 9741
rect 5608 9682 5662 9689
rect 5708 9767 5762 9940
rect 5802 9899 5868 9900
rect 5802 9847 5809 9899
rect 5861 9847 5868 9899
rect 5802 9846 5868 9847
rect 5708 9733 5718 9767
rect 5752 9733 5762 9767
rect 5508 9593 5518 9627
rect 5552 9593 5562 9627
rect 5308 9453 5318 9487
rect 5352 9453 5362 9487
rect 5108 9313 5118 9347
rect 5152 9313 5162 9347
rect 4908 9173 4918 9207
rect 4952 9173 4962 9207
rect 4708 9033 4718 9067
rect 4752 9033 4762 9067
rect 4508 8893 4518 8927
rect 4552 8893 4562 8927
rect 4308 8753 4318 8787
rect 4352 8753 4362 8787
rect 4202 8689 4268 8690
rect 4202 8637 4209 8689
rect 4261 8637 4268 8689
rect 4202 8636 4268 8637
rect 4108 8523 4118 8557
rect 4152 8523 4162 8557
rect 3908 8383 3918 8417
rect 3952 8383 3962 8417
rect 3708 8243 3718 8277
rect 3752 8243 3762 8277
rect 3508 8103 3518 8137
rect 3552 8103 3562 8137
rect 3308 7963 3318 7997
rect 3352 7963 3362 7997
rect 3108 7823 3118 7857
rect 3152 7823 3162 7857
rect 2908 7683 2918 7717
rect 2952 7683 2962 7717
rect 2708 7543 2718 7577
rect 2752 7543 2762 7577
rect 2602 7479 2668 7480
rect 2602 7427 2609 7479
rect 2661 7427 2668 7479
rect 2602 7426 2668 7427
rect 2508 7313 2518 7347
rect 2552 7313 2562 7347
rect 2308 7173 2318 7207
rect 2352 7173 2362 7207
rect 2108 7033 2118 7067
rect 2152 7033 2162 7067
rect 1908 6893 1918 6927
rect 1952 6893 1962 6927
rect 1708 6753 1718 6787
rect 1752 6753 1762 6787
rect 1508 6613 1518 6647
rect 1552 6613 1562 6647
rect 1308 6473 1318 6507
rect 1352 6473 1362 6507
rect 1108 6333 1118 6367
rect 1152 6333 1162 6367
rect 1002 6269 1068 6270
rect 1002 6217 1009 6269
rect 1061 6217 1068 6269
rect 1002 6216 1068 6217
rect 908 6103 918 6137
rect 952 6103 962 6137
rect 708 5963 718 5997
rect 752 5963 762 5997
rect 508 5823 518 5857
rect 552 5823 562 5857
rect 308 5683 318 5717
rect 352 5683 362 5717
rect 108 5543 118 5577
rect 152 5543 162 5577
rect 8 5437 62 5449
rect 8 5411 18 5437
rect 52 5411 62 5437
rect 8 5359 9 5411
rect 61 5359 62 5411
rect 8 5352 62 5359
rect 108 5437 162 5543
rect 208 5621 262 5628
rect 208 5569 209 5621
rect 261 5569 262 5621
rect 208 5543 218 5569
rect 252 5543 262 5569
rect 208 5531 262 5543
rect 308 5577 362 5683
rect 408 5717 462 5729
rect 408 5691 418 5717
rect 452 5691 462 5717
rect 408 5639 409 5691
rect 461 5639 462 5691
rect 408 5632 462 5639
rect 508 5717 562 5823
rect 608 5901 662 5908
rect 608 5849 609 5901
rect 661 5849 662 5901
rect 608 5823 618 5849
rect 652 5823 662 5849
rect 608 5811 662 5823
rect 708 5857 762 5963
rect 808 5997 862 6009
rect 808 5971 818 5997
rect 852 5971 862 5997
rect 808 5919 809 5971
rect 861 5919 862 5971
rect 808 5912 862 5919
rect 908 5997 962 6103
rect 1008 6181 1062 6188
rect 1008 6129 1009 6181
rect 1061 6129 1062 6181
rect 1008 6103 1018 6129
rect 1052 6103 1062 6129
rect 1008 6091 1062 6103
rect 1108 6137 1162 6333
rect 1208 6367 1262 6379
rect 1208 6341 1218 6367
rect 1252 6341 1262 6367
rect 1208 6289 1209 6341
rect 1261 6289 1262 6341
rect 1208 6282 1262 6289
rect 1308 6367 1362 6473
rect 1408 6551 1462 6558
rect 1408 6499 1409 6551
rect 1461 6499 1462 6551
rect 1408 6473 1418 6499
rect 1452 6473 1462 6499
rect 1408 6461 1462 6473
rect 1508 6507 1562 6613
rect 1608 6647 1662 6659
rect 1608 6621 1618 6647
rect 1652 6621 1662 6647
rect 1608 6569 1609 6621
rect 1661 6569 1662 6621
rect 1608 6562 1662 6569
rect 1708 6647 1762 6753
rect 1808 6831 1862 6838
rect 1808 6779 1809 6831
rect 1861 6779 1862 6831
rect 1808 6753 1818 6779
rect 1852 6753 1862 6779
rect 1808 6741 1862 6753
rect 1908 6787 1962 6893
rect 2008 6927 2062 6939
rect 2008 6901 2018 6927
rect 2052 6901 2062 6927
rect 2008 6849 2009 6901
rect 2061 6849 2062 6901
rect 2008 6842 2062 6849
rect 2108 6927 2162 7033
rect 2208 7111 2262 7118
rect 2208 7059 2209 7111
rect 2261 7059 2262 7111
rect 2208 7033 2218 7059
rect 2252 7033 2262 7059
rect 2208 7021 2262 7033
rect 2308 7067 2362 7173
rect 2408 7207 2462 7219
rect 2408 7181 2418 7207
rect 2452 7181 2462 7207
rect 2408 7129 2409 7181
rect 2461 7129 2462 7181
rect 2408 7122 2462 7129
rect 2508 7207 2562 7313
rect 2608 7391 2662 7398
rect 2608 7339 2609 7391
rect 2661 7339 2662 7391
rect 2608 7313 2618 7339
rect 2652 7313 2662 7339
rect 2608 7301 2662 7313
rect 2708 7347 2762 7543
rect 2808 7577 2862 7589
rect 2808 7551 2818 7577
rect 2852 7551 2862 7577
rect 2808 7499 2809 7551
rect 2861 7499 2862 7551
rect 2808 7492 2862 7499
rect 2908 7577 2962 7683
rect 3008 7761 3062 7768
rect 3008 7709 3009 7761
rect 3061 7709 3062 7761
rect 3008 7683 3018 7709
rect 3052 7683 3062 7709
rect 3008 7671 3062 7683
rect 3108 7717 3162 7823
rect 3208 7857 3262 7869
rect 3208 7831 3218 7857
rect 3252 7831 3262 7857
rect 3208 7779 3209 7831
rect 3261 7779 3262 7831
rect 3208 7772 3262 7779
rect 3308 7857 3362 7963
rect 3408 8041 3462 8048
rect 3408 7989 3409 8041
rect 3461 7989 3462 8041
rect 3408 7963 3418 7989
rect 3452 7963 3462 7989
rect 3408 7951 3462 7963
rect 3508 7997 3562 8103
rect 3608 8137 3662 8149
rect 3608 8111 3618 8137
rect 3652 8111 3662 8137
rect 3608 8059 3609 8111
rect 3661 8059 3662 8111
rect 3608 8052 3662 8059
rect 3708 8137 3762 8243
rect 3808 8321 3862 8328
rect 3808 8269 3809 8321
rect 3861 8269 3862 8321
rect 3808 8243 3818 8269
rect 3852 8243 3862 8269
rect 3808 8231 3862 8243
rect 3908 8277 3962 8383
rect 4008 8417 4062 8429
rect 4008 8391 4018 8417
rect 4052 8391 4062 8417
rect 4008 8339 4009 8391
rect 4061 8339 4062 8391
rect 4008 8332 4062 8339
rect 4108 8417 4162 8523
rect 4208 8601 4262 8608
rect 4208 8549 4209 8601
rect 4261 8549 4262 8601
rect 4208 8523 4218 8549
rect 4252 8523 4262 8549
rect 4208 8511 4262 8523
rect 4308 8557 4362 8753
rect 4408 8787 4462 8799
rect 4408 8761 4418 8787
rect 4452 8761 4462 8787
rect 4408 8709 4409 8761
rect 4461 8709 4462 8761
rect 4408 8702 4462 8709
rect 4508 8787 4562 8893
rect 4608 8971 4662 8978
rect 4608 8919 4609 8971
rect 4661 8919 4662 8971
rect 4608 8893 4618 8919
rect 4652 8893 4662 8919
rect 4608 8881 4662 8893
rect 4708 8927 4762 9033
rect 4808 9067 4862 9079
rect 4808 9041 4818 9067
rect 4852 9041 4862 9067
rect 4808 8989 4809 9041
rect 4861 8989 4862 9041
rect 4808 8982 4862 8989
rect 4908 9067 4962 9173
rect 5008 9251 5062 9258
rect 5008 9199 5009 9251
rect 5061 9199 5062 9251
rect 5008 9173 5018 9199
rect 5052 9173 5062 9199
rect 5008 9161 5062 9173
rect 5108 9207 5162 9313
rect 5208 9347 5262 9359
rect 5208 9321 5218 9347
rect 5252 9321 5262 9347
rect 5208 9269 5209 9321
rect 5261 9269 5262 9321
rect 5208 9262 5262 9269
rect 5308 9347 5362 9453
rect 5408 9531 5462 9538
rect 5408 9479 5409 9531
rect 5461 9479 5462 9531
rect 5408 9453 5418 9479
rect 5452 9453 5462 9479
rect 5408 9441 5462 9453
rect 5508 9487 5562 9593
rect 5608 9627 5662 9639
rect 5608 9601 5618 9627
rect 5652 9601 5662 9627
rect 5608 9549 5609 9601
rect 5661 9549 5662 9601
rect 5608 9542 5662 9549
rect 5708 9627 5762 9733
rect 5808 9811 5862 9818
rect 5808 9759 5809 9811
rect 5861 9759 5862 9811
rect 5808 9733 5818 9759
rect 5852 9733 5862 9759
rect 5808 9721 5862 9733
rect 5908 9767 5962 9940
rect 6002 9883 6068 9884
rect 6002 9831 6009 9883
rect 6061 9831 6068 9883
rect 6002 9830 6068 9831
rect 5908 9733 5918 9767
rect 5952 9733 5962 9767
rect 5708 9593 5718 9627
rect 5752 9593 5762 9627
rect 5508 9453 5518 9487
rect 5552 9453 5562 9487
rect 5308 9313 5318 9347
rect 5352 9313 5362 9347
rect 5108 9173 5118 9207
rect 5152 9173 5162 9207
rect 4908 9033 4918 9067
rect 4952 9033 4962 9067
rect 4708 8893 4718 8927
rect 4752 8893 4762 8927
rect 4508 8753 4518 8787
rect 4552 8753 4562 8787
rect 4402 8673 4468 8674
rect 4402 8621 4409 8673
rect 4461 8621 4468 8673
rect 4402 8620 4468 8621
rect 4308 8523 4318 8557
rect 4352 8523 4362 8557
rect 4108 8383 4118 8417
rect 4152 8383 4162 8417
rect 3908 8243 3918 8277
rect 3952 8243 3962 8277
rect 3708 8103 3718 8137
rect 3752 8103 3762 8137
rect 3508 7963 3518 7997
rect 3552 7963 3562 7997
rect 3308 7823 3318 7857
rect 3352 7823 3362 7857
rect 3108 7683 3118 7717
rect 3152 7683 3162 7717
rect 2908 7543 2918 7577
rect 2952 7543 2962 7577
rect 2802 7463 2868 7464
rect 2802 7411 2809 7463
rect 2861 7411 2868 7463
rect 2802 7410 2868 7411
rect 2708 7313 2718 7347
rect 2752 7313 2762 7347
rect 2508 7173 2518 7207
rect 2552 7173 2562 7207
rect 2308 7033 2318 7067
rect 2352 7033 2362 7067
rect 2108 6893 2118 6927
rect 2152 6893 2162 6927
rect 1908 6753 1918 6787
rect 1952 6753 1962 6787
rect 1708 6613 1718 6647
rect 1752 6613 1762 6647
rect 1508 6473 1518 6507
rect 1552 6473 1562 6507
rect 1308 6333 1318 6367
rect 1352 6333 1362 6367
rect 1202 6253 1268 6254
rect 1202 6201 1209 6253
rect 1261 6201 1268 6253
rect 1202 6200 1268 6201
rect 1108 6103 1118 6137
rect 1152 6103 1162 6137
rect 908 5963 918 5997
rect 952 5963 962 5997
rect 708 5823 718 5857
rect 752 5823 762 5857
rect 508 5683 518 5717
rect 552 5683 562 5717
rect 308 5543 318 5577
rect 352 5543 362 5577
rect 108 5403 118 5437
rect 152 5403 162 5437
rect 8 5297 62 5309
rect 8 5271 18 5297
rect 52 5271 62 5297
rect 8 5219 9 5271
rect 61 5219 62 5271
rect 8 5212 62 5219
rect 108 5297 162 5403
rect 208 5481 262 5488
rect 208 5429 209 5481
rect 261 5429 262 5481
rect 208 5403 218 5429
rect 252 5403 262 5429
rect 208 5391 262 5403
rect 308 5437 362 5543
rect 408 5577 462 5589
rect 408 5551 418 5577
rect 452 5551 462 5577
rect 408 5499 409 5551
rect 461 5499 462 5551
rect 408 5492 462 5499
rect 508 5577 562 5683
rect 608 5761 662 5768
rect 608 5709 609 5761
rect 661 5709 662 5761
rect 608 5683 618 5709
rect 652 5683 662 5709
rect 608 5671 662 5683
rect 708 5717 762 5823
rect 808 5857 862 5869
rect 808 5831 818 5857
rect 852 5831 862 5857
rect 808 5779 809 5831
rect 861 5779 862 5831
rect 808 5772 862 5779
rect 908 5857 962 5963
rect 1008 6041 1062 6048
rect 1008 5989 1009 6041
rect 1061 5989 1062 6041
rect 1008 5963 1018 5989
rect 1052 5963 1062 5989
rect 1008 5951 1062 5963
rect 1108 5997 1162 6103
rect 1208 6137 1262 6149
rect 1208 6111 1218 6137
rect 1252 6111 1262 6137
rect 1208 6059 1209 6111
rect 1261 6059 1262 6111
rect 1208 6052 1262 6059
rect 1308 6137 1362 6333
rect 1408 6411 1462 6418
rect 1408 6359 1409 6411
rect 1461 6359 1462 6411
rect 1408 6333 1418 6359
rect 1452 6333 1462 6359
rect 1408 6321 1462 6333
rect 1508 6367 1562 6473
rect 1608 6507 1662 6519
rect 1608 6481 1618 6507
rect 1652 6481 1662 6507
rect 1608 6429 1609 6481
rect 1661 6429 1662 6481
rect 1608 6422 1662 6429
rect 1708 6507 1762 6613
rect 1808 6691 1862 6698
rect 1808 6639 1809 6691
rect 1861 6639 1862 6691
rect 1808 6613 1818 6639
rect 1852 6613 1862 6639
rect 1808 6601 1862 6613
rect 1908 6647 1962 6753
rect 2008 6787 2062 6799
rect 2008 6761 2018 6787
rect 2052 6761 2062 6787
rect 2008 6709 2009 6761
rect 2061 6709 2062 6761
rect 2008 6702 2062 6709
rect 2108 6787 2162 6893
rect 2208 6971 2262 6978
rect 2208 6919 2209 6971
rect 2261 6919 2262 6971
rect 2208 6893 2218 6919
rect 2252 6893 2262 6919
rect 2208 6881 2262 6893
rect 2308 6927 2362 7033
rect 2408 7067 2462 7079
rect 2408 7041 2418 7067
rect 2452 7041 2462 7067
rect 2408 6989 2409 7041
rect 2461 6989 2462 7041
rect 2408 6982 2462 6989
rect 2508 7067 2562 7173
rect 2608 7251 2662 7258
rect 2608 7199 2609 7251
rect 2661 7199 2662 7251
rect 2608 7173 2618 7199
rect 2652 7173 2662 7199
rect 2608 7161 2662 7173
rect 2708 7207 2762 7313
rect 2808 7347 2862 7359
rect 2808 7321 2818 7347
rect 2852 7321 2862 7347
rect 2808 7269 2809 7321
rect 2861 7269 2862 7321
rect 2808 7262 2862 7269
rect 2908 7347 2962 7543
rect 3008 7621 3062 7628
rect 3008 7569 3009 7621
rect 3061 7569 3062 7621
rect 3008 7543 3018 7569
rect 3052 7543 3062 7569
rect 3008 7531 3062 7543
rect 3108 7577 3162 7683
rect 3208 7717 3262 7729
rect 3208 7691 3218 7717
rect 3252 7691 3262 7717
rect 3208 7639 3209 7691
rect 3261 7639 3262 7691
rect 3208 7632 3262 7639
rect 3308 7717 3362 7823
rect 3408 7901 3462 7908
rect 3408 7849 3409 7901
rect 3461 7849 3462 7901
rect 3408 7823 3418 7849
rect 3452 7823 3462 7849
rect 3408 7811 3462 7823
rect 3508 7857 3562 7963
rect 3608 7997 3662 8009
rect 3608 7971 3618 7997
rect 3652 7971 3662 7997
rect 3608 7919 3609 7971
rect 3661 7919 3662 7971
rect 3608 7912 3662 7919
rect 3708 7997 3762 8103
rect 3808 8181 3862 8188
rect 3808 8129 3809 8181
rect 3861 8129 3862 8181
rect 3808 8103 3818 8129
rect 3852 8103 3862 8129
rect 3808 8091 3862 8103
rect 3908 8137 3962 8243
rect 4008 8277 4062 8289
rect 4008 8251 4018 8277
rect 4052 8251 4062 8277
rect 4008 8199 4009 8251
rect 4061 8199 4062 8251
rect 4008 8192 4062 8199
rect 4108 8277 4162 8383
rect 4208 8461 4262 8468
rect 4208 8409 4209 8461
rect 4261 8409 4262 8461
rect 4208 8383 4218 8409
rect 4252 8383 4262 8409
rect 4208 8371 4262 8383
rect 4308 8417 4362 8523
rect 4408 8557 4462 8569
rect 4408 8531 4418 8557
rect 4452 8531 4462 8557
rect 4408 8479 4409 8531
rect 4461 8479 4462 8531
rect 4408 8472 4462 8479
rect 4508 8557 4562 8753
rect 4608 8831 4662 8838
rect 4608 8779 4609 8831
rect 4661 8779 4662 8831
rect 4608 8753 4618 8779
rect 4652 8753 4662 8779
rect 4608 8741 4662 8753
rect 4708 8787 4762 8893
rect 4808 8927 4862 8939
rect 4808 8901 4818 8927
rect 4852 8901 4862 8927
rect 4808 8849 4809 8901
rect 4861 8849 4862 8901
rect 4808 8842 4862 8849
rect 4908 8927 4962 9033
rect 5008 9111 5062 9118
rect 5008 9059 5009 9111
rect 5061 9059 5062 9111
rect 5008 9033 5018 9059
rect 5052 9033 5062 9059
rect 5008 9021 5062 9033
rect 5108 9067 5162 9173
rect 5208 9207 5262 9219
rect 5208 9181 5218 9207
rect 5252 9181 5262 9207
rect 5208 9129 5209 9181
rect 5261 9129 5262 9181
rect 5208 9122 5262 9129
rect 5308 9207 5362 9313
rect 5408 9391 5462 9398
rect 5408 9339 5409 9391
rect 5461 9339 5462 9391
rect 5408 9313 5418 9339
rect 5452 9313 5462 9339
rect 5408 9301 5462 9313
rect 5508 9347 5562 9453
rect 5608 9487 5662 9499
rect 5608 9461 5618 9487
rect 5652 9461 5662 9487
rect 5608 9409 5609 9461
rect 5661 9409 5662 9461
rect 5608 9402 5662 9409
rect 5708 9487 5762 9593
rect 5808 9671 5862 9678
rect 5808 9619 5809 9671
rect 5861 9619 5862 9671
rect 5808 9593 5818 9619
rect 5852 9593 5862 9619
rect 5808 9581 5862 9593
rect 5908 9627 5962 9733
rect 6008 9767 6062 9779
rect 6008 9741 6018 9767
rect 6052 9741 6062 9767
rect 6008 9689 6009 9741
rect 6061 9689 6062 9741
rect 6008 9682 6062 9689
rect 6108 9767 6162 9940
rect 6202 9899 6268 9900
rect 6202 9847 6209 9899
rect 6261 9847 6268 9899
rect 6202 9846 6268 9847
rect 6108 9733 6118 9767
rect 6152 9733 6162 9767
rect 5908 9593 5918 9627
rect 5952 9593 5962 9627
rect 5708 9453 5718 9487
rect 5752 9453 5762 9487
rect 5508 9313 5518 9347
rect 5552 9313 5562 9347
rect 5308 9173 5318 9207
rect 5352 9173 5362 9207
rect 5108 9033 5118 9067
rect 5152 9033 5162 9067
rect 4908 8893 4918 8927
rect 4952 8893 4962 8927
rect 4708 8753 4718 8787
rect 4752 8753 4762 8787
rect 4602 8689 4668 8690
rect 4602 8637 4609 8689
rect 4661 8637 4668 8689
rect 4602 8636 4668 8637
rect 4508 8523 4518 8557
rect 4552 8523 4562 8557
rect 4308 8383 4318 8417
rect 4352 8383 4362 8417
rect 4108 8243 4118 8277
rect 4152 8243 4162 8277
rect 3908 8103 3918 8137
rect 3952 8103 3962 8137
rect 3708 7963 3718 7997
rect 3752 7963 3762 7997
rect 3508 7823 3518 7857
rect 3552 7823 3562 7857
rect 3308 7683 3318 7717
rect 3352 7683 3362 7717
rect 3108 7543 3118 7577
rect 3152 7543 3162 7577
rect 3002 7479 3068 7480
rect 3002 7427 3009 7479
rect 3061 7427 3068 7479
rect 3002 7426 3068 7427
rect 2908 7313 2918 7347
rect 2952 7313 2962 7347
rect 2708 7173 2718 7207
rect 2752 7173 2762 7207
rect 2508 7033 2518 7067
rect 2552 7033 2562 7067
rect 2308 6893 2318 6927
rect 2352 6893 2362 6927
rect 2108 6753 2118 6787
rect 2152 6753 2162 6787
rect 1908 6613 1918 6647
rect 1952 6613 1962 6647
rect 1708 6473 1718 6507
rect 1752 6473 1762 6507
rect 1508 6333 1518 6367
rect 1552 6333 1562 6367
rect 1402 6269 1468 6270
rect 1402 6217 1409 6269
rect 1461 6217 1468 6269
rect 1402 6216 1468 6217
rect 1308 6103 1318 6137
rect 1352 6103 1362 6137
rect 1108 5963 1118 5997
rect 1152 5963 1162 5997
rect 908 5823 918 5857
rect 952 5823 962 5857
rect 708 5683 718 5717
rect 752 5683 762 5717
rect 508 5543 518 5577
rect 552 5543 562 5577
rect 308 5403 318 5437
rect 352 5403 362 5437
rect 108 5263 118 5297
rect 152 5263 162 5297
rect 8 5157 62 5169
rect 8 5131 18 5157
rect 52 5131 62 5157
rect 8 5079 9 5131
rect 61 5079 62 5131
rect 8 5072 62 5079
rect 108 5157 162 5263
rect 208 5341 262 5348
rect 208 5289 209 5341
rect 261 5289 262 5341
rect 208 5263 218 5289
rect 252 5263 262 5289
rect 208 5251 262 5263
rect 308 5297 362 5403
rect 408 5437 462 5449
rect 408 5411 418 5437
rect 452 5411 462 5437
rect 408 5359 409 5411
rect 461 5359 462 5411
rect 408 5352 462 5359
rect 508 5437 562 5543
rect 608 5621 662 5628
rect 608 5569 609 5621
rect 661 5569 662 5621
rect 608 5543 618 5569
rect 652 5543 662 5569
rect 608 5531 662 5543
rect 708 5577 762 5683
rect 808 5717 862 5729
rect 808 5691 818 5717
rect 852 5691 862 5717
rect 808 5639 809 5691
rect 861 5639 862 5691
rect 808 5632 862 5639
rect 908 5717 962 5823
rect 1008 5901 1062 5908
rect 1008 5849 1009 5901
rect 1061 5849 1062 5901
rect 1008 5823 1018 5849
rect 1052 5823 1062 5849
rect 1008 5811 1062 5823
rect 1108 5857 1162 5963
rect 1208 5997 1262 6009
rect 1208 5971 1218 5997
rect 1252 5971 1262 5997
rect 1208 5919 1209 5971
rect 1261 5919 1262 5971
rect 1208 5912 1262 5919
rect 1308 5997 1362 6103
rect 1408 6181 1462 6188
rect 1408 6129 1409 6181
rect 1461 6129 1462 6181
rect 1408 6103 1418 6129
rect 1452 6103 1462 6129
rect 1408 6091 1462 6103
rect 1508 6137 1562 6333
rect 1608 6367 1662 6379
rect 1608 6341 1618 6367
rect 1652 6341 1662 6367
rect 1608 6289 1609 6341
rect 1661 6289 1662 6341
rect 1608 6282 1662 6289
rect 1708 6367 1762 6473
rect 1808 6551 1862 6558
rect 1808 6499 1809 6551
rect 1861 6499 1862 6551
rect 1808 6473 1818 6499
rect 1852 6473 1862 6499
rect 1808 6461 1862 6473
rect 1908 6507 1962 6613
rect 2008 6647 2062 6659
rect 2008 6621 2018 6647
rect 2052 6621 2062 6647
rect 2008 6569 2009 6621
rect 2061 6569 2062 6621
rect 2008 6562 2062 6569
rect 2108 6647 2162 6753
rect 2208 6831 2262 6838
rect 2208 6779 2209 6831
rect 2261 6779 2262 6831
rect 2208 6753 2218 6779
rect 2252 6753 2262 6779
rect 2208 6741 2262 6753
rect 2308 6787 2362 6893
rect 2408 6927 2462 6939
rect 2408 6901 2418 6927
rect 2452 6901 2462 6927
rect 2408 6849 2409 6901
rect 2461 6849 2462 6901
rect 2408 6842 2462 6849
rect 2508 6927 2562 7033
rect 2608 7111 2662 7118
rect 2608 7059 2609 7111
rect 2661 7059 2662 7111
rect 2608 7033 2618 7059
rect 2652 7033 2662 7059
rect 2608 7021 2662 7033
rect 2708 7067 2762 7173
rect 2808 7207 2862 7219
rect 2808 7181 2818 7207
rect 2852 7181 2862 7207
rect 2808 7129 2809 7181
rect 2861 7129 2862 7181
rect 2808 7122 2862 7129
rect 2908 7207 2962 7313
rect 3008 7391 3062 7398
rect 3008 7339 3009 7391
rect 3061 7339 3062 7391
rect 3008 7313 3018 7339
rect 3052 7313 3062 7339
rect 3008 7301 3062 7313
rect 3108 7347 3162 7543
rect 3208 7577 3262 7589
rect 3208 7551 3218 7577
rect 3252 7551 3262 7577
rect 3208 7499 3209 7551
rect 3261 7499 3262 7551
rect 3208 7492 3262 7499
rect 3308 7577 3362 7683
rect 3408 7761 3462 7768
rect 3408 7709 3409 7761
rect 3461 7709 3462 7761
rect 3408 7683 3418 7709
rect 3452 7683 3462 7709
rect 3408 7671 3462 7683
rect 3508 7717 3562 7823
rect 3608 7857 3662 7869
rect 3608 7831 3618 7857
rect 3652 7831 3662 7857
rect 3608 7779 3609 7831
rect 3661 7779 3662 7831
rect 3608 7772 3662 7779
rect 3708 7857 3762 7963
rect 3808 8041 3862 8048
rect 3808 7989 3809 8041
rect 3861 7989 3862 8041
rect 3808 7963 3818 7989
rect 3852 7963 3862 7989
rect 3808 7951 3862 7963
rect 3908 7997 3962 8103
rect 4008 8137 4062 8149
rect 4008 8111 4018 8137
rect 4052 8111 4062 8137
rect 4008 8059 4009 8111
rect 4061 8059 4062 8111
rect 4008 8052 4062 8059
rect 4108 8137 4162 8243
rect 4208 8321 4262 8328
rect 4208 8269 4209 8321
rect 4261 8269 4262 8321
rect 4208 8243 4218 8269
rect 4252 8243 4262 8269
rect 4208 8231 4262 8243
rect 4308 8277 4362 8383
rect 4408 8417 4462 8429
rect 4408 8391 4418 8417
rect 4452 8391 4462 8417
rect 4408 8339 4409 8391
rect 4461 8339 4462 8391
rect 4408 8332 4462 8339
rect 4508 8417 4562 8523
rect 4608 8601 4662 8608
rect 4608 8549 4609 8601
rect 4661 8549 4662 8601
rect 4608 8523 4618 8549
rect 4652 8523 4662 8549
rect 4608 8511 4662 8523
rect 4708 8557 4762 8753
rect 4808 8787 4862 8799
rect 4808 8761 4818 8787
rect 4852 8761 4862 8787
rect 4808 8709 4809 8761
rect 4861 8709 4862 8761
rect 4808 8702 4862 8709
rect 4908 8787 4962 8893
rect 5008 8971 5062 8978
rect 5008 8919 5009 8971
rect 5061 8919 5062 8971
rect 5008 8893 5018 8919
rect 5052 8893 5062 8919
rect 5008 8881 5062 8893
rect 5108 8927 5162 9033
rect 5208 9067 5262 9079
rect 5208 9041 5218 9067
rect 5252 9041 5262 9067
rect 5208 8989 5209 9041
rect 5261 8989 5262 9041
rect 5208 8982 5262 8989
rect 5308 9067 5362 9173
rect 5408 9251 5462 9258
rect 5408 9199 5409 9251
rect 5461 9199 5462 9251
rect 5408 9173 5418 9199
rect 5452 9173 5462 9199
rect 5408 9161 5462 9173
rect 5508 9207 5562 9313
rect 5608 9347 5662 9359
rect 5608 9321 5618 9347
rect 5652 9321 5662 9347
rect 5608 9269 5609 9321
rect 5661 9269 5662 9321
rect 5608 9262 5662 9269
rect 5708 9347 5762 9453
rect 5808 9531 5862 9538
rect 5808 9479 5809 9531
rect 5861 9479 5862 9531
rect 5808 9453 5818 9479
rect 5852 9453 5862 9479
rect 5808 9441 5862 9453
rect 5908 9487 5962 9593
rect 6008 9627 6062 9639
rect 6008 9601 6018 9627
rect 6052 9601 6062 9627
rect 6008 9549 6009 9601
rect 6061 9549 6062 9601
rect 6008 9542 6062 9549
rect 6108 9627 6162 9733
rect 6208 9811 6262 9818
rect 6208 9759 6209 9811
rect 6261 9759 6262 9811
rect 6208 9733 6218 9759
rect 6252 9733 6262 9759
rect 6208 9721 6262 9733
rect 6308 9767 6362 9940
rect 6590 9877 6620 10050
rect 6504 9871 6620 9877
rect 6504 9837 6516 9871
rect 6550 9837 6620 9871
rect 6504 9831 6620 9837
rect 6506 9782 6560 9794
rect 6308 9733 6318 9767
rect 6352 9733 6362 9767
rect 6108 9593 6118 9627
rect 6152 9593 6162 9627
rect 5908 9453 5918 9487
rect 5952 9453 5962 9487
rect 5708 9313 5718 9347
rect 5752 9313 5762 9347
rect 5508 9173 5518 9207
rect 5552 9173 5562 9207
rect 5308 9033 5318 9067
rect 5352 9033 5362 9067
rect 5108 8893 5118 8927
rect 5152 8893 5162 8927
rect 4908 8753 4918 8787
rect 4952 8753 4962 8787
rect 4802 8673 4868 8674
rect 4802 8621 4809 8673
rect 4861 8621 4868 8673
rect 4802 8620 4868 8621
rect 4708 8523 4718 8557
rect 4752 8523 4762 8557
rect 4508 8383 4518 8417
rect 4552 8383 4562 8417
rect 4308 8243 4318 8277
rect 4352 8243 4362 8277
rect 4108 8103 4118 8137
rect 4152 8103 4162 8137
rect 3908 7963 3918 7997
rect 3952 7963 3962 7997
rect 3708 7823 3718 7857
rect 3752 7823 3762 7857
rect 3508 7683 3518 7717
rect 3552 7683 3562 7717
rect 3308 7543 3318 7577
rect 3352 7543 3362 7577
rect 3202 7463 3268 7464
rect 3202 7411 3209 7463
rect 3261 7411 3268 7463
rect 3202 7410 3268 7411
rect 3108 7313 3118 7347
rect 3152 7313 3162 7347
rect 2908 7173 2918 7207
rect 2952 7173 2962 7207
rect 2708 7033 2718 7067
rect 2752 7033 2762 7067
rect 2508 6893 2518 6927
rect 2552 6893 2562 6927
rect 2308 6753 2318 6787
rect 2352 6753 2362 6787
rect 2108 6613 2118 6647
rect 2152 6613 2162 6647
rect 1908 6473 1918 6507
rect 1952 6473 1962 6507
rect 1708 6333 1718 6367
rect 1752 6333 1762 6367
rect 1602 6253 1668 6254
rect 1602 6201 1609 6253
rect 1661 6201 1668 6253
rect 1602 6200 1668 6201
rect 1508 6103 1518 6137
rect 1552 6103 1562 6137
rect 1308 5963 1318 5997
rect 1352 5963 1362 5997
rect 1108 5823 1118 5857
rect 1152 5823 1162 5857
rect 908 5683 918 5717
rect 952 5683 962 5717
rect 708 5543 718 5577
rect 752 5543 762 5577
rect 508 5403 518 5437
rect 552 5403 562 5437
rect 308 5263 318 5297
rect 352 5263 362 5297
rect 108 5123 118 5157
rect 152 5123 162 5157
rect 108 5040 162 5123
rect 208 5201 262 5208
rect 208 5149 209 5201
rect 261 5149 262 5201
rect 208 5123 218 5149
rect 252 5123 262 5149
rect 208 5111 262 5123
rect 308 5157 362 5263
rect 408 5297 462 5309
rect 408 5271 418 5297
rect 452 5271 462 5297
rect 408 5219 409 5271
rect 461 5219 462 5271
rect 408 5212 462 5219
rect 508 5297 562 5403
rect 608 5481 662 5488
rect 608 5429 609 5481
rect 661 5429 662 5481
rect 608 5403 618 5429
rect 652 5403 662 5429
rect 608 5391 662 5403
rect 708 5437 762 5543
rect 808 5577 862 5589
rect 808 5551 818 5577
rect 852 5551 862 5577
rect 808 5499 809 5551
rect 861 5499 862 5551
rect 808 5492 862 5499
rect 908 5577 962 5683
rect 1008 5761 1062 5768
rect 1008 5709 1009 5761
rect 1061 5709 1062 5761
rect 1008 5683 1018 5709
rect 1052 5683 1062 5709
rect 1008 5671 1062 5683
rect 1108 5717 1162 5823
rect 1208 5857 1262 5869
rect 1208 5831 1218 5857
rect 1252 5831 1262 5857
rect 1208 5779 1209 5831
rect 1261 5779 1262 5831
rect 1208 5772 1262 5779
rect 1308 5857 1362 5963
rect 1408 6041 1462 6048
rect 1408 5989 1409 6041
rect 1461 5989 1462 6041
rect 1408 5963 1418 5989
rect 1452 5963 1462 5989
rect 1408 5951 1462 5963
rect 1508 5997 1562 6103
rect 1608 6137 1662 6149
rect 1608 6111 1618 6137
rect 1652 6111 1662 6137
rect 1608 6059 1609 6111
rect 1661 6059 1662 6111
rect 1608 6052 1662 6059
rect 1708 6137 1762 6333
rect 1808 6411 1862 6418
rect 1808 6359 1809 6411
rect 1861 6359 1862 6411
rect 1808 6333 1818 6359
rect 1852 6333 1862 6359
rect 1808 6321 1862 6333
rect 1908 6367 1962 6473
rect 2008 6507 2062 6519
rect 2008 6481 2018 6507
rect 2052 6481 2062 6507
rect 2008 6429 2009 6481
rect 2061 6429 2062 6481
rect 2008 6422 2062 6429
rect 2108 6507 2162 6613
rect 2208 6691 2262 6698
rect 2208 6639 2209 6691
rect 2261 6639 2262 6691
rect 2208 6613 2218 6639
rect 2252 6613 2262 6639
rect 2208 6601 2262 6613
rect 2308 6647 2362 6753
rect 2408 6787 2462 6799
rect 2408 6761 2418 6787
rect 2452 6761 2462 6787
rect 2408 6709 2409 6761
rect 2461 6709 2462 6761
rect 2408 6702 2462 6709
rect 2508 6787 2562 6893
rect 2608 6971 2662 6978
rect 2608 6919 2609 6971
rect 2661 6919 2662 6971
rect 2608 6893 2618 6919
rect 2652 6893 2662 6919
rect 2608 6881 2662 6893
rect 2708 6927 2762 7033
rect 2808 7067 2862 7079
rect 2808 7041 2818 7067
rect 2852 7041 2862 7067
rect 2808 6989 2809 7041
rect 2861 6989 2862 7041
rect 2808 6982 2862 6989
rect 2908 7067 2962 7173
rect 3008 7251 3062 7258
rect 3008 7199 3009 7251
rect 3061 7199 3062 7251
rect 3008 7173 3018 7199
rect 3052 7173 3062 7199
rect 3008 7161 3062 7173
rect 3108 7207 3162 7313
rect 3208 7347 3262 7359
rect 3208 7321 3218 7347
rect 3252 7321 3262 7347
rect 3208 7269 3209 7321
rect 3261 7269 3262 7321
rect 3208 7262 3262 7269
rect 3308 7347 3362 7543
rect 3408 7621 3462 7628
rect 3408 7569 3409 7621
rect 3461 7569 3462 7621
rect 3408 7543 3418 7569
rect 3452 7543 3462 7569
rect 3408 7531 3462 7543
rect 3508 7577 3562 7683
rect 3608 7717 3662 7729
rect 3608 7691 3618 7717
rect 3652 7691 3662 7717
rect 3608 7639 3609 7691
rect 3661 7639 3662 7691
rect 3608 7632 3662 7639
rect 3708 7717 3762 7823
rect 3808 7901 3862 7908
rect 3808 7849 3809 7901
rect 3861 7849 3862 7901
rect 3808 7823 3818 7849
rect 3852 7823 3862 7849
rect 3808 7811 3862 7823
rect 3908 7857 3962 7963
rect 4008 7997 4062 8009
rect 4008 7971 4018 7997
rect 4052 7971 4062 7997
rect 4008 7919 4009 7971
rect 4061 7919 4062 7971
rect 4008 7912 4062 7919
rect 4108 7997 4162 8103
rect 4208 8181 4262 8188
rect 4208 8129 4209 8181
rect 4261 8129 4262 8181
rect 4208 8103 4218 8129
rect 4252 8103 4262 8129
rect 4208 8091 4262 8103
rect 4308 8137 4362 8243
rect 4408 8277 4462 8289
rect 4408 8251 4418 8277
rect 4452 8251 4462 8277
rect 4408 8199 4409 8251
rect 4461 8199 4462 8251
rect 4408 8192 4462 8199
rect 4508 8277 4562 8383
rect 4608 8461 4662 8468
rect 4608 8409 4609 8461
rect 4661 8409 4662 8461
rect 4608 8383 4618 8409
rect 4652 8383 4662 8409
rect 4608 8371 4662 8383
rect 4708 8417 4762 8523
rect 4808 8557 4862 8569
rect 4808 8531 4818 8557
rect 4852 8531 4862 8557
rect 4808 8479 4809 8531
rect 4861 8479 4862 8531
rect 4808 8472 4862 8479
rect 4908 8557 4962 8753
rect 5008 8831 5062 8838
rect 5008 8779 5009 8831
rect 5061 8779 5062 8831
rect 5008 8753 5018 8779
rect 5052 8753 5062 8779
rect 5008 8741 5062 8753
rect 5108 8787 5162 8893
rect 5208 8927 5262 8939
rect 5208 8901 5218 8927
rect 5252 8901 5262 8927
rect 5208 8849 5209 8901
rect 5261 8849 5262 8901
rect 5208 8842 5262 8849
rect 5308 8927 5362 9033
rect 5408 9111 5462 9118
rect 5408 9059 5409 9111
rect 5461 9059 5462 9111
rect 5408 9033 5418 9059
rect 5452 9033 5462 9059
rect 5408 9021 5462 9033
rect 5508 9067 5562 9173
rect 5608 9207 5662 9219
rect 5608 9181 5618 9207
rect 5652 9181 5662 9207
rect 5608 9129 5609 9181
rect 5661 9129 5662 9181
rect 5608 9122 5662 9129
rect 5708 9207 5762 9313
rect 5808 9391 5862 9398
rect 5808 9339 5809 9391
rect 5861 9339 5862 9391
rect 5808 9313 5818 9339
rect 5852 9313 5862 9339
rect 5808 9301 5862 9313
rect 5908 9347 5962 9453
rect 6008 9487 6062 9499
rect 6008 9461 6018 9487
rect 6052 9461 6062 9487
rect 6008 9409 6009 9461
rect 6061 9409 6062 9461
rect 6008 9402 6062 9409
rect 6108 9487 6162 9593
rect 6208 9671 6262 9678
rect 6208 9619 6209 9671
rect 6261 9619 6262 9671
rect 6208 9593 6218 9619
rect 6252 9593 6262 9619
rect 6208 9581 6262 9593
rect 6308 9627 6362 9733
rect 6408 9767 6462 9779
rect 6408 9741 6418 9767
rect 6452 9741 6462 9767
rect 6408 9689 6409 9741
rect 6461 9689 6462 9741
rect 6408 9682 6462 9689
rect 6506 9748 6516 9782
rect 6550 9748 6560 9782
rect 6506 9741 6560 9748
rect 6506 9689 6507 9741
rect 6559 9689 6560 9741
rect 6506 9682 6560 9689
rect 6506 9642 6560 9654
rect 6308 9593 6318 9627
rect 6352 9593 6362 9627
rect 6108 9453 6118 9487
rect 6152 9453 6162 9487
rect 5908 9313 5918 9347
rect 5952 9313 5962 9347
rect 5708 9173 5718 9207
rect 5752 9173 5762 9207
rect 5508 9033 5518 9067
rect 5552 9033 5562 9067
rect 5308 8893 5318 8927
rect 5352 8893 5362 8927
rect 5108 8753 5118 8787
rect 5152 8753 5162 8787
rect 5002 8689 5068 8690
rect 5002 8637 5009 8689
rect 5061 8637 5068 8689
rect 5002 8636 5068 8637
rect 4908 8523 4918 8557
rect 4952 8523 4962 8557
rect 4708 8383 4718 8417
rect 4752 8383 4762 8417
rect 4508 8243 4518 8277
rect 4552 8243 4562 8277
rect 4308 8103 4318 8137
rect 4352 8103 4362 8137
rect 4108 7963 4118 7997
rect 4152 7963 4162 7997
rect 3908 7823 3918 7857
rect 3952 7823 3962 7857
rect 3708 7683 3718 7717
rect 3752 7683 3762 7717
rect 3508 7543 3518 7577
rect 3552 7543 3562 7577
rect 3402 7479 3468 7480
rect 3402 7427 3409 7479
rect 3461 7427 3468 7479
rect 3402 7426 3468 7427
rect 3308 7313 3318 7347
rect 3352 7313 3362 7347
rect 3108 7173 3118 7207
rect 3152 7173 3162 7207
rect 2908 7033 2918 7067
rect 2952 7033 2962 7067
rect 2708 6893 2718 6927
rect 2752 6893 2762 6927
rect 2508 6753 2518 6787
rect 2552 6753 2562 6787
rect 2308 6613 2318 6647
rect 2352 6613 2362 6647
rect 2108 6473 2118 6507
rect 2152 6473 2162 6507
rect 1908 6333 1918 6367
rect 1952 6333 1962 6367
rect 1802 6269 1868 6270
rect 1802 6217 1809 6269
rect 1861 6217 1868 6269
rect 1802 6216 1868 6217
rect 1708 6103 1718 6137
rect 1752 6103 1762 6137
rect 1508 5963 1518 5997
rect 1552 5963 1562 5997
rect 1308 5823 1318 5857
rect 1352 5823 1362 5857
rect 1108 5683 1118 5717
rect 1152 5683 1162 5717
rect 908 5543 918 5577
rect 952 5543 962 5577
rect 708 5403 718 5437
rect 752 5403 762 5437
rect 508 5263 518 5297
rect 552 5263 562 5297
rect 308 5123 318 5157
rect 352 5123 362 5157
rect 308 5040 362 5123
rect 408 5157 462 5169
rect 408 5131 418 5157
rect 452 5131 462 5157
rect 408 5079 409 5131
rect 461 5079 462 5131
rect 408 5072 462 5079
rect 508 5157 562 5263
rect 608 5341 662 5348
rect 608 5289 609 5341
rect 661 5289 662 5341
rect 608 5263 618 5289
rect 652 5263 662 5289
rect 608 5251 662 5263
rect 708 5297 762 5403
rect 808 5437 862 5449
rect 808 5411 818 5437
rect 852 5411 862 5437
rect 808 5359 809 5411
rect 861 5359 862 5411
rect 808 5352 862 5359
rect 908 5437 962 5543
rect 1008 5621 1062 5628
rect 1008 5569 1009 5621
rect 1061 5569 1062 5621
rect 1008 5543 1018 5569
rect 1052 5543 1062 5569
rect 1008 5531 1062 5543
rect 1108 5577 1162 5683
rect 1208 5717 1262 5729
rect 1208 5691 1218 5717
rect 1252 5691 1262 5717
rect 1208 5639 1209 5691
rect 1261 5639 1262 5691
rect 1208 5632 1262 5639
rect 1308 5717 1362 5823
rect 1408 5901 1462 5908
rect 1408 5849 1409 5901
rect 1461 5849 1462 5901
rect 1408 5823 1418 5849
rect 1452 5823 1462 5849
rect 1408 5811 1462 5823
rect 1508 5857 1562 5963
rect 1608 5997 1662 6009
rect 1608 5971 1618 5997
rect 1652 5971 1662 5997
rect 1608 5919 1609 5971
rect 1661 5919 1662 5971
rect 1608 5912 1662 5919
rect 1708 5997 1762 6103
rect 1808 6181 1862 6188
rect 1808 6129 1809 6181
rect 1861 6129 1862 6181
rect 1808 6103 1818 6129
rect 1852 6103 1862 6129
rect 1808 6091 1862 6103
rect 1908 6137 1962 6333
rect 2008 6367 2062 6379
rect 2008 6341 2018 6367
rect 2052 6341 2062 6367
rect 2008 6289 2009 6341
rect 2061 6289 2062 6341
rect 2008 6282 2062 6289
rect 2108 6367 2162 6473
rect 2208 6551 2262 6558
rect 2208 6499 2209 6551
rect 2261 6499 2262 6551
rect 2208 6473 2218 6499
rect 2252 6473 2262 6499
rect 2208 6461 2262 6473
rect 2308 6507 2362 6613
rect 2408 6647 2462 6659
rect 2408 6621 2418 6647
rect 2452 6621 2462 6647
rect 2408 6569 2409 6621
rect 2461 6569 2462 6621
rect 2408 6562 2462 6569
rect 2508 6647 2562 6753
rect 2608 6831 2662 6838
rect 2608 6779 2609 6831
rect 2661 6779 2662 6831
rect 2608 6753 2618 6779
rect 2652 6753 2662 6779
rect 2608 6741 2662 6753
rect 2708 6787 2762 6893
rect 2808 6927 2862 6939
rect 2808 6901 2818 6927
rect 2852 6901 2862 6927
rect 2808 6849 2809 6901
rect 2861 6849 2862 6901
rect 2808 6842 2862 6849
rect 2908 6927 2962 7033
rect 3008 7111 3062 7118
rect 3008 7059 3009 7111
rect 3061 7059 3062 7111
rect 3008 7033 3018 7059
rect 3052 7033 3062 7059
rect 3008 7021 3062 7033
rect 3108 7067 3162 7173
rect 3208 7207 3262 7219
rect 3208 7181 3218 7207
rect 3252 7181 3262 7207
rect 3208 7129 3209 7181
rect 3261 7129 3262 7181
rect 3208 7122 3262 7129
rect 3308 7207 3362 7313
rect 3408 7391 3462 7398
rect 3408 7339 3409 7391
rect 3461 7339 3462 7391
rect 3408 7313 3418 7339
rect 3452 7313 3462 7339
rect 3408 7301 3462 7313
rect 3508 7347 3562 7543
rect 3608 7577 3662 7589
rect 3608 7551 3618 7577
rect 3652 7551 3662 7577
rect 3608 7499 3609 7551
rect 3661 7499 3662 7551
rect 3608 7492 3662 7499
rect 3708 7577 3762 7683
rect 3808 7761 3862 7768
rect 3808 7709 3809 7761
rect 3861 7709 3862 7761
rect 3808 7683 3818 7709
rect 3852 7683 3862 7709
rect 3808 7671 3862 7683
rect 3908 7717 3962 7823
rect 4008 7857 4062 7869
rect 4008 7831 4018 7857
rect 4052 7831 4062 7857
rect 4008 7779 4009 7831
rect 4061 7779 4062 7831
rect 4008 7772 4062 7779
rect 4108 7857 4162 7963
rect 4208 8041 4262 8048
rect 4208 7989 4209 8041
rect 4261 7989 4262 8041
rect 4208 7963 4218 7989
rect 4252 7963 4262 7989
rect 4208 7951 4262 7963
rect 4308 7997 4362 8103
rect 4408 8137 4462 8149
rect 4408 8111 4418 8137
rect 4452 8111 4462 8137
rect 4408 8059 4409 8111
rect 4461 8059 4462 8111
rect 4408 8052 4462 8059
rect 4508 8137 4562 8243
rect 4608 8321 4662 8328
rect 4608 8269 4609 8321
rect 4661 8269 4662 8321
rect 4608 8243 4618 8269
rect 4652 8243 4662 8269
rect 4608 8231 4662 8243
rect 4708 8277 4762 8383
rect 4808 8417 4862 8429
rect 4808 8391 4818 8417
rect 4852 8391 4862 8417
rect 4808 8339 4809 8391
rect 4861 8339 4862 8391
rect 4808 8332 4862 8339
rect 4908 8417 4962 8523
rect 5008 8601 5062 8608
rect 5008 8549 5009 8601
rect 5061 8549 5062 8601
rect 5008 8523 5018 8549
rect 5052 8523 5062 8549
rect 5008 8511 5062 8523
rect 5108 8557 5162 8753
rect 5208 8787 5262 8799
rect 5208 8761 5218 8787
rect 5252 8761 5262 8787
rect 5208 8709 5209 8761
rect 5261 8709 5262 8761
rect 5208 8702 5262 8709
rect 5308 8787 5362 8893
rect 5408 8971 5462 8978
rect 5408 8919 5409 8971
rect 5461 8919 5462 8971
rect 5408 8893 5418 8919
rect 5452 8893 5462 8919
rect 5408 8881 5462 8893
rect 5508 8927 5562 9033
rect 5608 9067 5662 9079
rect 5608 9041 5618 9067
rect 5652 9041 5662 9067
rect 5608 8989 5609 9041
rect 5661 8989 5662 9041
rect 5608 8982 5662 8989
rect 5708 9067 5762 9173
rect 5808 9251 5862 9258
rect 5808 9199 5809 9251
rect 5861 9199 5862 9251
rect 5808 9173 5818 9199
rect 5852 9173 5862 9199
rect 5808 9161 5862 9173
rect 5908 9207 5962 9313
rect 6008 9347 6062 9359
rect 6008 9321 6018 9347
rect 6052 9321 6062 9347
rect 6008 9269 6009 9321
rect 6061 9269 6062 9321
rect 6008 9262 6062 9269
rect 6108 9347 6162 9453
rect 6208 9531 6262 9538
rect 6208 9479 6209 9531
rect 6261 9479 6262 9531
rect 6208 9453 6218 9479
rect 6252 9453 6262 9479
rect 6208 9441 6262 9453
rect 6308 9487 6362 9593
rect 6408 9627 6462 9639
rect 6408 9601 6418 9627
rect 6452 9601 6462 9627
rect 6408 9549 6409 9601
rect 6461 9549 6462 9601
rect 6408 9542 6462 9549
rect 6506 9608 6516 9642
rect 6550 9608 6560 9642
rect 6506 9601 6560 9608
rect 6506 9549 6507 9601
rect 6559 9549 6560 9601
rect 6506 9542 6560 9549
rect 6506 9502 6560 9514
rect 6308 9453 6318 9487
rect 6352 9453 6362 9487
rect 6108 9313 6118 9347
rect 6152 9313 6162 9347
rect 5908 9173 5918 9207
rect 5952 9173 5962 9207
rect 5708 9033 5718 9067
rect 5752 9033 5762 9067
rect 5508 8893 5518 8927
rect 5552 8893 5562 8927
rect 5308 8753 5318 8787
rect 5352 8753 5362 8787
rect 5202 8673 5268 8674
rect 5202 8621 5209 8673
rect 5261 8621 5268 8673
rect 5202 8620 5268 8621
rect 5108 8523 5118 8557
rect 5152 8523 5162 8557
rect 4908 8383 4918 8417
rect 4952 8383 4962 8417
rect 4708 8243 4718 8277
rect 4752 8243 4762 8277
rect 4508 8103 4518 8137
rect 4552 8103 4562 8137
rect 4308 7963 4318 7997
rect 4352 7963 4362 7997
rect 4108 7823 4118 7857
rect 4152 7823 4162 7857
rect 3908 7683 3918 7717
rect 3952 7683 3962 7717
rect 3708 7543 3718 7577
rect 3752 7543 3762 7577
rect 3602 7463 3668 7464
rect 3602 7411 3609 7463
rect 3661 7411 3668 7463
rect 3602 7410 3668 7411
rect 3508 7313 3518 7347
rect 3552 7313 3562 7347
rect 3308 7173 3318 7207
rect 3352 7173 3362 7207
rect 3108 7033 3118 7067
rect 3152 7033 3162 7067
rect 2908 6893 2918 6927
rect 2952 6893 2962 6927
rect 2708 6753 2718 6787
rect 2752 6753 2762 6787
rect 2508 6613 2518 6647
rect 2552 6613 2562 6647
rect 2308 6473 2318 6507
rect 2352 6473 2362 6507
rect 2108 6333 2118 6367
rect 2152 6333 2162 6367
rect 2002 6253 2068 6254
rect 2002 6201 2009 6253
rect 2061 6201 2068 6253
rect 2002 6200 2068 6201
rect 1908 6103 1918 6137
rect 1952 6103 1962 6137
rect 1708 5963 1718 5997
rect 1752 5963 1762 5997
rect 1508 5823 1518 5857
rect 1552 5823 1562 5857
rect 1308 5683 1318 5717
rect 1352 5683 1362 5717
rect 1108 5543 1118 5577
rect 1152 5543 1162 5577
rect 908 5403 918 5437
rect 952 5403 962 5437
rect 708 5263 718 5297
rect 752 5263 762 5297
rect 508 5123 518 5157
rect 552 5123 562 5157
rect 508 5040 562 5123
rect 608 5201 662 5208
rect 608 5149 609 5201
rect 661 5149 662 5201
rect 608 5123 618 5149
rect 652 5123 662 5149
rect 608 5111 662 5123
rect 708 5157 762 5263
rect 808 5297 862 5309
rect 808 5271 818 5297
rect 852 5271 862 5297
rect 808 5219 809 5271
rect 861 5219 862 5271
rect 808 5212 862 5219
rect 908 5297 962 5403
rect 1008 5481 1062 5488
rect 1008 5429 1009 5481
rect 1061 5429 1062 5481
rect 1008 5403 1018 5429
rect 1052 5403 1062 5429
rect 1008 5391 1062 5403
rect 1108 5437 1162 5543
rect 1208 5577 1262 5589
rect 1208 5551 1218 5577
rect 1252 5551 1262 5577
rect 1208 5499 1209 5551
rect 1261 5499 1262 5551
rect 1208 5492 1262 5499
rect 1308 5577 1362 5683
rect 1408 5761 1462 5768
rect 1408 5709 1409 5761
rect 1461 5709 1462 5761
rect 1408 5683 1418 5709
rect 1452 5683 1462 5709
rect 1408 5671 1462 5683
rect 1508 5717 1562 5823
rect 1608 5857 1662 5869
rect 1608 5831 1618 5857
rect 1652 5831 1662 5857
rect 1608 5779 1609 5831
rect 1661 5779 1662 5831
rect 1608 5772 1662 5779
rect 1708 5857 1762 5963
rect 1808 6041 1862 6048
rect 1808 5989 1809 6041
rect 1861 5989 1862 6041
rect 1808 5963 1818 5989
rect 1852 5963 1862 5989
rect 1808 5951 1862 5963
rect 1908 5997 1962 6103
rect 2008 6137 2062 6149
rect 2008 6111 2018 6137
rect 2052 6111 2062 6137
rect 2008 6059 2009 6111
rect 2061 6059 2062 6111
rect 2008 6052 2062 6059
rect 2108 6137 2162 6333
rect 2208 6411 2262 6418
rect 2208 6359 2209 6411
rect 2261 6359 2262 6411
rect 2208 6333 2218 6359
rect 2252 6333 2262 6359
rect 2208 6321 2262 6333
rect 2308 6367 2362 6473
rect 2408 6507 2462 6519
rect 2408 6481 2418 6507
rect 2452 6481 2462 6507
rect 2408 6429 2409 6481
rect 2461 6429 2462 6481
rect 2408 6422 2462 6429
rect 2508 6507 2562 6613
rect 2608 6691 2662 6698
rect 2608 6639 2609 6691
rect 2661 6639 2662 6691
rect 2608 6613 2618 6639
rect 2652 6613 2662 6639
rect 2608 6601 2662 6613
rect 2708 6647 2762 6753
rect 2808 6787 2862 6799
rect 2808 6761 2818 6787
rect 2852 6761 2862 6787
rect 2808 6709 2809 6761
rect 2861 6709 2862 6761
rect 2808 6702 2862 6709
rect 2908 6787 2962 6893
rect 3008 6971 3062 6978
rect 3008 6919 3009 6971
rect 3061 6919 3062 6971
rect 3008 6893 3018 6919
rect 3052 6893 3062 6919
rect 3008 6881 3062 6893
rect 3108 6927 3162 7033
rect 3208 7067 3262 7079
rect 3208 7041 3218 7067
rect 3252 7041 3262 7067
rect 3208 6989 3209 7041
rect 3261 6989 3262 7041
rect 3208 6982 3262 6989
rect 3308 7067 3362 7173
rect 3408 7251 3462 7258
rect 3408 7199 3409 7251
rect 3461 7199 3462 7251
rect 3408 7173 3418 7199
rect 3452 7173 3462 7199
rect 3408 7161 3462 7173
rect 3508 7207 3562 7313
rect 3608 7347 3662 7359
rect 3608 7321 3618 7347
rect 3652 7321 3662 7347
rect 3608 7269 3609 7321
rect 3661 7269 3662 7321
rect 3608 7262 3662 7269
rect 3708 7347 3762 7543
rect 3808 7621 3862 7628
rect 3808 7569 3809 7621
rect 3861 7569 3862 7621
rect 3808 7543 3818 7569
rect 3852 7543 3862 7569
rect 3808 7531 3862 7543
rect 3908 7577 3962 7683
rect 4008 7717 4062 7729
rect 4008 7691 4018 7717
rect 4052 7691 4062 7717
rect 4008 7639 4009 7691
rect 4061 7639 4062 7691
rect 4008 7632 4062 7639
rect 4108 7717 4162 7823
rect 4208 7901 4262 7908
rect 4208 7849 4209 7901
rect 4261 7849 4262 7901
rect 4208 7823 4218 7849
rect 4252 7823 4262 7849
rect 4208 7811 4262 7823
rect 4308 7857 4362 7963
rect 4408 7997 4462 8009
rect 4408 7971 4418 7997
rect 4452 7971 4462 7997
rect 4408 7919 4409 7971
rect 4461 7919 4462 7971
rect 4408 7912 4462 7919
rect 4508 7997 4562 8103
rect 4608 8181 4662 8188
rect 4608 8129 4609 8181
rect 4661 8129 4662 8181
rect 4608 8103 4618 8129
rect 4652 8103 4662 8129
rect 4608 8091 4662 8103
rect 4708 8137 4762 8243
rect 4808 8277 4862 8289
rect 4808 8251 4818 8277
rect 4852 8251 4862 8277
rect 4808 8199 4809 8251
rect 4861 8199 4862 8251
rect 4808 8192 4862 8199
rect 4908 8277 4962 8383
rect 5008 8461 5062 8468
rect 5008 8409 5009 8461
rect 5061 8409 5062 8461
rect 5008 8383 5018 8409
rect 5052 8383 5062 8409
rect 5008 8371 5062 8383
rect 5108 8417 5162 8523
rect 5208 8557 5262 8569
rect 5208 8531 5218 8557
rect 5252 8531 5262 8557
rect 5208 8479 5209 8531
rect 5261 8479 5262 8531
rect 5208 8472 5262 8479
rect 5308 8557 5362 8753
rect 5408 8831 5462 8838
rect 5408 8779 5409 8831
rect 5461 8779 5462 8831
rect 5408 8753 5418 8779
rect 5452 8753 5462 8779
rect 5408 8741 5462 8753
rect 5508 8787 5562 8893
rect 5608 8927 5662 8939
rect 5608 8901 5618 8927
rect 5652 8901 5662 8927
rect 5608 8849 5609 8901
rect 5661 8849 5662 8901
rect 5608 8842 5662 8849
rect 5708 8927 5762 9033
rect 5808 9111 5862 9118
rect 5808 9059 5809 9111
rect 5861 9059 5862 9111
rect 5808 9033 5818 9059
rect 5852 9033 5862 9059
rect 5808 9021 5862 9033
rect 5908 9067 5962 9173
rect 6008 9207 6062 9219
rect 6008 9181 6018 9207
rect 6052 9181 6062 9207
rect 6008 9129 6009 9181
rect 6061 9129 6062 9181
rect 6008 9122 6062 9129
rect 6108 9207 6162 9313
rect 6208 9391 6262 9398
rect 6208 9339 6209 9391
rect 6261 9339 6262 9391
rect 6208 9313 6218 9339
rect 6252 9313 6262 9339
rect 6208 9301 6262 9313
rect 6308 9347 6362 9453
rect 6408 9487 6462 9499
rect 6408 9461 6418 9487
rect 6452 9461 6462 9487
rect 6408 9409 6409 9461
rect 6461 9409 6462 9461
rect 6408 9402 6462 9409
rect 6506 9468 6516 9502
rect 6550 9468 6560 9502
rect 6506 9461 6560 9468
rect 6506 9409 6507 9461
rect 6559 9409 6560 9461
rect 6506 9402 6560 9409
rect 6506 9362 6560 9374
rect 6308 9313 6318 9347
rect 6352 9313 6362 9347
rect 6108 9173 6118 9207
rect 6152 9173 6162 9207
rect 5908 9033 5918 9067
rect 5952 9033 5962 9067
rect 5708 8893 5718 8927
rect 5752 8893 5762 8927
rect 5508 8753 5518 8787
rect 5552 8753 5562 8787
rect 5402 8689 5468 8690
rect 5402 8637 5409 8689
rect 5461 8637 5468 8689
rect 5402 8636 5468 8637
rect 5308 8523 5318 8557
rect 5352 8523 5362 8557
rect 5108 8383 5118 8417
rect 5152 8383 5162 8417
rect 4908 8243 4918 8277
rect 4952 8243 4962 8277
rect 4708 8103 4718 8137
rect 4752 8103 4762 8137
rect 4508 7963 4518 7997
rect 4552 7963 4562 7997
rect 4308 7823 4318 7857
rect 4352 7823 4362 7857
rect 4108 7683 4118 7717
rect 4152 7683 4162 7717
rect 3908 7543 3918 7577
rect 3952 7543 3962 7577
rect 3802 7479 3868 7480
rect 3802 7427 3809 7479
rect 3861 7427 3868 7479
rect 3802 7426 3868 7427
rect 3708 7313 3718 7347
rect 3752 7313 3762 7347
rect 3508 7173 3518 7207
rect 3552 7173 3562 7207
rect 3308 7033 3318 7067
rect 3352 7033 3362 7067
rect 3108 6893 3118 6927
rect 3152 6893 3162 6927
rect 2908 6753 2918 6787
rect 2952 6753 2962 6787
rect 2708 6613 2718 6647
rect 2752 6613 2762 6647
rect 2508 6473 2518 6507
rect 2552 6473 2562 6507
rect 2308 6333 2318 6367
rect 2352 6333 2362 6367
rect 2202 6269 2268 6270
rect 2202 6217 2209 6269
rect 2261 6217 2268 6269
rect 2202 6216 2268 6217
rect 2108 6103 2118 6137
rect 2152 6103 2162 6137
rect 1908 5963 1918 5997
rect 1952 5963 1962 5997
rect 1708 5823 1718 5857
rect 1752 5823 1762 5857
rect 1508 5683 1518 5717
rect 1552 5683 1562 5717
rect 1308 5543 1318 5577
rect 1352 5543 1362 5577
rect 1108 5403 1118 5437
rect 1152 5403 1162 5437
rect 908 5263 918 5297
rect 952 5263 962 5297
rect 708 5123 718 5157
rect 752 5123 762 5157
rect 708 5040 762 5123
rect 808 5157 862 5169
rect 808 5131 818 5157
rect 852 5131 862 5157
rect 808 5079 809 5131
rect 861 5079 862 5131
rect 808 5072 862 5079
rect 908 5157 962 5263
rect 1008 5341 1062 5348
rect 1008 5289 1009 5341
rect 1061 5289 1062 5341
rect 1008 5263 1018 5289
rect 1052 5263 1062 5289
rect 1008 5251 1062 5263
rect 1108 5297 1162 5403
rect 1208 5437 1262 5449
rect 1208 5411 1218 5437
rect 1252 5411 1262 5437
rect 1208 5359 1209 5411
rect 1261 5359 1262 5411
rect 1208 5352 1262 5359
rect 1308 5437 1362 5543
rect 1408 5621 1462 5628
rect 1408 5569 1409 5621
rect 1461 5569 1462 5621
rect 1408 5543 1418 5569
rect 1452 5543 1462 5569
rect 1408 5531 1462 5543
rect 1508 5577 1562 5683
rect 1608 5717 1662 5729
rect 1608 5691 1618 5717
rect 1652 5691 1662 5717
rect 1608 5639 1609 5691
rect 1661 5639 1662 5691
rect 1608 5632 1662 5639
rect 1708 5717 1762 5823
rect 1808 5901 1862 5908
rect 1808 5849 1809 5901
rect 1861 5849 1862 5901
rect 1808 5823 1818 5849
rect 1852 5823 1862 5849
rect 1808 5811 1862 5823
rect 1908 5857 1962 5963
rect 2008 5997 2062 6009
rect 2008 5971 2018 5997
rect 2052 5971 2062 5997
rect 2008 5919 2009 5971
rect 2061 5919 2062 5971
rect 2008 5912 2062 5919
rect 2108 5997 2162 6103
rect 2208 6181 2262 6188
rect 2208 6129 2209 6181
rect 2261 6129 2262 6181
rect 2208 6103 2218 6129
rect 2252 6103 2262 6129
rect 2208 6091 2262 6103
rect 2308 6137 2362 6333
rect 2408 6367 2462 6379
rect 2408 6341 2418 6367
rect 2452 6341 2462 6367
rect 2408 6289 2409 6341
rect 2461 6289 2462 6341
rect 2408 6282 2462 6289
rect 2508 6367 2562 6473
rect 2608 6551 2662 6558
rect 2608 6499 2609 6551
rect 2661 6499 2662 6551
rect 2608 6473 2618 6499
rect 2652 6473 2662 6499
rect 2608 6461 2662 6473
rect 2708 6507 2762 6613
rect 2808 6647 2862 6659
rect 2808 6621 2818 6647
rect 2852 6621 2862 6647
rect 2808 6569 2809 6621
rect 2861 6569 2862 6621
rect 2808 6562 2862 6569
rect 2908 6647 2962 6753
rect 3008 6831 3062 6838
rect 3008 6779 3009 6831
rect 3061 6779 3062 6831
rect 3008 6753 3018 6779
rect 3052 6753 3062 6779
rect 3008 6741 3062 6753
rect 3108 6787 3162 6893
rect 3208 6927 3262 6939
rect 3208 6901 3218 6927
rect 3252 6901 3262 6927
rect 3208 6849 3209 6901
rect 3261 6849 3262 6901
rect 3208 6842 3262 6849
rect 3308 6927 3362 7033
rect 3408 7111 3462 7118
rect 3408 7059 3409 7111
rect 3461 7059 3462 7111
rect 3408 7033 3418 7059
rect 3452 7033 3462 7059
rect 3408 7021 3462 7033
rect 3508 7067 3562 7173
rect 3608 7207 3662 7219
rect 3608 7181 3618 7207
rect 3652 7181 3662 7207
rect 3608 7129 3609 7181
rect 3661 7129 3662 7181
rect 3608 7122 3662 7129
rect 3708 7207 3762 7313
rect 3808 7391 3862 7398
rect 3808 7339 3809 7391
rect 3861 7339 3862 7391
rect 3808 7313 3818 7339
rect 3852 7313 3862 7339
rect 3808 7301 3862 7313
rect 3908 7347 3962 7543
rect 4008 7577 4062 7589
rect 4008 7551 4018 7577
rect 4052 7551 4062 7577
rect 4008 7499 4009 7551
rect 4061 7499 4062 7551
rect 4008 7492 4062 7499
rect 4108 7577 4162 7683
rect 4208 7761 4262 7768
rect 4208 7709 4209 7761
rect 4261 7709 4262 7761
rect 4208 7683 4218 7709
rect 4252 7683 4262 7709
rect 4208 7671 4262 7683
rect 4308 7717 4362 7823
rect 4408 7857 4462 7869
rect 4408 7831 4418 7857
rect 4452 7831 4462 7857
rect 4408 7779 4409 7831
rect 4461 7779 4462 7831
rect 4408 7772 4462 7779
rect 4508 7857 4562 7963
rect 4608 8041 4662 8048
rect 4608 7989 4609 8041
rect 4661 7989 4662 8041
rect 4608 7963 4618 7989
rect 4652 7963 4662 7989
rect 4608 7951 4662 7963
rect 4708 7997 4762 8103
rect 4808 8137 4862 8149
rect 4808 8111 4818 8137
rect 4852 8111 4862 8137
rect 4808 8059 4809 8111
rect 4861 8059 4862 8111
rect 4808 8052 4862 8059
rect 4908 8137 4962 8243
rect 5008 8321 5062 8328
rect 5008 8269 5009 8321
rect 5061 8269 5062 8321
rect 5008 8243 5018 8269
rect 5052 8243 5062 8269
rect 5008 8231 5062 8243
rect 5108 8277 5162 8383
rect 5208 8417 5262 8429
rect 5208 8391 5218 8417
rect 5252 8391 5262 8417
rect 5208 8339 5209 8391
rect 5261 8339 5262 8391
rect 5208 8332 5262 8339
rect 5308 8417 5362 8523
rect 5408 8601 5462 8608
rect 5408 8549 5409 8601
rect 5461 8549 5462 8601
rect 5408 8523 5418 8549
rect 5452 8523 5462 8549
rect 5408 8511 5462 8523
rect 5508 8557 5562 8753
rect 5608 8787 5662 8799
rect 5608 8761 5618 8787
rect 5652 8761 5662 8787
rect 5608 8709 5609 8761
rect 5661 8709 5662 8761
rect 5608 8702 5662 8709
rect 5708 8787 5762 8893
rect 5808 8971 5862 8978
rect 5808 8919 5809 8971
rect 5861 8919 5862 8971
rect 5808 8893 5818 8919
rect 5852 8893 5862 8919
rect 5808 8881 5862 8893
rect 5908 8927 5962 9033
rect 6008 9067 6062 9079
rect 6008 9041 6018 9067
rect 6052 9041 6062 9067
rect 6008 8989 6009 9041
rect 6061 8989 6062 9041
rect 6008 8982 6062 8989
rect 6108 9067 6162 9173
rect 6208 9251 6262 9258
rect 6208 9199 6209 9251
rect 6261 9199 6262 9251
rect 6208 9173 6218 9199
rect 6252 9173 6262 9199
rect 6208 9161 6262 9173
rect 6308 9207 6362 9313
rect 6408 9347 6462 9359
rect 6408 9321 6418 9347
rect 6452 9321 6462 9347
rect 6408 9269 6409 9321
rect 6461 9269 6462 9321
rect 6408 9262 6462 9269
rect 6506 9328 6516 9362
rect 6550 9328 6560 9362
rect 6506 9321 6560 9328
rect 6506 9269 6507 9321
rect 6559 9269 6560 9321
rect 6506 9262 6560 9269
rect 6506 9222 6560 9234
rect 6308 9173 6318 9207
rect 6352 9173 6362 9207
rect 6108 9033 6118 9067
rect 6152 9033 6162 9067
rect 5908 8893 5918 8927
rect 5952 8893 5962 8927
rect 5708 8753 5718 8787
rect 5752 8753 5762 8787
rect 5602 8673 5668 8674
rect 5602 8621 5609 8673
rect 5661 8621 5668 8673
rect 5602 8620 5668 8621
rect 5508 8523 5518 8557
rect 5552 8523 5562 8557
rect 5308 8383 5318 8417
rect 5352 8383 5362 8417
rect 5108 8243 5118 8277
rect 5152 8243 5162 8277
rect 4908 8103 4918 8137
rect 4952 8103 4962 8137
rect 4708 7963 4718 7997
rect 4752 7963 4762 7997
rect 4508 7823 4518 7857
rect 4552 7823 4562 7857
rect 4308 7683 4318 7717
rect 4352 7683 4362 7717
rect 4108 7543 4118 7577
rect 4152 7543 4162 7577
rect 4002 7463 4068 7464
rect 4002 7411 4009 7463
rect 4061 7411 4068 7463
rect 4002 7410 4068 7411
rect 3908 7313 3918 7347
rect 3952 7313 3962 7347
rect 3708 7173 3718 7207
rect 3752 7173 3762 7207
rect 3508 7033 3518 7067
rect 3552 7033 3562 7067
rect 3308 6893 3318 6927
rect 3352 6893 3362 6927
rect 3108 6753 3118 6787
rect 3152 6753 3162 6787
rect 2908 6613 2918 6647
rect 2952 6613 2962 6647
rect 2708 6473 2718 6507
rect 2752 6473 2762 6507
rect 2508 6333 2518 6367
rect 2552 6333 2562 6367
rect 2402 6253 2468 6254
rect 2402 6201 2409 6253
rect 2461 6201 2468 6253
rect 2402 6200 2468 6201
rect 2308 6103 2318 6137
rect 2352 6103 2362 6137
rect 2108 5963 2118 5997
rect 2152 5963 2162 5997
rect 1908 5823 1918 5857
rect 1952 5823 1962 5857
rect 1708 5683 1718 5717
rect 1752 5683 1762 5717
rect 1508 5543 1518 5577
rect 1552 5543 1562 5577
rect 1308 5403 1318 5437
rect 1352 5403 1362 5437
rect 1108 5263 1118 5297
rect 1152 5263 1162 5297
rect 908 5123 918 5157
rect 952 5123 962 5157
rect 908 5040 962 5123
rect 1008 5201 1062 5208
rect 1008 5149 1009 5201
rect 1061 5149 1062 5201
rect 1008 5123 1018 5149
rect 1052 5123 1062 5149
rect 1008 5111 1062 5123
rect 1108 5157 1162 5263
rect 1208 5297 1262 5309
rect 1208 5271 1218 5297
rect 1252 5271 1262 5297
rect 1208 5219 1209 5271
rect 1261 5219 1262 5271
rect 1208 5212 1262 5219
rect 1308 5297 1362 5403
rect 1408 5481 1462 5488
rect 1408 5429 1409 5481
rect 1461 5429 1462 5481
rect 1408 5403 1418 5429
rect 1452 5403 1462 5429
rect 1408 5391 1462 5403
rect 1508 5437 1562 5543
rect 1608 5577 1662 5589
rect 1608 5551 1618 5577
rect 1652 5551 1662 5577
rect 1608 5499 1609 5551
rect 1661 5499 1662 5551
rect 1608 5492 1662 5499
rect 1708 5577 1762 5683
rect 1808 5761 1862 5768
rect 1808 5709 1809 5761
rect 1861 5709 1862 5761
rect 1808 5683 1818 5709
rect 1852 5683 1862 5709
rect 1808 5671 1862 5683
rect 1908 5717 1962 5823
rect 2008 5857 2062 5869
rect 2008 5831 2018 5857
rect 2052 5831 2062 5857
rect 2008 5779 2009 5831
rect 2061 5779 2062 5831
rect 2008 5772 2062 5779
rect 2108 5857 2162 5963
rect 2208 6041 2262 6048
rect 2208 5989 2209 6041
rect 2261 5989 2262 6041
rect 2208 5963 2218 5989
rect 2252 5963 2262 5989
rect 2208 5951 2262 5963
rect 2308 5997 2362 6103
rect 2408 6137 2462 6149
rect 2408 6111 2418 6137
rect 2452 6111 2462 6137
rect 2408 6059 2409 6111
rect 2461 6059 2462 6111
rect 2408 6052 2462 6059
rect 2508 6137 2562 6333
rect 2608 6411 2662 6418
rect 2608 6359 2609 6411
rect 2661 6359 2662 6411
rect 2608 6333 2618 6359
rect 2652 6333 2662 6359
rect 2608 6321 2662 6333
rect 2708 6367 2762 6473
rect 2808 6507 2862 6519
rect 2808 6481 2818 6507
rect 2852 6481 2862 6507
rect 2808 6429 2809 6481
rect 2861 6429 2862 6481
rect 2808 6422 2862 6429
rect 2908 6507 2962 6613
rect 3008 6691 3062 6698
rect 3008 6639 3009 6691
rect 3061 6639 3062 6691
rect 3008 6613 3018 6639
rect 3052 6613 3062 6639
rect 3008 6601 3062 6613
rect 3108 6647 3162 6753
rect 3208 6787 3262 6799
rect 3208 6761 3218 6787
rect 3252 6761 3262 6787
rect 3208 6709 3209 6761
rect 3261 6709 3262 6761
rect 3208 6702 3262 6709
rect 3308 6787 3362 6893
rect 3408 6971 3462 6978
rect 3408 6919 3409 6971
rect 3461 6919 3462 6971
rect 3408 6893 3418 6919
rect 3452 6893 3462 6919
rect 3408 6881 3462 6893
rect 3508 6927 3562 7033
rect 3608 7067 3662 7079
rect 3608 7041 3618 7067
rect 3652 7041 3662 7067
rect 3608 6989 3609 7041
rect 3661 6989 3662 7041
rect 3608 6982 3662 6989
rect 3708 7067 3762 7173
rect 3808 7251 3862 7258
rect 3808 7199 3809 7251
rect 3861 7199 3862 7251
rect 3808 7173 3818 7199
rect 3852 7173 3862 7199
rect 3808 7161 3862 7173
rect 3908 7207 3962 7313
rect 4008 7347 4062 7359
rect 4008 7321 4018 7347
rect 4052 7321 4062 7347
rect 4008 7269 4009 7321
rect 4061 7269 4062 7321
rect 4008 7262 4062 7269
rect 4108 7347 4162 7543
rect 4208 7621 4262 7628
rect 4208 7569 4209 7621
rect 4261 7569 4262 7621
rect 4208 7543 4218 7569
rect 4252 7543 4262 7569
rect 4208 7531 4262 7543
rect 4308 7577 4362 7683
rect 4408 7717 4462 7729
rect 4408 7691 4418 7717
rect 4452 7691 4462 7717
rect 4408 7639 4409 7691
rect 4461 7639 4462 7691
rect 4408 7632 4462 7639
rect 4508 7717 4562 7823
rect 4608 7901 4662 7908
rect 4608 7849 4609 7901
rect 4661 7849 4662 7901
rect 4608 7823 4618 7849
rect 4652 7823 4662 7849
rect 4608 7811 4662 7823
rect 4708 7857 4762 7963
rect 4808 7997 4862 8009
rect 4808 7971 4818 7997
rect 4852 7971 4862 7997
rect 4808 7919 4809 7971
rect 4861 7919 4862 7971
rect 4808 7912 4862 7919
rect 4908 7997 4962 8103
rect 5008 8181 5062 8188
rect 5008 8129 5009 8181
rect 5061 8129 5062 8181
rect 5008 8103 5018 8129
rect 5052 8103 5062 8129
rect 5008 8091 5062 8103
rect 5108 8137 5162 8243
rect 5208 8277 5262 8289
rect 5208 8251 5218 8277
rect 5252 8251 5262 8277
rect 5208 8199 5209 8251
rect 5261 8199 5262 8251
rect 5208 8192 5262 8199
rect 5308 8277 5362 8383
rect 5408 8461 5462 8468
rect 5408 8409 5409 8461
rect 5461 8409 5462 8461
rect 5408 8383 5418 8409
rect 5452 8383 5462 8409
rect 5408 8371 5462 8383
rect 5508 8417 5562 8523
rect 5608 8557 5662 8569
rect 5608 8531 5618 8557
rect 5652 8531 5662 8557
rect 5608 8479 5609 8531
rect 5661 8479 5662 8531
rect 5608 8472 5662 8479
rect 5708 8557 5762 8753
rect 5808 8831 5862 8838
rect 5808 8779 5809 8831
rect 5861 8779 5862 8831
rect 5808 8753 5818 8779
rect 5852 8753 5862 8779
rect 5808 8741 5862 8753
rect 5908 8787 5962 8893
rect 6008 8927 6062 8939
rect 6008 8901 6018 8927
rect 6052 8901 6062 8927
rect 6008 8849 6009 8901
rect 6061 8849 6062 8901
rect 6008 8842 6062 8849
rect 6108 8927 6162 9033
rect 6208 9111 6262 9118
rect 6208 9059 6209 9111
rect 6261 9059 6262 9111
rect 6208 9033 6218 9059
rect 6252 9033 6262 9059
rect 6208 9021 6262 9033
rect 6308 9067 6362 9173
rect 6408 9207 6462 9219
rect 6408 9181 6418 9207
rect 6452 9181 6462 9207
rect 6408 9129 6409 9181
rect 6461 9129 6462 9181
rect 6408 9122 6462 9129
rect 6506 9188 6516 9222
rect 6550 9188 6560 9222
rect 6506 9181 6560 9188
rect 6506 9129 6507 9181
rect 6559 9129 6560 9181
rect 6506 9122 6560 9129
rect 6506 9082 6560 9094
rect 6308 9033 6318 9067
rect 6352 9033 6362 9067
rect 6108 8893 6118 8927
rect 6152 8893 6162 8927
rect 5908 8753 5918 8787
rect 5952 8753 5962 8787
rect 5802 8689 5868 8690
rect 5802 8637 5809 8689
rect 5861 8637 5868 8689
rect 5802 8636 5868 8637
rect 5708 8523 5718 8557
rect 5752 8523 5762 8557
rect 5508 8383 5518 8417
rect 5552 8383 5562 8417
rect 5308 8243 5318 8277
rect 5352 8243 5362 8277
rect 5108 8103 5118 8137
rect 5152 8103 5162 8137
rect 4908 7963 4918 7997
rect 4952 7963 4962 7997
rect 4708 7823 4718 7857
rect 4752 7823 4762 7857
rect 4508 7683 4518 7717
rect 4552 7683 4562 7717
rect 4308 7543 4318 7577
rect 4352 7543 4362 7577
rect 4202 7479 4268 7480
rect 4202 7427 4209 7479
rect 4261 7427 4268 7479
rect 4202 7426 4268 7427
rect 4108 7313 4118 7347
rect 4152 7313 4162 7347
rect 3908 7173 3918 7207
rect 3952 7173 3962 7207
rect 3708 7033 3718 7067
rect 3752 7033 3762 7067
rect 3508 6893 3518 6927
rect 3552 6893 3562 6927
rect 3308 6753 3318 6787
rect 3352 6753 3362 6787
rect 3108 6613 3118 6647
rect 3152 6613 3162 6647
rect 2908 6473 2918 6507
rect 2952 6473 2962 6507
rect 2708 6333 2718 6367
rect 2752 6333 2762 6367
rect 2602 6269 2668 6270
rect 2602 6217 2609 6269
rect 2661 6217 2668 6269
rect 2602 6216 2668 6217
rect 2508 6103 2518 6137
rect 2552 6103 2562 6137
rect 2308 5963 2318 5997
rect 2352 5963 2362 5997
rect 2108 5823 2118 5857
rect 2152 5823 2162 5857
rect 1908 5683 1918 5717
rect 1952 5683 1962 5717
rect 1708 5543 1718 5577
rect 1752 5543 1762 5577
rect 1508 5403 1518 5437
rect 1552 5403 1562 5437
rect 1308 5263 1318 5297
rect 1352 5263 1362 5297
rect 1108 5123 1118 5157
rect 1152 5123 1162 5157
rect 1108 5040 1162 5123
rect 1208 5157 1262 5169
rect 1208 5131 1218 5157
rect 1252 5131 1262 5157
rect 1208 5079 1209 5131
rect 1261 5079 1262 5131
rect 1208 5072 1262 5079
rect 1308 5157 1362 5263
rect 1408 5341 1462 5348
rect 1408 5289 1409 5341
rect 1461 5289 1462 5341
rect 1408 5263 1418 5289
rect 1452 5263 1462 5289
rect 1408 5251 1462 5263
rect 1508 5297 1562 5403
rect 1608 5437 1662 5449
rect 1608 5411 1618 5437
rect 1652 5411 1662 5437
rect 1608 5359 1609 5411
rect 1661 5359 1662 5411
rect 1608 5352 1662 5359
rect 1708 5437 1762 5543
rect 1808 5621 1862 5628
rect 1808 5569 1809 5621
rect 1861 5569 1862 5621
rect 1808 5543 1818 5569
rect 1852 5543 1862 5569
rect 1808 5531 1862 5543
rect 1908 5577 1962 5683
rect 2008 5717 2062 5729
rect 2008 5691 2018 5717
rect 2052 5691 2062 5717
rect 2008 5639 2009 5691
rect 2061 5639 2062 5691
rect 2008 5632 2062 5639
rect 2108 5717 2162 5823
rect 2208 5901 2262 5908
rect 2208 5849 2209 5901
rect 2261 5849 2262 5901
rect 2208 5823 2218 5849
rect 2252 5823 2262 5849
rect 2208 5811 2262 5823
rect 2308 5857 2362 5963
rect 2408 5997 2462 6009
rect 2408 5971 2418 5997
rect 2452 5971 2462 5997
rect 2408 5919 2409 5971
rect 2461 5919 2462 5971
rect 2408 5912 2462 5919
rect 2508 5997 2562 6103
rect 2608 6181 2662 6188
rect 2608 6129 2609 6181
rect 2661 6129 2662 6181
rect 2608 6103 2618 6129
rect 2652 6103 2662 6129
rect 2608 6091 2662 6103
rect 2708 6137 2762 6333
rect 2808 6367 2862 6379
rect 2808 6341 2818 6367
rect 2852 6341 2862 6367
rect 2808 6289 2809 6341
rect 2861 6289 2862 6341
rect 2808 6282 2862 6289
rect 2908 6367 2962 6473
rect 3008 6551 3062 6558
rect 3008 6499 3009 6551
rect 3061 6499 3062 6551
rect 3008 6473 3018 6499
rect 3052 6473 3062 6499
rect 3008 6461 3062 6473
rect 3108 6507 3162 6613
rect 3208 6647 3262 6659
rect 3208 6621 3218 6647
rect 3252 6621 3262 6647
rect 3208 6569 3209 6621
rect 3261 6569 3262 6621
rect 3208 6562 3262 6569
rect 3308 6647 3362 6753
rect 3408 6831 3462 6838
rect 3408 6779 3409 6831
rect 3461 6779 3462 6831
rect 3408 6753 3418 6779
rect 3452 6753 3462 6779
rect 3408 6741 3462 6753
rect 3508 6787 3562 6893
rect 3608 6927 3662 6939
rect 3608 6901 3618 6927
rect 3652 6901 3662 6927
rect 3608 6849 3609 6901
rect 3661 6849 3662 6901
rect 3608 6842 3662 6849
rect 3708 6927 3762 7033
rect 3808 7111 3862 7118
rect 3808 7059 3809 7111
rect 3861 7059 3862 7111
rect 3808 7033 3818 7059
rect 3852 7033 3862 7059
rect 3808 7021 3862 7033
rect 3908 7067 3962 7173
rect 4008 7207 4062 7219
rect 4008 7181 4018 7207
rect 4052 7181 4062 7207
rect 4008 7129 4009 7181
rect 4061 7129 4062 7181
rect 4008 7122 4062 7129
rect 4108 7207 4162 7313
rect 4208 7391 4262 7398
rect 4208 7339 4209 7391
rect 4261 7339 4262 7391
rect 4208 7313 4218 7339
rect 4252 7313 4262 7339
rect 4208 7301 4262 7313
rect 4308 7347 4362 7543
rect 4408 7577 4462 7589
rect 4408 7551 4418 7577
rect 4452 7551 4462 7577
rect 4408 7499 4409 7551
rect 4461 7499 4462 7551
rect 4408 7492 4462 7499
rect 4508 7577 4562 7683
rect 4608 7761 4662 7768
rect 4608 7709 4609 7761
rect 4661 7709 4662 7761
rect 4608 7683 4618 7709
rect 4652 7683 4662 7709
rect 4608 7671 4662 7683
rect 4708 7717 4762 7823
rect 4808 7857 4862 7869
rect 4808 7831 4818 7857
rect 4852 7831 4862 7857
rect 4808 7779 4809 7831
rect 4861 7779 4862 7831
rect 4808 7772 4862 7779
rect 4908 7857 4962 7963
rect 5008 8041 5062 8048
rect 5008 7989 5009 8041
rect 5061 7989 5062 8041
rect 5008 7963 5018 7989
rect 5052 7963 5062 7989
rect 5008 7951 5062 7963
rect 5108 7997 5162 8103
rect 5208 8137 5262 8149
rect 5208 8111 5218 8137
rect 5252 8111 5262 8137
rect 5208 8059 5209 8111
rect 5261 8059 5262 8111
rect 5208 8052 5262 8059
rect 5308 8137 5362 8243
rect 5408 8321 5462 8328
rect 5408 8269 5409 8321
rect 5461 8269 5462 8321
rect 5408 8243 5418 8269
rect 5452 8243 5462 8269
rect 5408 8231 5462 8243
rect 5508 8277 5562 8383
rect 5608 8417 5662 8429
rect 5608 8391 5618 8417
rect 5652 8391 5662 8417
rect 5608 8339 5609 8391
rect 5661 8339 5662 8391
rect 5608 8332 5662 8339
rect 5708 8417 5762 8523
rect 5808 8601 5862 8608
rect 5808 8549 5809 8601
rect 5861 8549 5862 8601
rect 5808 8523 5818 8549
rect 5852 8523 5862 8549
rect 5808 8511 5862 8523
rect 5908 8557 5962 8753
rect 6008 8787 6062 8799
rect 6008 8761 6018 8787
rect 6052 8761 6062 8787
rect 6008 8709 6009 8761
rect 6061 8709 6062 8761
rect 6008 8702 6062 8709
rect 6108 8787 6162 8893
rect 6208 8971 6262 8978
rect 6208 8919 6209 8971
rect 6261 8919 6262 8971
rect 6208 8893 6218 8919
rect 6252 8893 6262 8919
rect 6208 8881 6262 8893
rect 6308 8927 6362 9033
rect 6408 9067 6462 9079
rect 6408 9041 6418 9067
rect 6452 9041 6462 9067
rect 6408 8989 6409 9041
rect 6461 8989 6462 9041
rect 6408 8982 6462 8989
rect 6506 9048 6516 9082
rect 6550 9048 6560 9082
rect 6506 9041 6560 9048
rect 6506 8989 6507 9041
rect 6559 8989 6560 9041
rect 6506 8982 6560 8989
rect 6506 8942 6560 8954
rect 6308 8893 6318 8927
rect 6352 8893 6362 8927
rect 6108 8753 6118 8787
rect 6152 8753 6162 8787
rect 6002 8673 6068 8674
rect 6002 8621 6009 8673
rect 6061 8621 6068 8673
rect 6002 8620 6068 8621
rect 5908 8523 5918 8557
rect 5952 8523 5962 8557
rect 5708 8383 5718 8417
rect 5752 8383 5762 8417
rect 5508 8243 5518 8277
rect 5552 8243 5562 8277
rect 5308 8103 5318 8137
rect 5352 8103 5362 8137
rect 5108 7963 5118 7997
rect 5152 7963 5162 7997
rect 4908 7823 4918 7857
rect 4952 7823 4962 7857
rect 4708 7683 4718 7717
rect 4752 7683 4762 7717
rect 4508 7543 4518 7577
rect 4552 7543 4562 7577
rect 4402 7463 4468 7464
rect 4402 7411 4409 7463
rect 4461 7411 4468 7463
rect 4402 7410 4468 7411
rect 4308 7313 4318 7347
rect 4352 7313 4362 7347
rect 4108 7173 4118 7207
rect 4152 7173 4162 7207
rect 3908 7033 3918 7067
rect 3952 7033 3962 7067
rect 3708 6893 3718 6927
rect 3752 6893 3762 6927
rect 3508 6753 3518 6787
rect 3552 6753 3562 6787
rect 3308 6613 3318 6647
rect 3352 6613 3362 6647
rect 3108 6473 3118 6507
rect 3152 6473 3162 6507
rect 2908 6333 2918 6367
rect 2952 6333 2962 6367
rect 2802 6253 2868 6254
rect 2802 6201 2809 6253
rect 2861 6201 2868 6253
rect 2802 6200 2868 6201
rect 2708 6103 2718 6137
rect 2752 6103 2762 6137
rect 2508 5963 2518 5997
rect 2552 5963 2562 5997
rect 2308 5823 2318 5857
rect 2352 5823 2362 5857
rect 2108 5683 2118 5717
rect 2152 5683 2162 5717
rect 1908 5543 1918 5577
rect 1952 5543 1962 5577
rect 1708 5403 1718 5437
rect 1752 5403 1762 5437
rect 1508 5263 1518 5297
rect 1552 5263 1562 5297
rect 1308 5123 1318 5157
rect 1352 5123 1362 5157
rect 1308 5040 1362 5123
rect 1408 5201 1462 5208
rect 1408 5149 1409 5201
rect 1461 5149 1462 5201
rect 1408 5123 1418 5149
rect 1452 5123 1462 5149
rect 1408 5111 1462 5123
rect 1508 5157 1562 5263
rect 1608 5297 1662 5309
rect 1608 5271 1618 5297
rect 1652 5271 1662 5297
rect 1608 5219 1609 5271
rect 1661 5219 1662 5271
rect 1608 5212 1662 5219
rect 1708 5297 1762 5403
rect 1808 5481 1862 5488
rect 1808 5429 1809 5481
rect 1861 5429 1862 5481
rect 1808 5403 1818 5429
rect 1852 5403 1862 5429
rect 1808 5391 1862 5403
rect 1908 5437 1962 5543
rect 2008 5577 2062 5589
rect 2008 5551 2018 5577
rect 2052 5551 2062 5577
rect 2008 5499 2009 5551
rect 2061 5499 2062 5551
rect 2008 5492 2062 5499
rect 2108 5577 2162 5683
rect 2208 5761 2262 5768
rect 2208 5709 2209 5761
rect 2261 5709 2262 5761
rect 2208 5683 2218 5709
rect 2252 5683 2262 5709
rect 2208 5671 2262 5683
rect 2308 5717 2362 5823
rect 2408 5857 2462 5869
rect 2408 5831 2418 5857
rect 2452 5831 2462 5857
rect 2408 5779 2409 5831
rect 2461 5779 2462 5831
rect 2408 5772 2462 5779
rect 2508 5857 2562 5963
rect 2608 6041 2662 6048
rect 2608 5989 2609 6041
rect 2661 5989 2662 6041
rect 2608 5963 2618 5989
rect 2652 5963 2662 5989
rect 2608 5951 2662 5963
rect 2708 5997 2762 6103
rect 2808 6137 2862 6149
rect 2808 6111 2818 6137
rect 2852 6111 2862 6137
rect 2808 6059 2809 6111
rect 2861 6059 2862 6111
rect 2808 6052 2862 6059
rect 2908 6137 2962 6333
rect 3008 6411 3062 6418
rect 3008 6359 3009 6411
rect 3061 6359 3062 6411
rect 3008 6333 3018 6359
rect 3052 6333 3062 6359
rect 3008 6321 3062 6333
rect 3108 6367 3162 6473
rect 3208 6507 3262 6519
rect 3208 6481 3218 6507
rect 3252 6481 3262 6507
rect 3208 6429 3209 6481
rect 3261 6429 3262 6481
rect 3208 6422 3262 6429
rect 3308 6507 3362 6613
rect 3408 6691 3462 6698
rect 3408 6639 3409 6691
rect 3461 6639 3462 6691
rect 3408 6613 3418 6639
rect 3452 6613 3462 6639
rect 3408 6601 3462 6613
rect 3508 6647 3562 6753
rect 3608 6787 3662 6799
rect 3608 6761 3618 6787
rect 3652 6761 3662 6787
rect 3608 6709 3609 6761
rect 3661 6709 3662 6761
rect 3608 6702 3662 6709
rect 3708 6787 3762 6893
rect 3808 6971 3862 6978
rect 3808 6919 3809 6971
rect 3861 6919 3862 6971
rect 3808 6893 3818 6919
rect 3852 6893 3862 6919
rect 3808 6881 3862 6893
rect 3908 6927 3962 7033
rect 4008 7067 4062 7079
rect 4008 7041 4018 7067
rect 4052 7041 4062 7067
rect 4008 6989 4009 7041
rect 4061 6989 4062 7041
rect 4008 6982 4062 6989
rect 4108 7067 4162 7173
rect 4208 7251 4262 7258
rect 4208 7199 4209 7251
rect 4261 7199 4262 7251
rect 4208 7173 4218 7199
rect 4252 7173 4262 7199
rect 4208 7161 4262 7173
rect 4308 7207 4362 7313
rect 4408 7347 4462 7359
rect 4408 7321 4418 7347
rect 4452 7321 4462 7347
rect 4408 7269 4409 7321
rect 4461 7269 4462 7321
rect 4408 7262 4462 7269
rect 4508 7347 4562 7543
rect 4608 7621 4662 7628
rect 4608 7569 4609 7621
rect 4661 7569 4662 7621
rect 4608 7543 4618 7569
rect 4652 7543 4662 7569
rect 4608 7531 4662 7543
rect 4708 7577 4762 7683
rect 4808 7717 4862 7729
rect 4808 7691 4818 7717
rect 4852 7691 4862 7717
rect 4808 7639 4809 7691
rect 4861 7639 4862 7691
rect 4808 7632 4862 7639
rect 4908 7717 4962 7823
rect 5008 7901 5062 7908
rect 5008 7849 5009 7901
rect 5061 7849 5062 7901
rect 5008 7823 5018 7849
rect 5052 7823 5062 7849
rect 5008 7811 5062 7823
rect 5108 7857 5162 7963
rect 5208 7997 5262 8009
rect 5208 7971 5218 7997
rect 5252 7971 5262 7997
rect 5208 7919 5209 7971
rect 5261 7919 5262 7971
rect 5208 7912 5262 7919
rect 5308 7997 5362 8103
rect 5408 8181 5462 8188
rect 5408 8129 5409 8181
rect 5461 8129 5462 8181
rect 5408 8103 5418 8129
rect 5452 8103 5462 8129
rect 5408 8091 5462 8103
rect 5508 8137 5562 8243
rect 5608 8277 5662 8289
rect 5608 8251 5618 8277
rect 5652 8251 5662 8277
rect 5608 8199 5609 8251
rect 5661 8199 5662 8251
rect 5608 8192 5662 8199
rect 5708 8277 5762 8383
rect 5808 8461 5862 8468
rect 5808 8409 5809 8461
rect 5861 8409 5862 8461
rect 5808 8383 5818 8409
rect 5852 8383 5862 8409
rect 5808 8371 5862 8383
rect 5908 8417 5962 8523
rect 6008 8557 6062 8569
rect 6008 8531 6018 8557
rect 6052 8531 6062 8557
rect 6008 8479 6009 8531
rect 6061 8479 6062 8531
rect 6008 8472 6062 8479
rect 6108 8557 6162 8753
rect 6208 8831 6262 8838
rect 6208 8779 6209 8831
rect 6261 8779 6262 8831
rect 6208 8753 6218 8779
rect 6252 8753 6262 8779
rect 6208 8741 6262 8753
rect 6308 8787 6362 8893
rect 6408 8927 6462 8939
rect 6408 8901 6418 8927
rect 6452 8901 6462 8927
rect 6408 8849 6409 8901
rect 6461 8849 6462 8901
rect 6408 8842 6462 8849
rect 6506 8908 6516 8942
rect 6550 8908 6560 8942
rect 6506 8901 6560 8908
rect 6506 8849 6507 8901
rect 6559 8849 6560 8901
rect 6506 8842 6560 8849
rect 6506 8802 6560 8814
rect 6308 8753 6318 8787
rect 6352 8753 6362 8787
rect 6202 8689 6268 8690
rect 6202 8637 6209 8689
rect 6261 8637 6268 8689
rect 6202 8636 6268 8637
rect 6108 8523 6118 8557
rect 6152 8523 6162 8557
rect 5908 8383 5918 8417
rect 5952 8383 5962 8417
rect 5708 8243 5718 8277
rect 5752 8243 5762 8277
rect 5508 8103 5518 8137
rect 5552 8103 5562 8137
rect 5308 7963 5318 7997
rect 5352 7963 5362 7997
rect 5108 7823 5118 7857
rect 5152 7823 5162 7857
rect 4908 7683 4918 7717
rect 4952 7683 4962 7717
rect 4708 7543 4718 7577
rect 4752 7543 4762 7577
rect 4602 7479 4668 7480
rect 4602 7427 4609 7479
rect 4661 7427 4668 7479
rect 4602 7426 4668 7427
rect 4508 7313 4518 7347
rect 4552 7313 4562 7347
rect 4308 7173 4318 7207
rect 4352 7173 4362 7207
rect 4108 7033 4118 7067
rect 4152 7033 4162 7067
rect 3908 6893 3918 6927
rect 3952 6893 3962 6927
rect 3708 6753 3718 6787
rect 3752 6753 3762 6787
rect 3508 6613 3518 6647
rect 3552 6613 3562 6647
rect 3308 6473 3318 6507
rect 3352 6473 3362 6507
rect 3108 6333 3118 6367
rect 3152 6333 3162 6367
rect 3002 6269 3068 6270
rect 3002 6217 3009 6269
rect 3061 6217 3068 6269
rect 3002 6216 3068 6217
rect 2908 6103 2918 6137
rect 2952 6103 2962 6137
rect 2708 5963 2718 5997
rect 2752 5963 2762 5997
rect 2508 5823 2518 5857
rect 2552 5823 2562 5857
rect 2308 5683 2318 5717
rect 2352 5683 2362 5717
rect 2108 5543 2118 5577
rect 2152 5543 2162 5577
rect 1908 5403 1918 5437
rect 1952 5403 1962 5437
rect 1708 5263 1718 5297
rect 1752 5263 1762 5297
rect 1508 5123 1518 5157
rect 1552 5123 1562 5157
rect 1508 5040 1562 5123
rect 1608 5157 1662 5169
rect 1608 5131 1618 5157
rect 1652 5131 1662 5157
rect 1608 5079 1609 5131
rect 1661 5079 1662 5131
rect 1608 5072 1662 5079
rect 1708 5157 1762 5263
rect 1808 5341 1862 5348
rect 1808 5289 1809 5341
rect 1861 5289 1862 5341
rect 1808 5263 1818 5289
rect 1852 5263 1862 5289
rect 1808 5251 1862 5263
rect 1908 5297 1962 5403
rect 2008 5437 2062 5449
rect 2008 5411 2018 5437
rect 2052 5411 2062 5437
rect 2008 5359 2009 5411
rect 2061 5359 2062 5411
rect 2008 5352 2062 5359
rect 2108 5437 2162 5543
rect 2208 5621 2262 5628
rect 2208 5569 2209 5621
rect 2261 5569 2262 5621
rect 2208 5543 2218 5569
rect 2252 5543 2262 5569
rect 2208 5531 2262 5543
rect 2308 5577 2362 5683
rect 2408 5717 2462 5729
rect 2408 5691 2418 5717
rect 2452 5691 2462 5717
rect 2408 5639 2409 5691
rect 2461 5639 2462 5691
rect 2408 5632 2462 5639
rect 2508 5717 2562 5823
rect 2608 5901 2662 5908
rect 2608 5849 2609 5901
rect 2661 5849 2662 5901
rect 2608 5823 2618 5849
rect 2652 5823 2662 5849
rect 2608 5811 2662 5823
rect 2708 5857 2762 5963
rect 2808 5997 2862 6009
rect 2808 5971 2818 5997
rect 2852 5971 2862 5997
rect 2808 5919 2809 5971
rect 2861 5919 2862 5971
rect 2808 5912 2862 5919
rect 2908 5997 2962 6103
rect 3008 6181 3062 6188
rect 3008 6129 3009 6181
rect 3061 6129 3062 6181
rect 3008 6103 3018 6129
rect 3052 6103 3062 6129
rect 3008 6091 3062 6103
rect 3108 6137 3162 6333
rect 3208 6367 3262 6379
rect 3208 6341 3218 6367
rect 3252 6341 3262 6367
rect 3208 6289 3209 6341
rect 3261 6289 3262 6341
rect 3208 6282 3262 6289
rect 3308 6367 3362 6473
rect 3408 6551 3462 6558
rect 3408 6499 3409 6551
rect 3461 6499 3462 6551
rect 3408 6473 3418 6499
rect 3452 6473 3462 6499
rect 3408 6461 3462 6473
rect 3508 6507 3562 6613
rect 3608 6647 3662 6659
rect 3608 6621 3618 6647
rect 3652 6621 3662 6647
rect 3608 6569 3609 6621
rect 3661 6569 3662 6621
rect 3608 6562 3662 6569
rect 3708 6647 3762 6753
rect 3808 6831 3862 6838
rect 3808 6779 3809 6831
rect 3861 6779 3862 6831
rect 3808 6753 3818 6779
rect 3852 6753 3862 6779
rect 3808 6741 3862 6753
rect 3908 6787 3962 6893
rect 4008 6927 4062 6939
rect 4008 6901 4018 6927
rect 4052 6901 4062 6927
rect 4008 6849 4009 6901
rect 4061 6849 4062 6901
rect 4008 6842 4062 6849
rect 4108 6927 4162 7033
rect 4208 7111 4262 7118
rect 4208 7059 4209 7111
rect 4261 7059 4262 7111
rect 4208 7033 4218 7059
rect 4252 7033 4262 7059
rect 4208 7021 4262 7033
rect 4308 7067 4362 7173
rect 4408 7207 4462 7219
rect 4408 7181 4418 7207
rect 4452 7181 4462 7207
rect 4408 7129 4409 7181
rect 4461 7129 4462 7181
rect 4408 7122 4462 7129
rect 4508 7207 4562 7313
rect 4608 7391 4662 7398
rect 4608 7339 4609 7391
rect 4661 7339 4662 7391
rect 4608 7313 4618 7339
rect 4652 7313 4662 7339
rect 4608 7301 4662 7313
rect 4708 7347 4762 7543
rect 4808 7577 4862 7589
rect 4808 7551 4818 7577
rect 4852 7551 4862 7577
rect 4808 7499 4809 7551
rect 4861 7499 4862 7551
rect 4808 7492 4862 7499
rect 4908 7577 4962 7683
rect 5008 7761 5062 7768
rect 5008 7709 5009 7761
rect 5061 7709 5062 7761
rect 5008 7683 5018 7709
rect 5052 7683 5062 7709
rect 5008 7671 5062 7683
rect 5108 7717 5162 7823
rect 5208 7857 5262 7869
rect 5208 7831 5218 7857
rect 5252 7831 5262 7857
rect 5208 7779 5209 7831
rect 5261 7779 5262 7831
rect 5208 7772 5262 7779
rect 5308 7857 5362 7963
rect 5408 8041 5462 8048
rect 5408 7989 5409 8041
rect 5461 7989 5462 8041
rect 5408 7963 5418 7989
rect 5452 7963 5462 7989
rect 5408 7951 5462 7963
rect 5508 7997 5562 8103
rect 5608 8137 5662 8149
rect 5608 8111 5618 8137
rect 5652 8111 5662 8137
rect 5608 8059 5609 8111
rect 5661 8059 5662 8111
rect 5608 8052 5662 8059
rect 5708 8137 5762 8243
rect 5808 8321 5862 8328
rect 5808 8269 5809 8321
rect 5861 8269 5862 8321
rect 5808 8243 5818 8269
rect 5852 8243 5862 8269
rect 5808 8231 5862 8243
rect 5908 8277 5962 8383
rect 6008 8417 6062 8429
rect 6008 8391 6018 8417
rect 6052 8391 6062 8417
rect 6008 8339 6009 8391
rect 6061 8339 6062 8391
rect 6008 8332 6062 8339
rect 6108 8417 6162 8523
rect 6208 8601 6262 8608
rect 6208 8549 6209 8601
rect 6261 8549 6262 8601
rect 6208 8523 6218 8549
rect 6252 8523 6262 8549
rect 6208 8511 6262 8523
rect 6308 8557 6362 8753
rect 6408 8787 6462 8799
rect 6408 8761 6418 8787
rect 6452 8761 6462 8787
rect 6408 8709 6409 8761
rect 6461 8709 6462 8761
rect 6408 8702 6462 8709
rect 6506 8768 6516 8802
rect 6550 8768 6560 8802
rect 6506 8761 6560 8768
rect 6506 8709 6507 8761
rect 6559 8709 6560 8761
rect 6506 8702 6560 8709
rect 6590 8667 6620 9831
rect 6504 8661 6620 8667
rect 6504 8627 6516 8661
rect 6550 8627 6620 8661
rect 6504 8621 6620 8627
rect 6506 8572 6560 8584
rect 6308 8523 6318 8557
rect 6352 8523 6362 8557
rect 6108 8383 6118 8417
rect 6152 8383 6162 8417
rect 5908 8243 5918 8277
rect 5952 8243 5962 8277
rect 5708 8103 5718 8137
rect 5752 8103 5762 8137
rect 5508 7963 5518 7997
rect 5552 7963 5562 7997
rect 5308 7823 5318 7857
rect 5352 7823 5362 7857
rect 5108 7683 5118 7717
rect 5152 7683 5162 7717
rect 4908 7543 4918 7577
rect 4952 7543 4962 7577
rect 4802 7463 4868 7464
rect 4802 7411 4809 7463
rect 4861 7411 4868 7463
rect 4802 7410 4868 7411
rect 4708 7313 4718 7347
rect 4752 7313 4762 7347
rect 4508 7173 4518 7207
rect 4552 7173 4562 7207
rect 4308 7033 4318 7067
rect 4352 7033 4362 7067
rect 4108 6893 4118 6927
rect 4152 6893 4162 6927
rect 3908 6753 3918 6787
rect 3952 6753 3962 6787
rect 3708 6613 3718 6647
rect 3752 6613 3762 6647
rect 3508 6473 3518 6507
rect 3552 6473 3562 6507
rect 3308 6333 3318 6367
rect 3352 6333 3362 6367
rect 3202 6253 3268 6254
rect 3202 6201 3209 6253
rect 3261 6201 3268 6253
rect 3202 6200 3268 6201
rect 3108 6103 3118 6137
rect 3152 6103 3162 6137
rect 2908 5963 2918 5997
rect 2952 5963 2962 5997
rect 2708 5823 2718 5857
rect 2752 5823 2762 5857
rect 2508 5683 2518 5717
rect 2552 5683 2562 5717
rect 2308 5543 2318 5577
rect 2352 5543 2362 5577
rect 2108 5403 2118 5437
rect 2152 5403 2162 5437
rect 1908 5263 1918 5297
rect 1952 5263 1962 5297
rect 1708 5123 1718 5157
rect 1752 5123 1762 5157
rect 1708 5040 1762 5123
rect 1808 5201 1862 5208
rect 1808 5149 1809 5201
rect 1861 5149 1862 5201
rect 1808 5123 1818 5149
rect 1852 5123 1862 5149
rect 1808 5111 1862 5123
rect 1908 5157 1962 5263
rect 2008 5297 2062 5309
rect 2008 5271 2018 5297
rect 2052 5271 2062 5297
rect 2008 5219 2009 5271
rect 2061 5219 2062 5271
rect 2008 5212 2062 5219
rect 2108 5297 2162 5403
rect 2208 5481 2262 5488
rect 2208 5429 2209 5481
rect 2261 5429 2262 5481
rect 2208 5403 2218 5429
rect 2252 5403 2262 5429
rect 2208 5391 2262 5403
rect 2308 5437 2362 5543
rect 2408 5577 2462 5589
rect 2408 5551 2418 5577
rect 2452 5551 2462 5577
rect 2408 5499 2409 5551
rect 2461 5499 2462 5551
rect 2408 5492 2462 5499
rect 2508 5577 2562 5683
rect 2608 5761 2662 5768
rect 2608 5709 2609 5761
rect 2661 5709 2662 5761
rect 2608 5683 2618 5709
rect 2652 5683 2662 5709
rect 2608 5671 2662 5683
rect 2708 5717 2762 5823
rect 2808 5857 2862 5869
rect 2808 5831 2818 5857
rect 2852 5831 2862 5857
rect 2808 5779 2809 5831
rect 2861 5779 2862 5831
rect 2808 5772 2862 5779
rect 2908 5857 2962 5963
rect 3008 6041 3062 6048
rect 3008 5989 3009 6041
rect 3061 5989 3062 6041
rect 3008 5963 3018 5989
rect 3052 5963 3062 5989
rect 3008 5951 3062 5963
rect 3108 5997 3162 6103
rect 3208 6137 3262 6149
rect 3208 6111 3218 6137
rect 3252 6111 3262 6137
rect 3208 6059 3209 6111
rect 3261 6059 3262 6111
rect 3208 6052 3262 6059
rect 3308 6137 3362 6333
rect 3408 6411 3462 6418
rect 3408 6359 3409 6411
rect 3461 6359 3462 6411
rect 3408 6333 3418 6359
rect 3452 6333 3462 6359
rect 3408 6321 3462 6333
rect 3508 6367 3562 6473
rect 3608 6507 3662 6519
rect 3608 6481 3618 6507
rect 3652 6481 3662 6507
rect 3608 6429 3609 6481
rect 3661 6429 3662 6481
rect 3608 6422 3662 6429
rect 3708 6507 3762 6613
rect 3808 6691 3862 6698
rect 3808 6639 3809 6691
rect 3861 6639 3862 6691
rect 3808 6613 3818 6639
rect 3852 6613 3862 6639
rect 3808 6601 3862 6613
rect 3908 6647 3962 6753
rect 4008 6787 4062 6799
rect 4008 6761 4018 6787
rect 4052 6761 4062 6787
rect 4008 6709 4009 6761
rect 4061 6709 4062 6761
rect 4008 6702 4062 6709
rect 4108 6787 4162 6893
rect 4208 6971 4262 6978
rect 4208 6919 4209 6971
rect 4261 6919 4262 6971
rect 4208 6893 4218 6919
rect 4252 6893 4262 6919
rect 4208 6881 4262 6893
rect 4308 6927 4362 7033
rect 4408 7067 4462 7079
rect 4408 7041 4418 7067
rect 4452 7041 4462 7067
rect 4408 6989 4409 7041
rect 4461 6989 4462 7041
rect 4408 6982 4462 6989
rect 4508 7067 4562 7173
rect 4608 7251 4662 7258
rect 4608 7199 4609 7251
rect 4661 7199 4662 7251
rect 4608 7173 4618 7199
rect 4652 7173 4662 7199
rect 4608 7161 4662 7173
rect 4708 7207 4762 7313
rect 4808 7347 4862 7359
rect 4808 7321 4818 7347
rect 4852 7321 4862 7347
rect 4808 7269 4809 7321
rect 4861 7269 4862 7321
rect 4808 7262 4862 7269
rect 4908 7347 4962 7543
rect 5008 7621 5062 7628
rect 5008 7569 5009 7621
rect 5061 7569 5062 7621
rect 5008 7543 5018 7569
rect 5052 7543 5062 7569
rect 5008 7531 5062 7543
rect 5108 7577 5162 7683
rect 5208 7717 5262 7729
rect 5208 7691 5218 7717
rect 5252 7691 5262 7717
rect 5208 7639 5209 7691
rect 5261 7639 5262 7691
rect 5208 7632 5262 7639
rect 5308 7717 5362 7823
rect 5408 7901 5462 7908
rect 5408 7849 5409 7901
rect 5461 7849 5462 7901
rect 5408 7823 5418 7849
rect 5452 7823 5462 7849
rect 5408 7811 5462 7823
rect 5508 7857 5562 7963
rect 5608 7997 5662 8009
rect 5608 7971 5618 7997
rect 5652 7971 5662 7997
rect 5608 7919 5609 7971
rect 5661 7919 5662 7971
rect 5608 7912 5662 7919
rect 5708 7997 5762 8103
rect 5808 8181 5862 8188
rect 5808 8129 5809 8181
rect 5861 8129 5862 8181
rect 5808 8103 5818 8129
rect 5852 8103 5862 8129
rect 5808 8091 5862 8103
rect 5908 8137 5962 8243
rect 6008 8277 6062 8289
rect 6008 8251 6018 8277
rect 6052 8251 6062 8277
rect 6008 8199 6009 8251
rect 6061 8199 6062 8251
rect 6008 8192 6062 8199
rect 6108 8277 6162 8383
rect 6208 8461 6262 8468
rect 6208 8409 6209 8461
rect 6261 8409 6262 8461
rect 6208 8383 6218 8409
rect 6252 8383 6262 8409
rect 6208 8371 6262 8383
rect 6308 8417 6362 8523
rect 6408 8557 6462 8569
rect 6408 8531 6418 8557
rect 6452 8531 6462 8557
rect 6408 8479 6409 8531
rect 6461 8479 6462 8531
rect 6408 8472 6462 8479
rect 6506 8538 6516 8572
rect 6550 8538 6560 8572
rect 6506 8531 6560 8538
rect 6506 8479 6507 8531
rect 6559 8479 6560 8531
rect 6506 8472 6560 8479
rect 6506 8432 6560 8444
rect 6308 8383 6318 8417
rect 6352 8383 6362 8417
rect 6108 8243 6118 8277
rect 6152 8243 6162 8277
rect 5908 8103 5918 8137
rect 5952 8103 5962 8137
rect 5708 7963 5718 7997
rect 5752 7963 5762 7997
rect 5508 7823 5518 7857
rect 5552 7823 5562 7857
rect 5308 7683 5318 7717
rect 5352 7683 5362 7717
rect 5108 7543 5118 7577
rect 5152 7543 5162 7577
rect 5002 7479 5068 7480
rect 5002 7427 5009 7479
rect 5061 7427 5068 7479
rect 5002 7426 5068 7427
rect 4908 7313 4918 7347
rect 4952 7313 4962 7347
rect 4708 7173 4718 7207
rect 4752 7173 4762 7207
rect 4508 7033 4518 7067
rect 4552 7033 4562 7067
rect 4308 6893 4318 6927
rect 4352 6893 4362 6927
rect 4108 6753 4118 6787
rect 4152 6753 4162 6787
rect 3908 6613 3918 6647
rect 3952 6613 3962 6647
rect 3708 6473 3718 6507
rect 3752 6473 3762 6507
rect 3508 6333 3518 6367
rect 3552 6333 3562 6367
rect 3402 6269 3468 6270
rect 3402 6217 3409 6269
rect 3461 6217 3468 6269
rect 3402 6216 3468 6217
rect 3308 6103 3318 6137
rect 3352 6103 3362 6137
rect 3108 5963 3118 5997
rect 3152 5963 3162 5997
rect 2908 5823 2918 5857
rect 2952 5823 2962 5857
rect 2708 5683 2718 5717
rect 2752 5683 2762 5717
rect 2508 5543 2518 5577
rect 2552 5543 2562 5577
rect 2308 5403 2318 5437
rect 2352 5403 2362 5437
rect 2108 5263 2118 5297
rect 2152 5263 2162 5297
rect 1908 5123 1918 5157
rect 1952 5123 1962 5157
rect 1908 5040 1962 5123
rect 2008 5157 2062 5169
rect 2008 5131 2018 5157
rect 2052 5131 2062 5157
rect 2008 5079 2009 5131
rect 2061 5079 2062 5131
rect 2008 5072 2062 5079
rect 2108 5157 2162 5263
rect 2208 5341 2262 5348
rect 2208 5289 2209 5341
rect 2261 5289 2262 5341
rect 2208 5263 2218 5289
rect 2252 5263 2262 5289
rect 2208 5251 2262 5263
rect 2308 5297 2362 5403
rect 2408 5437 2462 5449
rect 2408 5411 2418 5437
rect 2452 5411 2462 5437
rect 2408 5359 2409 5411
rect 2461 5359 2462 5411
rect 2408 5352 2462 5359
rect 2508 5437 2562 5543
rect 2608 5621 2662 5628
rect 2608 5569 2609 5621
rect 2661 5569 2662 5621
rect 2608 5543 2618 5569
rect 2652 5543 2662 5569
rect 2608 5531 2662 5543
rect 2708 5577 2762 5683
rect 2808 5717 2862 5729
rect 2808 5691 2818 5717
rect 2852 5691 2862 5717
rect 2808 5639 2809 5691
rect 2861 5639 2862 5691
rect 2808 5632 2862 5639
rect 2908 5717 2962 5823
rect 3008 5901 3062 5908
rect 3008 5849 3009 5901
rect 3061 5849 3062 5901
rect 3008 5823 3018 5849
rect 3052 5823 3062 5849
rect 3008 5811 3062 5823
rect 3108 5857 3162 5963
rect 3208 5997 3262 6009
rect 3208 5971 3218 5997
rect 3252 5971 3262 5997
rect 3208 5919 3209 5971
rect 3261 5919 3262 5971
rect 3208 5912 3262 5919
rect 3308 5997 3362 6103
rect 3408 6181 3462 6188
rect 3408 6129 3409 6181
rect 3461 6129 3462 6181
rect 3408 6103 3418 6129
rect 3452 6103 3462 6129
rect 3408 6091 3462 6103
rect 3508 6137 3562 6333
rect 3608 6367 3662 6379
rect 3608 6341 3618 6367
rect 3652 6341 3662 6367
rect 3608 6289 3609 6341
rect 3661 6289 3662 6341
rect 3608 6282 3662 6289
rect 3708 6367 3762 6473
rect 3808 6551 3862 6558
rect 3808 6499 3809 6551
rect 3861 6499 3862 6551
rect 3808 6473 3818 6499
rect 3852 6473 3862 6499
rect 3808 6461 3862 6473
rect 3908 6507 3962 6613
rect 4008 6647 4062 6659
rect 4008 6621 4018 6647
rect 4052 6621 4062 6647
rect 4008 6569 4009 6621
rect 4061 6569 4062 6621
rect 4008 6562 4062 6569
rect 4108 6647 4162 6753
rect 4208 6831 4262 6838
rect 4208 6779 4209 6831
rect 4261 6779 4262 6831
rect 4208 6753 4218 6779
rect 4252 6753 4262 6779
rect 4208 6741 4262 6753
rect 4308 6787 4362 6893
rect 4408 6927 4462 6939
rect 4408 6901 4418 6927
rect 4452 6901 4462 6927
rect 4408 6849 4409 6901
rect 4461 6849 4462 6901
rect 4408 6842 4462 6849
rect 4508 6927 4562 7033
rect 4608 7111 4662 7118
rect 4608 7059 4609 7111
rect 4661 7059 4662 7111
rect 4608 7033 4618 7059
rect 4652 7033 4662 7059
rect 4608 7021 4662 7033
rect 4708 7067 4762 7173
rect 4808 7207 4862 7219
rect 4808 7181 4818 7207
rect 4852 7181 4862 7207
rect 4808 7129 4809 7181
rect 4861 7129 4862 7181
rect 4808 7122 4862 7129
rect 4908 7207 4962 7313
rect 5008 7391 5062 7398
rect 5008 7339 5009 7391
rect 5061 7339 5062 7391
rect 5008 7313 5018 7339
rect 5052 7313 5062 7339
rect 5008 7301 5062 7313
rect 5108 7347 5162 7543
rect 5208 7577 5262 7589
rect 5208 7551 5218 7577
rect 5252 7551 5262 7577
rect 5208 7499 5209 7551
rect 5261 7499 5262 7551
rect 5208 7492 5262 7499
rect 5308 7577 5362 7683
rect 5408 7761 5462 7768
rect 5408 7709 5409 7761
rect 5461 7709 5462 7761
rect 5408 7683 5418 7709
rect 5452 7683 5462 7709
rect 5408 7671 5462 7683
rect 5508 7717 5562 7823
rect 5608 7857 5662 7869
rect 5608 7831 5618 7857
rect 5652 7831 5662 7857
rect 5608 7779 5609 7831
rect 5661 7779 5662 7831
rect 5608 7772 5662 7779
rect 5708 7857 5762 7963
rect 5808 8041 5862 8048
rect 5808 7989 5809 8041
rect 5861 7989 5862 8041
rect 5808 7963 5818 7989
rect 5852 7963 5862 7989
rect 5808 7951 5862 7963
rect 5908 7997 5962 8103
rect 6008 8137 6062 8149
rect 6008 8111 6018 8137
rect 6052 8111 6062 8137
rect 6008 8059 6009 8111
rect 6061 8059 6062 8111
rect 6008 8052 6062 8059
rect 6108 8137 6162 8243
rect 6208 8321 6262 8328
rect 6208 8269 6209 8321
rect 6261 8269 6262 8321
rect 6208 8243 6218 8269
rect 6252 8243 6262 8269
rect 6208 8231 6262 8243
rect 6308 8277 6362 8383
rect 6408 8417 6462 8429
rect 6408 8391 6418 8417
rect 6452 8391 6462 8417
rect 6408 8339 6409 8391
rect 6461 8339 6462 8391
rect 6408 8332 6462 8339
rect 6506 8398 6516 8432
rect 6550 8398 6560 8432
rect 6506 8391 6560 8398
rect 6506 8339 6507 8391
rect 6559 8339 6560 8391
rect 6506 8332 6560 8339
rect 6506 8292 6560 8304
rect 6308 8243 6318 8277
rect 6352 8243 6362 8277
rect 6108 8103 6118 8137
rect 6152 8103 6162 8137
rect 5908 7963 5918 7997
rect 5952 7963 5962 7997
rect 5708 7823 5718 7857
rect 5752 7823 5762 7857
rect 5508 7683 5518 7717
rect 5552 7683 5562 7717
rect 5308 7543 5318 7577
rect 5352 7543 5362 7577
rect 5202 7463 5268 7464
rect 5202 7411 5209 7463
rect 5261 7411 5268 7463
rect 5202 7410 5268 7411
rect 5108 7313 5118 7347
rect 5152 7313 5162 7347
rect 4908 7173 4918 7207
rect 4952 7173 4962 7207
rect 4708 7033 4718 7067
rect 4752 7033 4762 7067
rect 4508 6893 4518 6927
rect 4552 6893 4562 6927
rect 4308 6753 4318 6787
rect 4352 6753 4362 6787
rect 4108 6613 4118 6647
rect 4152 6613 4162 6647
rect 3908 6473 3918 6507
rect 3952 6473 3962 6507
rect 3708 6333 3718 6367
rect 3752 6333 3762 6367
rect 3602 6253 3668 6254
rect 3602 6201 3609 6253
rect 3661 6201 3668 6253
rect 3602 6200 3668 6201
rect 3508 6103 3518 6137
rect 3552 6103 3562 6137
rect 3308 5963 3318 5997
rect 3352 5963 3362 5997
rect 3108 5823 3118 5857
rect 3152 5823 3162 5857
rect 2908 5683 2918 5717
rect 2952 5683 2962 5717
rect 2708 5543 2718 5577
rect 2752 5543 2762 5577
rect 2508 5403 2518 5437
rect 2552 5403 2562 5437
rect 2308 5263 2318 5297
rect 2352 5263 2362 5297
rect 2108 5123 2118 5157
rect 2152 5123 2162 5157
rect 2108 5040 2162 5123
rect 2208 5201 2262 5208
rect 2208 5149 2209 5201
rect 2261 5149 2262 5201
rect 2208 5123 2218 5149
rect 2252 5123 2262 5149
rect 2208 5111 2262 5123
rect 2308 5157 2362 5263
rect 2408 5297 2462 5309
rect 2408 5271 2418 5297
rect 2452 5271 2462 5297
rect 2408 5219 2409 5271
rect 2461 5219 2462 5271
rect 2408 5212 2462 5219
rect 2508 5297 2562 5403
rect 2608 5481 2662 5488
rect 2608 5429 2609 5481
rect 2661 5429 2662 5481
rect 2608 5403 2618 5429
rect 2652 5403 2662 5429
rect 2608 5391 2662 5403
rect 2708 5437 2762 5543
rect 2808 5577 2862 5589
rect 2808 5551 2818 5577
rect 2852 5551 2862 5577
rect 2808 5499 2809 5551
rect 2861 5499 2862 5551
rect 2808 5492 2862 5499
rect 2908 5577 2962 5683
rect 3008 5761 3062 5768
rect 3008 5709 3009 5761
rect 3061 5709 3062 5761
rect 3008 5683 3018 5709
rect 3052 5683 3062 5709
rect 3008 5671 3062 5683
rect 3108 5717 3162 5823
rect 3208 5857 3262 5869
rect 3208 5831 3218 5857
rect 3252 5831 3262 5857
rect 3208 5779 3209 5831
rect 3261 5779 3262 5831
rect 3208 5772 3262 5779
rect 3308 5857 3362 5963
rect 3408 6041 3462 6048
rect 3408 5989 3409 6041
rect 3461 5989 3462 6041
rect 3408 5963 3418 5989
rect 3452 5963 3462 5989
rect 3408 5951 3462 5963
rect 3508 5997 3562 6103
rect 3608 6137 3662 6149
rect 3608 6111 3618 6137
rect 3652 6111 3662 6137
rect 3608 6059 3609 6111
rect 3661 6059 3662 6111
rect 3608 6052 3662 6059
rect 3708 6137 3762 6333
rect 3808 6411 3862 6418
rect 3808 6359 3809 6411
rect 3861 6359 3862 6411
rect 3808 6333 3818 6359
rect 3852 6333 3862 6359
rect 3808 6321 3862 6333
rect 3908 6367 3962 6473
rect 4008 6507 4062 6519
rect 4008 6481 4018 6507
rect 4052 6481 4062 6507
rect 4008 6429 4009 6481
rect 4061 6429 4062 6481
rect 4008 6422 4062 6429
rect 4108 6507 4162 6613
rect 4208 6691 4262 6698
rect 4208 6639 4209 6691
rect 4261 6639 4262 6691
rect 4208 6613 4218 6639
rect 4252 6613 4262 6639
rect 4208 6601 4262 6613
rect 4308 6647 4362 6753
rect 4408 6787 4462 6799
rect 4408 6761 4418 6787
rect 4452 6761 4462 6787
rect 4408 6709 4409 6761
rect 4461 6709 4462 6761
rect 4408 6702 4462 6709
rect 4508 6787 4562 6893
rect 4608 6971 4662 6978
rect 4608 6919 4609 6971
rect 4661 6919 4662 6971
rect 4608 6893 4618 6919
rect 4652 6893 4662 6919
rect 4608 6881 4662 6893
rect 4708 6927 4762 7033
rect 4808 7067 4862 7079
rect 4808 7041 4818 7067
rect 4852 7041 4862 7067
rect 4808 6989 4809 7041
rect 4861 6989 4862 7041
rect 4808 6982 4862 6989
rect 4908 7067 4962 7173
rect 5008 7251 5062 7258
rect 5008 7199 5009 7251
rect 5061 7199 5062 7251
rect 5008 7173 5018 7199
rect 5052 7173 5062 7199
rect 5008 7161 5062 7173
rect 5108 7207 5162 7313
rect 5208 7347 5262 7359
rect 5208 7321 5218 7347
rect 5252 7321 5262 7347
rect 5208 7269 5209 7321
rect 5261 7269 5262 7321
rect 5208 7262 5262 7269
rect 5308 7347 5362 7543
rect 5408 7621 5462 7628
rect 5408 7569 5409 7621
rect 5461 7569 5462 7621
rect 5408 7543 5418 7569
rect 5452 7543 5462 7569
rect 5408 7531 5462 7543
rect 5508 7577 5562 7683
rect 5608 7717 5662 7729
rect 5608 7691 5618 7717
rect 5652 7691 5662 7717
rect 5608 7639 5609 7691
rect 5661 7639 5662 7691
rect 5608 7632 5662 7639
rect 5708 7717 5762 7823
rect 5808 7901 5862 7908
rect 5808 7849 5809 7901
rect 5861 7849 5862 7901
rect 5808 7823 5818 7849
rect 5852 7823 5862 7849
rect 5808 7811 5862 7823
rect 5908 7857 5962 7963
rect 6008 7997 6062 8009
rect 6008 7971 6018 7997
rect 6052 7971 6062 7997
rect 6008 7919 6009 7971
rect 6061 7919 6062 7971
rect 6008 7912 6062 7919
rect 6108 7997 6162 8103
rect 6208 8181 6262 8188
rect 6208 8129 6209 8181
rect 6261 8129 6262 8181
rect 6208 8103 6218 8129
rect 6252 8103 6262 8129
rect 6208 8091 6262 8103
rect 6308 8137 6362 8243
rect 6408 8277 6462 8289
rect 6408 8251 6418 8277
rect 6452 8251 6462 8277
rect 6408 8199 6409 8251
rect 6461 8199 6462 8251
rect 6408 8192 6462 8199
rect 6506 8258 6516 8292
rect 6550 8258 6560 8292
rect 6506 8251 6560 8258
rect 6506 8199 6507 8251
rect 6559 8199 6560 8251
rect 6506 8192 6560 8199
rect 6506 8152 6560 8164
rect 6308 8103 6318 8137
rect 6352 8103 6362 8137
rect 6108 7963 6118 7997
rect 6152 7963 6162 7997
rect 5908 7823 5918 7857
rect 5952 7823 5962 7857
rect 5708 7683 5718 7717
rect 5752 7683 5762 7717
rect 5508 7543 5518 7577
rect 5552 7543 5562 7577
rect 5402 7479 5468 7480
rect 5402 7427 5409 7479
rect 5461 7427 5468 7479
rect 5402 7426 5468 7427
rect 5308 7313 5318 7347
rect 5352 7313 5362 7347
rect 5108 7173 5118 7207
rect 5152 7173 5162 7207
rect 4908 7033 4918 7067
rect 4952 7033 4962 7067
rect 4708 6893 4718 6927
rect 4752 6893 4762 6927
rect 4508 6753 4518 6787
rect 4552 6753 4562 6787
rect 4308 6613 4318 6647
rect 4352 6613 4362 6647
rect 4108 6473 4118 6507
rect 4152 6473 4162 6507
rect 3908 6333 3918 6367
rect 3952 6333 3962 6367
rect 3802 6269 3868 6270
rect 3802 6217 3809 6269
rect 3861 6217 3868 6269
rect 3802 6216 3868 6217
rect 3708 6103 3718 6137
rect 3752 6103 3762 6137
rect 3508 5963 3518 5997
rect 3552 5963 3562 5997
rect 3308 5823 3318 5857
rect 3352 5823 3362 5857
rect 3108 5683 3118 5717
rect 3152 5683 3162 5717
rect 2908 5543 2918 5577
rect 2952 5543 2962 5577
rect 2708 5403 2718 5437
rect 2752 5403 2762 5437
rect 2508 5263 2518 5297
rect 2552 5263 2562 5297
rect 2308 5123 2318 5157
rect 2352 5123 2362 5157
rect 2308 5040 2362 5123
rect 2408 5157 2462 5169
rect 2408 5131 2418 5157
rect 2452 5131 2462 5157
rect 2408 5079 2409 5131
rect 2461 5079 2462 5131
rect 2408 5072 2462 5079
rect 2508 5157 2562 5263
rect 2608 5341 2662 5348
rect 2608 5289 2609 5341
rect 2661 5289 2662 5341
rect 2608 5263 2618 5289
rect 2652 5263 2662 5289
rect 2608 5251 2662 5263
rect 2708 5297 2762 5403
rect 2808 5437 2862 5449
rect 2808 5411 2818 5437
rect 2852 5411 2862 5437
rect 2808 5359 2809 5411
rect 2861 5359 2862 5411
rect 2808 5352 2862 5359
rect 2908 5437 2962 5543
rect 3008 5621 3062 5628
rect 3008 5569 3009 5621
rect 3061 5569 3062 5621
rect 3008 5543 3018 5569
rect 3052 5543 3062 5569
rect 3008 5531 3062 5543
rect 3108 5577 3162 5683
rect 3208 5717 3262 5729
rect 3208 5691 3218 5717
rect 3252 5691 3262 5717
rect 3208 5639 3209 5691
rect 3261 5639 3262 5691
rect 3208 5632 3262 5639
rect 3308 5717 3362 5823
rect 3408 5901 3462 5908
rect 3408 5849 3409 5901
rect 3461 5849 3462 5901
rect 3408 5823 3418 5849
rect 3452 5823 3462 5849
rect 3408 5811 3462 5823
rect 3508 5857 3562 5963
rect 3608 5997 3662 6009
rect 3608 5971 3618 5997
rect 3652 5971 3662 5997
rect 3608 5919 3609 5971
rect 3661 5919 3662 5971
rect 3608 5912 3662 5919
rect 3708 5997 3762 6103
rect 3808 6181 3862 6188
rect 3808 6129 3809 6181
rect 3861 6129 3862 6181
rect 3808 6103 3818 6129
rect 3852 6103 3862 6129
rect 3808 6091 3862 6103
rect 3908 6137 3962 6333
rect 4008 6367 4062 6379
rect 4008 6341 4018 6367
rect 4052 6341 4062 6367
rect 4008 6289 4009 6341
rect 4061 6289 4062 6341
rect 4008 6282 4062 6289
rect 4108 6367 4162 6473
rect 4208 6551 4262 6558
rect 4208 6499 4209 6551
rect 4261 6499 4262 6551
rect 4208 6473 4218 6499
rect 4252 6473 4262 6499
rect 4208 6461 4262 6473
rect 4308 6507 4362 6613
rect 4408 6647 4462 6659
rect 4408 6621 4418 6647
rect 4452 6621 4462 6647
rect 4408 6569 4409 6621
rect 4461 6569 4462 6621
rect 4408 6562 4462 6569
rect 4508 6647 4562 6753
rect 4608 6831 4662 6838
rect 4608 6779 4609 6831
rect 4661 6779 4662 6831
rect 4608 6753 4618 6779
rect 4652 6753 4662 6779
rect 4608 6741 4662 6753
rect 4708 6787 4762 6893
rect 4808 6927 4862 6939
rect 4808 6901 4818 6927
rect 4852 6901 4862 6927
rect 4808 6849 4809 6901
rect 4861 6849 4862 6901
rect 4808 6842 4862 6849
rect 4908 6927 4962 7033
rect 5008 7111 5062 7118
rect 5008 7059 5009 7111
rect 5061 7059 5062 7111
rect 5008 7033 5018 7059
rect 5052 7033 5062 7059
rect 5008 7021 5062 7033
rect 5108 7067 5162 7173
rect 5208 7207 5262 7219
rect 5208 7181 5218 7207
rect 5252 7181 5262 7207
rect 5208 7129 5209 7181
rect 5261 7129 5262 7181
rect 5208 7122 5262 7129
rect 5308 7207 5362 7313
rect 5408 7391 5462 7398
rect 5408 7339 5409 7391
rect 5461 7339 5462 7391
rect 5408 7313 5418 7339
rect 5452 7313 5462 7339
rect 5408 7301 5462 7313
rect 5508 7347 5562 7543
rect 5608 7577 5662 7589
rect 5608 7551 5618 7577
rect 5652 7551 5662 7577
rect 5608 7499 5609 7551
rect 5661 7499 5662 7551
rect 5608 7492 5662 7499
rect 5708 7577 5762 7683
rect 5808 7761 5862 7768
rect 5808 7709 5809 7761
rect 5861 7709 5862 7761
rect 5808 7683 5818 7709
rect 5852 7683 5862 7709
rect 5808 7671 5862 7683
rect 5908 7717 5962 7823
rect 6008 7857 6062 7869
rect 6008 7831 6018 7857
rect 6052 7831 6062 7857
rect 6008 7779 6009 7831
rect 6061 7779 6062 7831
rect 6008 7772 6062 7779
rect 6108 7857 6162 7963
rect 6208 8041 6262 8048
rect 6208 7989 6209 8041
rect 6261 7989 6262 8041
rect 6208 7963 6218 7989
rect 6252 7963 6262 7989
rect 6208 7951 6262 7963
rect 6308 7997 6362 8103
rect 6408 8137 6462 8149
rect 6408 8111 6418 8137
rect 6452 8111 6462 8137
rect 6408 8059 6409 8111
rect 6461 8059 6462 8111
rect 6408 8052 6462 8059
rect 6506 8118 6516 8152
rect 6550 8118 6560 8152
rect 6506 8111 6560 8118
rect 6506 8059 6507 8111
rect 6559 8059 6560 8111
rect 6506 8052 6560 8059
rect 6506 8012 6560 8024
rect 6308 7963 6318 7997
rect 6352 7963 6362 7997
rect 6108 7823 6118 7857
rect 6152 7823 6162 7857
rect 5908 7683 5918 7717
rect 5952 7683 5962 7717
rect 5708 7543 5718 7577
rect 5752 7543 5762 7577
rect 5602 7463 5668 7464
rect 5602 7411 5609 7463
rect 5661 7411 5668 7463
rect 5602 7410 5668 7411
rect 5508 7313 5518 7347
rect 5552 7313 5562 7347
rect 5308 7173 5318 7207
rect 5352 7173 5362 7207
rect 5108 7033 5118 7067
rect 5152 7033 5162 7067
rect 4908 6893 4918 6927
rect 4952 6893 4962 6927
rect 4708 6753 4718 6787
rect 4752 6753 4762 6787
rect 4508 6613 4518 6647
rect 4552 6613 4562 6647
rect 4308 6473 4318 6507
rect 4352 6473 4362 6507
rect 4108 6333 4118 6367
rect 4152 6333 4162 6367
rect 4002 6253 4068 6254
rect 4002 6201 4009 6253
rect 4061 6201 4068 6253
rect 4002 6200 4068 6201
rect 3908 6103 3918 6137
rect 3952 6103 3962 6137
rect 3708 5963 3718 5997
rect 3752 5963 3762 5997
rect 3508 5823 3518 5857
rect 3552 5823 3562 5857
rect 3308 5683 3318 5717
rect 3352 5683 3362 5717
rect 3108 5543 3118 5577
rect 3152 5543 3162 5577
rect 2908 5403 2918 5437
rect 2952 5403 2962 5437
rect 2708 5263 2718 5297
rect 2752 5263 2762 5297
rect 2508 5123 2518 5157
rect 2552 5123 2562 5157
rect 2508 5040 2562 5123
rect 2608 5201 2662 5208
rect 2608 5149 2609 5201
rect 2661 5149 2662 5201
rect 2608 5123 2618 5149
rect 2652 5123 2662 5149
rect 2608 5111 2662 5123
rect 2708 5157 2762 5263
rect 2808 5297 2862 5309
rect 2808 5271 2818 5297
rect 2852 5271 2862 5297
rect 2808 5219 2809 5271
rect 2861 5219 2862 5271
rect 2808 5212 2862 5219
rect 2908 5297 2962 5403
rect 3008 5481 3062 5488
rect 3008 5429 3009 5481
rect 3061 5429 3062 5481
rect 3008 5403 3018 5429
rect 3052 5403 3062 5429
rect 3008 5391 3062 5403
rect 3108 5437 3162 5543
rect 3208 5577 3262 5589
rect 3208 5551 3218 5577
rect 3252 5551 3262 5577
rect 3208 5499 3209 5551
rect 3261 5499 3262 5551
rect 3208 5492 3262 5499
rect 3308 5577 3362 5683
rect 3408 5761 3462 5768
rect 3408 5709 3409 5761
rect 3461 5709 3462 5761
rect 3408 5683 3418 5709
rect 3452 5683 3462 5709
rect 3408 5671 3462 5683
rect 3508 5717 3562 5823
rect 3608 5857 3662 5869
rect 3608 5831 3618 5857
rect 3652 5831 3662 5857
rect 3608 5779 3609 5831
rect 3661 5779 3662 5831
rect 3608 5772 3662 5779
rect 3708 5857 3762 5963
rect 3808 6041 3862 6048
rect 3808 5989 3809 6041
rect 3861 5989 3862 6041
rect 3808 5963 3818 5989
rect 3852 5963 3862 5989
rect 3808 5951 3862 5963
rect 3908 5997 3962 6103
rect 4008 6137 4062 6149
rect 4008 6111 4018 6137
rect 4052 6111 4062 6137
rect 4008 6059 4009 6111
rect 4061 6059 4062 6111
rect 4008 6052 4062 6059
rect 4108 6137 4162 6333
rect 4208 6411 4262 6418
rect 4208 6359 4209 6411
rect 4261 6359 4262 6411
rect 4208 6333 4218 6359
rect 4252 6333 4262 6359
rect 4208 6321 4262 6333
rect 4308 6367 4362 6473
rect 4408 6507 4462 6519
rect 4408 6481 4418 6507
rect 4452 6481 4462 6507
rect 4408 6429 4409 6481
rect 4461 6429 4462 6481
rect 4408 6422 4462 6429
rect 4508 6507 4562 6613
rect 4608 6691 4662 6698
rect 4608 6639 4609 6691
rect 4661 6639 4662 6691
rect 4608 6613 4618 6639
rect 4652 6613 4662 6639
rect 4608 6601 4662 6613
rect 4708 6647 4762 6753
rect 4808 6787 4862 6799
rect 4808 6761 4818 6787
rect 4852 6761 4862 6787
rect 4808 6709 4809 6761
rect 4861 6709 4862 6761
rect 4808 6702 4862 6709
rect 4908 6787 4962 6893
rect 5008 6971 5062 6978
rect 5008 6919 5009 6971
rect 5061 6919 5062 6971
rect 5008 6893 5018 6919
rect 5052 6893 5062 6919
rect 5008 6881 5062 6893
rect 5108 6927 5162 7033
rect 5208 7067 5262 7079
rect 5208 7041 5218 7067
rect 5252 7041 5262 7067
rect 5208 6989 5209 7041
rect 5261 6989 5262 7041
rect 5208 6982 5262 6989
rect 5308 7067 5362 7173
rect 5408 7251 5462 7258
rect 5408 7199 5409 7251
rect 5461 7199 5462 7251
rect 5408 7173 5418 7199
rect 5452 7173 5462 7199
rect 5408 7161 5462 7173
rect 5508 7207 5562 7313
rect 5608 7347 5662 7359
rect 5608 7321 5618 7347
rect 5652 7321 5662 7347
rect 5608 7269 5609 7321
rect 5661 7269 5662 7321
rect 5608 7262 5662 7269
rect 5708 7347 5762 7543
rect 5808 7621 5862 7628
rect 5808 7569 5809 7621
rect 5861 7569 5862 7621
rect 5808 7543 5818 7569
rect 5852 7543 5862 7569
rect 5808 7531 5862 7543
rect 5908 7577 5962 7683
rect 6008 7717 6062 7729
rect 6008 7691 6018 7717
rect 6052 7691 6062 7717
rect 6008 7639 6009 7691
rect 6061 7639 6062 7691
rect 6008 7632 6062 7639
rect 6108 7717 6162 7823
rect 6208 7901 6262 7908
rect 6208 7849 6209 7901
rect 6261 7849 6262 7901
rect 6208 7823 6218 7849
rect 6252 7823 6262 7849
rect 6208 7811 6262 7823
rect 6308 7857 6362 7963
rect 6408 7997 6462 8009
rect 6408 7971 6418 7997
rect 6452 7971 6462 7997
rect 6408 7919 6409 7971
rect 6461 7919 6462 7971
rect 6408 7912 6462 7919
rect 6506 7978 6516 8012
rect 6550 7978 6560 8012
rect 6506 7971 6560 7978
rect 6506 7919 6507 7971
rect 6559 7919 6560 7971
rect 6506 7912 6560 7919
rect 6506 7872 6560 7884
rect 6308 7823 6318 7857
rect 6352 7823 6362 7857
rect 6108 7683 6118 7717
rect 6152 7683 6162 7717
rect 5908 7543 5918 7577
rect 5952 7543 5962 7577
rect 5802 7479 5868 7480
rect 5802 7427 5809 7479
rect 5861 7427 5868 7479
rect 5802 7426 5868 7427
rect 5708 7313 5718 7347
rect 5752 7313 5762 7347
rect 5508 7173 5518 7207
rect 5552 7173 5562 7207
rect 5308 7033 5318 7067
rect 5352 7033 5362 7067
rect 5108 6893 5118 6927
rect 5152 6893 5162 6927
rect 4908 6753 4918 6787
rect 4952 6753 4962 6787
rect 4708 6613 4718 6647
rect 4752 6613 4762 6647
rect 4508 6473 4518 6507
rect 4552 6473 4562 6507
rect 4308 6333 4318 6367
rect 4352 6333 4362 6367
rect 4202 6269 4268 6270
rect 4202 6217 4209 6269
rect 4261 6217 4268 6269
rect 4202 6216 4268 6217
rect 4108 6103 4118 6137
rect 4152 6103 4162 6137
rect 3908 5963 3918 5997
rect 3952 5963 3962 5997
rect 3708 5823 3718 5857
rect 3752 5823 3762 5857
rect 3508 5683 3518 5717
rect 3552 5683 3562 5717
rect 3308 5543 3318 5577
rect 3352 5543 3362 5577
rect 3108 5403 3118 5437
rect 3152 5403 3162 5437
rect 2908 5263 2918 5297
rect 2952 5263 2962 5297
rect 2708 5123 2718 5157
rect 2752 5123 2762 5157
rect 2708 5040 2762 5123
rect 2808 5157 2862 5169
rect 2808 5131 2818 5157
rect 2852 5131 2862 5157
rect 2808 5079 2809 5131
rect 2861 5079 2862 5131
rect 2808 5072 2862 5079
rect 2908 5157 2962 5263
rect 3008 5341 3062 5348
rect 3008 5289 3009 5341
rect 3061 5289 3062 5341
rect 3008 5263 3018 5289
rect 3052 5263 3062 5289
rect 3008 5251 3062 5263
rect 3108 5297 3162 5403
rect 3208 5437 3262 5449
rect 3208 5411 3218 5437
rect 3252 5411 3262 5437
rect 3208 5359 3209 5411
rect 3261 5359 3262 5411
rect 3208 5352 3262 5359
rect 3308 5437 3362 5543
rect 3408 5621 3462 5628
rect 3408 5569 3409 5621
rect 3461 5569 3462 5621
rect 3408 5543 3418 5569
rect 3452 5543 3462 5569
rect 3408 5531 3462 5543
rect 3508 5577 3562 5683
rect 3608 5717 3662 5729
rect 3608 5691 3618 5717
rect 3652 5691 3662 5717
rect 3608 5639 3609 5691
rect 3661 5639 3662 5691
rect 3608 5632 3662 5639
rect 3708 5717 3762 5823
rect 3808 5901 3862 5908
rect 3808 5849 3809 5901
rect 3861 5849 3862 5901
rect 3808 5823 3818 5849
rect 3852 5823 3862 5849
rect 3808 5811 3862 5823
rect 3908 5857 3962 5963
rect 4008 5997 4062 6009
rect 4008 5971 4018 5997
rect 4052 5971 4062 5997
rect 4008 5919 4009 5971
rect 4061 5919 4062 5971
rect 4008 5912 4062 5919
rect 4108 5997 4162 6103
rect 4208 6181 4262 6188
rect 4208 6129 4209 6181
rect 4261 6129 4262 6181
rect 4208 6103 4218 6129
rect 4252 6103 4262 6129
rect 4208 6091 4262 6103
rect 4308 6137 4362 6333
rect 4408 6367 4462 6379
rect 4408 6341 4418 6367
rect 4452 6341 4462 6367
rect 4408 6289 4409 6341
rect 4461 6289 4462 6341
rect 4408 6282 4462 6289
rect 4508 6367 4562 6473
rect 4608 6551 4662 6558
rect 4608 6499 4609 6551
rect 4661 6499 4662 6551
rect 4608 6473 4618 6499
rect 4652 6473 4662 6499
rect 4608 6461 4662 6473
rect 4708 6507 4762 6613
rect 4808 6647 4862 6659
rect 4808 6621 4818 6647
rect 4852 6621 4862 6647
rect 4808 6569 4809 6621
rect 4861 6569 4862 6621
rect 4808 6562 4862 6569
rect 4908 6647 4962 6753
rect 5008 6831 5062 6838
rect 5008 6779 5009 6831
rect 5061 6779 5062 6831
rect 5008 6753 5018 6779
rect 5052 6753 5062 6779
rect 5008 6741 5062 6753
rect 5108 6787 5162 6893
rect 5208 6927 5262 6939
rect 5208 6901 5218 6927
rect 5252 6901 5262 6927
rect 5208 6849 5209 6901
rect 5261 6849 5262 6901
rect 5208 6842 5262 6849
rect 5308 6927 5362 7033
rect 5408 7111 5462 7118
rect 5408 7059 5409 7111
rect 5461 7059 5462 7111
rect 5408 7033 5418 7059
rect 5452 7033 5462 7059
rect 5408 7021 5462 7033
rect 5508 7067 5562 7173
rect 5608 7207 5662 7219
rect 5608 7181 5618 7207
rect 5652 7181 5662 7207
rect 5608 7129 5609 7181
rect 5661 7129 5662 7181
rect 5608 7122 5662 7129
rect 5708 7207 5762 7313
rect 5808 7391 5862 7398
rect 5808 7339 5809 7391
rect 5861 7339 5862 7391
rect 5808 7313 5818 7339
rect 5852 7313 5862 7339
rect 5808 7301 5862 7313
rect 5908 7347 5962 7543
rect 6008 7577 6062 7589
rect 6008 7551 6018 7577
rect 6052 7551 6062 7577
rect 6008 7499 6009 7551
rect 6061 7499 6062 7551
rect 6008 7492 6062 7499
rect 6108 7577 6162 7683
rect 6208 7761 6262 7768
rect 6208 7709 6209 7761
rect 6261 7709 6262 7761
rect 6208 7683 6218 7709
rect 6252 7683 6262 7709
rect 6208 7671 6262 7683
rect 6308 7717 6362 7823
rect 6408 7857 6462 7869
rect 6408 7831 6418 7857
rect 6452 7831 6462 7857
rect 6408 7779 6409 7831
rect 6461 7779 6462 7831
rect 6408 7772 6462 7779
rect 6506 7838 6516 7872
rect 6550 7838 6560 7872
rect 6506 7831 6560 7838
rect 6506 7779 6507 7831
rect 6559 7779 6560 7831
rect 6506 7772 6560 7779
rect 6506 7732 6560 7744
rect 6308 7683 6318 7717
rect 6352 7683 6362 7717
rect 6108 7543 6118 7577
rect 6152 7543 6162 7577
rect 6002 7463 6068 7464
rect 6002 7411 6009 7463
rect 6061 7411 6068 7463
rect 6002 7410 6068 7411
rect 5908 7313 5918 7347
rect 5952 7313 5962 7347
rect 5708 7173 5718 7207
rect 5752 7173 5762 7207
rect 5508 7033 5518 7067
rect 5552 7033 5562 7067
rect 5308 6893 5318 6927
rect 5352 6893 5362 6927
rect 5108 6753 5118 6787
rect 5152 6753 5162 6787
rect 4908 6613 4918 6647
rect 4952 6613 4962 6647
rect 4708 6473 4718 6507
rect 4752 6473 4762 6507
rect 4508 6333 4518 6367
rect 4552 6333 4562 6367
rect 4402 6253 4468 6254
rect 4402 6201 4409 6253
rect 4461 6201 4468 6253
rect 4402 6200 4468 6201
rect 4308 6103 4318 6137
rect 4352 6103 4362 6137
rect 4108 5963 4118 5997
rect 4152 5963 4162 5997
rect 3908 5823 3918 5857
rect 3952 5823 3962 5857
rect 3708 5683 3718 5717
rect 3752 5683 3762 5717
rect 3508 5543 3518 5577
rect 3552 5543 3562 5577
rect 3308 5403 3318 5437
rect 3352 5403 3362 5437
rect 3108 5263 3118 5297
rect 3152 5263 3162 5297
rect 2908 5123 2918 5157
rect 2952 5123 2962 5157
rect 2908 5040 2962 5123
rect 3008 5201 3062 5208
rect 3008 5149 3009 5201
rect 3061 5149 3062 5201
rect 3008 5123 3018 5149
rect 3052 5123 3062 5149
rect 3008 5111 3062 5123
rect 3108 5157 3162 5263
rect 3208 5297 3262 5309
rect 3208 5271 3218 5297
rect 3252 5271 3262 5297
rect 3208 5219 3209 5271
rect 3261 5219 3262 5271
rect 3208 5212 3262 5219
rect 3308 5297 3362 5403
rect 3408 5481 3462 5488
rect 3408 5429 3409 5481
rect 3461 5429 3462 5481
rect 3408 5403 3418 5429
rect 3452 5403 3462 5429
rect 3408 5391 3462 5403
rect 3508 5437 3562 5543
rect 3608 5577 3662 5589
rect 3608 5551 3618 5577
rect 3652 5551 3662 5577
rect 3608 5499 3609 5551
rect 3661 5499 3662 5551
rect 3608 5492 3662 5499
rect 3708 5577 3762 5683
rect 3808 5761 3862 5768
rect 3808 5709 3809 5761
rect 3861 5709 3862 5761
rect 3808 5683 3818 5709
rect 3852 5683 3862 5709
rect 3808 5671 3862 5683
rect 3908 5717 3962 5823
rect 4008 5857 4062 5869
rect 4008 5831 4018 5857
rect 4052 5831 4062 5857
rect 4008 5779 4009 5831
rect 4061 5779 4062 5831
rect 4008 5772 4062 5779
rect 4108 5857 4162 5963
rect 4208 6041 4262 6048
rect 4208 5989 4209 6041
rect 4261 5989 4262 6041
rect 4208 5963 4218 5989
rect 4252 5963 4262 5989
rect 4208 5951 4262 5963
rect 4308 5997 4362 6103
rect 4408 6137 4462 6149
rect 4408 6111 4418 6137
rect 4452 6111 4462 6137
rect 4408 6059 4409 6111
rect 4461 6059 4462 6111
rect 4408 6052 4462 6059
rect 4508 6137 4562 6333
rect 4608 6411 4662 6418
rect 4608 6359 4609 6411
rect 4661 6359 4662 6411
rect 4608 6333 4618 6359
rect 4652 6333 4662 6359
rect 4608 6321 4662 6333
rect 4708 6367 4762 6473
rect 4808 6507 4862 6519
rect 4808 6481 4818 6507
rect 4852 6481 4862 6507
rect 4808 6429 4809 6481
rect 4861 6429 4862 6481
rect 4808 6422 4862 6429
rect 4908 6507 4962 6613
rect 5008 6691 5062 6698
rect 5008 6639 5009 6691
rect 5061 6639 5062 6691
rect 5008 6613 5018 6639
rect 5052 6613 5062 6639
rect 5008 6601 5062 6613
rect 5108 6647 5162 6753
rect 5208 6787 5262 6799
rect 5208 6761 5218 6787
rect 5252 6761 5262 6787
rect 5208 6709 5209 6761
rect 5261 6709 5262 6761
rect 5208 6702 5262 6709
rect 5308 6787 5362 6893
rect 5408 6971 5462 6978
rect 5408 6919 5409 6971
rect 5461 6919 5462 6971
rect 5408 6893 5418 6919
rect 5452 6893 5462 6919
rect 5408 6881 5462 6893
rect 5508 6927 5562 7033
rect 5608 7067 5662 7079
rect 5608 7041 5618 7067
rect 5652 7041 5662 7067
rect 5608 6989 5609 7041
rect 5661 6989 5662 7041
rect 5608 6982 5662 6989
rect 5708 7067 5762 7173
rect 5808 7251 5862 7258
rect 5808 7199 5809 7251
rect 5861 7199 5862 7251
rect 5808 7173 5818 7199
rect 5852 7173 5862 7199
rect 5808 7161 5862 7173
rect 5908 7207 5962 7313
rect 6008 7347 6062 7359
rect 6008 7321 6018 7347
rect 6052 7321 6062 7347
rect 6008 7269 6009 7321
rect 6061 7269 6062 7321
rect 6008 7262 6062 7269
rect 6108 7347 6162 7543
rect 6208 7621 6262 7628
rect 6208 7569 6209 7621
rect 6261 7569 6262 7621
rect 6208 7543 6218 7569
rect 6252 7543 6262 7569
rect 6208 7531 6262 7543
rect 6308 7577 6362 7683
rect 6408 7717 6462 7729
rect 6408 7691 6418 7717
rect 6452 7691 6462 7717
rect 6408 7639 6409 7691
rect 6461 7639 6462 7691
rect 6408 7632 6462 7639
rect 6506 7698 6516 7732
rect 6550 7698 6560 7732
rect 6506 7691 6560 7698
rect 6506 7639 6507 7691
rect 6559 7639 6560 7691
rect 6506 7632 6560 7639
rect 6506 7592 6560 7604
rect 6308 7543 6318 7577
rect 6352 7543 6362 7577
rect 6202 7479 6268 7480
rect 6202 7427 6209 7479
rect 6261 7427 6268 7479
rect 6202 7426 6268 7427
rect 6108 7313 6118 7347
rect 6152 7313 6162 7347
rect 5908 7173 5918 7207
rect 5952 7173 5962 7207
rect 5708 7033 5718 7067
rect 5752 7033 5762 7067
rect 5508 6893 5518 6927
rect 5552 6893 5562 6927
rect 5308 6753 5318 6787
rect 5352 6753 5362 6787
rect 5108 6613 5118 6647
rect 5152 6613 5162 6647
rect 4908 6473 4918 6507
rect 4952 6473 4962 6507
rect 4708 6333 4718 6367
rect 4752 6333 4762 6367
rect 4602 6269 4668 6270
rect 4602 6217 4609 6269
rect 4661 6217 4668 6269
rect 4602 6216 4668 6217
rect 4508 6103 4518 6137
rect 4552 6103 4562 6137
rect 4308 5963 4318 5997
rect 4352 5963 4362 5997
rect 4108 5823 4118 5857
rect 4152 5823 4162 5857
rect 3908 5683 3918 5717
rect 3952 5683 3962 5717
rect 3708 5543 3718 5577
rect 3752 5543 3762 5577
rect 3508 5403 3518 5437
rect 3552 5403 3562 5437
rect 3308 5263 3318 5297
rect 3352 5263 3362 5297
rect 3108 5123 3118 5157
rect 3152 5123 3162 5157
rect 3108 5040 3162 5123
rect 3208 5157 3262 5169
rect 3208 5131 3218 5157
rect 3252 5131 3262 5157
rect 3208 5079 3209 5131
rect 3261 5079 3262 5131
rect 3208 5072 3262 5079
rect 3308 5157 3362 5263
rect 3408 5341 3462 5348
rect 3408 5289 3409 5341
rect 3461 5289 3462 5341
rect 3408 5263 3418 5289
rect 3452 5263 3462 5289
rect 3408 5251 3462 5263
rect 3508 5297 3562 5403
rect 3608 5437 3662 5449
rect 3608 5411 3618 5437
rect 3652 5411 3662 5437
rect 3608 5359 3609 5411
rect 3661 5359 3662 5411
rect 3608 5352 3662 5359
rect 3708 5437 3762 5543
rect 3808 5621 3862 5628
rect 3808 5569 3809 5621
rect 3861 5569 3862 5621
rect 3808 5543 3818 5569
rect 3852 5543 3862 5569
rect 3808 5531 3862 5543
rect 3908 5577 3962 5683
rect 4008 5717 4062 5729
rect 4008 5691 4018 5717
rect 4052 5691 4062 5717
rect 4008 5639 4009 5691
rect 4061 5639 4062 5691
rect 4008 5632 4062 5639
rect 4108 5717 4162 5823
rect 4208 5901 4262 5908
rect 4208 5849 4209 5901
rect 4261 5849 4262 5901
rect 4208 5823 4218 5849
rect 4252 5823 4262 5849
rect 4208 5811 4262 5823
rect 4308 5857 4362 5963
rect 4408 5997 4462 6009
rect 4408 5971 4418 5997
rect 4452 5971 4462 5997
rect 4408 5919 4409 5971
rect 4461 5919 4462 5971
rect 4408 5912 4462 5919
rect 4508 5997 4562 6103
rect 4608 6181 4662 6188
rect 4608 6129 4609 6181
rect 4661 6129 4662 6181
rect 4608 6103 4618 6129
rect 4652 6103 4662 6129
rect 4608 6091 4662 6103
rect 4708 6137 4762 6333
rect 4808 6367 4862 6379
rect 4808 6341 4818 6367
rect 4852 6341 4862 6367
rect 4808 6289 4809 6341
rect 4861 6289 4862 6341
rect 4808 6282 4862 6289
rect 4908 6367 4962 6473
rect 5008 6551 5062 6558
rect 5008 6499 5009 6551
rect 5061 6499 5062 6551
rect 5008 6473 5018 6499
rect 5052 6473 5062 6499
rect 5008 6461 5062 6473
rect 5108 6507 5162 6613
rect 5208 6647 5262 6659
rect 5208 6621 5218 6647
rect 5252 6621 5262 6647
rect 5208 6569 5209 6621
rect 5261 6569 5262 6621
rect 5208 6562 5262 6569
rect 5308 6647 5362 6753
rect 5408 6831 5462 6838
rect 5408 6779 5409 6831
rect 5461 6779 5462 6831
rect 5408 6753 5418 6779
rect 5452 6753 5462 6779
rect 5408 6741 5462 6753
rect 5508 6787 5562 6893
rect 5608 6927 5662 6939
rect 5608 6901 5618 6927
rect 5652 6901 5662 6927
rect 5608 6849 5609 6901
rect 5661 6849 5662 6901
rect 5608 6842 5662 6849
rect 5708 6927 5762 7033
rect 5808 7111 5862 7118
rect 5808 7059 5809 7111
rect 5861 7059 5862 7111
rect 5808 7033 5818 7059
rect 5852 7033 5862 7059
rect 5808 7021 5862 7033
rect 5908 7067 5962 7173
rect 6008 7207 6062 7219
rect 6008 7181 6018 7207
rect 6052 7181 6062 7207
rect 6008 7129 6009 7181
rect 6061 7129 6062 7181
rect 6008 7122 6062 7129
rect 6108 7207 6162 7313
rect 6208 7391 6262 7398
rect 6208 7339 6209 7391
rect 6261 7339 6262 7391
rect 6208 7313 6218 7339
rect 6252 7313 6262 7339
rect 6208 7301 6262 7313
rect 6308 7347 6362 7543
rect 6408 7577 6462 7589
rect 6408 7551 6418 7577
rect 6452 7551 6462 7577
rect 6408 7499 6409 7551
rect 6461 7499 6462 7551
rect 6408 7492 6462 7499
rect 6506 7558 6516 7592
rect 6550 7558 6560 7592
rect 6506 7551 6560 7558
rect 6506 7499 6507 7551
rect 6559 7499 6560 7551
rect 6506 7492 6560 7499
rect 6590 7457 6620 8621
rect 6504 7451 6620 7457
rect 6504 7417 6516 7451
rect 6550 7417 6620 7451
rect 6504 7411 6620 7417
rect 6506 7362 6560 7374
rect 6308 7313 6318 7347
rect 6352 7313 6362 7347
rect 6108 7173 6118 7207
rect 6152 7173 6162 7207
rect 5908 7033 5918 7067
rect 5952 7033 5962 7067
rect 5708 6893 5718 6927
rect 5752 6893 5762 6927
rect 5508 6753 5518 6787
rect 5552 6753 5562 6787
rect 5308 6613 5318 6647
rect 5352 6613 5362 6647
rect 5108 6473 5118 6507
rect 5152 6473 5162 6507
rect 4908 6333 4918 6367
rect 4952 6333 4962 6367
rect 4802 6253 4868 6254
rect 4802 6201 4809 6253
rect 4861 6201 4868 6253
rect 4802 6200 4868 6201
rect 4708 6103 4718 6137
rect 4752 6103 4762 6137
rect 4508 5963 4518 5997
rect 4552 5963 4562 5997
rect 4308 5823 4318 5857
rect 4352 5823 4362 5857
rect 4108 5683 4118 5717
rect 4152 5683 4162 5717
rect 3908 5543 3918 5577
rect 3952 5543 3962 5577
rect 3708 5403 3718 5437
rect 3752 5403 3762 5437
rect 3508 5263 3518 5297
rect 3552 5263 3562 5297
rect 3308 5123 3318 5157
rect 3352 5123 3362 5157
rect 3308 5040 3362 5123
rect 3408 5201 3462 5208
rect 3408 5149 3409 5201
rect 3461 5149 3462 5201
rect 3408 5123 3418 5149
rect 3452 5123 3462 5149
rect 3408 5111 3462 5123
rect 3508 5157 3562 5263
rect 3608 5297 3662 5309
rect 3608 5271 3618 5297
rect 3652 5271 3662 5297
rect 3608 5219 3609 5271
rect 3661 5219 3662 5271
rect 3608 5212 3662 5219
rect 3708 5297 3762 5403
rect 3808 5481 3862 5488
rect 3808 5429 3809 5481
rect 3861 5429 3862 5481
rect 3808 5403 3818 5429
rect 3852 5403 3862 5429
rect 3808 5391 3862 5403
rect 3908 5437 3962 5543
rect 4008 5577 4062 5589
rect 4008 5551 4018 5577
rect 4052 5551 4062 5577
rect 4008 5499 4009 5551
rect 4061 5499 4062 5551
rect 4008 5492 4062 5499
rect 4108 5577 4162 5683
rect 4208 5761 4262 5768
rect 4208 5709 4209 5761
rect 4261 5709 4262 5761
rect 4208 5683 4218 5709
rect 4252 5683 4262 5709
rect 4208 5671 4262 5683
rect 4308 5717 4362 5823
rect 4408 5857 4462 5869
rect 4408 5831 4418 5857
rect 4452 5831 4462 5857
rect 4408 5779 4409 5831
rect 4461 5779 4462 5831
rect 4408 5772 4462 5779
rect 4508 5857 4562 5963
rect 4608 6041 4662 6048
rect 4608 5989 4609 6041
rect 4661 5989 4662 6041
rect 4608 5963 4618 5989
rect 4652 5963 4662 5989
rect 4608 5951 4662 5963
rect 4708 5997 4762 6103
rect 4808 6137 4862 6149
rect 4808 6111 4818 6137
rect 4852 6111 4862 6137
rect 4808 6059 4809 6111
rect 4861 6059 4862 6111
rect 4808 6052 4862 6059
rect 4908 6137 4962 6333
rect 5008 6411 5062 6418
rect 5008 6359 5009 6411
rect 5061 6359 5062 6411
rect 5008 6333 5018 6359
rect 5052 6333 5062 6359
rect 5008 6321 5062 6333
rect 5108 6367 5162 6473
rect 5208 6507 5262 6519
rect 5208 6481 5218 6507
rect 5252 6481 5262 6507
rect 5208 6429 5209 6481
rect 5261 6429 5262 6481
rect 5208 6422 5262 6429
rect 5308 6507 5362 6613
rect 5408 6691 5462 6698
rect 5408 6639 5409 6691
rect 5461 6639 5462 6691
rect 5408 6613 5418 6639
rect 5452 6613 5462 6639
rect 5408 6601 5462 6613
rect 5508 6647 5562 6753
rect 5608 6787 5662 6799
rect 5608 6761 5618 6787
rect 5652 6761 5662 6787
rect 5608 6709 5609 6761
rect 5661 6709 5662 6761
rect 5608 6702 5662 6709
rect 5708 6787 5762 6893
rect 5808 6971 5862 6978
rect 5808 6919 5809 6971
rect 5861 6919 5862 6971
rect 5808 6893 5818 6919
rect 5852 6893 5862 6919
rect 5808 6881 5862 6893
rect 5908 6927 5962 7033
rect 6008 7067 6062 7079
rect 6008 7041 6018 7067
rect 6052 7041 6062 7067
rect 6008 6989 6009 7041
rect 6061 6989 6062 7041
rect 6008 6982 6062 6989
rect 6108 7067 6162 7173
rect 6208 7251 6262 7258
rect 6208 7199 6209 7251
rect 6261 7199 6262 7251
rect 6208 7173 6218 7199
rect 6252 7173 6262 7199
rect 6208 7161 6262 7173
rect 6308 7207 6362 7313
rect 6408 7347 6462 7359
rect 6408 7321 6418 7347
rect 6452 7321 6462 7347
rect 6408 7269 6409 7321
rect 6461 7269 6462 7321
rect 6408 7262 6462 7269
rect 6506 7328 6516 7362
rect 6550 7328 6560 7362
rect 6506 7321 6560 7328
rect 6506 7269 6507 7321
rect 6559 7269 6560 7321
rect 6506 7262 6560 7269
rect 6506 7222 6560 7234
rect 6308 7173 6318 7207
rect 6352 7173 6362 7207
rect 6108 7033 6118 7067
rect 6152 7033 6162 7067
rect 5908 6893 5918 6927
rect 5952 6893 5962 6927
rect 5708 6753 5718 6787
rect 5752 6753 5762 6787
rect 5508 6613 5518 6647
rect 5552 6613 5562 6647
rect 5308 6473 5318 6507
rect 5352 6473 5362 6507
rect 5108 6333 5118 6367
rect 5152 6333 5162 6367
rect 5002 6269 5068 6270
rect 5002 6217 5009 6269
rect 5061 6217 5068 6269
rect 5002 6216 5068 6217
rect 4908 6103 4918 6137
rect 4952 6103 4962 6137
rect 4708 5963 4718 5997
rect 4752 5963 4762 5997
rect 4508 5823 4518 5857
rect 4552 5823 4562 5857
rect 4308 5683 4318 5717
rect 4352 5683 4362 5717
rect 4108 5543 4118 5577
rect 4152 5543 4162 5577
rect 3908 5403 3918 5437
rect 3952 5403 3962 5437
rect 3708 5263 3718 5297
rect 3752 5263 3762 5297
rect 3508 5123 3518 5157
rect 3552 5123 3562 5157
rect 3508 5040 3562 5123
rect 3608 5157 3662 5169
rect 3608 5131 3618 5157
rect 3652 5131 3662 5157
rect 3608 5079 3609 5131
rect 3661 5079 3662 5131
rect 3608 5072 3662 5079
rect 3708 5157 3762 5263
rect 3808 5341 3862 5348
rect 3808 5289 3809 5341
rect 3861 5289 3862 5341
rect 3808 5263 3818 5289
rect 3852 5263 3862 5289
rect 3808 5251 3862 5263
rect 3908 5297 3962 5403
rect 4008 5437 4062 5449
rect 4008 5411 4018 5437
rect 4052 5411 4062 5437
rect 4008 5359 4009 5411
rect 4061 5359 4062 5411
rect 4008 5352 4062 5359
rect 4108 5437 4162 5543
rect 4208 5621 4262 5628
rect 4208 5569 4209 5621
rect 4261 5569 4262 5621
rect 4208 5543 4218 5569
rect 4252 5543 4262 5569
rect 4208 5531 4262 5543
rect 4308 5577 4362 5683
rect 4408 5717 4462 5729
rect 4408 5691 4418 5717
rect 4452 5691 4462 5717
rect 4408 5639 4409 5691
rect 4461 5639 4462 5691
rect 4408 5632 4462 5639
rect 4508 5717 4562 5823
rect 4608 5901 4662 5908
rect 4608 5849 4609 5901
rect 4661 5849 4662 5901
rect 4608 5823 4618 5849
rect 4652 5823 4662 5849
rect 4608 5811 4662 5823
rect 4708 5857 4762 5963
rect 4808 5997 4862 6009
rect 4808 5971 4818 5997
rect 4852 5971 4862 5997
rect 4808 5919 4809 5971
rect 4861 5919 4862 5971
rect 4808 5912 4862 5919
rect 4908 5997 4962 6103
rect 5008 6181 5062 6188
rect 5008 6129 5009 6181
rect 5061 6129 5062 6181
rect 5008 6103 5018 6129
rect 5052 6103 5062 6129
rect 5008 6091 5062 6103
rect 5108 6137 5162 6333
rect 5208 6367 5262 6379
rect 5208 6341 5218 6367
rect 5252 6341 5262 6367
rect 5208 6289 5209 6341
rect 5261 6289 5262 6341
rect 5208 6282 5262 6289
rect 5308 6367 5362 6473
rect 5408 6551 5462 6558
rect 5408 6499 5409 6551
rect 5461 6499 5462 6551
rect 5408 6473 5418 6499
rect 5452 6473 5462 6499
rect 5408 6461 5462 6473
rect 5508 6507 5562 6613
rect 5608 6647 5662 6659
rect 5608 6621 5618 6647
rect 5652 6621 5662 6647
rect 5608 6569 5609 6621
rect 5661 6569 5662 6621
rect 5608 6562 5662 6569
rect 5708 6647 5762 6753
rect 5808 6831 5862 6838
rect 5808 6779 5809 6831
rect 5861 6779 5862 6831
rect 5808 6753 5818 6779
rect 5852 6753 5862 6779
rect 5808 6741 5862 6753
rect 5908 6787 5962 6893
rect 6008 6927 6062 6939
rect 6008 6901 6018 6927
rect 6052 6901 6062 6927
rect 6008 6849 6009 6901
rect 6061 6849 6062 6901
rect 6008 6842 6062 6849
rect 6108 6927 6162 7033
rect 6208 7111 6262 7118
rect 6208 7059 6209 7111
rect 6261 7059 6262 7111
rect 6208 7033 6218 7059
rect 6252 7033 6262 7059
rect 6208 7021 6262 7033
rect 6308 7067 6362 7173
rect 6408 7207 6462 7219
rect 6408 7181 6418 7207
rect 6452 7181 6462 7207
rect 6408 7129 6409 7181
rect 6461 7129 6462 7181
rect 6408 7122 6462 7129
rect 6506 7188 6516 7222
rect 6550 7188 6560 7222
rect 6506 7181 6560 7188
rect 6506 7129 6507 7181
rect 6559 7129 6560 7181
rect 6506 7122 6560 7129
rect 6506 7082 6560 7094
rect 6308 7033 6318 7067
rect 6352 7033 6362 7067
rect 6108 6893 6118 6927
rect 6152 6893 6162 6927
rect 5908 6753 5918 6787
rect 5952 6753 5962 6787
rect 5708 6613 5718 6647
rect 5752 6613 5762 6647
rect 5508 6473 5518 6507
rect 5552 6473 5562 6507
rect 5308 6333 5318 6367
rect 5352 6333 5362 6367
rect 5202 6253 5268 6254
rect 5202 6201 5209 6253
rect 5261 6201 5268 6253
rect 5202 6200 5268 6201
rect 5108 6103 5118 6137
rect 5152 6103 5162 6137
rect 4908 5963 4918 5997
rect 4952 5963 4962 5997
rect 4708 5823 4718 5857
rect 4752 5823 4762 5857
rect 4508 5683 4518 5717
rect 4552 5683 4562 5717
rect 4308 5543 4318 5577
rect 4352 5543 4362 5577
rect 4108 5403 4118 5437
rect 4152 5403 4162 5437
rect 3908 5263 3918 5297
rect 3952 5263 3962 5297
rect 3708 5123 3718 5157
rect 3752 5123 3762 5157
rect 3708 5040 3762 5123
rect 3808 5201 3862 5208
rect 3808 5149 3809 5201
rect 3861 5149 3862 5201
rect 3808 5123 3818 5149
rect 3852 5123 3862 5149
rect 3808 5111 3862 5123
rect 3908 5157 3962 5263
rect 4008 5297 4062 5309
rect 4008 5271 4018 5297
rect 4052 5271 4062 5297
rect 4008 5219 4009 5271
rect 4061 5219 4062 5271
rect 4008 5212 4062 5219
rect 4108 5297 4162 5403
rect 4208 5481 4262 5488
rect 4208 5429 4209 5481
rect 4261 5429 4262 5481
rect 4208 5403 4218 5429
rect 4252 5403 4262 5429
rect 4208 5391 4262 5403
rect 4308 5437 4362 5543
rect 4408 5577 4462 5589
rect 4408 5551 4418 5577
rect 4452 5551 4462 5577
rect 4408 5499 4409 5551
rect 4461 5499 4462 5551
rect 4408 5492 4462 5499
rect 4508 5577 4562 5683
rect 4608 5761 4662 5768
rect 4608 5709 4609 5761
rect 4661 5709 4662 5761
rect 4608 5683 4618 5709
rect 4652 5683 4662 5709
rect 4608 5671 4662 5683
rect 4708 5717 4762 5823
rect 4808 5857 4862 5869
rect 4808 5831 4818 5857
rect 4852 5831 4862 5857
rect 4808 5779 4809 5831
rect 4861 5779 4862 5831
rect 4808 5772 4862 5779
rect 4908 5857 4962 5963
rect 5008 6041 5062 6048
rect 5008 5989 5009 6041
rect 5061 5989 5062 6041
rect 5008 5963 5018 5989
rect 5052 5963 5062 5989
rect 5008 5951 5062 5963
rect 5108 5997 5162 6103
rect 5208 6137 5262 6149
rect 5208 6111 5218 6137
rect 5252 6111 5262 6137
rect 5208 6059 5209 6111
rect 5261 6059 5262 6111
rect 5208 6052 5262 6059
rect 5308 6137 5362 6333
rect 5408 6411 5462 6418
rect 5408 6359 5409 6411
rect 5461 6359 5462 6411
rect 5408 6333 5418 6359
rect 5452 6333 5462 6359
rect 5408 6321 5462 6333
rect 5508 6367 5562 6473
rect 5608 6507 5662 6519
rect 5608 6481 5618 6507
rect 5652 6481 5662 6507
rect 5608 6429 5609 6481
rect 5661 6429 5662 6481
rect 5608 6422 5662 6429
rect 5708 6507 5762 6613
rect 5808 6691 5862 6698
rect 5808 6639 5809 6691
rect 5861 6639 5862 6691
rect 5808 6613 5818 6639
rect 5852 6613 5862 6639
rect 5808 6601 5862 6613
rect 5908 6647 5962 6753
rect 6008 6787 6062 6799
rect 6008 6761 6018 6787
rect 6052 6761 6062 6787
rect 6008 6709 6009 6761
rect 6061 6709 6062 6761
rect 6008 6702 6062 6709
rect 6108 6787 6162 6893
rect 6208 6971 6262 6978
rect 6208 6919 6209 6971
rect 6261 6919 6262 6971
rect 6208 6893 6218 6919
rect 6252 6893 6262 6919
rect 6208 6881 6262 6893
rect 6308 6927 6362 7033
rect 6408 7067 6462 7079
rect 6408 7041 6418 7067
rect 6452 7041 6462 7067
rect 6408 6989 6409 7041
rect 6461 6989 6462 7041
rect 6408 6982 6462 6989
rect 6506 7048 6516 7082
rect 6550 7048 6560 7082
rect 6506 7041 6560 7048
rect 6506 6989 6507 7041
rect 6559 6989 6560 7041
rect 6506 6982 6560 6989
rect 6506 6942 6560 6954
rect 6308 6893 6318 6927
rect 6352 6893 6362 6927
rect 6108 6753 6118 6787
rect 6152 6753 6162 6787
rect 5908 6613 5918 6647
rect 5952 6613 5962 6647
rect 5708 6473 5718 6507
rect 5752 6473 5762 6507
rect 5508 6333 5518 6367
rect 5552 6333 5562 6367
rect 5402 6269 5468 6270
rect 5402 6217 5409 6269
rect 5461 6217 5468 6269
rect 5402 6216 5468 6217
rect 5308 6103 5318 6137
rect 5352 6103 5362 6137
rect 5108 5963 5118 5997
rect 5152 5963 5162 5997
rect 4908 5823 4918 5857
rect 4952 5823 4962 5857
rect 4708 5683 4718 5717
rect 4752 5683 4762 5717
rect 4508 5543 4518 5577
rect 4552 5543 4562 5577
rect 4308 5403 4318 5437
rect 4352 5403 4362 5437
rect 4108 5263 4118 5297
rect 4152 5263 4162 5297
rect 3908 5123 3918 5157
rect 3952 5123 3962 5157
rect 3908 5040 3962 5123
rect 4008 5157 4062 5169
rect 4008 5131 4018 5157
rect 4052 5131 4062 5157
rect 4008 5079 4009 5131
rect 4061 5079 4062 5131
rect 4008 5072 4062 5079
rect 4108 5157 4162 5263
rect 4208 5341 4262 5348
rect 4208 5289 4209 5341
rect 4261 5289 4262 5341
rect 4208 5263 4218 5289
rect 4252 5263 4262 5289
rect 4208 5251 4262 5263
rect 4308 5297 4362 5403
rect 4408 5437 4462 5449
rect 4408 5411 4418 5437
rect 4452 5411 4462 5437
rect 4408 5359 4409 5411
rect 4461 5359 4462 5411
rect 4408 5352 4462 5359
rect 4508 5437 4562 5543
rect 4608 5621 4662 5628
rect 4608 5569 4609 5621
rect 4661 5569 4662 5621
rect 4608 5543 4618 5569
rect 4652 5543 4662 5569
rect 4608 5531 4662 5543
rect 4708 5577 4762 5683
rect 4808 5717 4862 5729
rect 4808 5691 4818 5717
rect 4852 5691 4862 5717
rect 4808 5639 4809 5691
rect 4861 5639 4862 5691
rect 4808 5632 4862 5639
rect 4908 5717 4962 5823
rect 5008 5901 5062 5908
rect 5008 5849 5009 5901
rect 5061 5849 5062 5901
rect 5008 5823 5018 5849
rect 5052 5823 5062 5849
rect 5008 5811 5062 5823
rect 5108 5857 5162 5963
rect 5208 5997 5262 6009
rect 5208 5971 5218 5997
rect 5252 5971 5262 5997
rect 5208 5919 5209 5971
rect 5261 5919 5262 5971
rect 5208 5912 5262 5919
rect 5308 5997 5362 6103
rect 5408 6181 5462 6188
rect 5408 6129 5409 6181
rect 5461 6129 5462 6181
rect 5408 6103 5418 6129
rect 5452 6103 5462 6129
rect 5408 6091 5462 6103
rect 5508 6137 5562 6333
rect 5608 6367 5662 6379
rect 5608 6341 5618 6367
rect 5652 6341 5662 6367
rect 5608 6289 5609 6341
rect 5661 6289 5662 6341
rect 5608 6282 5662 6289
rect 5708 6367 5762 6473
rect 5808 6551 5862 6558
rect 5808 6499 5809 6551
rect 5861 6499 5862 6551
rect 5808 6473 5818 6499
rect 5852 6473 5862 6499
rect 5808 6461 5862 6473
rect 5908 6507 5962 6613
rect 6008 6647 6062 6659
rect 6008 6621 6018 6647
rect 6052 6621 6062 6647
rect 6008 6569 6009 6621
rect 6061 6569 6062 6621
rect 6008 6562 6062 6569
rect 6108 6647 6162 6753
rect 6208 6831 6262 6838
rect 6208 6779 6209 6831
rect 6261 6779 6262 6831
rect 6208 6753 6218 6779
rect 6252 6753 6262 6779
rect 6208 6741 6262 6753
rect 6308 6787 6362 6893
rect 6408 6927 6462 6939
rect 6408 6901 6418 6927
rect 6452 6901 6462 6927
rect 6408 6849 6409 6901
rect 6461 6849 6462 6901
rect 6408 6842 6462 6849
rect 6506 6908 6516 6942
rect 6550 6908 6560 6942
rect 6506 6901 6560 6908
rect 6506 6849 6507 6901
rect 6559 6849 6560 6901
rect 6506 6842 6560 6849
rect 6506 6802 6560 6814
rect 6308 6753 6318 6787
rect 6352 6753 6362 6787
rect 6108 6613 6118 6647
rect 6152 6613 6162 6647
rect 5908 6473 5918 6507
rect 5952 6473 5962 6507
rect 5708 6333 5718 6367
rect 5752 6333 5762 6367
rect 5602 6253 5668 6254
rect 5602 6201 5609 6253
rect 5661 6201 5668 6253
rect 5602 6200 5668 6201
rect 5508 6103 5518 6137
rect 5552 6103 5562 6137
rect 5308 5963 5318 5997
rect 5352 5963 5362 5997
rect 5108 5823 5118 5857
rect 5152 5823 5162 5857
rect 4908 5683 4918 5717
rect 4952 5683 4962 5717
rect 4708 5543 4718 5577
rect 4752 5543 4762 5577
rect 4508 5403 4518 5437
rect 4552 5403 4562 5437
rect 4308 5263 4318 5297
rect 4352 5263 4362 5297
rect 4108 5123 4118 5157
rect 4152 5123 4162 5157
rect 4108 5040 4162 5123
rect 4208 5201 4262 5208
rect 4208 5149 4209 5201
rect 4261 5149 4262 5201
rect 4208 5123 4218 5149
rect 4252 5123 4262 5149
rect 4208 5111 4262 5123
rect 4308 5157 4362 5263
rect 4408 5297 4462 5309
rect 4408 5271 4418 5297
rect 4452 5271 4462 5297
rect 4408 5219 4409 5271
rect 4461 5219 4462 5271
rect 4408 5212 4462 5219
rect 4508 5297 4562 5403
rect 4608 5481 4662 5488
rect 4608 5429 4609 5481
rect 4661 5429 4662 5481
rect 4608 5403 4618 5429
rect 4652 5403 4662 5429
rect 4608 5391 4662 5403
rect 4708 5437 4762 5543
rect 4808 5577 4862 5589
rect 4808 5551 4818 5577
rect 4852 5551 4862 5577
rect 4808 5499 4809 5551
rect 4861 5499 4862 5551
rect 4808 5492 4862 5499
rect 4908 5577 4962 5683
rect 5008 5761 5062 5768
rect 5008 5709 5009 5761
rect 5061 5709 5062 5761
rect 5008 5683 5018 5709
rect 5052 5683 5062 5709
rect 5008 5671 5062 5683
rect 5108 5717 5162 5823
rect 5208 5857 5262 5869
rect 5208 5831 5218 5857
rect 5252 5831 5262 5857
rect 5208 5779 5209 5831
rect 5261 5779 5262 5831
rect 5208 5772 5262 5779
rect 5308 5857 5362 5963
rect 5408 6041 5462 6048
rect 5408 5989 5409 6041
rect 5461 5989 5462 6041
rect 5408 5963 5418 5989
rect 5452 5963 5462 5989
rect 5408 5951 5462 5963
rect 5508 5997 5562 6103
rect 5608 6137 5662 6149
rect 5608 6111 5618 6137
rect 5652 6111 5662 6137
rect 5608 6059 5609 6111
rect 5661 6059 5662 6111
rect 5608 6052 5662 6059
rect 5708 6137 5762 6333
rect 5808 6411 5862 6418
rect 5808 6359 5809 6411
rect 5861 6359 5862 6411
rect 5808 6333 5818 6359
rect 5852 6333 5862 6359
rect 5808 6321 5862 6333
rect 5908 6367 5962 6473
rect 6008 6507 6062 6519
rect 6008 6481 6018 6507
rect 6052 6481 6062 6507
rect 6008 6429 6009 6481
rect 6061 6429 6062 6481
rect 6008 6422 6062 6429
rect 6108 6507 6162 6613
rect 6208 6691 6262 6698
rect 6208 6639 6209 6691
rect 6261 6639 6262 6691
rect 6208 6613 6218 6639
rect 6252 6613 6262 6639
rect 6208 6601 6262 6613
rect 6308 6647 6362 6753
rect 6408 6787 6462 6799
rect 6408 6761 6418 6787
rect 6452 6761 6462 6787
rect 6408 6709 6409 6761
rect 6461 6709 6462 6761
rect 6408 6702 6462 6709
rect 6506 6768 6516 6802
rect 6550 6768 6560 6802
rect 6506 6761 6560 6768
rect 6506 6709 6507 6761
rect 6559 6709 6560 6761
rect 6506 6702 6560 6709
rect 6506 6662 6560 6674
rect 6308 6613 6318 6647
rect 6352 6613 6362 6647
rect 6108 6473 6118 6507
rect 6152 6473 6162 6507
rect 5908 6333 5918 6367
rect 5952 6333 5962 6367
rect 5802 6269 5868 6270
rect 5802 6217 5809 6269
rect 5861 6217 5868 6269
rect 5802 6216 5868 6217
rect 5708 6103 5718 6137
rect 5752 6103 5762 6137
rect 5508 5963 5518 5997
rect 5552 5963 5562 5997
rect 5308 5823 5318 5857
rect 5352 5823 5362 5857
rect 5108 5683 5118 5717
rect 5152 5683 5162 5717
rect 4908 5543 4918 5577
rect 4952 5543 4962 5577
rect 4708 5403 4718 5437
rect 4752 5403 4762 5437
rect 4508 5263 4518 5297
rect 4552 5263 4562 5297
rect 4308 5123 4318 5157
rect 4352 5123 4362 5157
rect 4308 5040 4362 5123
rect 4408 5157 4462 5169
rect 4408 5131 4418 5157
rect 4452 5131 4462 5157
rect 4408 5079 4409 5131
rect 4461 5079 4462 5131
rect 4408 5072 4462 5079
rect 4508 5157 4562 5263
rect 4608 5341 4662 5348
rect 4608 5289 4609 5341
rect 4661 5289 4662 5341
rect 4608 5263 4618 5289
rect 4652 5263 4662 5289
rect 4608 5251 4662 5263
rect 4708 5297 4762 5403
rect 4808 5437 4862 5449
rect 4808 5411 4818 5437
rect 4852 5411 4862 5437
rect 4808 5359 4809 5411
rect 4861 5359 4862 5411
rect 4808 5352 4862 5359
rect 4908 5437 4962 5543
rect 5008 5621 5062 5628
rect 5008 5569 5009 5621
rect 5061 5569 5062 5621
rect 5008 5543 5018 5569
rect 5052 5543 5062 5569
rect 5008 5531 5062 5543
rect 5108 5577 5162 5683
rect 5208 5717 5262 5729
rect 5208 5691 5218 5717
rect 5252 5691 5262 5717
rect 5208 5639 5209 5691
rect 5261 5639 5262 5691
rect 5208 5632 5262 5639
rect 5308 5717 5362 5823
rect 5408 5901 5462 5908
rect 5408 5849 5409 5901
rect 5461 5849 5462 5901
rect 5408 5823 5418 5849
rect 5452 5823 5462 5849
rect 5408 5811 5462 5823
rect 5508 5857 5562 5963
rect 5608 5997 5662 6009
rect 5608 5971 5618 5997
rect 5652 5971 5662 5997
rect 5608 5919 5609 5971
rect 5661 5919 5662 5971
rect 5608 5912 5662 5919
rect 5708 5997 5762 6103
rect 5808 6181 5862 6188
rect 5808 6129 5809 6181
rect 5861 6129 5862 6181
rect 5808 6103 5818 6129
rect 5852 6103 5862 6129
rect 5808 6091 5862 6103
rect 5908 6137 5962 6333
rect 6008 6367 6062 6379
rect 6008 6341 6018 6367
rect 6052 6341 6062 6367
rect 6008 6289 6009 6341
rect 6061 6289 6062 6341
rect 6008 6282 6062 6289
rect 6108 6367 6162 6473
rect 6208 6551 6262 6558
rect 6208 6499 6209 6551
rect 6261 6499 6262 6551
rect 6208 6473 6218 6499
rect 6252 6473 6262 6499
rect 6208 6461 6262 6473
rect 6308 6507 6362 6613
rect 6408 6647 6462 6659
rect 6408 6621 6418 6647
rect 6452 6621 6462 6647
rect 6408 6569 6409 6621
rect 6461 6569 6462 6621
rect 6408 6562 6462 6569
rect 6506 6628 6516 6662
rect 6550 6628 6560 6662
rect 6506 6621 6560 6628
rect 6506 6569 6507 6621
rect 6559 6569 6560 6621
rect 6506 6562 6560 6569
rect 6506 6522 6560 6534
rect 6308 6473 6318 6507
rect 6352 6473 6362 6507
rect 6108 6333 6118 6367
rect 6152 6333 6162 6367
rect 6002 6253 6068 6254
rect 6002 6201 6009 6253
rect 6061 6201 6068 6253
rect 6002 6200 6068 6201
rect 5908 6103 5918 6137
rect 5952 6103 5962 6137
rect 5708 5963 5718 5997
rect 5752 5963 5762 5997
rect 5508 5823 5518 5857
rect 5552 5823 5562 5857
rect 5308 5683 5318 5717
rect 5352 5683 5362 5717
rect 5108 5543 5118 5577
rect 5152 5543 5162 5577
rect 4908 5403 4918 5437
rect 4952 5403 4962 5437
rect 4708 5263 4718 5297
rect 4752 5263 4762 5297
rect 4508 5123 4518 5157
rect 4552 5123 4562 5157
rect 4508 5040 4562 5123
rect 4608 5201 4662 5208
rect 4608 5149 4609 5201
rect 4661 5149 4662 5201
rect 4608 5123 4618 5149
rect 4652 5123 4662 5149
rect 4608 5111 4662 5123
rect 4708 5157 4762 5263
rect 4808 5297 4862 5309
rect 4808 5271 4818 5297
rect 4852 5271 4862 5297
rect 4808 5219 4809 5271
rect 4861 5219 4862 5271
rect 4808 5212 4862 5219
rect 4908 5297 4962 5403
rect 5008 5481 5062 5488
rect 5008 5429 5009 5481
rect 5061 5429 5062 5481
rect 5008 5403 5018 5429
rect 5052 5403 5062 5429
rect 5008 5391 5062 5403
rect 5108 5437 5162 5543
rect 5208 5577 5262 5589
rect 5208 5551 5218 5577
rect 5252 5551 5262 5577
rect 5208 5499 5209 5551
rect 5261 5499 5262 5551
rect 5208 5492 5262 5499
rect 5308 5577 5362 5683
rect 5408 5761 5462 5768
rect 5408 5709 5409 5761
rect 5461 5709 5462 5761
rect 5408 5683 5418 5709
rect 5452 5683 5462 5709
rect 5408 5671 5462 5683
rect 5508 5717 5562 5823
rect 5608 5857 5662 5869
rect 5608 5831 5618 5857
rect 5652 5831 5662 5857
rect 5608 5779 5609 5831
rect 5661 5779 5662 5831
rect 5608 5772 5662 5779
rect 5708 5857 5762 5963
rect 5808 6041 5862 6048
rect 5808 5989 5809 6041
rect 5861 5989 5862 6041
rect 5808 5963 5818 5989
rect 5852 5963 5862 5989
rect 5808 5951 5862 5963
rect 5908 5997 5962 6103
rect 6008 6137 6062 6149
rect 6008 6111 6018 6137
rect 6052 6111 6062 6137
rect 6008 6059 6009 6111
rect 6061 6059 6062 6111
rect 6008 6052 6062 6059
rect 6108 6137 6162 6333
rect 6208 6411 6262 6418
rect 6208 6359 6209 6411
rect 6261 6359 6262 6411
rect 6208 6333 6218 6359
rect 6252 6333 6262 6359
rect 6208 6321 6262 6333
rect 6308 6367 6362 6473
rect 6408 6507 6462 6519
rect 6408 6481 6418 6507
rect 6452 6481 6462 6507
rect 6408 6429 6409 6481
rect 6461 6429 6462 6481
rect 6408 6422 6462 6429
rect 6506 6488 6516 6522
rect 6550 6488 6560 6522
rect 6506 6481 6560 6488
rect 6506 6429 6507 6481
rect 6559 6429 6560 6481
rect 6506 6422 6560 6429
rect 6506 6382 6560 6394
rect 6308 6333 6318 6367
rect 6352 6333 6362 6367
rect 6202 6269 6268 6270
rect 6202 6217 6209 6269
rect 6261 6217 6268 6269
rect 6202 6216 6268 6217
rect 6108 6103 6118 6137
rect 6152 6103 6162 6137
rect 5908 5963 5918 5997
rect 5952 5963 5962 5997
rect 5708 5823 5718 5857
rect 5752 5823 5762 5857
rect 5508 5683 5518 5717
rect 5552 5683 5562 5717
rect 5308 5543 5318 5577
rect 5352 5543 5362 5577
rect 5108 5403 5118 5437
rect 5152 5403 5162 5437
rect 4908 5263 4918 5297
rect 4952 5263 4962 5297
rect 4708 5123 4718 5157
rect 4752 5123 4762 5157
rect 4708 5040 4762 5123
rect 4808 5157 4862 5169
rect 4808 5131 4818 5157
rect 4852 5131 4862 5157
rect 4808 5079 4809 5131
rect 4861 5079 4862 5131
rect 4808 5072 4862 5079
rect 4908 5157 4962 5263
rect 5008 5341 5062 5348
rect 5008 5289 5009 5341
rect 5061 5289 5062 5341
rect 5008 5263 5018 5289
rect 5052 5263 5062 5289
rect 5008 5251 5062 5263
rect 5108 5297 5162 5403
rect 5208 5437 5262 5449
rect 5208 5411 5218 5437
rect 5252 5411 5262 5437
rect 5208 5359 5209 5411
rect 5261 5359 5262 5411
rect 5208 5352 5262 5359
rect 5308 5437 5362 5543
rect 5408 5621 5462 5628
rect 5408 5569 5409 5621
rect 5461 5569 5462 5621
rect 5408 5543 5418 5569
rect 5452 5543 5462 5569
rect 5408 5531 5462 5543
rect 5508 5577 5562 5683
rect 5608 5717 5662 5729
rect 5608 5691 5618 5717
rect 5652 5691 5662 5717
rect 5608 5639 5609 5691
rect 5661 5639 5662 5691
rect 5608 5632 5662 5639
rect 5708 5717 5762 5823
rect 5808 5901 5862 5908
rect 5808 5849 5809 5901
rect 5861 5849 5862 5901
rect 5808 5823 5818 5849
rect 5852 5823 5862 5849
rect 5808 5811 5862 5823
rect 5908 5857 5962 5963
rect 6008 5997 6062 6009
rect 6008 5971 6018 5997
rect 6052 5971 6062 5997
rect 6008 5919 6009 5971
rect 6061 5919 6062 5971
rect 6008 5912 6062 5919
rect 6108 5997 6162 6103
rect 6208 6181 6262 6188
rect 6208 6129 6209 6181
rect 6261 6129 6262 6181
rect 6208 6103 6218 6129
rect 6252 6103 6262 6129
rect 6208 6091 6262 6103
rect 6308 6137 6362 6333
rect 6408 6367 6462 6379
rect 6408 6341 6418 6367
rect 6452 6341 6462 6367
rect 6408 6289 6409 6341
rect 6461 6289 6462 6341
rect 6408 6282 6462 6289
rect 6506 6348 6516 6382
rect 6550 6348 6560 6382
rect 6506 6341 6560 6348
rect 6506 6289 6507 6341
rect 6559 6289 6560 6341
rect 6506 6282 6560 6289
rect 6590 6247 6620 7411
rect 6504 6241 6620 6247
rect 6504 6207 6516 6241
rect 6550 6207 6620 6241
rect 6504 6201 6620 6207
rect 6506 6152 6560 6164
rect 6308 6103 6318 6137
rect 6352 6103 6362 6137
rect 6108 5963 6118 5997
rect 6152 5963 6162 5997
rect 5908 5823 5918 5857
rect 5952 5823 5962 5857
rect 5708 5683 5718 5717
rect 5752 5683 5762 5717
rect 5508 5543 5518 5577
rect 5552 5543 5562 5577
rect 5308 5403 5318 5437
rect 5352 5403 5362 5437
rect 5108 5263 5118 5297
rect 5152 5263 5162 5297
rect 4908 5123 4918 5157
rect 4952 5123 4962 5157
rect 4908 5040 4962 5123
rect 5008 5201 5062 5208
rect 5008 5149 5009 5201
rect 5061 5149 5062 5201
rect 5008 5123 5018 5149
rect 5052 5123 5062 5149
rect 5008 5111 5062 5123
rect 5108 5157 5162 5263
rect 5208 5297 5262 5309
rect 5208 5271 5218 5297
rect 5252 5271 5262 5297
rect 5208 5219 5209 5271
rect 5261 5219 5262 5271
rect 5208 5212 5262 5219
rect 5308 5297 5362 5403
rect 5408 5481 5462 5488
rect 5408 5429 5409 5481
rect 5461 5429 5462 5481
rect 5408 5403 5418 5429
rect 5452 5403 5462 5429
rect 5408 5391 5462 5403
rect 5508 5437 5562 5543
rect 5608 5577 5662 5589
rect 5608 5551 5618 5577
rect 5652 5551 5662 5577
rect 5608 5499 5609 5551
rect 5661 5499 5662 5551
rect 5608 5492 5662 5499
rect 5708 5577 5762 5683
rect 5808 5761 5862 5768
rect 5808 5709 5809 5761
rect 5861 5709 5862 5761
rect 5808 5683 5818 5709
rect 5852 5683 5862 5709
rect 5808 5671 5862 5683
rect 5908 5717 5962 5823
rect 6008 5857 6062 5869
rect 6008 5831 6018 5857
rect 6052 5831 6062 5857
rect 6008 5779 6009 5831
rect 6061 5779 6062 5831
rect 6008 5772 6062 5779
rect 6108 5857 6162 5963
rect 6208 6041 6262 6048
rect 6208 5989 6209 6041
rect 6261 5989 6262 6041
rect 6208 5963 6218 5989
rect 6252 5963 6262 5989
rect 6208 5951 6262 5963
rect 6308 5997 6362 6103
rect 6408 6137 6462 6149
rect 6408 6111 6418 6137
rect 6452 6111 6462 6137
rect 6408 6059 6409 6111
rect 6461 6059 6462 6111
rect 6408 6052 6462 6059
rect 6506 6118 6516 6152
rect 6550 6118 6560 6152
rect 6506 6111 6560 6118
rect 6506 6059 6507 6111
rect 6559 6059 6560 6111
rect 6506 6052 6560 6059
rect 6506 6012 6560 6024
rect 6308 5963 6318 5997
rect 6352 5963 6362 5997
rect 6108 5823 6118 5857
rect 6152 5823 6162 5857
rect 5908 5683 5918 5717
rect 5952 5683 5962 5717
rect 5708 5543 5718 5577
rect 5752 5543 5762 5577
rect 5508 5403 5518 5437
rect 5552 5403 5562 5437
rect 5308 5263 5318 5297
rect 5352 5263 5362 5297
rect 5108 5123 5118 5157
rect 5152 5123 5162 5157
rect 5108 5040 5162 5123
rect 5208 5157 5262 5169
rect 5208 5131 5218 5157
rect 5252 5131 5262 5157
rect 5208 5079 5209 5131
rect 5261 5079 5262 5131
rect 5208 5072 5262 5079
rect 5308 5157 5362 5263
rect 5408 5341 5462 5348
rect 5408 5289 5409 5341
rect 5461 5289 5462 5341
rect 5408 5263 5418 5289
rect 5452 5263 5462 5289
rect 5408 5251 5462 5263
rect 5508 5297 5562 5403
rect 5608 5437 5662 5449
rect 5608 5411 5618 5437
rect 5652 5411 5662 5437
rect 5608 5359 5609 5411
rect 5661 5359 5662 5411
rect 5608 5352 5662 5359
rect 5708 5437 5762 5543
rect 5808 5621 5862 5628
rect 5808 5569 5809 5621
rect 5861 5569 5862 5621
rect 5808 5543 5818 5569
rect 5852 5543 5862 5569
rect 5808 5531 5862 5543
rect 5908 5577 5962 5683
rect 6008 5717 6062 5729
rect 6008 5691 6018 5717
rect 6052 5691 6062 5717
rect 6008 5639 6009 5691
rect 6061 5639 6062 5691
rect 6008 5632 6062 5639
rect 6108 5717 6162 5823
rect 6208 5901 6262 5908
rect 6208 5849 6209 5901
rect 6261 5849 6262 5901
rect 6208 5823 6218 5849
rect 6252 5823 6262 5849
rect 6208 5811 6262 5823
rect 6308 5857 6362 5963
rect 6408 5997 6462 6009
rect 6408 5971 6418 5997
rect 6452 5971 6462 5997
rect 6408 5919 6409 5971
rect 6461 5919 6462 5971
rect 6408 5912 6462 5919
rect 6506 5978 6516 6012
rect 6550 5978 6560 6012
rect 6506 5971 6560 5978
rect 6506 5919 6507 5971
rect 6559 5919 6560 5971
rect 6506 5912 6560 5919
rect 6506 5872 6560 5884
rect 6308 5823 6318 5857
rect 6352 5823 6362 5857
rect 6108 5683 6118 5717
rect 6152 5683 6162 5717
rect 5908 5543 5918 5577
rect 5952 5543 5962 5577
rect 5708 5403 5718 5437
rect 5752 5403 5762 5437
rect 5508 5263 5518 5297
rect 5552 5263 5562 5297
rect 5308 5123 5318 5157
rect 5352 5123 5362 5157
rect 5308 5040 5362 5123
rect 5408 5201 5462 5208
rect 5408 5149 5409 5201
rect 5461 5149 5462 5201
rect 5408 5123 5418 5149
rect 5452 5123 5462 5149
rect 5408 5111 5462 5123
rect 5508 5157 5562 5263
rect 5608 5297 5662 5309
rect 5608 5271 5618 5297
rect 5652 5271 5662 5297
rect 5608 5219 5609 5271
rect 5661 5219 5662 5271
rect 5608 5212 5662 5219
rect 5708 5297 5762 5403
rect 5808 5481 5862 5488
rect 5808 5429 5809 5481
rect 5861 5429 5862 5481
rect 5808 5403 5818 5429
rect 5852 5403 5862 5429
rect 5808 5391 5862 5403
rect 5908 5437 5962 5543
rect 6008 5577 6062 5589
rect 6008 5551 6018 5577
rect 6052 5551 6062 5577
rect 6008 5499 6009 5551
rect 6061 5499 6062 5551
rect 6008 5492 6062 5499
rect 6108 5577 6162 5683
rect 6208 5761 6262 5768
rect 6208 5709 6209 5761
rect 6261 5709 6262 5761
rect 6208 5683 6218 5709
rect 6252 5683 6262 5709
rect 6208 5671 6262 5683
rect 6308 5717 6362 5823
rect 6408 5857 6462 5869
rect 6408 5831 6418 5857
rect 6452 5831 6462 5857
rect 6408 5779 6409 5831
rect 6461 5779 6462 5831
rect 6408 5772 6462 5779
rect 6506 5838 6516 5872
rect 6550 5838 6560 5872
rect 6506 5831 6560 5838
rect 6506 5779 6507 5831
rect 6559 5779 6560 5831
rect 6506 5772 6560 5779
rect 6506 5732 6560 5744
rect 6308 5683 6318 5717
rect 6352 5683 6362 5717
rect 6108 5543 6118 5577
rect 6152 5543 6162 5577
rect 5908 5403 5918 5437
rect 5952 5403 5962 5437
rect 5708 5263 5718 5297
rect 5752 5263 5762 5297
rect 5508 5123 5518 5157
rect 5552 5123 5562 5157
rect 5508 5040 5562 5123
rect 5608 5157 5662 5169
rect 5608 5131 5618 5157
rect 5652 5131 5662 5157
rect 5608 5079 5609 5131
rect 5661 5079 5662 5131
rect 5608 5072 5662 5079
rect 5708 5157 5762 5263
rect 5808 5341 5862 5348
rect 5808 5289 5809 5341
rect 5861 5289 5862 5341
rect 5808 5263 5818 5289
rect 5852 5263 5862 5289
rect 5808 5251 5862 5263
rect 5908 5297 5962 5403
rect 6008 5437 6062 5449
rect 6008 5411 6018 5437
rect 6052 5411 6062 5437
rect 6008 5359 6009 5411
rect 6061 5359 6062 5411
rect 6008 5352 6062 5359
rect 6108 5437 6162 5543
rect 6208 5621 6262 5628
rect 6208 5569 6209 5621
rect 6261 5569 6262 5621
rect 6208 5543 6218 5569
rect 6252 5543 6262 5569
rect 6208 5531 6262 5543
rect 6308 5577 6362 5683
rect 6408 5717 6462 5729
rect 6408 5691 6418 5717
rect 6452 5691 6462 5717
rect 6408 5639 6409 5691
rect 6461 5639 6462 5691
rect 6408 5632 6462 5639
rect 6506 5698 6516 5732
rect 6550 5698 6560 5732
rect 6506 5691 6560 5698
rect 6506 5639 6507 5691
rect 6559 5639 6560 5691
rect 6506 5632 6560 5639
rect 6506 5592 6560 5604
rect 6308 5543 6318 5577
rect 6352 5543 6362 5577
rect 6108 5403 6118 5437
rect 6152 5403 6162 5437
rect 5908 5263 5918 5297
rect 5952 5263 5962 5297
rect 5708 5123 5718 5157
rect 5752 5123 5762 5157
rect 5708 5040 5762 5123
rect 5808 5201 5862 5208
rect 5808 5149 5809 5201
rect 5861 5149 5862 5201
rect 5808 5123 5818 5149
rect 5852 5123 5862 5149
rect 5808 5111 5862 5123
rect 5908 5157 5962 5263
rect 6008 5297 6062 5309
rect 6008 5271 6018 5297
rect 6052 5271 6062 5297
rect 6008 5219 6009 5271
rect 6061 5219 6062 5271
rect 6008 5212 6062 5219
rect 6108 5297 6162 5403
rect 6208 5481 6262 5488
rect 6208 5429 6209 5481
rect 6261 5429 6262 5481
rect 6208 5403 6218 5429
rect 6252 5403 6262 5429
rect 6208 5391 6262 5403
rect 6308 5437 6362 5543
rect 6408 5577 6462 5589
rect 6408 5551 6418 5577
rect 6452 5551 6462 5577
rect 6408 5499 6409 5551
rect 6461 5499 6462 5551
rect 6408 5492 6462 5499
rect 6506 5558 6516 5592
rect 6550 5558 6560 5592
rect 6506 5551 6560 5558
rect 6506 5499 6507 5551
rect 6559 5499 6560 5551
rect 6506 5492 6560 5499
rect 6506 5452 6560 5464
rect 6308 5403 6318 5437
rect 6352 5403 6362 5437
rect 6108 5263 6118 5297
rect 6152 5263 6162 5297
rect 5908 5123 5918 5157
rect 5952 5123 5962 5157
rect 5908 5040 5962 5123
rect 6008 5157 6062 5169
rect 6008 5131 6018 5157
rect 6052 5131 6062 5157
rect 6008 5079 6009 5131
rect 6061 5079 6062 5131
rect 6008 5072 6062 5079
rect 6108 5157 6162 5263
rect 6208 5341 6262 5348
rect 6208 5289 6209 5341
rect 6261 5289 6262 5341
rect 6208 5263 6218 5289
rect 6252 5263 6262 5289
rect 6208 5251 6262 5263
rect 6308 5297 6362 5403
rect 6408 5437 6462 5449
rect 6408 5411 6418 5437
rect 6452 5411 6462 5437
rect 6408 5359 6409 5411
rect 6461 5359 6462 5411
rect 6408 5352 6462 5359
rect 6506 5418 6516 5452
rect 6550 5418 6560 5452
rect 6506 5411 6560 5418
rect 6506 5359 6507 5411
rect 6559 5359 6560 5411
rect 6506 5352 6560 5359
rect 6506 5312 6560 5324
rect 6308 5263 6318 5297
rect 6352 5263 6362 5297
rect 6108 5123 6118 5157
rect 6152 5123 6162 5157
rect 6108 5040 6162 5123
rect 6208 5201 6262 5208
rect 6208 5149 6209 5201
rect 6261 5149 6262 5201
rect 6208 5123 6218 5149
rect 6252 5123 6262 5149
rect 6208 5111 6262 5123
rect 6308 5157 6362 5263
rect 6408 5297 6462 5309
rect 6408 5271 6418 5297
rect 6452 5271 6462 5297
rect 6408 5219 6409 5271
rect 6461 5219 6462 5271
rect 6408 5212 6462 5219
rect 6506 5278 6516 5312
rect 6550 5278 6560 5312
rect 6506 5271 6560 5278
rect 6506 5219 6507 5271
rect 6559 5219 6560 5271
rect 6506 5212 6560 5219
rect 6506 5172 6560 5184
rect 6308 5123 6318 5157
rect 6352 5123 6362 5157
rect 6308 5040 6362 5123
rect 6408 5157 6462 5169
rect 6408 5131 6418 5157
rect 6452 5131 6462 5157
rect 6408 5079 6409 5131
rect 6461 5079 6462 5131
rect 6408 5072 6462 5079
rect 6506 5138 6516 5172
rect 6550 5138 6560 5172
rect 6506 5131 6560 5138
rect 6506 5079 6507 5131
rect 6559 5079 6560 5131
rect 6506 5072 6560 5079
rect 35 5017 6435 5040
rect 35 4983 118 5017
rect 152 4983 318 5017
rect 352 4983 518 5017
rect 552 4983 718 5017
rect 752 4983 918 5017
rect 952 4983 1118 5017
rect 1152 4983 1318 5017
rect 1352 4983 1518 5017
rect 1552 4983 1718 5017
rect 1752 4983 1918 5017
rect 1952 4983 2118 5017
rect 2152 4983 2318 5017
rect 2352 4983 2518 5017
rect 2552 4983 2718 5017
rect 2752 4983 2918 5017
rect 2952 4983 3118 5017
rect 3152 4983 3318 5017
rect 3352 4983 3518 5017
rect 3552 4983 3718 5017
rect 3752 4983 3918 5017
rect 3952 4983 4118 5017
rect 4152 4983 4318 5017
rect 4352 4983 4518 5017
rect 4552 4983 4718 5017
rect 4752 4983 4918 5017
rect 4952 4983 5118 5017
rect 5152 4983 5318 5017
rect 5352 4983 5518 5017
rect 5552 4983 5718 5017
rect 5752 4983 5918 5017
rect 5952 4983 6118 5017
rect 6152 4983 6318 5017
rect 6352 4983 6435 5017
rect 35 4960 6435 4983
rect 2 4903 68 4904
rect 2 4851 9 4903
rect 61 4851 68 4903
rect 2 4850 68 4851
rect 8 4787 62 4799
rect 8 4761 18 4787
rect 52 4761 62 4787
rect 8 4709 9 4761
rect 61 4709 62 4761
rect 8 4702 62 4709
rect 108 4787 162 4960
rect 202 4919 268 4920
rect 202 4867 209 4919
rect 261 4867 268 4919
rect 202 4866 268 4867
rect 108 4753 118 4787
rect 152 4753 162 4787
rect 8 4647 62 4659
rect 8 4621 18 4647
rect 52 4621 62 4647
rect 8 4569 9 4621
rect 61 4569 62 4621
rect 8 4562 62 4569
rect 108 4647 162 4753
rect 208 4831 262 4838
rect 208 4779 209 4831
rect 261 4779 262 4831
rect 208 4753 218 4779
rect 252 4753 262 4779
rect 208 4741 262 4753
rect 308 4787 362 4960
rect 402 4903 468 4904
rect 402 4851 409 4903
rect 461 4851 468 4903
rect 402 4850 468 4851
rect 308 4753 318 4787
rect 352 4753 362 4787
rect 108 4613 118 4647
rect 152 4613 162 4647
rect 8 4507 62 4519
rect 8 4481 18 4507
rect 52 4481 62 4507
rect 8 4429 9 4481
rect 61 4429 62 4481
rect 8 4422 62 4429
rect 108 4507 162 4613
rect 208 4691 262 4698
rect 208 4639 209 4691
rect 261 4639 262 4691
rect 208 4613 218 4639
rect 252 4613 262 4639
rect 208 4601 262 4613
rect 308 4647 362 4753
rect 408 4787 462 4799
rect 408 4761 418 4787
rect 452 4761 462 4787
rect 408 4709 409 4761
rect 461 4709 462 4761
rect 408 4702 462 4709
rect 508 4787 562 4960
rect 602 4919 668 4920
rect 602 4867 609 4919
rect 661 4867 668 4919
rect 602 4866 668 4867
rect 508 4753 518 4787
rect 552 4753 562 4787
rect 308 4613 318 4647
rect 352 4613 362 4647
rect 108 4473 118 4507
rect 152 4473 162 4507
rect 8 4367 62 4379
rect 8 4341 18 4367
rect 52 4341 62 4367
rect 8 4289 9 4341
rect 61 4289 62 4341
rect 8 4282 62 4289
rect 108 4367 162 4473
rect 208 4551 262 4558
rect 208 4499 209 4551
rect 261 4499 262 4551
rect 208 4473 218 4499
rect 252 4473 262 4499
rect 208 4461 262 4473
rect 308 4507 362 4613
rect 408 4647 462 4659
rect 408 4621 418 4647
rect 452 4621 462 4647
rect 408 4569 409 4621
rect 461 4569 462 4621
rect 408 4562 462 4569
rect 508 4647 562 4753
rect 608 4831 662 4838
rect 608 4779 609 4831
rect 661 4779 662 4831
rect 608 4753 618 4779
rect 652 4753 662 4779
rect 608 4741 662 4753
rect 708 4787 762 4960
rect 802 4903 868 4904
rect 802 4851 809 4903
rect 861 4851 868 4903
rect 802 4850 868 4851
rect 708 4753 718 4787
rect 752 4753 762 4787
rect 508 4613 518 4647
rect 552 4613 562 4647
rect 308 4473 318 4507
rect 352 4473 362 4507
rect 108 4333 118 4367
rect 152 4333 162 4367
rect 8 4227 62 4239
rect 8 4201 18 4227
rect 52 4201 62 4227
rect 8 4149 9 4201
rect 61 4149 62 4201
rect 8 4142 62 4149
rect 108 4227 162 4333
rect 208 4411 262 4418
rect 208 4359 209 4411
rect 261 4359 262 4411
rect 208 4333 218 4359
rect 252 4333 262 4359
rect 208 4321 262 4333
rect 308 4367 362 4473
rect 408 4507 462 4519
rect 408 4481 418 4507
rect 452 4481 462 4507
rect 408 4429 409 4481
rect 461 4429 462 4481
rect 408 4422 462 4429
rect 508 4507 562 4613
rect 608 4691 662 4698
rect 608 4639 609 4691
rect 661 4639 662 4691
rect 608 4613 618 4639
rect 652 4613 662 4639
rect 608 4601 662 4613
rect 708 4647 762 4753
rect 808 4787 862 4799
rect 808 4761 818 4787
rect 852 4761 862 4787
rect 808 4709 809 4761
rect 861 4709 862 4761
rect 808 4702 862 4709
rect 908 4787 962 4960
rect 1002 4919 1068 4920
rect 1002 4867 1009 4919
rect 1061 4867 1068 4919
rect 1002 4866 1068 4867
rect 908 4753 918 4787
rect 952 4753 962 4787
rect 708 4613 718 4647
rect 752 4613 762 4647
rect 508 4473 518 4507
rect 552 4473 562 4507
rect 308 4333 318 4367
rect 352 4333 362 4367
rect 108 4193 118 4227
rect 152 4193 162 4227
rect 8 4087 62 4099
rect 8 4061 18 4087
rect 52 4061 62 4087
rect 8 4009 9 4061
rect 61 4009 62 4061
rect 8 4002 62 4009
rect 108 4087 162 4193
rect 208 4271 262 4278
rect 208 4219 209 4271
rect 261 4219 262 4271
rect 208 4193 218 4219
rect 252 4193 262 4219
rect 208 4181 262 4193
rect 308 4227 362 4333
rect 408 4367 462 4379
rect 408 4341 418 4367
rect 452 4341 462 4367
rect 408 4289 409 4341
rect 461 4289 462 4341
rect 408 4282 462 4289
rect 508 4367 562 4473
rect 608 4551 662 4558
rect 608 4499 609 4551
rect 661 4499 662 4551
rect 608 4473 618 4499
rect 652 4473 662 4499
rect 608 4461 662 4473
rect 708 4507 762 4613
rect 808 4647 862 4659
rect 808 4621 818 4647
rect 852 4621 862 4647
rect 808 4569 809 4621
rect 861 4569 862 4621
rect 808 4562 862 4569
rect 908 4647 962 4753
rect 1008 4831 1062 4838
rect 1008 4779 1009 4831
rect 1061 4779 1062 4831
rect 1008 4753 1018 4779
rect 1052 4753 1062 4779
rect 1008 4741 1062 4753
rect 1108 4787 1162 4960
rect 1202 4903 1268 4904
rect 1202 4851 1209 4903
rect 1261 4851 1268 4903
rect 1202 4850 1268 4851
rect 1108 4753 1118 4787
rect 1152 4753 1162 4787
rect 908 4613 918 4647
rect 952 4613 962 4647
rect 708 4473 718 4507
rect 752 4473 762 4507
rect 508 4333 518 4367
rect 552 4333 562 4367
rect 308 4193 318 4227
rect 352 4193 362 4227
rect 108 4053 118 4087
rect 152 4053 162 4087
rect 8 3947 62 3959
rect 8 3921 18 3947
rect 52 3921 62 3947
rect 8 3869 9 3921
rect 61 3869 62 3921
rect 8 3862 62 3869
rect 108 3947 162 4053
rect 208 4131 262 4138
rect 208 4079 209 4131
rect 261 4079 262 4131
rect 208 4053 218 4079
rect 252 4053 262 4079
rect 208 4041 262 4053
rect 308 4087 362 4193
rect 408 4227 462 4239
rect 408 4201 418 4227
rect 452 4201 462 4227
rect 408 4149 409 4201
rect 461 4149 462 4201
rect 408 4142 462 4149
rect 508 4227 562 4333
rect 608 4411 662 4418
rect 608 4359 609 4411
rect 661 4359 662 4411
rect 608 4333 618 4359
rect 652 4333 662 4359
rect 608 4321 662 4333
rect 708 4367 762 4473
rect 808 4507 862 4519
rect 808 4481 818 4507
rect 852 4481 862 4507
rect 808 4429 809 4481
rect 861 4429 862 4481
rect 808 4422 862 4429
rect 908 4507 962 4613
rect 1008 4691 1062 4698
rect 1008 4639 1009 4691
rect 1061 4639 1062 4691
rect 1008 4613 1018 4639
rect 1052 4613 1062 4639
rect 1008 4601 1062 4613
rect 1108 4647 1162 4753
rect 1208 4787 1262 4799
rect 1208 4761 1218 4787
rect 1252 4761 1262 4787
rect 1208 4709 1209 4761
rect 1261 4709 1262 4761
rect 1208 4702 1262 4709
rect 1308 4787 1362 4960
rect 1402 4919 1468 4920
rect 1402 4867 1409 4919
rect 1461 4867 1468 4919
rect 1402 4866 1468 4867
rect 1308 4753 1318 4787
rect 1352 4753 1362 4787
rect 1108 4613 1118 4647
rect 1152 4613 1162 4647
rect 908 4473 918 4507
rect 952 4473 962 4507
rect 708 4333 718 4367
rect 752 4333 762 4367
rect 508 4193 518 4227
rect 552 4193 562 4227
rect 308 4053 318 4087
rect 352 4053 362 4087
rect 108 3913 118 3947
rect 152 3913 162 3947
rect 8 3807 62 3819
rect 8 3781 18 3807
rect 52 3781 62 3807
rect 8 3729 9 3781
rect 61 3729 62 3781
rect 8 3722 62 3729
rect 108 3807 162 3913
rect 208 3991 262 3998
rect 208 3939 209 3991
rect 261 3939 262 3991
rect 208 3913 218 3939
rect 252 3913 262 3939
rect 208 3901 262 3913
rect 308 3947 362 4053
rect 408 4087 462 4099
rect 408 4061 418 4087
rect 452 4061 462 4087
rect 408 4009 409 4061
rect 461 4009 462 4061
rect 408 4002 462 4009
rect 508 4087 562 4193
rect 608 4271 662 4278
rect 608 4219 609 4271
rect 661 4219 662 4271
rect 608 4193 618 4219
rect 652 4193 662 4219
rect 608 4181 662 4193
rect 708 4227 762 4333
rect 808 4367 862 4379
rect 808 4341 818 4367
rect 852 4341 862 4367
rect 808 4289 809 4341
rect 861 4289 862 4341
rect 808 4282 862 4289
rect 908 4367 962 4473
rect 1008 4551 1062 4558
rect 1008 4499 1009 4551
rect 1061 4499 1062 4551
rect 1008 4473 1018 4499
rect 1052 4473 1062 4499
rect 1008 4461 1062 4473
rect 1108 4507 1162 4613
rect 1208 4647 1262 4659
rect 1208 4621 1218 4647
rect 1252 4621 1262 4647
rect 1208 4569 1209 4621
rect 1261 4569 1262 4621
rect 1208 4562 1262 4569
rect 1308 4647 1362 4753
rect 1408 4831 1462 4838
rect 1408 4779 1409 4831
rect 1461 4779 1462 4831
rect 1408 4753 1418 4779
rect 1452 4753 1462 4779
rect 1408 4741 1462 4753
rect 1508 4787 1562 4960
rect 1602 4903 1668 4904
rect 1602 4851 1609 4903
rect 1661 4851 1668 4903
rect 1602 4850 1668 4851
rect 1508 4753 1518 4787
rect 1552 4753 1562 4787
rect 1308 4613 1318 4647
rect 1352 4613 1362 4647
rect 1108 4473 1118 4507
rect 1152 4473 1162 4507
rect 908 4333 918 4367
rect 952 4333 962 4367
rect 708 4193 718 4227
rect 752 4193 762 4227
rect 508 4053 518 4087
rect 552 4053 562 4087
rect 308 3913 318 3947
rect 352 3913 362 3947
rect 108 3773 118 3807
rect 152 3773 162 3807
rect 2 3693 68 3694
rect 2 3641 9 3693
rect 61 3641 68 3693
rect 2 3640 68 3641
rect 8 3577 62 3589
rect 8 3551 18 3577
rect 52 3551 62 3577
rect 8 3499 9 3551
rect 61 3499 62 3551
rect 8 3492 62 3499
rect 108 3577 162 3773
rect 208 3851 262 3858
rect 208 3799 209 3851
rect 261 3799 262 3851
rect 208 3773 218 3799
rect 252 3773 262 3799
rect 208 3761 262 3773
rect 308 3807 362 3913
rect 408 3947 462 3959
rect 408 3921 418 3947
rect 452 3921 462 3947
rect 408 3869 409 3921
rect 461 3869 462 3921
rect 408 3862 462 3869
rect 508 3947 562 4053
rect 608 4131 662 4138
rect 608 4079 609 4131
rect 661 4079 662 4131
rect 608 4053 618 4079
rect 652 4053 662 4079
rect 608 4041 662 4053
rect 708 4087 762 4193
rect 808 4227 862 4239
rect 808 4201 818 4227
rect 852 4201 862 4227
rect 808 4149 809 4201
rect 861 4149 862 4201
rect 808 4142 862 4149
rect 908 4227 962 4333
rect 1008 4411 1062 4418
rect 1008 4359 1009 4411
rect 1061 4359 1062 4411
rect 1008 4333 1018 4359
rect 1052 4333 1062 4359
rect 1008 4321 1062 4333
rect 1108 4367 1162 4473
rect 1208 4507 1262 4519
rect 1208 4481 1218 4507
rect 1252 4481 1262 4507
rect 1208 4429 1209 4481
rect 1261 4429 1262 4481
rect 1208 4422 1262 4429
rect 1308 4507 1362 4613
rect 1408 4691 1462 4698
rect 1408 4639 1409 4691
rect 1461 4639 1462 4691
rect 1408 4613 1418 4639
rect 1452 4613 1462 4639
rect 1408 4601 1462 4613
rect 1508 4647 1562 4753
rect 1608 4787 1662 4799
rect 1608 4761 1618 4787
rect 1652 4761 1662 4787
rect 1608 4709 1609 4761
rect 1661 4709 1662 4761
rect 1608 4702 1662 4709
rect 1708 4787 1762 4960
rect 1802 4919 1868 4920
rect 1802 4867 1809 4919
rect 1861 4867 1868 4919
rect 1802 4866 1868 4867
rect 1708 4753 1718 4787
rect 1752 4753 1762 4787
rect 1508 4613 1518 4647
rect 1552 4613 1562 4647
rect 1308 4473 1318 4507
rect 1352 4473 1362 4507
rect 1108 4333 1118 4367
rect 1152 4333 1162 4367
rect 908 4193 918 4227
rect 952 4193 962 4227
rect 708 4053 718 4087
rect 752 4053 762 4087
rect 508 3913 518 3947
rect 552 3913 562 3947
rect 308 3773 318 3807
rect 352 3773 362 3807
rect 202 3709 268 3710
rect 202 3657 209 3709
rect 261 3657 268 3709
rect 202 3656 268 3657
rect 108 3543 118 3577
rect 152 3543 162 3577
rect 8 3437 62 3449
rect 8 3411 18 3437
rect 52 3411 62 3437
rect 8 3359 9 3411
rect 61 3359 62 3411
rect 8 3352 62 3359
rect 108 3437 162 3543
rect 208 3621 262 3628
rect 208 3569 209 3621
rect 261 3569 262 3621
rect 208 3543 218 3569
rect 252 3543 262 3569
rect 208 3531 262 3543
rect 308 3577 362 3773
rect 408 3807 462 3819
rect 408 3781 418 3807
rect 452 3781 462 3807
rect 408 3729 409 3781
rect 461 3729 462 3781
rect 408 3722 462 3729
rect 508 3807 562 3913
rect 608 3991 662 3998
rect 608 3939 609 3991
rect 661 3939 662 3991
rect 608 3913 618 3939
rect 652 3913 662 3939
rect 608 3901 662 3913
rect 708 3947 762 4053
rect 808 4087 862 4099
rect 808 4061 818 4087
rect 852 4061 862 4087
rect 808 4009 809 4061
rect 861 4009 862 4061
rect 808 4002 862 4009
rect 908 4087 962 4193
rect 1008 4271 1062 4278
rect 1008 4219 1009 4271
rect 1061 4219 1062 4271
rect 1008 4193 1018 4219
rect 1052 4193 1062 4219
rect 1008 4181 1062 4193
rect 1108 4227 1162 4333
rect 1208 4367 1262 4379
rect 1208 4341 1218 4367
rect 1252 4341 1262 4367
rect 1208 4289 1209 4341
rect 1261 4289 1262 4341
rect 1208 4282 1262 4289
rect 1308 4367 1362 4473
rect 1408 4551 1462 4558
rect 1408 4499 1409 4551
rect 1461 4499 1462 4551
rect 1408 4473 1418 4499
rect 1452 4473 1462 4499
rect 1408 4461 1462 4473
rect 1508 4507 1562 4613
rect 1608 4647 1662 4659
rect 1608 4621 1618 4647
rect 1652 4621 1662 4647
rect 1608 4569 1609 4621
rect 1661 4569 1662 4621
rect 1608 4562 1662 4569
rect 1708 4647 1762 4753
rect 1808 4831 1862 4838
rect 1808 4779 1809 4831
rect 1861 4779 1862 4831
rect 1808 4753 1818 4779
rect 1852 4753 1862 4779
rect 1808 4741 1862 4753
rect 1908 4787 1962 4960
rect 2002 4903 2068 4904
rect 2002 4851 2009 4903
rect 2061 4851 2068 4903
rect 2002 4850 2068 4851
rect 1908 4753 1918 4787
rect 1952 4753 1962 4787
rect 1708 4613 1718 4647
rect 1752 4613 1762 4647
rect 1508 4473 1518 4507
rect 1552 4473 1562 4507
rect 1308 4333 1318 4367
rect 1352 4333 1362 4367
rect 1108 4193 1118 4227
rect 1152 4193 1162 4227
rect 908 4053 918 4087
rect 952 4053 962 4087
rect 708 3913 718 3947
rect 752 3913 762 3947
rect 508 3773 518 3807
rect 552 3773 562 3807
rect 402 3693 468 3694
rect 402 3641 409 3693
rect 461 3641 468 3693
rect 402 3640 468 3641
rect 308 3543 318 3577
rect 352 3543 362 3577
rect 108 3403 118 3437
rect 152 3403 162 3437
rect 8 3297 62 3309
rect 8 3271 18 3297
rect 52 3271 62 3297
rect 8 3219 9 3271
rect 61 3219 62 3271
rect 8 3212 62 3219
rect 108 3297 162 3403
rect 208 3481 262 3488
rect 208 3429 209 3481
rect 261 3429 262 3481
rect 208 3403 218 3429
rect 252 3403 262 3429
rect 208 3391 262 3403
rect 308 3437 362 3543
rect 408 3577 462 3589
rect 408 3551 418 3577
rect 452 3551 462 3577
rect 408 3499 409 3551
rect 461 3499 462 3551
rect 408 3492 462 3499
rect 508 3577 562 3773
rect 608 3851 662 3858
rect 608 3799 609 3851
rect 661 3799 662 3851
rect 608 3773 618 3799
rect 652 3773 662 3799
rect 608 3761 662 3773
rect 708 3807 762 3913
rect 808 3947 862 3959
rect 808 3921 818 3947
rect 852 3921 862 3947
rect 808 3869 809 3921
rect 861 3869 862 3921
rect 808 3862 862 3869
rect 908 3947 962 4053
rect 1008 4131 1062 4138
rect 1008 4079 1009 4131
rect 1061 4079 1062 4131
rect 1008 4053 1018 4079
rect 1052 4053 1062 4079
rect 1008 4041 1062 4053
rect 1108 4087 1162 4193
rect 1208 4227 1262 4239
rect 1208 4201 1218 4227
rect 1252 4201 1262 4227
rect 1208 4149 1209 4201
rect 1261 4149 1262 4201
rect 1208 4142 1262 4149
rect 1308 4227 1362 4333
rect 1408 4411 1462 4418
rect 1408 4359 1409 4411
rect 1461 4359 1462 4411
rect 1408 4333 1418 4359
rect 1452 4333 1462 4359
rect 1408 4321 1462 4333
rect 1508 4367 1562 4473
rect 1608 4507 1662 4519
rect 1608 4481 1618 4507
rect 1652 4481 1662 4507
rect 1608 4429 1609 4481
rect 1661 4429 1662 4481
rect 1608 4422 1662 4429
rect 1708 4507 1762 4613
rect 1808 4691 1862 4698
rect 1808 4639 1809 4691
rect 1861 4639 1862 4691
rect 1808 4613 1818 4639
rect 1852 4613 1862 4639
rect 1808 4601 1862 4613
rect 1908 4647 1962 4753
rect 2008 4787 2062 4799
rect 2008 4761 2018 4787
rect 2052 4761 2062 4787
rect 2008 4709 2009 4761
rect 2061 4709 2062 4761
rect 2008 4702 2062 4709
rect 2108 4787 2162 4960
rect 2202 4919 2268 4920
rect 2202 4867 2209 4919
rect 2261 4867 2268 4919
rect 2202 4866 2268 4867
rect 2108 4753 2118 4787
rect 2152 4753 2162 4787
rect 1908 4613 1918 4647
rect 1952 4613 1962 4647
rect 1708 4473 1718 4507
rect 1752 4473 1762 4507
rect 1508 4333 1518 4367
rect 1552 4333 1562 4367
rect 1308 4193 1318 4227
rect 1352 4193 1362 4227
rect 1108 4053 1118 4087
rect 1152 4053 1162 4087
rect 908 3913 918 3947
rect 952 3913 962 3947
rect 708 3773 718 3807
rect 752 3773 762 3807
rect 602 3709 668 3710
rect 602 3657 609 3709
rect 661 3657 668 3709
rect 602 3656 668 3657
rect 508 3543 518 3577
rect 552 3543 562 3577
rect 308 3403 318 3437
rect 352 3403 362 3437
rect 108 3263 118 3297
rect 152 3263 162 3297
rect 8 3157 62 3169
rect 8 3131 18 3157
rect 52 3131 62 3157
rect 8 3079 9 3131
rect 61 3079 62 3131
rect 8 3072 62 3079
rect 108 3157 162 3263
rect 208 3341 262 3348
rect 208 3289 209 3341
rect 261 3289 262 3341
rect 208 3263 218 3289
rect 252 3263 262 3289
rect 208 3251 262 3263
rect 308 3297 362 3403
rect 408 3437 462 3449
rect 408 3411 418 3437
rect 452 3411 462 3437
rect 408 3359 409 3411
rect 461 3359 462 3411
rect 408 3352 462 3359
rect 508 3437 562 3543
rect 608 3621 662 3628
rect 608 3569 609 3621
rect 661 3569 662 3621
rect 608 3543 618 3569
rect 652 3543 662 3569
rect 608 3531 662 3543
rect 708 3577 762 3773
rect 808 3807 862 3819
rect 808 3781 818 3807
rect 852 3781 862 3807
rect 808 3729 809 3781
rect 861 3729 862 3781
rect 808 3722 862 3729
rect 908 3807 962 3913
rect 1008 3991 1062 3998
rect 1008 3939 1009 3991
rect 1061 3939 1062 3991
rect 1008 3913 1018 3939
rect 1052 3913 1062 3939
rect 1008 3901 1062 3913
rect 1108 3947 1162 4053
rect 1208 4087 1262 4099
rect 1208 4061 1218 4087
rect 1252 4061 1262 4087
rect 1208 4009 1209 4061
rect 1261 4009 1262 4061
rect 1208 4002 1262 4009
rect 1308 4087 1362 4193
rect 1408 4271 1462 4278
rect 1408 4219 1409 4271
rect 1461 4219 1462 4271
rect 1408 4193 1418 4219
rect 1452 4193 1462 4219
rect 1408 4181 1462 4193
rect 1508 4227 1562 4333
rect 1608 4367 1662 4379
rect 1608 4341 1618 4367
rect 1652 4341 1662 4367
rect 1608 4289 1609 4341
rect 1661 4289 1662 4341
rect 1608 4282 1662 4289
rect 1708 4367 1762 4473
rect 1808 4551 1862 4558
rect 1808 4499 1809 4551
rect 1861 4499 1862 4551
rect 1808 4473 1818 4499
rect 1852 4473 1862 4499
rect 1808 4461 1862 4473
rect 1908 4507 1962 4613
rect 2008 4647 2062 4659
rect 2008 4621 2018 4647
rect 2052 4621 2062 4647
rect 2008 4569 2009 4621
rect 2061 4569 2062 4621
rect 2008 4562 2062 4569
rect 2108 4647 2162 4753
rect 2208 4831 2262 4838
rect 2208 4779 2209 4831
rect 2261 4779 2262 4831
rect 2208 4753 2218 4779
rect 2252 4753 2262 4779
rect 2208 4741 2262 4753
rect 2308 4787 2362 4960
rect 2402 4903 2468 4904
rect 2402 4851 2409 4903
rect 2461 4851 2468 4903
rect 2402 4850 2468 4851
rect 2308 4753 2318 4787
rect 2352 4753 2362 4787
rect 2108 4613 2118 4647
rect 2152 4613 2162 4647
rect 1908 4473 1918 4507
rect 1952 4473 1962 4507
rect 1708 4333 1718 4367
rect 1752 4333 1762 4367
rect 1508 4193 1518 4227
rect 1552 4193 1562 4227
rect 1308 4053 1318 4087
rect 1352 4053 1362 4087
rect 1108 3913 1118 3947
rect 1152 3913 1162 3947
rect 908 3773 918 3807
rect 952 3773 962 3807
rect 802 3693 868 3694
rect 802 3641 809 3693
rect 861 3641 868 3693
rect 802 3640 868 3641
rect 708 3543 718 3577
rect 752 3543 762 3577
rect 508 3403 518 3437
rect 552 3403 562 3437
rect 308 3263 318 3297
rect 352 3263 362 3297
rect 108 3123 118 3157
rect 152 3123 162 3157
rect 8 3017 62 3029
rect 8 2991 18 3017
rect 52 2991 62 3017
rect 8 2939 9 2991
rect 61 2939 62 2991
rect 8 2932 62 2939
rect 108 3017 162 3123
rect 208 3201 262 3208
rect 208 3149 209 3201
rect 261 3149 262 3201
rect 208 3123 218 3149
rect 252 3123 262 3149
rect 208 3111 262 3123
rect 308 3157 362 3263
rect 408 3297 462 3309
rect 408 3271 418 3297
rect 452 3271 462 3297
rect 408 3219 409 3271
rect 461 3219 462 3271
rect 408 3212 462 3219
rect 508 3297 562 3403
rect 608 3481 662 3488
rect 608 3429 609 3481
rect 661 3429 662 3481
rect 608 3403 618 3429
rect 652 3403 662 3429
rect 608 3391 662 3403
rect 708 3437 762 3543
rect 808 3577 862 3589
rect 808 3551 818 3577
rect 852 3551 862 3577
rect 808 3499 809 3551
rect 861 3499 862 3551
rect 808 3492 862 3499
rect 908 3577 962 3773
rect 1008 3851 1062 3858
rect 1008 3799 1009 3851
rect 1061 3799 1062 3851
rect 1008 3773 1018 3799
rect 1052 3773 1062 3799
rect 1008 3761 1062 3773
rect 1108 3807 1162 3913
rect 1208 3947 1262 3959
rect 1208 3921 1218 3947
rect 1252 3921 1262 3947
rect 1208 3869 1209 3921
rect 1261 3869 1262 3921
rect 1208 3862 1262 3869
rect 1308 3947 1362 4053
rect 1408 4131 1462 4138
rect 1408 4079 1409 4131
rect 1461 4079 1462 4131
rect 1408 4053 1418 4079
rect 1452 4053 1462 4079
rect 1408 4041 1462 4053
rect 1508 4087 1562 4193
rect 1608 4227 1662 4239
rect 1608 4201 1618 4227
rect 1652 4201 1662 4227
rect 1608 4149 1609 4201
rect 1661 4149 1662 4201
rect 1608 4142 1662 4149
rect 1708 4227 1762 4333
rect 1808 4411 1862 4418
rect 1808 4359 1809 4411
rect 1861 4359 1862 4411
rect 1808 4333 1818 4359
rect 1852 4333 1862 4359
rect 1808 4321 1862 4333
rect 1908 4367 1962 4473
rect 2008 4507 2062 4519
rect 2008 4481 2018 4507
rect 2052 4481 2062 4507
rect 2008 4429 2009 4481
rect 2061 4429 2062 4481
rect 2008 4422 2062 4429
rect 2108 4507 2162 4613
rect 2208 4691 2262 4698
rect 2208 4639 2209 4691
rect 2261 4639 2262 4691
rect 2208 4613 2218 4639
rect 2252 4613 2262 4639
rect 2208 4601 2262 4613
rect 2308 4647 2362 4753
rect 2408 4787 2462 4799
rect 2408 4761 2418 4787
rect 2452 4761 2462 4787
rect 2408 4709 2409 4761
rect 2461 4709 2462 4761
rect 2408 4702 2462 4709
rect 2508 4787 2562 4960
rect 2602 4919 2668 4920
rect 2602 4867 2609 4919
rect 2661 4867 2668 4919
rect 2602 4866 2668 4867
rect 2508 4753 2518 4787
rect 2552 4753 2562 4787
rect 2308 4613 2318 4647
rect 2352 4613 2362 4647
rect 2108 4473 2118 4507
rect 2152 4473 2162 4507
rect 1908 4333 1918 4367
rect 1952 4333 1962 4367
rect 1708 4193 1718 4227
rect 1752 4193 1762 4227
rect 1508 4053 1518 4087
rect 1552 4053 1562 4087
rect 1308 3913 1318 3947
rect 1352 3913 1362 3947
rect 1108 3773 1118 3807
rect 1152 3773 1162 3807
rect 1002 3709 1068 3710
rect 1002 3657 1009 3709
rect 1061 3657 1068 3709
rect 1002 3656 1068 3657
rect 908 3543 918 3577
rect 952 3543 962 3577
rect 708 3403 718 3437
rect 752 3403 762 3437
rect 508 3263 518 3297
rect 552 3263 562 3297
rect 308 3123 318 3157
rect 352 3123 362 3157
rect 108 2983 118 3017
rect 152 2983 162 3017
rect 8 2877 62 2889
rect 8 2851 18 2877
rect 52 2851 62 2877
rect 8 2799 9 2851
rect 61 2799 62 2851
rect 8 2792 62 2799
rect 108 2877 162 2983
rect 208 3061 262 3068
rect 208 3009 209 3061
rect 261 3009 262 3061
rect 208 2983 218 3009
rect 252 2983 262 3009
rect 208 2971 262 2983
rect 308 3017 362 3123
rect 408 3157 462 3169
rect 408 3131 418 3157
rect 452 3131 462 3157
rect 408 3079 409 3131
rect 461 3079 462 3131
rect 408 3072 462 3079
rect 508 3157 562 3263
rect 608 3341 662 3348
rect 608 3289 609 3341
rect 661 3289 662 3341
rect 608 3263 618 3289
rect 652 3263 662 3289
rect 608 3251 662 3263
rect 708 3297 762 3403
rect 808 3437 862 3449
rect 808 3411 818 3437
rect 852 3411 862 3437
rect 808 3359 809 3411
rect 861 3359 862 3411
rect 808 3352 862 3359
rect 908 3437 962 3543
rect 1008 3621 1062 3628
rect 1008 3569 1009 3621
rect 1061 3569 1062 3621
rect 1008 3543 1018 3569
rect 1052 3543 1062 3569
rect 1008 3531 1062 3543
rect 1108 3577 1162 3773
rect 1208 3807 1262 3819
rect 1208 3781 1218 3807
rect 1252 3781 1262 3807
rect 1208 3729 1209 3781
rect 1261 3729 1262 3781
rect 1208 3722 1262 3729
rect 1308 3807 1362 3913
rect 1408 3991 1462 3998
rect 1408 3939 1409 3991
rect 1461 3939 1462 3991
rect 1408 3913 1418 3939
rect 1452 3913 1462 3939
rect 1408 3901 1462 3913
rect 1508 3947 1562 4053
rect 1608 4087 1662 4099
rect 1608 4061 1618 4087
rect 1652 4061 1662 4087
rect 1608 4009 1609 4061
rect 1661 4009 1662 4061
rect 1608 4002 1662 4009
rect 1708 4087 1762 4193
rect 1808 4271 1862 4278
rect 1808 4219 1809 4271
rect 1861 4219 1862 4271
rect 1808 4193 1818 4219
rect 1852 4193 1862 4219
rect 1808 4181 1862 4193
rect 1908 4227 1962 4333
rect 2008 4367 2062 4379
rect 2008 4341 2018 4367
rect 2052 4341 2062 4367
rect 2008 4289 2009 4341
rect 2061 4289 2062 4341
rect 2008 4282 2062 4289
rect 2108 4367 2162 4473
rect 2208 4551 2262 4558
rect 2208 4499 2209 4551
rect 2261 4499 2262 4551
rect 2208 4473 2218 4499
rect 2252 4473 2262 4499
rect 2208 4461 2262 4473
rect 2308 4507 2362 4613
rect 2408 4647 2462 4659
rect 2408 4621 2418 4647
rect 2452 4621 2462 4647
rect 2408 4569 2409 4621
rect 2461 4569 2462 4621
rect 2408 4562 2462 4569
rect 2508 4647 2562 4753
rect 2608 4831 2662 4838
rect 2608 4779 2609 4831
rect 2661 4779 2662 4831
rect 2608 4753 2618 4779
rect 2652 4753 2662 4779
rect 2608 4741 2662 4753
rect 2708 4787 2762 4960
rect 2802 4903 2868 4904
rect 2802 4851 2809 4903
rect 2861 4851 2868 4903
rect 2802 4850 2868 4851
rect 2708 4753 2718 4787
rect 2752 4753 2762 4787
rect 2508 4613 2518 4647
rect 2552 4613 2562 4647
rect 2308 4473 2318 4507
rect 2352 4473 2362 4507
rect 2108 4333 2118 4367
rect 2152 4333 2162 4367
rect 1908 4193 1918 4227
rect 1952 4193 1962 4227
rect 1708 4053 1718 4087
rect 1752 4053 1762 4087
rect 1508 3913 1518 3947
rect 1552 3913 1562 3947
rect 1308 3773 1318 3807
rect 1352 3773 1362 3807
rect 1202 3693 1268 3694
rect 1202 3641 1209 3693
rect 1261 3641 1268 3693
rect 1202 3640 1268 3641
rect 1108 3543 1118 3577
rect 1152 3543 1162 3577
rect 908 3403 918 3437
rect 952 3403 962 3437
rect 708 3263 718 3297
rect 752 3263 762 3297
rect 508 3123 518 3157
rect 552 3123 562 3157
rect 308 2983 318 3017
rect 352 2983 362 3017
rect 108 2843 118 2877
rect 152 2843 162 2877
rect 8 2737 62 2749
rect 8 2711 18 2737
rect 52 2711 62 2737
rect 8 2659 9 2711
rect 61 2659 62 2711
rect 8 2652 62 2659
rect 108 2737 162 2843
rect 208 2921 262 2928
rect 208 2869 209 2921
rect 261 2869 262 2921
rect 208 2843 218 2869
rect 252 2843 262 2869
rect 208 2831 262 2843
rect 308 2877 362 2983
rect 408 3017 462 3029
rect 408 2991 418 3017
rect 452 2991 462 3017
rect 408 2939 409 2991
rect 461 2939 462 2991
rect 408 2932 462 2939
rect 508 3017 562 3123
rect 608 3201 662 3208
rect 608 3149 609 3201
rect 661 3149 662 3201
rect 608 3123 618 3149
rect 652 3123 662 3149
rect 608 3111 662 3123
rect 708 3157 762 3263
rect 808 3297 862 3309
rect 808 3271 818 3297
rect 852 3271 862 3297
rect 808 3219 809 3271
rect 861 3219 862 3271
rect 808 3212 862 3219
rect 908 3297 962 3403
rect 1008 3481 1062 3488
rect 1008 3429 1009 3481
rect 1061 3429 1062 3481
rect 1008 3403 1018 3429
rect 1052 3403 1062 3429
rect 1008 3391 1062 3403
rect 1108 3437 1162 3543
rect 1208 3577 1262 3589
rect 1208 3551 1218 3577
rect 1252 3551 1262 3577
rect 1208 3499 1209 3551
rect 1261 3499 1262 3551
rect 1208 3492 1262 3499
rect 1308 3577 1362 3773
rect 1408 3851 1462 3858
rect 1408 3799 1409 3851
rect 1461 3799 1462 3851
rect 1408 3773 1418 3799
rect 1452 3773 1462 3799
rect 1408 3761 1462 3773
rect 1508 3807 1562 3913
rect 1608 3947 1662 3959
rect 1608 3921 1618 3947
rect 1652 3921 1662 3947
rect 1608 3869 1609 3921
rect 1661 3869 1662 3921
rect 1608 3862 1662 3869
rect 1708 3947 1762 4053
rect 1808 4131 1862 4138
rect 1808 4079 1809 4131
rect 1861 4079 1862 4131
rect 1808 4053 1818 4079
rect 1852 4053 1862 4079
rect 1808 4041 1862 4053
rect 1908 4087 1962 4193
rect 2008 4227 2062 4239
rect 2008 4201 2018 4227
rect 2052 4201 2062 4227
rect 2008 4149 2009 4201
rect 2061 4149 2062 4201
rect 2008 4142 2062 4149
rect 2108 4227 2162 4333
rect 2208 4411 2262 4418
rect 2208 4359 2209 4411
rect 2261 4359 2262 4411
rect 2208 4333 2218 4359
rect 2252 4333 2262 4359
rect 2208 4321 2262 4333
rect 2308 4367 2362 4473
rect 2408 4507 2462 4519
rect 2408 4481 2418 4507
rect 2452 4481 2462 4507
rect 2408 4429 2409 4481
rect 2461 4429 2462 4481
rect 2408 4422 2462 4429
rect 2508 4507 2562 4613
rect 2608 4691 2662 4698
rect 2608 4639 2609 4691
rect 2661 4639 2662 4691
rect 2608 4613 2618 4639
rect 2652 4613 2662 4639
rect 2608 4601 2662 4613
rect 2708 4647 2762 4753
rect 2808 4787 2862 4799
rect 2808 4761 2818 4787
rect 2852 4761 2862 4787
rect 2808 4709 2809 4761
rect 2861 4709 2862 4761
rect 2808 4702 2862 4709
rect 2908 4787 2962 4960
rect 3002 4919 3068 4920
rect 3002 4867 3009 4919
rect 3061 4867 3068 4919
rect 3002 4866 3068 4867
rect 2908 4753 2918 4787
rect 2952 4753 2962 4787
rect 2708 4613 2718 4647
rect 2752 4613 2762 4647
rect 2508 4473 2518 4507
rect 2552 4473 2562 4507
rect 2308 4333 2318 4367
rect 2352 4333 2362 4367
rect 2108 4193 2118 4227
rect 2152 4193 2162 4227
rect 1908 4053 1918 4087
rect 1952 4053 1962 4087
rect 1708 3913 1718 3947
rect 1752 3913 1762 3947
rect 1508 3773 1518 3807
rect 1552 3773 1562 3807
rect 1402 3709 1468 3710
rect 1402 3657 1409 3709
rect 1461 3657 1468 3709
rect 1402 3656 1468 3657
rect 1308 3543 1318 3577
rect 1352 3543 1362 3577
rect 1108 3403 1118 3437
rect 1152 3403 1162 3437
rect 908 3263 918 3297
rect 952 3263 962 3297
rect 708 3123 718 3157
rect 752 3123 762 3157
rect 508 2983 518 3017
rect 552 2983 562 3017
rect 308 2843 318 2877
rect 352 2843 362 2877
rect 108 2703 118 2737
rect 152 2703 162 2737
rect 8 2597 62 2609
rect 8 2571 18 2597
rect 52 2571 62 2597
rect 8 2519 9 2571
rect 61 2519 62 2571
rect 8 2512 62 2519
rect 108 2597 162 2703
rect 208 2781 262 2788
rect 208 2729 209 2781
rect 261 2729 262 2781
rect 208 2703 218 2729
rect 252 2703 262 2729
rect 208 2691 262 2703
rect 308 2737 362 2843
rect 408 2877 462 2889
rect 408 2851 418 2877
rect 452 2851 462 2877
rect 408 2799 409 2851
rect 461 2799 462 2851
rect 408 2792 462 2799
rect 508 2877 562 2983
rect 608 3061 662 3068
rect 608 3009 609 3061
rect 661 3009 662 3061
rect 608 2983 618 3009
rect 652 2983 662 3009
rect 608 2971 662 2983
rect 708 3017 762 3123
rect 808 3157 862 3169
rect 808 3131 818 3157
rect 852 3131 862 3157
rect 808 3079 809 3131
rect 861 3079 862 3131
rect 808 3072 862 3079
rect 908 3157 962 3263
rect 1008 3341 1062 3348
rect 1008 3289 1009 3341
rect 1061 3289 1062 3341
rect 1008 3263 1018 3289
rect 1052 3263 1062 3289
rect 1008 3251 1062 3263
rect 1108 3297 1162 3403
rect 1208 3437 1262 3449
rect 1208 3411 1218 3437
rect 1252 3411 1262 3437
rect 1208 3359 1209 3411
rect 1261 3359 1262 3411
rect 1208 3352 1262 3359
rect 1308 3437 1362 3543
rect 1408 3621 1462 3628
rect 1408 3569 1409 3621
rect 1461 3569 1462 3621
rect 1408 3543 1418 3569
rect 1452 3543 1462 3569
rect 1408 3531 1462 3543
rect 1508 3577 1562 3773
rect 1608 3807 1662 3819
rect 1608 3781 1618 3807
rect 1652 3781 1662 3807
rect 1608 3729 1609 3781
rect 1661 3729 1662 3781
rect 1608 3722 1662 3729
rect 1708 3807 1762 3913
rect 1808 3991 1862 3998
rect 1808 3939 1809 3991
rect 1861 3939 1862 3991
rect 1808 3913 1818 3939
rect 1852 3913 1862 3939
rect 1808 3901 1862 3913
rect 1908 3947 1962 4053
rect 2008 4087 2062 4099
rect 2008 4061 2018 4087
rect 2052 4061 2062 4087
rect 2008 4009 2009 4061
rect 2061 4009 2062 4061
rect 2008 4002 2062 4009
rect 2108 4087 2162 4193
rect 2208 4271 2262 4278
rect 2208 4219 2209 4271
rect 2261 4219 2262 4271
rect 2208 4193 2218 4219
rect 2252 4193 2262 4219
rect 2208 4181 2262 4193
rect 2308 4227 2362 4333
rect 2408 4367 2462 4379
rect 2408 4341 2418 4367
rect 2452 4341 2462 4367
rect 2408 4289 2409 4341
rect 2461 4289 2462 4341
rect 2408 4282 2462 4289
rect 2508 4367 2562 4473
rect 2608 4551 2662 4558
rect 2608 4499 2609 4551
rect 2661 4499 2662 4551
rect 2608 4473 2618 4499
rect 2652 4473 2662 4499
rect 2608 4461 2662 4473
rect 2708 4507 2762 4613
rect 2808 4647 2862 4659
rect 2808 4621 2818 4647
rect 2852 4621 2862 4647
rect 2808 4569 2809 4621
rect 2861 4569 2862 4621
rect 2808 4562 2862 4569
rect 2908 4647 2962 4753
rect 3008 4831 3062 4838
rect 3008 4779 3009 4831
rect 3061 4779 3062 4831
rect 3008 4753 3018 4779
rect 3052 4753 3062 4779
rect 3008 4741 3062 4753
rect 3108 4787 3162 4960
rect 3202 4903 3268 4904
rect 3202 4851 3209 4903
rect 3261 4851 3268 4903
rect 3202 4850 3268 4851
rect 3108 4753 3118 4787
rect 3152 4753 3162 4787
rect 2908 4613 2918 4647
rect 2952 4613 2962 4647
rect 2708 4473 2718 4507
rect 2752 4473 2762 4507
rect 2508 4333 2518 4367
rect 2552 4333 2562 4367
rect 2308 4193 2318 4227
rect 2352 4193 2362 4227
rect 2108 4053 2118 4087
rect 2152 4053 2162 4087
rect 1908 3913 1918 3947
rect 1952 3913 1962 3947
rect 1708 3773 1718 3807
rect 1752 3773 1762 3807
rect 1602 3693 1668 3694
rect 1602 3641 1609 3693
rect 1661 3641 1668 3693
rect 1602 3640 1668 3641
rect 1508 3543 1518 3577
rect 1552 3543 1562 3577
rect 1308 3403 1318 3437
rect 1352 3403 1362 3437
rect 1108 3263 1118 3297
rect 1152 3263 1162 3297
rect 908 3123 918 3157
rect 952 3123 962 3157
rect 708 2983 718 3017
rect 752 2983 762 3017
rect 508 2843 518 2877
rect 552 2843 562 2877
rect 308 2703 318 2737
rect 352 2703 362 2737
rect 108 2563 118 2597
rect 152 2563 162 2597
rect 2 2483 68 2484
rect 2 2431 9 2483
rect 61 2431 68 2483
rect 2 2430 68 2431
rect 8 2367 62 2379
rect 8 2341 18 2367
rect 52 2341 62 2367
rect 8 2289 9 2341
rect 61 2289 62 2341
rect 8 2282 62 2289
rect 108 2367 162 2563
rect 208 2641 262 2648
rect 208 2589 209 2641
rect 261 2589 262 2641
rect 208 2563 218 2589
rect 252 2563 262 2589
rect 208 2551 262 2563
rect 308 2597 362 2703
rect 408 2737 462 2749
rect 408 2711 418 2737
rect 452 2711 462 2737
rect 408 2659 409 2711
rect 461 2659 462 2711
rect 408 2652 462 2659
rect 508 2737 562 2843
rect 608 2921 662 2928
rect 608 2869 609 2921
rect 661 2869 662 2921
rect 608 2843 618 2869
rect 652 2843 662 2869
rect 608 2831 662 2843
rect 708 2877 762 2983
rect 808 3017 862 3029
rect 808 2991 818 3017
rect 852 2991 862 3017
rect 808 2939 809 2991
rect 861 2939 862 2991
rect 808 2932 862 2939
rect 908 3017 962 3123
rect 1008 3201 1062 3208
rect 1008 3149 1009 3201
rect 1061 3149 1062 3201
rect 1008 3123 1018 3149
rect 1052 3123 1062 3149
rect 1008 3111 1062 3123
rect 1108 3157 1162 3263
rect 1208 3297 1262 3309
rect 1208 3271 1218 3297
rect 1252 3271 1262 3297
rect 1208 3219 1209 3271
rect 1261 3219 1262 3271
rect 1208 3212 1262 3219
rect 1308 3297 1362 3403
rect 1408 3481 1462 3488
rect 1408 3429 1409 3481
rect 1461 3429 1462 3481
rect 1408 3403 1418 3429
rect 1452 3403 1462 3429
rect 1408 3391 1462 3403
rect 1508 3437 1562 3543
rect 1608 3577 1662 3589
rect 1608 3551 1618 3577
rect 1652 3551 1662 3577
rect 1608 3499 1609 3551
rect 1661 3499 1662 3551
rect 1608 3492 1662 3499
rect 1708 3577 1762 3773
rect 1808 3851 1862 3858
rect 1808 3799 1809 3851
rect 1861 3799 1862 3851
rect 1808 3773 1818 3799
rect 1852 3773 1862 3799
rect 1808 3761 1862 3773
rect 1908 3807 1962 3913
rect 2008 3947 2062 3959
rect 2008 3921 2018 3947
rect 2052 3921 2062 3947
rect 2008 3869 2009 3921
rect 2061 3869 2062 3921
rect 2008 3862 2062 3869
rect 2108 3947 2162 4053
rect 2208 4131 2262 4138
rect 2208 4079 2209 4131
rect 2261 4079 2262 4131
rect 2208 4053 2218 4079
rect 2252 4053 2262 4079
rect 2208 4041 2262 4053
rect 2308 4087 2362 4193
rect 2408 4227 2462 4239
rect 2408 4201 2418 4227
rect 2452 4201 2462 4227
rect 2408 4149 2409 4201
rect 2461 4149 2462 4201
rect 2408 4142 2462 4149
rect 2508 4227 2562 4333
rect 2608 4411 2662 4418
rect 2608 4359 2609 4411
rect 2661 4359 2662 4411
rect 2608 4333 2618 4359
rect 2652 4333 2662 4359
rect 2608 4321 2662 4333
rect 2708 4367 2762 4473
rect 2808 4507 2862 4519
rect 2808 4481 2818 4507
rect 2852 4481 2862 4507
rect 2808 4429 2809 4481
rect 2861 4429 2862 4481
rect 2808 4422 2862 4429
rect 2908 4507 2962 4613
rect 3008 4691 3062 4698
rect 3008 4639 3009 4691
rect 3061 4639 3062 4691
rect 3008 4613 3018 4639
rect 3052 4613 3062 4639
rect 3008 4601 3062 4613
rect 3108 4647 3162 4753
rect 3208 4787 3262 4799
rect 3208 4761 3218 4787
rect 3252 4761 3262 4787
rect 3208 4709 3209 4761
rect 3261 4709 3262 4761
rect 3208 4702 3262 4709
rect 3308 4787 3362 4960
rect 3402 4919 3468 4920
rect 3402 4867 3409 4919
rect 3461 4867 3468 4919
rect 3402 4866 3468 4867
rect 3308 4753 3318 4787
rect 3352 4753 3362 4787
rect 3108 4613 3118 4647
rect 3152 4613 3162 4647
rect 2908 4473 2918 4507
rect 2952 4473 2962 4507
rect 2708 4333 2718 4367
rect 2752 4333 2762 4367
rect 2508 4193 2518 4227
rect 2552 4193 2562 4227
rect 2308 4053 2318 4087
rect 2352 4053 2362 4087
rect 2108 3913 2118 3947
rect 2152 3913 2162 3947
rect 1908 3773 1918 3807
rect 1952 3773 1962 3807
rect 1802 3709 1868 3710
rect 1802 3657 1809 3709
rect 1861 3657 1868 3709
rect 1802 3656 1868 3657
rect 1708 3543 1718 3577
rect 1752 3543 1762 3577
rect 1508 3403 1518 3437
rect 1552 3403 1562 3437
rect 1308 3263 1318 3297
rect 1352 3263 1362 3297
rect 1108 3123 1118 3157
rect 1152 3123 1162 3157
rect 908 2983 918 3017
rect 952 2983 962 3017
rect 708 2843 718 2877
rect 752 2843 762 2877
rect 508 2703 518 2737
rect 552 2703 562 2737
rect 308 2563 318 2597
rect 352 2563 362 2597
rect 202 2499 268 2500
rect 202 2447 209 2499
rect 261 2447 268 2499
rect 202 2446 268 2447
rect 108 2333 118 2367
rect 152 2333 162 2367
rect 8 2227 62 2239
rect 8 2201 18 2227
rect 52 2201 62 2227
rect 8 2149 9 2201
rect 61 2149 62 2201
rect 8 2142 62 2149
rect 108 2227 162 2333
rect 208 2411 262 2418
rect 208 2359 209 2411
rect 261 2359 262 2411
rect 208 2333 218 2359
rect 252 2333 262 2359
rect 208 2321 262 2333
rect 308 2367 362 2563
rect 408 2597 462 2609
rect 408 2571 418 2597
rect 452 2571 462 2597
rect 408 2519 409 2571
rect 461 2519 462 2571
rect 408 2512 462 2519
rect 508 2597 562 2703
rect 608 2781 662 2788
rect 608 2729 609 2781
rect 661 2729 662 2781
rect 608 2703 618 2729
rect 652 2703 662 2729
rect 608 2691 662 2703
rect 708 2737 762 2843
rect 808 2877 862 2889
rect 808 2851 818 2877
rect 852 2851 862 2877
rect 808 2799 809 2851
rect 861 2799 862 2851
rect 808 2792 862 2799
rect 908 2877 962 2983
rect 1008 3061 1062 3068
rect 1008 3009 1009 3061
rect 1061 3009 1062 3061
rect 1008 2983 1018 3009
rect 1052 2983 1062 3009
rect 1008 2971 1062 2983
rect 1108 3017 1162 3123
rect 1208 3157 1262 3169
rect 1208 3131 1218 3157
rect 1252 3131 1262 3157
rect 1208 3079 1209 3131
rect 1261 3079 1262 3131
rect 1208 3072 1262 3079
rect 1308 3157 1362 3263
rect 1408 3341 1462 3348
rect 1408 3289 1409 3341
rect 1461 3289 1462 3341
rect 1408 3263 1418 3289
rect 1452 3263 1462 3289
rect 1408 3251 1462 3263
rect 1508 3297 1562 3403
rect 1608 3437 1662 3449
rect 1608 3411 1618 3437
rect 1652 3411 1662 3437
rect 1608 3359 1609 3411
rect 1661 3359 1662 3411
rect 1608 3352 1662 3359
rect 1708 3437 1762 3543
rect 1808 3621 1862 3628
rect 1808 3569 1809 3621
rect 1861 3569 1862 3621
rect 1808 3543 1818 3569
rect 1852 3543 1862 3569
rect 1808 3531 1862 3543
rect 1908 3577 1962 3773
rect 2008 3807 2062 3819
rect 2008 3781 2018 3807
rect 2052 3781 2062 3807
rect 2008 3729 2009 3781
rect 2061 3729 2062 3781
rect 2008 3722 2062 3729
rect 2108 3807 2162 3913
rect 2208 3991 2262 3998
rect 2208 3939 2209 3991
rect 2261 3939 2262 3991
rect 2208 3913 2218 3939
rect 2252 3913 2262 3939
rect 2208 3901 2262 3913
rect 2308 3947 2362 4053
rect 2408 4087 2462 4099
rect 2408 4061 2418 4087
rect 2452 4061 2462 4087
rect 2408 4009 2409 4061
rect 2461 4009 2462 4061
rect 2408 4002 2462 4009
rect 2508 4087 2562 4193
rect 2608 4271 2662 4278
rect 2608 4219 2609 4271
rect 2661 4219 2662 4271
rect 2608 4193 2618 4219
rect 2652 4193 2662 4219
rect 2608 4181 2662 4193
rect 2708 4227 2762 4333
rect 2808 4367 2862 4379
rect 2808 4341 2818 4367
rect 2852 4341 2862 4367
rect 2808 4289 2809 4341
rect 2861 4289 2862 4341
rect 2808 4282 2862 4289
rect 2908 4367 2962 4473
rect 3008 4551 3062 4558
rect 3008 4499 3009 4551
rect 3061 4499 3062 4551
rect 3008 4473 3018 4499
rect 3052 4473 3062 4499
rect 3008 4461 3062 4473
rect 3108 4507 3162 4613
rect 3208 4647 3262 4659
rect 3208 4621 3218 4647
rect 3252 4621 3262 4647
rect 3208 4569 3209 4621
rect 3261 4569 3262 4621
rect 3208 4562 3262 4569
rect 3308 4647 3362 4753
rect 3408 4831 3462 4838
rect 3408 4779 3409 4831
rect 3461 4779 3462 4831
rect 3408 4753 3418 4779
rect 3452 4753 3462 4779
rect 3408 4741 3462 4753
rect 3508 4787 3562 4960
rect 3602 4903 3668 4904
rect 3602 4851 3609 4903
rect 3661 4851 3668 4903
rect 3602 4850 3668 4851
rect 3508 4753 3518 4787
rect 3552 4753 3562 4787
rect 3308 4613 3318 4647
rect 3352 4613 3362 4647
rect 3108 4473 3118 4507
rect 3152 4473 3162 4507
rect 2908 4333 2918 4367
rect 2952 4333 2962 4367
rect 2708 4193 2718 4227
rect 2752 4193 2762 4227
rect 2508 4053 2518 4087
rect 2552 4053 2562 4087
rect 2308 3913 2318 3947
rect 2352 3913 2362 3947
rect 2108 3773 2118 3807
rect 2152 3773 2162 3807
rect 2002 3693 2068 3694
rect 2002 3641 2009 3693
rect 2061 3641 2068 3693
rect 2002 3640 2068 3641
rect 1908 3543 1918 3577
rect 1952 3543 1962 3577
rect 1708 3403 1718 3437
rect 1752 3403 1762 3437
rect 1508 3263 1518 3297
rect 1552 3263 1562 3297
rect 1308 3123 1318 3157
rect 1352 3123 1362 3157
rect 1108 2983 1118 3017
rect 1152 2983 1162 3017
rect 908 2843 918 2877
rect 952 2843 962 2877
rect 708 2703 718 2737
rect 752 2703 762 2737
rect 508 2563 518 2597
rect 552 2563 562 2597
rect 402 2483 468 2484
rect 402 2431 409 2483
rect 461 2431 468 2483
rect 402 2430 468 2431
rect 308 2333 318 2367
rect 352 2333 362 2367
rect 108 2193 118 2227
rect 152 2193 162 2227
rect 8 2087 62 2099
rect 8 2061 18 2087
rect 52 2061 62 2087
rect 8 2009 9 2061
rect 61 2009 62 2061
rect 8 2002 62 2009
rect 108 2087 162 2193
rect 208 2271 262 2278
rect 208 2219 209 2271
rect 261 2219 262 2271
rect 208 2193 218 2219
rect 252 2193 262 2219
rect 208 2181 262 2193
rect 308 2227 362 2333
rect 408 2367 462 2379
rect 408 2341 418 2367
rect 452 2341 462 2367
rect 408 2289 409 2341
rect 461 2289 462 2341
rect 408 2282 462 2289
rect 508 2367 562 2563
rect 608 2641 662 2648
rect 608 2589 609 2641
rect 661 2589 662 2641
rect 608 2563 618 2589
rect 652 2563 662 2589
rect 608 2551 662 2563
rect 708 2597 762 2703
rect 808 2737 862 2749
rect 808 2711 818 2737
rect 852 2711 862 2737
rect 808 2659 809 2711
rect 861 2659 862 2711
rect 808 2652 862 2659
rect 908 2737 962 2843
rect 1008 2921 1062 2928
rect 1008 2869 1009 2921
rect 1061 2869 1062 2921
rect 1008 2843 1018 2869
rect 1052 2843 1062 2869
rect 1008 2831 1062 2843
rect 1108 2877 1162 2983
rect 1208 3017 1262 3029
rect 1208 2991 1218 3017
rect 1252 2991 1262 3017
rect 1208 2939 1209 2991
rect 1261 2939 1262 2991
rect 1208 2932 1262 2939
rect 1308 3017 1362 3123
rect 1408 3201 1462 3208
rect 1408 3149 1409 3201
rect 1461 3149 1462 3201
rect 1408 3123 1418 3149
rect 1452 3123 1462 3149
rect 1408 3111 1462 3123
rect 1508 3157 1562 3263
rect 1608 3297 1662 3309
rect 1608 3271 1618 3297
rect 1652 3271 1662 3297
rect 1608 3219 1609 3271
rect 1661 3219 1662 3271
rect 1608 3212 1662 3219
rect 1708 3297 1762 3403
rect 1808 3481 1862 3488
rect 1808 3429 1809 3481
rect 1861 3429 1862 3481
rect 1808 3403 1818 3429
rect 1852 3403 1862 3429
rect 1808 3391 1862 3403
rect 1908 3437 1962 3543
rect 2008 3577 2062 3589
rect 2008 3551 2018 3577
rect 2052 3551 2062 3577
rect 2008 3499 2009 3551
rect 2061 3499 2062 3551
rect 2008 3492 2062 3499
rect 2108 3577 2162 3773
rect 2208 3851 2262 3858
rect 2208 3799 2209 3851
rect 2261 3799 2262 3851
rect 2208 3773 2218 3799
rect 2252 3773 2262 3799
rect 2208 3761 2262 3773
rect 2308 3807 2362 3913
rect 2408 3947 2462 3959
rect 2408 3921 2418 3947
rect 2452 3921 2462 3947
rect 2408 3869 2409 3921
rect 2461 3869 2462 3921
rect 2408 3862 2462 3869
rect 2508 3947 2562 4053
rect 2608 4131 2662 4138
rect 2608 4079 2609 4131
rect 2661 4079 2662 4131
rect 2608 4053 2618 4079
rect 2652 4053 2662 4079
rect 2608 4041 2662 4053
rect 2708 4087 2762 4193
rect 2808 4227 2862 4239
rect 2808 4201 2818 4227
rect 2852 4201 2862 4227
rect 2808 4149 2809 4201
rect 2861 4149 2862 4201
rect 2808 4142 2862 4149
rect 2908 4227 2962 4333
rect 3008 4411 3062 4418
rect 3008 4359 3009 4411
rect 3061 4359 3062 4411
rect 3008 4333 3018 4359
rect 3052 4333 3062 4359
rect 3008 4321 3062 4333
rect 3108 4367 3162 4473
rect 3208 4507 3262 4519
rect 3208 4481 3218 4507
rect 3252 4481 3262 4507
rect 3208 4429 3209 4481
rect 3261 4429 3262 4481
rect 3208 4422 3262 4429
rect 3308 4507 3362 4613
rect 3408 4691 3462 4698
rect 3408 4639 3409 4691
rect 3461 4639 3462 4691
rect 3408 4613 3418 4639
rect 3452 4613 3462 4639
rect 3408 4601 3462 4613
rect 3508 4647 3562 4753
rect 3608 4787 3662 4799
rect 3608 4761 3618 4787
rect 3652 4761 3662 4787
rect 3608 4709 3609 4761
rect 3661 4709 3662 4761
rect 3608 4702 3662 4709
rect 3708 4787 3762 4960
rect 3802 4919 3868 4920
rect 3802 4867 3809 4919
rect 3861 4867 3868 4919
rect 3802 4866 3868 4867
rect 3708 4753 3718 4787
rect 3752 4753 3762 4787
rect 3508 4613 3518 4647
rect 3552 4613 3562 4647
rect 3308 4473 3318 4507
rect 3352 4473 3362 4507
rect 3108 4333 3118 4367
rect 3152 4333 3162 4367
rect 2908 4193 2918 4227
rect 2952 4193 2962 4227
rect 2708 4053 2718 4087
rect 2752 4053 2762 4087
rect 2508 3913 2518 3947
rect 2552 3913 2562 3947
rect 2308 3773 2318 3807
rect 2352 3773 2362 3807
rect 2202 3709 2268 3710
rect 2202 3657 2209 3709
rect 2261 3657 2268 3709
rect 2202 3656 2268 3657
rect 2108 3543 2118 3577
rect 2152 3543 2162 3577
rect 1908 3403 1918 3437
rect 1952 3403 1962 3437
rect 1708 3263 1718 3297
rect 1752 3263 1762 3297
rect 1508 3123 1518 3157
rect 1552 3123 1562 3157
rect 1308 2983 1318 3017
rect 1352 2983 1362 3017
rect 1108 2843 1118 2877
rect 1152 2843 1162 2877
rect 908 2703 918 2737
rect 952 2703 962 2737
rect 708 2563 718 2597
rect 752 2563 762 2597
rect 602 2499 668 2500
rect 602 2447 609 2499
rect 661 2447 668 2499
rect 602 2446 668 2447
rect 508 2333 518 2367
rect 552 2333 562 2367
rect 308 2193 318 2227
rect 352 2193 362 2227
rect 108 2053 118 2087
rect 152 2053 162 2087
rect 8 1947 62 1959
rect 8 1921 18 1947
rect 52 1921 62 1947
rect 8 1869 9 1921
rect 61 1869 62 1921
rect 8 1862 62 1869
rect 108 1947 162 2053
rect 208 2131 262 2138
rect 208 2079 209 2131
rect 261 2079 262 2131
rect 208 2053 218 2079
rect 252 2053 262 2079
rect 208 2041 262 2053
rect 308 2087 362 2193
rect 408 2227 462 2239
rect 408 2201 418 2227
rect 452 2201 462 2227
rect 408 2149 409 2201
rect 461 2149 462 2201
rect 408 2142 462 2149
rect 508 2227 562 2333
rect 608 2411 662 2418
rect 608 2359 609 2411
rect 661 2359 662 2411
rect 608 2333 618 2359
rect 652 2333 662 2359
rect 608 2321 662 2333
rect 708 2367 762 2563
rect 808 2597 862 2609
rect 808 2571 818 2597
rect 852 2571 862 2597
rect 808 2519 809 2571
rect 861 2519 862 2571
rect 808 2512 862 2519
rect 908 2597 962 2703
rect 1008 2781 1062 2788
rect 1008 2729 1009 2781
rect 1061 2729 1062 2781
rect 1008 2703 1018 2729
rect 1052 2703 1062 2729
rect 1008 2691 1062 2703
rect 1108 2737 1162 2843
rect 1208 2877 1262 2889
rect 1208 2851 1218 2877
rect 1252 2851 1262 2877
rect 1208 2799 1209 2851
rect 1261 2799 1262 2851
rect 1208 2792 1262 2799
rect 1308 2877 1362 2983
rect 1408 3061 1462 3068
rect 1408 3009 1409 3061
rect 1461 3009 1462 3061
rect 1408 2983 1418 3009
rect 1452 2983 1462 3009
rect 1408 2971 1462 2983
rect 1508 3017 1562 3123
rect 1608 3157 1662 3169
rect 1608 3131 1618 3157
rect 1652 3131 1662 3157
rect 1608 3079 1609 3131
rect 1661 3079 1662 3131
rect 1608 3072 1662 3079
rect 1708 3157 1762 3263
rect 1808 3341 1862 3348
rect 1808 3289 1809 3341
rect 1861 3289 1862 3341
rect 1808 3263 1818 3289
rect 1852 3263 1862 3289
rect 1808 3251 1862 3263
rect 1908 3297 1962 3403
rect 2008 3437 2062 3449
rect 2008 3411 2018 3437
rect 2052 3411 2062 3437
rect 2008 3359 2009 3411
rect 2061 3359 2062 3411
rect 2008 3352 2062 3359
rect 2108 3437 2162 3543
rect 2208 3621 2262 3628
rect 2208 3569 2209 3621
rect 2261 3569 2262 3621
rect 2208 3543 2218 3569
rect 2252 3543 2262 3569
rect 2208 3531 2262 3543
rect 2308 3577 2362 3773
rect 2408 3807 2462 3819
rect 2408 3781 2418 3807
rect 2452 3781 2462 3807
rect 2408 3729 2409 3781
rect 2461 3729 2462 3781
rect 2408 3722 2462 3729
rect 2508 3807 2562 3913
rect 2608 3991 2662 3998
rect 2608 3939 2609 3991
rect 2661 3939 2662 3991
rect 2608 3913 2618 3939
rect 2652 3913 2662 3939
rect 2608 3901 2662 3913
rect 2708 3947 2762 4053
rect 2808 4087 2862 4099
rect 2808 4061 2818 4087
rect 2852 4061 2862 4087
rect 2808 4009 2809 4061
rect 2861 4009 2862 4061
rect 2808 4002 2862 4009
rect 2908 4087 2962 4193
rect 3008 4271 3062 4278
rect 3008 4219 3009 4271
rect 3061 4219 3062 4271
rect 3008 4193 3018 4219
rect 3052 4193 3062 4219
rect 3008 4181 3062 4193
rect 3108 4227 3162 4333
rect 3208 4367 3262 4379
rect 3208 4341 3218 4367
rect 3252 4341 3262 4367
rect 3208 4289 3209 4341
rect 3261 4289 3262 4341
rect 3208 4282 3262 4289
rect 3308 4367 3362 4473
rect 3408 4551 3462 4558
rect 3408 4499 3409 4551
rect 3461 4499 3462 4551
rect 3408 4473 3418 4499
rect 3452 4473 3462 4499
rect 3408 4461 3462 4473
rect 3508 4507 3562 4613
rect 3608 4647 3662 4659
rect 3608 4621 3618 4647
rect 3652 4621 3662 4647
rect 3608 4569 3609 4621
rect 3661 4569 3662 4621
rect 3608 4562 3662 4569
rect 3708 4647 3762 4753
rect 3808 4831 3862 4838
rect 3808 4779 3809 4831
rect 3861 4779 3862 4831
rect 3808 4753 3818 4779
rect 3852 4753 3862 4779
rect 3808 4741 3862 4753
rect 3908 4787 3962 4960
rect 4002 4903 4068 4904
rect 4002 4851 4009 4903
rect 4061 4851 4068 4903
rect 4002 4850 4068 4851
rect 3908 4753 3918 4787
rect 3952 4753 3962 4787
rect 3708 4613 3718 4647
rect 3752 4613 3762 4647
rect 3508 4473 3518 4507
rect 3552 4473 3562 4507
rect 3308 4333 3318 4367
rect 3352 4333 3362 4367
rect 3108 4193 3118 4227
rect 3152 4193 3162 4227
rect 2908 4053 2918 4087
rect 2952 4053 2962 4087
rect 2708 3913 2718 3947
rect 2752 3913 2762 3947
rect 2508 3773 2518 3807
rect 2552 3773 2562 3807
rect 2402 3693 2468 3694
rect 2402 3641 2409 3693
rect 2461 3641 2468 3693
rect 2402 3640 2468 3641
rect 2308 3543 2318 3577
rect 2352 3543 2362 3577
rect 2108 3403 2118 3437
rect 2152 3403 2162 3437
rect 1908 3263 1918 3297
rect 1952 3263 1962 3297
rect 1708 3123 1718 3157
rect 1752 3123 1762 3157
rect 1508 2983 1518 3017
rect 1552 2983 1562 3017
rect 1308 2843 1318 2877
rect 1352 2843 1362 2877
rect 1108 2703 1118 2737
rect 1152 2703 1162 2737
rect 908 2563 918 2597
rect 952 2563 962 2597
rect 802 2483 868 2484
rect 802 2431 809 2483
rect 861 2431 868 2483
rect 802 2430 868 2431
rect 708 2333 718 2367
rect 752 2333 762 2367
rect 508 2193 518 2227
rect 552 2193 562 2227
rect 308 2053 318 2087
rect 352 2053 362 2087
rect 108 1913 118 1947
rect 152 1913 162 1947
rect 8 1807 62 1819
rect 8 1781 18 1807
rect 52 1781 62 1807
rect 8 1729 9 1781
rect 61 1729 62 1781
rect 8 1722 62 1729
rect 108 1807 162 1913
rect 208 1991 262 1998
rect 208 1939 209 1991
rect 261 1939 262 1991
rect 208 1913 218 1939
rect 252 1913 262 1939
rect 208 1901 262 1913
rect 308 1947 362 2053
rect 408 2087 462 2099
rect 408 2061 418 2087
rect 452 2061 462 2087
rect 408 2009 409 2061
rect 461 2009 462 2061
rect 408 2002 462 2009
rect 508 2087 562 2193
rect 608 2271 662 2278
rect 608 2219 609 2271
rect 661 2219 662 2271
rect 608 2193 618 2219
rect 652 2193 662 2219
rect 608 2181 662 2193
rect 708 2227 762 2333
rect 808 2367 862 2379
rect 808 2341 818 2367
rect 852 2341 862 2367
rect 808 2289 809 2341
rect 861 2289 862 2341
rect 808 2282 862 2289
rect 908 2367 962 2563
rect 1008 2641 1062 2648
rect 1008 2589 1009 2641
rect 1061 2589 1062 2641
rect 1008 2563 1018 2589
rect 1052 2563 1062 2589
rect 1008 2551 1062 2563
rect 1108 2597 1162 2703
rect 1208 2737 1262 2749
rect 1208 2711 1218 2737
rect 1252 2711 1262 2737
rect 1208 2659 1209 2711
rect 1261 2659 1262 2711
rect 1208 2652 1262 2659
rect 1308 2737 1362 2843
rect 1408 2921 1462 2928
rect 1408 2869 1409 2921
rect 1461 2869 1462 2921
rect 1408 2843 1418 2869
rect 1452 2843 1462 2869
rect 1408 2831 1462 2843
rect 1508 2877 1562 2983
rect 1608 3017 1662 3029
rect 1608 2991 1618 3017
rect 1652 2991 1662 3017
rect 1608 2939 1609 2991
rect 1661 2939 1662 2991
rect 1608 2932 1662 2939
rect 1708 3017 1762 3123
rect 1808 3201 1862 3208
rect 1808 3149 1809 3201
rect 1861 3149 1862 3201
rect 1808 3123 1818 3149
rect 1852 3123 1862 3149
rect 1808 3111 1862 3123
rect 1908 3157 1962 3263
rect 2008 3297 2062 3309
rect 2008 3271 2018 3297
rect 2052 3271 2062 3297
rect 2008 3219 2009 3271
rect 2061 3219 2062 3271
rect 2008 3212 2062 3219
rect 2108 3297 2162 3403
rect 2208 3481 2262 3488
rect 2208 3429 2209 3481
rect 2261 3429 2262 3481
rect 2208 3403 2218 3429
rect 2252 3403 2262 3429
rect 2208 3391 2262 3403
rect 2308 3437 2362 3543
rect 2408 3577 2462 3589
rect 2408 3551 2418 3577
rect 2452 3551 2462 3577
rect 2408 3499 2409 3551
rect 2461 3499 2462 3551
rect 2408 3492 2462 3499
rect 2508 3577 2562 3773
rect 2608 3851 2662 3858
rect 2608 3799 2609 3851
rect 2661 3799 2662 3851
rect 2608 3773 2618 3799
rect 2652 3773 2662 3799
rect 2608 3761 2662 3773
rect 2708 3807 2762 3913
rect 2808 3947 2862 3959
rect 2808 3921 2818 3947
rect 2852 3921 2862 3947
rect 2808 3869 2809 3921
rect 2861 3869 2862 3921
rect 2808 3862 2862 3869
rect 2908 3947 2962 4053
rect 3008 4131 3062 4138
rect 3008 4079 3009 4131
rect 3061 4079 3062 4131
rect 3008 4053 3018 4079
rect 3052 4053 3062 4079
rect 3008 4041 3062 4053
rect 3108 4087 3162 4193
rect 3208 4227 3262 4239
rect 3208 4201 3218 4227
rect 3252 4201 3262 4227
rect 3208 4149 3209 4201
rect 3261 4149 3262 4201
rect 3208 4142 3262 4149
rect 3308 4227 3362 4333
rect 3408 4411 3462 4418
rect 3408 4359 3409 4411
rect 3461 4359 3462 4411
rect 3408 4333 3418 4359
rect 3452 4333 3462 4359
rect 3408 4321 3462 4333
rect 3508 4367 3562 4473
rect 3608 4507 3662 4519
rect 3608 4481 3618 4507
rect 3652 4481 3662 4507
rect 3608 4429 3609 4481
rect 3661 4429 3662 4481
rect 3608 4422 3662 4429
rect 3708 4507 3762 4613
rect 3808 4691 3862 4698
rect 3808 4639 3809 4691
rect 3861 4639 3862 4691
rect 3808 4613 3818 4639
rect 3852 4613 3862 4639
rect 3808 4601 3862 4613
rect 3908 4647 3962 4753
rect 4008 4787 4062 4799
rect 4008 4761 4018 4787
rect 4052 4761 4062 4787
rect 4008 4709 4009 4761
rect 4061 4709 4062 4761
rect 4008 4702 4062 4709
rect 4108 4787 4162 4960
rect 4202 4919 4268 4920
rect 4202 4867 4209 4919
rect 4261 4867 4268 4919
rect 4202 4866 4268 4867
rect 4108 4753 4118 4787
rect 4152 4753 4162 4787
rect 3908 4613 3918 4647
rect 3952 4613 3962 4647
rect 3708 4473 3718 4507
rect 3752 4473 3762 4507
rect 3508 4333 3518 4367
rect 3552 4333 3562 4367
rect 3308 4193 3318 4227
rect 3352 4193 3362 4227
rect 3108 4053 3118 4087
rect 3152 4053 3162 4087
rect 2908 3913 2918 3947
rect 2952 3913 2962 3947
rect 2708 3773 2718 3807
rect 2752 3773 2762 3807
rect 2602 3709 2668 3710
rect 2602 3657 2609 3709
rect 2661 3657 2668 3709
rect 2602 3656 2668 3657
rect 2508 3543 2518 3577
rect 2552 3543 2562 3577
rect 2308 3403 2318 3437
rect 2352 3403 2362 3437
rect 2108 3263 2118 3297
rect 2152 3263 2162 3297
rect 1908 3123 1918 3157
rect 1952 3123 1962 3157
rect 1708 2983 1718 3017
rect 1752 2983 1762 3017
rect 1508 2843 1518 2877
rect 1552 2843 1562 2877
rect 1308 2703 1318 2737
rect 1352 2703 1362 2737
rect 1108 2563 1118 2597
rect 1152 2563 1162 2597
rect 1002 2499 1068 2500
rect 1002 2447 1009 2499
rect 1061 2447 1068 2499
rect 1002 2446 1068 2447
rect 908 2333 918 2367
rect 952 2333 962 2367
rect 708 2193 718 2227
rect 752 2193 762 2227
rect 508 2053 518 2087
rect 552 2053 562 2087
rect 308 1913 318 1947
rect 352 1913 362 1947
rect 108 1773 118 1807
rect 152 1773 162 1807
rect 8 1667 62 1679
rect 8 1641 18 1667
rect 52 1641 62 1667
rect 8 1589 9 1641
rect 61 1589 62 1641
rect 8 1582 62 1589
rect 108 1667 162 1773
rect 208 1851 262 1858
rect 208 1799 209 1851
rect 261 1799 262 1851
rect 208 1773 218 1799
rect 252 1773 262 1799
rect 208 1761 262 1773
rect 308 1807 362 1913
rect 408 1947 462 1959
rect 408 1921 418 1947
rect 452 1921 462 1947
rect 408 1869 409 1921
rect 461 1869 462 1921
rect 408 1862 462 1869
rect 508 1947 562 2053
rect 608 2131 662 2138
rect 608 2079 609 2131
rect 661 2079 662 2131
rect 608 2053 618 2079
rect 652 2053 662 2079
rect 608 2041 662 2053
rect 708 2087 762 2193
rect 808 2227 862 2239
rect 808 2201 818 2227
rect 852 2201 862 2227
rect 808 2149 809 2201
rect 861 2149 862 2201
rect 808 2142 862 2149
rect 908 2227 962 2333
rect 1008 2411 1062 2418
rect 1008 2359 1009 2411
rect 1061 2359 1062 2411
rect 1008 2333 1018 2359
rect 1052 2333 1062 2359
rect 1008 2321 1062 2333
rect 1108 2367 1162 2563
rect 1208 2597 1262 2609
rect 1208 2571 1218 2597
rect 1252 2571 1262 2597
rect 1208 2519 1209 2571
rect 1261 2519 1262 2571
rect 1208 2512 1262 2519
rect 1308 2597 1362 2703
rect 1408 2781 1462 2788
rect 1408 2729 1409 2781
rect 1461 2729 1462 2781
rect 1408 2703 1418 2729
rect 1452 2703 1462 2729
rect 1408 2691 1462 2703
rect 1508 2737 1562 2843
rect 1608 2877 1662 2889
rect 1608 2851 1618 2877
rect 1652 2851 1662 2877
rect 1608 2799 1609 2851
rect 1661 2799 1662 2851
rect 1608 2792 1662 2799
rect 1708 2877 1762 2983
rect 1808 3061 1862 3068
rect 1808 3009 1809 3061
rect 1861 3009 1862 3061
rect 1808 2983 1818 3009
rect 1852 2983 1862 3009
rect 1808 2971 1862 2983
rect 1908 3017 1962 3123
rect 2008 3157 2062 3169
rect 2008 3131 2018 3157
rect 2052 3131 2062 3157
rect 2008 3079 2009 3131
rect 2061 3079 2062 3131
rect 2008 3072 2062 3079
rect 2108 3157 2162 3263
rect 2208 3341 2262 3348
rect 2208 3289 2209 3341
rect 2261 3289 2262 3341
rect 2208 3263 2218 3289
rect 2252 3263 2262 3289
rect 2208 3251 2262 3263
rect 2308 3297 2362 3403
rect 2408 3437 2462 3449
rect 2408 3411 2418 3437
rect 2452 3411 2462 3437
rect 2408 3359 2409 3411
rect 2461 3359 2462 3411
rect 2408 3352 2462 3359
rect 2508 3437 2562 3543
rect 2608 3621 2662 3628
rect 2608 3569 2609 3621
rect 2661 3569 2662 3621
rect 2608 3543 2618 3569
rect 2652 3543 2662 3569
rect 2608 3531 2662 3543
rect 2708 3577 2762 3773
rect 2808 3807 2862 3819
rect 2808 3781 2818 3807
rect 2852 3781 2862 3807
rect 2808 3729 2809 3781
rect 2861 3729 2862 3781
rect 2808 3722 2862 3729
rect 2908 3807 2962 3913
rect 3008 3991 3062 3998
rect 3008 3939 3009 3991
rect 3061 3939 3062 3991
rect 3008 3913 3018 3939
rect 3052 3913 3062 3939
rect 3008 3901 3062 3913
rect 3108 3947 3162 4053
rect 3208 4087 3262 4099
rect 3208 4061 3218 4087
rect 3252 4061 3262 4087
rect 3208 4009 3209 4061
rect 3261 4009 3262 4061
rect 3208 4002 3262 4009
rect 3308 4087 3362 4193
rect 3408 4271 3462 4278
rect 3408 4219 3409 4271
rect 3461 4219 3462 4271
rect 3408 4193 3418 4219
rect 3452 4193 3462 4219
rect 3408 4181 3462 4193
rect 3508 4227 3562 4333
rect 3608 4367 3662 4379
rect 3608 4341 3618 4367
rect 3652 4341 3662 4367
rect 3608 4289 3609 4341
rect 3661 4289 3662 4341
rect 3608 4282 3662 4289
rect 3708 4367 3762 4473
rect 3808 4551 3862 4558
rect 3808 4499 3809 4551
rect 3861 4499 3862 4551
rect 3808 4473 3818 4499
rect 3852 4473 3862 4499
rect 3808 4461 3862 4473
rect 3908 4507 3962 4613
rect 4008 4647 4062 4659
rect 4008 4621 4018 4647
rect 4052 4621 4062 4647
rect 4008 4569 4009 4621
rect 4061 4569 4062 4621
rect 4008 4562 4062 4569
rect 4108 4647 4162 4753
rect 4208 4831 4262 4838
rect 4208 4779 4209 4831
rect 4261 4779 4262 4831
rect 4208 4753 4218 4779
rect 4252 4753 4262 4779
rect 4208 4741 4262 4753
rect 4308 4787 4362 4960
rect 4402 4903 4468 4904
rect 4402 4851 4409 4903
rect 4461 4851 4468 4903
rect 4402 4850 4468 4851
rect 4308 4753 4318 4787
rect 4352 4753 4362 4787
rect 4108 4613 4118 4647
rect 4152 4613 4162 4647
rect 3908 4473 3918 4507
rect 3952 4473 3962 4507
rect 3708 4333 3718 4367
rect 3752 4333 3762 4367
rect 3508 4193 3518 4227
rect 3552 4193 3562 4227
rect 3308 4053 3318 4087
rect 3352 4053 3362 4087
rect 3108 3913 3118 3947
rect 3152 3913 3162 3947
rect 2908 3773 2918 3807
rect 2952 3773 2962 3807
rect 2802 3693 2868 3694
rect 2802 3641 2809 3693
rect 2861 3641 2868 3693
rect 2802 3640 2868 3641
rect 2708 3543 2718 3577
rect 2752 3543 2762 3577
rect 2508 3403 2518 3437
rect 2552 3403 2562 3437
rect 2308 3263 2318 3297
rect 2352 3263 2362 3297
rect 2108 3123 2118 3157
rect 2152 3123 2162 3157
rect 1908 2983 1918 3017
rect 1952 2983 1962 3017
rect 1708 2843 1718 2877
rect 1752 2843 1762 2877
rect 1508 2703 1518 2737
rect 1552 2703 1562 2737
rect 1308 2563 1318 2597
rect 1352 2563 1362 2597
rect 1202 2483 1268 2484
rect 1202 2431 1209 2483
rect 1261 2431 1268 2483
rect 1202 2430 1268 2431
rect 1108 2333 1118 2367
rect 1152 2333 1162 2367
rect 908 2193 918 2227
rect 952 2193 962 2227
rect 708 2053 718 2087
rect 752 2053 762 2087
rect 508 1913 518 1947
rect 552 1913 562 1947
rect 308 1773 318 1807
rect 352 1773 362 1807
rect 108 1633 118 1667
rect 152 1633 162 1667
rect 8 1527 62 1539
rect 8 1501 18 1527
rect 52 1501 62 1527
rect 8 1449 9 1501
rect 61 1449 62 1501
rect 8 1442 62 1449
rect 108 1527 162 1633
rect 208 1711 262 1718
rect 208 1659 209 1711
rect 261 1659 262 1711
rect 208 1633 218 1659
rect 252 1633 262 1659
rect 208 1621 262 1633
rect 308 1667 362 1773
rect 408 1807 462 1819
rect 408 1781 418 1807
rect 452 1781 462 1807
rect 408 1729 409 1781
rect 461 1729 462 1781
rect 408 1722 462 1729
rect 508 1807 562 1913
rect 608 1991 662 1998
rect 608 1939 609 1991
rect 661 1939 662 1991
rect 608 1913 618 1939
rect 652 1913 662 1939
rect 608 1901 662 1913
rect 708 1947 762 2053
rect 808 2087 862 2099
rect 808 2061 818 2087
rect 852 2061 862 2087
rect 808 2009 809 2061
rect 861 2009 862 2061
rect 808 2002 862 2009
rect 908 2087 962 2193
rect 1008 2271 1062 2278
rect 1008 2219 1009 2271
rect 1061 2219 1062 2271
rect 1008 2193 1018 2219
rect 1052 2193 1062 2219
rect 1008 2181 1062 2193
rect 1108 2227 1162 2333
rect 1208 2367 1262 2379
rect 1208 2341 1218 2367
rect 1252 2341 1262 2367
rect 1208 2289 1209 2341
rect 1261 2289 1262 2341
rect 1208 2282 1262 2289
rect 1308 2367 1362 2563
rect 1408 2641 1462 2648
rect 1408 2589 1409 2641
rect 1461 2589 1462 2641
rect 1408 2563 1418 2589
rect 1452 2563 1462 2589
rect 1408 2551 1462 2563
rect 1508 2597 1562 2703
rect 1608 2737 1662 2749
rect 1608 2711 1618 2737
rect 1652 2711 1662 2737
rect 1608 2659 1609 2711
rect 1661 2659 1662 2711
rect 1608 2652 1662 2659
rect 1708 2737 1762 2843
rect 1808 2921 1862 2928
rect 1808 2869 1809 2921
rect 1861 2869 1862 2921
rect 1808 2843 1818 2869
rect 1852 2843 1862 2869
rect 1808 2831 1862 2843
rect 1908 2877 1962 2983
rect 2008 3017 2062 3029
rect 2008 2991 2018 3017
rect 2052 2991 2062 3017
rect 2008 2939 2009 2991
rect 2061 2939 2062 2991
rect 2008 2932 2062 2939
rect 2108 3017 2162 3123
rect 2208 3201 2262 3208
rect 2208 3149 2209 3201
rect 2261 3149 2262 3201
rect 2208 3123 2218 3149
rect 2252 3123 2262 3149
rect 2208 3111 2262 3123
rect 2308 3157 2362 3263
rect 2408 3297 2462 3309
rect 2408 3271 2418 3297
rect 2452 3271 2462 3297
rect 2408 3219 2409 3271
rect 2461 3219 2462 3271
rect 2408 3212 2462 3219
rect 2508 3297 2562 3403
rect 2608 3481 2662 3488
rect 2608 3429 2609 3481
rect 2661 3429 2662 3481
rect 2608 3403 2618 3429
rect 2652 3403 2662 3429
rect 2608 3391 2662 3403
rect 2708 3437 2762 3543
rect 2808 3577 2862 3589
rect 2808 3551 2818 3577
rect 2852 3551 2862 3577
rect 2808 3499 2809 3551
rect 2861 3499 2862 3551
rect 2808 3492 2862 3499
rect 2908 3577 2962 3773
rect 3008 3851 3062 3858
rect 3008 3799 3009 3851
rect 3061 3799 3062 3851
rect 3008 3773 3018 3799
rect 3052 3773 3062 3799
rect 3008 3761 3062 3773
rect 3108 3807 3162 3913
rect 3208 3947 3262 3959
rect 3208 3921 3218 3947
rect 3252 3921 3262 3947
rect 3208 3869 3209 3921
rect 3261 3869 3262 3921
rect 3208 3862 3262 3869
rect 3308 3947 3362 4053
rect 3408 4131 3462 4138
rect 3408 4079 3409 4131
rect 3461 4079 3462 4131
rect 3408 4053 3418 4079
rect 3452 4053 3462 4079
rect 3408 4041 3462 4053
rect 3508 4087 3562 4193
rect 3608 4227 3662 4239
rect 3608 4201 3618 4227
rect 3652 4201 3662 4227
rect 3608 4149 3609 4201
rect 3661 4149 3662 4201
rect 3608 4142 3662 4149
rect 3708 4227 3762 4333
rect 3808 4411 3862 4418
rect 3808 4359 3809 4411
rect 3861 4359 3862 4411
rect 3808 4333 3818 4359
rect 3852 4333 3862 4359
rect 3808 4321 3862 4333
rect 3908 4367 3962 4473
rect 4008 4507 4062 4519
rect 4008 4481 4018 4507
rect 4052 4481 4062 4507
rect 4008 4429 4009 4481
rect 4061 4429 4062 4481
rect 4008 4422 4062 4429
rect 4108 4507 4162 4613
rect 4208 4691 4262 4698
rect 4208 4639 4209 4691
rect 4261 4639 4262 4691
rect 4208 4613 4218 4639
rect 4252 4613 4262 4639
rect 4208 4601 4262 4613
rect 4308 4647 4362 4753
rect 4408 4787 4462 4799
rect 4408 4761 4418 4787
rect 4452 4761 4462 4787
rect 4408 4709 4409 4761
rect 4461 4709 4462 4761
rect 4408 4702 4462 4709
rect 4508 4787 4562 4960
rect 4602 4919 4668 4920
rect 4602 4867 4609 4919
rect 4661 4867 4668 4919
rect 4602 4866 4668 4867
rect 4508 4753 4518 4787
rect 4552 4753 4562 4787
rect 4308 4613 4318 4647
rect 4352 4613 4362 4647
rect 4108 4473 4118 4507
rect 4152 4473 4162 4507
rect 3908 4333 3918 4367
rect 3952 4333 3962 4367
rect 3708 4193 3718 4227
rect 3752 4193 3762 4227
rect 3508 4053 3518 4087
rect 3552 4053 3562 4087
rect 3308 3913 3318 3947
rect 3352 3913 3362 3947
rect 3108 3773 3118 3807
rect 3152 3773 3162 3807
rect 3002 3709 3068 3710
rect 3002 3657 3009 3709
rect 3061 3657 3068 3709
rect 3002 3656 3068 3657
rect 2908 3543 2918 3577
rect 2952 3543 2962 3577
rect 2708 3403 2718 3437
rect 2752 3403 2762 3437
rect 2508 3263 2518 3297
rect 2552 3263 2562 3297
rect 2308 3123 2318 3157
rect 2352 3123 2362 3157
rect 2108 2983 2118 3017
rect 2152 2983 2162 3017
rect 1908 2843 1918 2877
rect 1952 2843 1962 2877
rect 1708 2703 1718 2737
rect 1752 2703 1762 2737
rect 1508 2563 1518 2597
rect 1552 2563 1562 2597
rect 1402 2499 1468 2500
rect 1402 2447 1409 2499
rect 1461 2447 1468 2499
rect 1402 2446 1468 2447
rect 1308 2333 1318 2367
rect 1352 2333 1362 2367
rect 1108 2193 1118 2227
rect 1152 2193 1162 2227
rect 908 2053 918 2087
rect 952 2053 962 2087
rect 708 1913 718 1947
rect 752 1913 762 1947
rect 508 1773 518 1807
rect 552 1773 562 1807
rect 308 1633 318 1667
rect 352 1633 362 1667
rect 108 1493 118 1527
rect 152 1493 162 1527
rect 8 1387 62 1399
rect 8 1361 18 1387
rect 52 1361 62 1387
rect 8 1309 9 1361
rect 61 1309 62 1361
rect 8 1302 62 1309
rect 108 1387 162 1493
rect 208 1571 262 1578
rect 208 1519 209 1571
rect 261 1519 262 1571
rect 208 1493 218 1519
rect 252 1493 262 1519
rect 208 1481 262 1493
rect 308 1527 362 1633
rect 408 1667 462 1679
rect 408 1641 418 1667
rect 452 1641 462 1667
rect 408 1589 409 1641
rect 461 1589 462 1641
rect 408 1582 462 1589
rect 508 1667 562 1773
rect 608 1851 662 1858
rect 608 1799 609 1851
rect 661 1799 662 1851
rect 608 1773 618 1799
rect 652 1773 662 1799
rect 608 1761 662 1773
rect 708 1807 762 1913
rect 808 1947 862 1959
rect 808 1921 818 1947
rect 852 1921 862 1947
rect 808 1869 809 1921
rect 861 1869 862 1921
rect 808 1862 862 1869
rect 908 1947 962 2053
rect 1008 2131 1062 2138
rect 1008 2079 1009 2131
rect 1061 2079 1062 2131
rect 1008 2053 1018 2079
rect 1052 2053 1062 2079
rect 1008 2041 1062 2053
rect 1108 2087 1162 2193
rect 1208 2227 1262 2239
rect 1208 2201 1218 2227
rect 1252 2201 1262 2227
rect 1208 2149 1209 2201
rect 1261 2149 1262 2201
rect 1208 2142 1262 2149
rect 1308 2227 1362 2333
rect 1408 2411 1462 2418
rect 1408 2359 1409 2411
rect 1461 2359 1462 2411
rect 1408 2333 1418 2359
rect 1452 2333 1462 2359
rect 1408 2321 1462 2333
rect 1508 2367 1562 2563
rect 1608 2597 1662 2609
rect 1608 2571 1618 2597
rect 1652 2571 1662 2597
rect 1608 2519 1609 2571
rect 1661 2519 1662 2571
rect 1608 2512 1662 2519
rect 1708 2597 1762 2703
rect 1808 2781 1862 2788
rect 1808 2729 1809 2781
rect 1861 2729 1862 2781
rect 1808 2703 1818 2729
rect 1852 2703 1862 2729
rect 1808 2691 1862 2703
rect 1908 2737 1962 2843
rect 2008 2877 2062 2889
rect 2008 2851 2018 2877
rect 2052 2851 2062 2877
rect 2008 2799 2009 2851
rect 2061 2799 2062 2851
rect 2008 2792 2062 2799
rect 2108 2877 2162 2983
rect 2208 3061 2262 3068
rect 2208 3009 2209 3061
rect 2261 3009 2262 3061
rect 2208 2983 2218 3009
rect 2252 2983 2262 3009
rect 2208 2971 2262 2983
rect 2308 3017 2362 3123
rect 2408 3157 2462 3169
rect 2408 3131 2418 3157
rect 2452 3131 2462 3157
rect 2408 3079 2409 3131
rect 2461 3079 2462 3131
rect 2408 3072 2462 3079
rect 2508 3157 2562 3263
rect 2608 3341 2662 3348
rect 2608 3289 2609 3341
rect 2661 3289 2662 3341
rect 2608 3263 2618 3289
rect 2652 3263 2662 3289
rect 2608 3251 2662 3263
rect 2708 3297 2762 3403
rect 2808 3437 2862 3449
rect 2808 3411 2818 3437
rect 2852 3411 2862 3437
rect 2808 3359 2809 3411
rect 2861 3359 2862 3411
rect 2808 3352 2862 3359
rect 2908 3437 2962 3543
rect 3008 3621 3062 3628
rect 3008 3569 3009 3621
rect 3061 3569 3062 3621
rect 3008 3543 3018 3569
rect 3052 3543 3062 3569
rect 3008 3531 3062 3543
rect 3108 3577 3162 3773
rect 3208 3807 3262 3819
rect 3208 3781 3218 3807
rect 3252 3781 3262 3807
rect 3208 3729 3209 3781
rect 3261 3729 3262 3781
rect 3208 3722 3262 3729
rect 3308 3807 3362 3913
rect 3408 3991 3462 3998
rect 3408 3939 3409 3991
rect 3461 3939 3462 3991
rect 3408 3913 3418 3939
rect 3452 3913 3462 3939
rect 3408 3901 3462 3913
rect 3508 3947 3562 4053
rect 3608 4087 3662 4099
rect 3608 4061 3618 4087
rect 3652 4061 3662 4087
rect 3608 4009 3609 4061
rect 3661 4009 3662 4061
rect 3608 4002 3662 4009
rect 3708 4087 3762 4193
rect 3808 4271 3862 4278
rect 3808 4219 3809 4271
rect 3861 4219 3862 4271
rect 3808 4193 3818 4219
rect 3852 4193 3862 4219
rect 3808 4181 3862 4193
rect 3908 4227 3962 4333
rect 4008 4367 4062 4379
rect 4008 4341 4018 4367
rect 4052 4341 4062 4367
rect 4008 4289 4009 4341
rect 4061 4289 4062 4341
rect 4008 4282 4062 4289
rect 4108 4367 4162 4473
rect 4208 4551 4262 4558
rect 4208 4499 4209 4551
rect 4261 4499 4262 4551
rect 4208 4473 4218 4499
rect 4252 4473 4262 4499
rect 4208 4461 4262 4473
rect 4308 4507 4362 4613
rect 4408 4647 4462 4659
rect 4408 4621 4418 4647
rect 4452 4621 4462 4647
rect 4408 4569 4409 4621
rect 4461 4569 4462 4621
rect 4408 4562 4462 4569
rect 4508 4647 4562 4753
rect 4608 4831 4662 4838
rect 4608 4779 4609 4831
rect 4661 4779 4662 4831
rect 4608 4753 4618 4779
rect 4652 4753 4662 4779
rect 4608 4741 4662 4753
rect 4708 4787 4762 4960
rect 4802 4903 4868 4904
rect 4802 4851 4809 4903
rect 4861 4851 4868 4903
rect 4802 4850 4868 4851
rect 4708 4753 4718 4787
rect 4752 4753 4762 4787
rect 4508 4613 4518 4647
rect 4552 4613 4562 4647
rect 4308 4473 4318 4507
rect 4352 4473 4362 4507
rect 4108 4333 4118 4367
rect 4152 4333 4162 4367
rect 3908 4193 3918 4227
rect 3952 4193 3962 4227
rect 3708 4053 3718 4087
rect 3752 4053 3762 4087
rect 3508 3913 3518 3947
rect 3552 3913 3562 3947
rect 3308 3773 3318 3807
rect 3352 3773 3362 3807
rect 3202 3693 3268 3694
rect 3202 3641 3209 3693
rect 3261 3641 3268 3693
rect 3202 3640 3268 3641
rect 3108 3543 3118 3577
rect 3152 3543 3162 3577
rect 2908 3403 2918 3437
rect 2952 3403 2962 3437
rect 2708 3263 2718 3297
rect 2752 3263 2762 3297
rect 2508 3123 2518 3157
rect 2552 3123 2562 3157
rect 2308 2983 2318 3017
rect 2352 2983 2362 3017
rect 2108 2843 2118 2877
rect 2152 2843 2162 2877
rect 1908 2703 1918 2737
rect 1952 2703 1962 2737
rect 1708 2563 1718 2597
rect 1752 2563 1762 2597
rect 1602 2483 1668 2484
rect 1602 2431 1609 2483
rect 1661 2431 1668 2483
rect 1602 2430 1668 2431
rect 1508 2333 1518 2367
rect 1552 2333 1562 2367
rect 1308 2193 1318 2227
rect 1352 2193 1362 2227
rect 1108 2053 1118 2087
rect 1152 2053 1162 2087
rect 908 1913 918 1947
rect 952 1913 962 1947
rect 708 1773 718 1807
rect 752 1773 762 1807
rect 508 1633 518 1667
rect 552 1633 562 1667
rect 308 1493 318 1527
rect 352 1493 362 1527
rect 108 1353 118 1387
rect 152 1353 162 1387
rect 2 1273 68 1274
rect 2 1221 9 1273
rect 61 1221 68 1273
rect 2 1220 68 1221
rect 8 1157 62 1169
rect 8 1131 18 1157
rect 52 1131 62 1157
rect 8 1079 9 1131
rect 61 1079 62 1131
rect 8 1072 62 1079
rect 108 1157 162 1353
rect 208 1431 262 1438
rect 208 1379 209 1431
rect 261 1379 262 1431
rect 208 1353 218 1379
rect 252 1353 262 1379
rect 208 1341 262 1353
rect 308 1387 362 1493
rect 408 1527 462 1539
rect 408 1501 418 1527
rect 452 1501 462 1527
rect 408 1449 409 1501
rect 461 1449 462 1501
rect 408 1442 462 1449
rect 508 1527 562 1633
rect 608 1711 662 1718
rect 608 1659 609 1711
rect 661 1659 662 1711
rect 608 1633 618 1659
rect 652 1633 662 1659
rect 608 1621 662 1633
rect 708 1667 762 1773
rect 808 1807 862 1819
rect 808 1781 818 1807
rect 852 1781 862 1807
rect 808 1729 809 1781
rect 861 1729 862 1781
rect 808 1722 862 1729
rect 908 1807 962 1913
rect 1008 1991 1062 1998
rect 1008 1939 1009 1991
rect 1061 1939 1062 1991
rect 1008 1913 1018 1939
rect 1052 1913 1062 1939
rect 1008 1901 1062 1913
rect 1108 1947 1162 2053
rect 1208 2087 1262 2099
rect 1208 2061 1218 2087
rect 1252 2061 1262 2087
rect 1208 2009 1209 2061
rect 1261 2009 1262 2061
rect 1208 2002 1262 2009
rect 1308 2087 1362 2193
rect 1408 2271 1462 2278
rect 1408 2219 1409 2271
rect 1461 2219 1462 2271
rect 1408 2193 1418 2219
rect 1452 2193 1462 2219
rect 1408 2181 1462 2193
rect 1508 2227 1562 2333
rect 1608 2367 1662 2379
rect 1608 2341 1618 2367
rect 1652 2341 1662 2367
rect 1608 2289 1609 2341
rect 1661 2289 1662 2341
rect 1608 2282 1662 2289
rect 1708 2367 1762 2563
rect 1808 2641 1862 2648
rect 1808 2589 1809 2641
rect 1861 2589 1862 2641
rect 1808 2563 1818 2589
rect 1852 2563 1862 2589
rect 1808 2551 1862 2563
rect 1908 2597 1962 2703
rect 2008 2737 2062 2749
rect 2008 2711 2018 2737
rect 2052 2711 2062 2737
rect 2008 2659 2009 2711
rect 2061 2659 2062 2711
rect 2008 2652 2062 2659
rect 2108 2737 2162 2843
rect 2208 2921 2262 2928
rect 2208 2869 2209 2921
rect 2261 2869 2262 2921
rect 2208 2843 2218 2869
rect 2252 2843 2262 2869
rect 2208 2831 2262 2843
rect 2308 2877 2362 2983
rect 2408 3017 2462 3029
rect 2408 2991 2418 3017
rect 2452 2991 2462 3017
rect 2408 2939 2409 2991
rect 2461 2939 2462 2991
rect 2408 2932 2462 2939
rect 2508 3017 2562 3123
rect 2608 3201 2662 3208
rect 2608 3149 2609 3201
rect 2661 3149 2662 3201
rect 2608 3123 2618 3149
rect 2652 3123 2662 3149
rect 2608 3111 2662 3123
rect 2708 3157 2762 3263
rect 2808 3297 2862 3309
rect 2808 3271 2818 3297
rect 2852 3271 2862 3297
rect 2808 3219 2809 3271
rect 2861 3219 2862 3271
rect 2808 3212 2862 3219
rect 2908 3297 2962 3403
rect 3008 3481 3062 3488
rect 3008 3429 3009 3481
rect 3061 3429 3062 3481
rect 3008 3403 3018 3429
rect 3052 3403 3062 3429
rect 3008 3391 3062 3403
rect 3108 3437 3162 3543
rect 3208 3577 3262 3589
rect 3208 3551 3218 3577
rect 3252 3551 3262 3577
rect 3208 3499 3209 3551
rect 3261 3499 3262 3551
rect 3208 3492 3262 3499
rect 3308 3577 3362 3773
rect 3408 3851 3462 3858
rect 3408 3799 3409 3851
rect 3461 3799 3462 3851
rect 3408 3773 3418 3799
rect 3452 3773 3462 3799
rect 3408 3761 3462 3773
rect 3508 3807 3562 3913
rect 3608 3947 3662 3959
rect 3608 3921 3618 3947
rect 3652 3921 3662 3947
rect 3608 3869 3609 3921
rect 3661 3869 3662 3921
rect 3608 3862 3662 3869
rect 3708 3947 3762 4053
rect 3808 4131 3862 4138
rect 3808 4079 3809 4131
rect 3861 4079 3862 4131
rect 3808 4053 3818 4079
rect 3852 4053 3862 4079
rect 3808 4041 3862 4053
rect 3908 4087 3962 4193
rect 4008 4227 4062 4239
rect 4008 4201 4018 4227
rect 4052 4201 4062 4227
rect 4008 4149 4009 4201
rect 4061 4149 4062 4201
rect 4008 4142 4062 4149
rect 4108 4227 4162 4333
rect 4208 4411 4262 4418
rect 4208 4359 4209 4411
rect 4261 4359 4262 4411
rect 4208 4333 4218 4359
rect 4252 4333 4262 4359
rect 4208 4321 4262 4333
rect 4308 4367 4362 4473
rect 4408 4507 4462 4519
rect 4408 4481 4418 4507
rect 4452 4481 4462 4507
rect 4408 4429 4409 4481
rect 4461 4429 4462 4481
rect 4408 4422 4462 4429
rect 4508 4507 4562 4613
rect 4608 4691 4662 4698
rect 4608 4639 4609 4691
rect 4661 4639 4662 4691
rect 4608 4613 4618 4639
rect 4652 4613 4662 4639
rect 4608 4601 4662 4613
rect 4708 4647 4762 4753
rect 4808 4787 4862 4799
rect 4808 4761 4818 4787
rect 4852 4761 4862 4787
rect 4808 4709 4809 4761
rect 4861 4709 4862 4761
rect 4808 4702 4862 4709
rect 4908 4787 4962 4960
rect 5002 4919 5068 4920
rect 5002 4867 5009 4919
rect 5061 4867 5068 4919
rect 5002 4866 5068 4867
rect 4908 4753 4918 4787
rect 4952 4753 4962 4787
rect 4708 4613 4718 4647
rect 4752 4613 4762 4647
rect 4508 4473 4518 4507
rect 4552 4473 4562 4507
rect 4308 4333 4318 4367
rect 4352 4333 4362 4367
rect 4108 4193 4118 4227
rect 4152 4193 4162 4227
rect 3908 4053 3918 4087
rect 3952 4053 3962 4087
rect 3708 3913 3718 3947
rect 3752 3913 3762 3947
rect 3508 3773 3518 3807
rect 3552 3773 3562 3807
rect 3402 3709 3468 3710
rect 3402 3657 3409 3709
rect 3461 3657 3468 3709
rect 3402 3656 3468 3657
rect 3308 3543 3318 3577
rect 3352 3543 3362 3577
rect 3108 3403 3118 3437
rect 3152 3403 3162 3437
rect 2908 3263 2918 3297
rect 2952 3263 2962 3297
rect 2708 3123 2718 3157
rect 2752 3123 2762 3157
rect 2508 2983 2518 3017
rect 2552 2983 2562 3017
rect 2308 2843 2318 2877
rect 2352 2843 2362 2877
rect 2108 2703 2118 2737
rect 2152 2703 2162 2737
rect 1908 2563 1918 2597
rect 1952 2563 1962 2597
rect 1802 2499 1868 2500
rect 1802 2447 1809 2499
rect 1861 2447 1868 2499
rect 1802 2446 1868 2447
rect 1708 2333 1718 2367
rect 1752 2333 1762 2367
rect 1508 2193 1518 2227
rect 1552 2193 1562 2227
rect 1308 2053 1318 2087
rect 1352 2053 1362 2087
rect 1108 1913 1118 1947
rect 1152 1913 1162 1947
rect 908 1773 918 1807
rect 952 1773 962 1807
rect 708 1633 718 1667
rect 752 1633 762 1667
rect 508 1493 518 1527
rect 552 1493 562 1527
rect 308 1353 318 1387
rect 352 1353 362 1387
rect 202 1289 268 1290
rect 202 1237 209 1289
rect 261 1237 268 1289
rect 202 1236 268 1237
rect 108 1123 118 1157
rect 152 1123 162 1157
rect 8 1017 62 1029
rect 8 991 18 1017
rect 52 991 62 1017
rect 8 939 9 991
rect 61 939 62 991
rect 8 932 62 939
rect 108 1017 162 1123
rect 208 1201 262 1208
rect 208 1149 209 1201
rect 261 1149 262 1201
rect 208 1123 218 1149
rect 252 1123 262 1149
rect 208 1111 262 1123
rect 308 1157 362 1353
rect 408 1387 462 1399
rect 408 1361 418 1387
rect 452 1361 462 1387
rect 408 1309 409 1361
rect 461 1309 462 1361
rect 408 1302 462 1309
rect 508 1387 562 1493
rect 608 1571 662 1578
rect 608 1519 609 1571
rect 661 1519 662 1571
rect 608 1493 618 1519
rect 652 1493 662 1519
rect 608 1481 662 1493
rect 708 1527 762 1633
rect 808 1667 862 1679
rect 808 1641 818 1667
rect 852 1641 862 1667
rect 808 1589 809 1641
rect 861 1589 862 1641
rect 808 1582 862 1589
rect 908 1667 962 1773
rect 1008 1851 1062 1858
rect 1008 1799 1009 1851
rect 1061 1799 1062 1851
rect 1008 1773 1018 1799
rect 1052 1773 1062 1799
rect 1008 1761 1062 1773
rect 1108 1807 1162 1913
rect 1208 1947 1262 1959
rect 1208 1921 1218 1947
rect 1252 1921 1262 1947
rect 1208 1869 1209 1921
rect 1261 1869 1262 1921
rect 1208 1862 1262 1869
rect 1308 1947 1362 2053
rect 1408 2131 1462 2138
rect 1408 2079 1409 2131
rect 1461 2079 1462 2131
rect 1408 2053 1418 2079
rect 1452 2053 1462 2079
rect 1408 2041 1462 2053
rect 1508 2087 1562 2193
rect 1608 2227 1662 2239
rect 1608 2201 1618 2227
rect 1652 2201 1662 2227
rect 1608 2149 1609 2201
rect 1661 2149 1662 2201
rect 1608 2142 1662 2149
rect 1708 2227 1762 2333
rect 1808 2411 1862 2418
rect 1808 2359 1809 2411
rect 1861 2359 1862 2411
rect 1808 2333 1818 2359
rect 1852 2333 1862 2359
rect 1808 2321 1862 2333
rect 1908 2367 1962 2563
rect 2008 2597 2062 2609
rect 2008 2571 2018 2597
rect 2052 2571 2062 2597
rect 2008 2519 2009 2571
rect 2061 2519 2062 2571
rect 2008 2512 2062 2519
rect 2108 2597 2162 2703
rect 2208 2781 2262 2788
rect 2208 2729 2209 2781
rect 2261 2729 2262 2781
rect 2208 2703 2218 2729
rect 2252 2703 2262 2729
rect 2208 2691 2262 2703
rect 2308 2737 2362 2843
rect 2408 2877 2462 2889
rect 2408 2851 2418 2877
rect 2452 2851 2462 2877
rect 2408 2799 2409 2851
rect 2461 2799 2462 2851
rect 2408 2792 2462 2799
rect 2508 2877 2562 2983
rect 2608 3061 2662 3068
rect 2608 3009 2609 3061
rect 2661 3009 2662 3061
rect 2608 2983 2618 3009
rect 2652 2983 2662 3009
rect 2608 2971 2662 2983
rect 2708 3017 2762 3123
rect 2808 3157 2862 3169
rect 2808 3131 2818 3157
rect 2852 3131 2862 3157
rect 2808 3079 2809 3131
rect 2861 3079 2862 3131
rect 2808 3072 2862 3079
rect 2908 3157 2962 3263
rect 3008 3341 3062 3348
rect 3008 3289 3009 3341
rect 3061 3289 3062 3341
rect 3008 3263 3018 3289
rect 3052 3263 3062 3289
rect 3008 3251 3062 3263
rect 3108 3297 3162 3403
rect 3208 3437 3262 3449
rect 3208 3411 3218 3437
rect 3252 3411 3262 3437
rect 3208 3359 3209 3411
rect 3261 3359 3262 3411
rect 3208 3352 3262 3359
rect 3308 3437 3362 3543
rect 3408 3621 3462 3628
rect 3408 3569 3409 3621
rect 3461 3569 3462 3621
rect 3408 3543 3418 3569
rect 3452 3543 3462 3569
rect 3408 3531 3462 3543
rect 3508 3577 3562 3773
rect 3608 3807 3662 3819
rect 3608 3781 3618 3807
rect 3652 3781 3662 3807
rect 3608 3729 3609 3781
rect 3661 3729 3662 3781
rect 3608 3722 3662 3729
rect 3708 3807 3762 3913
rect 3808 3991 3862 3998
rect 3808 3939 3809 3991
rect 3861 3939 3862 3991
rect 3808 3913 3818 3939
rect 3852 3913 3862 3939
rect 3808 3901 3862 3913
rect 3908 3947 3962 4053
rect 4008 4087 4062 4099
rect 4008 4061 4018 4087
rect 4052 4061 4062 4087
rect 4008 4009 4009 4061
rect 4061 4009 4062 4061
rect 4008 4002 4062 4009
rect 4108 4087 4162 4193
rect 4208 4271 4262 4278
rect 4208 4219 4209 4271
rect 4261 4219 4262 4271
rect 4208 4193 4218 4219
rect 4252 4193 4262 4219
rect 4208 4181 4262 4193
rect 4308 4227 4362 4333
rect 4408 4367 4462 4379
rect 4408 4341 4418 4367
rect 4452 4341 4462 4367
rect 4408 4289 4409 4341
rect 4461 4289 4462 4341
rect 4408 4282 4462 4289
rect 4508 4367 4562 4473
rect 4608 4551 4662 4558
rect 4608 4499 4609 4551
rect 4661 4499 4662 4551
rect 4608 4473 4618 4499
rect 4652 4473 4662 4499
rect 4608 4461 4662 4473
rect 4708 4507 4762 4613
rect 4808 4647 4862 4659
rect 4808 4621 4818 4647
rect 4852 4621 4862 4647
rect 4808 4569 4809 4621
rect 4861 4569 4862 4621
rect 4808 4562 4862 4569
rect 4908 4647 4962 4753
rect 5008 4831 5062 4838
rect 5008 4779 5009 4831
rect 5061 4779 5062 4831
rect 5008 4753 5018 4779
rect 5052 4753 5062 4779
rect 5008 4741 5062 4753
rect 5108 4787 5162 4960
rect 5202 4903 5268 4904
rect 5202 4851 5209 4903
rect 5261 4851 5268 4903
rect 5202 4850 5268 4851
rect 5108 4753 5118 4787
rect 5152 4753 5162 4787
rect 4908 4613 4918 4647
rect 4952 4613 4962 4647
rect 4708 4473 4718 4507
rect 4752 4473 4762 4507
rect 4508 4333 4518 4367
rect 4552 4333 4562 4367
rect 4308 4193 4318 4227
rect 4352 4193 4362 4227
rect 4108 4053 4118 4087
rect 4152 4053 4162 4087
rect 3908 3913 3918 3947
rect 3952 3913 3962 3947
rect 3708 3773 3718 3807
rect 3752 3773 3762 3807
rect 3602 3693 3668 3694
rect 3602 3641 3609 3693
rect 3661 3641 3668 3693
rect 3602 3640 3668 3641
rect 3508 3543 3518 3577
rect 3552 3543 3562 3577
rect 3308 3403 3318 3437
rect 3352 3403 3362 3437
rect 3108 3263 3118 3297
rect 3152 3263 3162 3297
rect 2908 3123 2918 3157
rect 2952 3123 2962 3157
rect 2708 2983 2718 3017
rect 2752 2983 2762 3017
rect 2508 2843 2518 2877
rect 2552 2843 2562 2877
rect 2308 2703 2318 2737
rect 2352 2703 2362 2737
rect 2108 2563 2118 2597
rect 2152 2563 2162 2597
rect 2002 2483 2068 2484
rect 2002 2431 2009 2483
rect 2061 2431 2068 2483
rect 2002 2430 2068 2431
rect 1908 2333 1918 2367
rect 1952 2333 1962 2367
rect 1708 2193 1718 2227
rect 1752 2193 1762 2227
rect 1508 2053 1518 2087
rect 1552 2053 1562 2087
rect 1308 1913 1318 1947
rect 1352 1913 1362 1947
rect 1108 1773 1118 1807
rect 1152 1773 1162 1807
rect 908 1633 918 1667
rect 952 1633 962 1667
rect 708 1493 718 1527
rect 752 1493 762 1527
rect 508 1353 518 1387
rect 552 1353 562 1387
rect 402 1273 468 1274
rect 402 1221 409 1273
rect 461 1221 468 1273
rect 402 1220 468 1221
rect 308 1123 318 1157
rect 352 1123 362 1157
rect 108 983 118 1017
rect 152 983 162 1017
rect 8 877 62 889
rect 8 851 18 877
rect 52 851 62 877
rect 8 799 9 851
rect 61 799 62 851
rect 8 792 62 799
rect 108 877 162 983
rect 208 1061 262 1068
rect 208 1009 209 1061
rect 261 1009 262 1061
rect 208 983 218 1009
rect 252 983 262 1009
rect 208 971 262 983
rect 308 1017 362 1123
rect 408 1157 462 1169
rect 408 1131 418 1157
rect 452 1131 462 1157
rect 408 1079 409 1131
rect 461 1079 462 1131
rect 408 1072 462 1079
rect 508 1157 562 1353
rect 608 1431 662 1438
rect 608 1379 609 1431
rect 661 1379 662 1431
rect 608 1353 618 1379
rect 652 1353 662 1379
rect 608 1341 662 1353
rect 708 1387 762 1493
rect 808 1527 862 1539
rect 808 1501 818 1527
rect 852 1501 862 1527
rect 808 1449 809 1501
rect 861 1449 862 1501
rect 808 1442 862 1449
rect 908 1527 962 1633
rect 1008 1711 1062 1718
rect 1008 1659 1009 1711
rect 1061 1659 1062 1711
rect 1008 1633 1018 1659
rect 1052 1633 1062 1659
rect 1008 1621 1062 1633
rect 1108 1667 1162 1773
rect 1208 1807 1262 1819
rect 1208 1781 1218 1807
rect 1252 1781 1262 1807
rect 1208 1729 1209 1781
rect 1261 1729 1262 1781
rect 1208 1722 1262 1729
rect 1308 1807 1362 1913
rect 1408 1991 1462 1998
rect 1408 1939 1409 1991
rect 1461 1939 1462 1991
rect 1408 1913 1418 1939
rect 1452 1913 1462 1939
rect 1408 1901 1462 1913
rect 1508 1947 1562 2053
rect 1608 2087 1662 2099
rect 1608 2061 1618 2087
rect 1652 2061 1662 2087
rect 1608 2009 1609 2061
rect 1661 2009 1662 2061
rect 1608 2002 1662 2009
rect 1708 2087 1762 2193
rect 1808 2271 1862 2278
rect 1808 2219 1809 2271
rect 1861 2219 1862 2271
rect 1808 2193 1818 2219
rect 1852 2193 1862 2219
rect 1808 2181 1862 2193
rect 1908 2227 1962 2333
rect 2008 2367 2062 2379
rect 2008 2341 2018 2367
rect 2052 2341 2062 2367
rect 2008 2289 2009 2341
rect 2061 2289 2062 2341
rect 2008 2282 2062 2289
rect 2108 2367 2162 2563
rect 2208 2641 2262 2648
rect 2208 2589 2209 2641
rect 2261 2589 2262 2641
rect 2208 2563 2218 2589
rect 2252 2563 2262 2589
rect 2208 2551 2262 2563
rect 2308 2597 2362 2703
rect 2408 2737 2462 2749
rect 2408 2711 2418 2737
rect 2452 2711 2462 2737
rect 2408 2659 2409 2711
rect 2461 2659 2462 2711
rect 2408 2652 2462 2659
rect 2508 2737 2562 2843
rect 2608 2921 2662 2928
rect 2608 2869 2609 2921
rect 2661 2869 2662 2921
rect 2608 2843 2618 2869
rect 2652 2843 2662 2869
rect 2608 2831 2662 2843
rect 2708 2877 2762 2983
rect 2808 3017 2862 3029
rect 2808 2991 2818 3017
rect 2852 2991 2862 3017
rect 2808 2939 2809 2991
rect 2861 2939 2862 2991
rect 2808 2932 2862 2939
rect 2908 3017 2962 3123
rect 3008 3201 3062 3208
rect 3008 3149 3009 3201
rect 3061 3149 3062 3201
rect 3008 3123 3018 3149
rect 3052 3123 3062 3149
rect 3008 3111 3062 3123
rect 3108 3157 3162 3263
rect 3208 3297 3262 3309
rect 3208 3271 3218 3297
rect 3252 3271 3262 3297
rect 3208 3219 3209 3271
rect 3261 3219 3262 3271
rect 3208 3212 3262 3219
rect 3308 3297 3362 3403
rect 3408 3481 3462 3488
rect 3408 3429 3409 3481
rect 3461 3429 3462 3481
rect 3408 3403 3418 3429
rect 3452 3403 3462 3429
rect 3408 3391 3462 3403
rect 3508 3437 3562 3543
rect 3608 3577 3662 3589
rect 3608 3551 3618 3577
rect 3652 3551 3662 3577
rect 3608 3499 3609 3551
rect 3661 3499 3662 3551
rect 3608 3492 3662 3499
rect 3708 3577 3762 3773
rect 3808 3851 3862 3858
rect 3808 3799 3809 3851
rect 3861 3799 3862 3851
rect 3808 3773 3818 3799
rect 3852 3773 3862 3799
rect 3808 3761 3862 3773
rect 3908 3807 3962 3913
rect 4008 3947 4062 3959
rect 4008 3921 4018 3947
rect 4052 3921 4062 3947
rect 4008 3869 4009 3921
rect 4061 3869 4062 3921
rect 4008 3862 4062 3869
rect 4108 3947 4162 4053
rect 4208 4131 4262 4138
rect 4208 4079 4209 4131
rect 4261 4079 4262 4131
rect 4208 4053 4218 4079
rect 4252 4053 4262 4079
rect 4208 4041 4262 4053
rect 4308 4087 4362 4193
rect 4408 4227 4462 4239
rect 4408 4201 4418 4227
rect 4452 4201 4462 4227
rect 4408 4149 4409 4201
rect 4461 4149 4462 4201
rect 4408 4142 4462 4149
rect 4508 4227 4562 4333
rect 4608 4411 4662 4418
rect 4608 4359 4609 4411
rect 4661 4359 4662 4411
rect 4608 4333 4618 4359
rect 4652 4333 4662 4359
rect 4608 4321 4662 4333
rect 4708 4367 4762 4473
rect 4808 4507 4862 4519
rect 4808 4481 4818 4507
rect 4852 4481 4862 4507
rect 4808 4429 4809 4481
rect 4861 4429 4862 4481
rect 4808 4422 4862 4429
rect 4908 4507 4962 4613
rect 5008 4691 5062 4698
rect 5008 4639 5009 4691
rect 5061 4639 5062 4691
rect 5008 4613 5018 4639
rect 5052 4613 5062 4639
rect 5008 4601 5062 4613
rect 5108 4647 5162 4753
rect 5208 4787 5262 4799
rect 5208 4761 5218 4787
rect 5252 4761 5262 4787
rect 5208 4709 5209 4761
rect 5261 4709 5262 4761
rect 5208 4702 5262 4709
rect 5308 4787 5362 4960
rect 5402 4919 5468 4920
rect 5402 4867 5409 4919
rect 5461 4867 5468 4919
rect 5402 4866 5468 4867
rect 5308 4753 5318 4787
rect 5352 4753 5362 4787
rect 5108 4613 5118 4647
rect 5152 4613 5162 4647
rect 4908 4473 4918 4507
rect 4952 4473 4962 4507
rect 4708 4333 4718 4367
rect 4752 4333 4762 4367
rect 4508 4193 4518 4227
rect 4552 4193 4562 4227
rect 4308 4053 4318 4087
rect 4352 4053 4362 4087
rect 4108 3913 4118 3947
rect 4152 3913 4162 3947
rect 3908 3773 3918 3807
rect 3952 3773 3962 3807
rect 3802 3709 3868 3710
rect 3802 3657 3809 3709
rect 3861 3657 3868 3709
rect 3802 3656 3868 3657
rect 3708 3543 3718 3577
rect 3752 3543 3762 3577
rect 3508 3403 3518 3437
rect 3552 3403 3562 3437
rect 3308 3263 3318 3297
rect 3352 3263 3362 3297
rect 3108 3123 3118 3157
rect 3152 3123 3162 3157
rect 2908 2983 2918 3017
rect 2952 2983 2962 3017
rect 2708 2843 2718 2877
rect 2752 2843 2762 2877
rect 2508 2703 2518 2737
rect 2552 2703 2562 2737
rect 2308 2563 2318 2597
rect 2352 2563 2362 2597
rect 2202 2499 2268 2500
rect 2202 2447 2209 2499
rect 2261 2447 2268 2499
rect 2202 2446 2268 2447
rect 2108 2333 2118 2367
rect 2152 2333 2162 2367
rect 1908 2193 1918 2227
rect 1952 2193 1962 2227
rect 1708 2053 1718 2087
rect 1752 2053 1762 2087
rect 1508 1913 1518 1947
rect 1552 1913 1562 1947
rect 1308 1773 1318 1807
rect 1352 1773 1362 1807
rect 1108 1633 1118 1667
rect 1152 1633 1162 1667
rect 908 1493 918 1527
rect 952 1493 962 1527
rect 708 1353 718 1387
rect 752 1353 762 1387
rect 602 1289 668 1290
rect 602 1237 609 1289
rect 661 1237 668 1289
rect 602 1236 668 1237
rect 508 1123 518 1157
rect 552 1123 562 1157
rect 308 983 318 1017
rect 352 983 362 1017
rect 108 843 118 877
rect 152 843 162 877
rect 8 737 62 749
rect 8 711 18 737
rect 52 711 62 737
rect 8 659 9 711
rect 61 659 62 711
rect 8 652 62 659
rect 108 737 162 843
rect 208 921 262 928
rect 208 869 209 921
rect 261 869 262 921
rect 208 843 218 869
rect 252 843 262 869
rect 208 831 262 843
rect 308 877 362 983
rect 408 1017 462 1029
rect 408 991 418 1017
rect 452 991 462 1017
rect 408 939 409 991
rect 461 939 462 991
rect 408 932 462 939
rect 508 1017 562 1123
rect 608 1201 662 1208
rect 608 1149 609 1201
rect 661 1149 662 1201
rect 608 1123 618 1149
rect 652 1123 662 1149
rect 608 1111 662 1123
rect 708 1157 762 1353
rect 808 1387 862 1399
rect 808 1361 818 1387
rect 852 1361 862 1387
rect 808 1309 809 1361
rect 861 1309 862 1361
rect 808 1302 862 1309
rect 908 1387 962 1493
rect 1008 1571 1062 1578
rect 1008 1519 1009 1571
rect 1061 1519 1062 1571
rect 1008 1493 1018 1519
rect 1052 1493 1062 1519
rect 1008 1481 1062 1493
rect 1108 1527 1162 1633
rect 1208 1667 1262 1679
rect 1208 1641 1218 1667
rect 1252 1641 1262 1667
rect 1208 1589 1209 1641
rect 1261 1589 1262 1641
rect 1208 1582 1262 1589
rect 1308 1667 1362 1773
rect 1408 1851 1462 1858
rect 1408 1799 1409 1851
rect 1461 1799 1462 1851
rect 1408 1773 1418 1799
rect 1452 1773 1462 1799
rect 1408 1761 1462 1773
rect 1508 1807 1562 1913
rect 1608 1947 1662 1959
rect 1608 1921 1618 1947
rect 1652 1921 1662 1947
rect 1608 1869 1609 1921
rect 1661 1869 1662 1921
rect 1608 1862 1662 1869
rect 1708 1947 1762 2053
rect 1808 2131 1862 2138
rect 1808 2079 1809 2131
rect 1861 2079 1862 2131
rect 1808 2053 1818 2079
rect 1852 2053 1862 2079
rect 1808 2041 1862 2053
rect 1908 2087 1962 2193
rect 2008 2227 2062 2239
rect 2008 2201 2018 2227
rect 2052 2201 2062 2227
rect 2008 2149 2009 2201
rect 2061 2149 2062 2201
rect 2008 2142 2062 2149
rect 2108 2227 2162 2333
rect 2208 2411 2262 2418
rect 2208 2359 2209 2411
rect 2261 2359 2262 2411
rect 2208 2333 2218 2359
rect 2252 2333 2262 2359
rect 2208 2321 2262 2333
rect 2308 2367 2362 2563
rect 2408 2597 2462 2609
rect 2408 2571 2418 2597
rect 2452 2571 2462 2597
rect 2408 2519 2409 2571
rect 2461 2519 2462 2571
rect 2408 2512 2462 2519
rect 2508 2597 2562 2703
rect 2608 2781 2662 2788
rect 2608 2729 2609 2781
rect 2661 2729 2662 2781
rect 2608 2703 2618 2729
rect 2652 2703 2662 2729
rect 2608 2691 2662 2703
rect 2708 2737 2762 2843
rect 2808 2877 2862 2889
rect 2808 2851 2818 2877
rect 2852 2851 2862 2877
rect 2808 2799 2809 2851
rect 2861 2799 2862 2851
rect 2808 2792 2862 2799
rect 2908 2877 2962 2983
rect 3008 3061 3062 3068
rect 3008 3009 3009 3061
rect 3061 3009 3062 3061
rect 3008 2983 3018 3009
rect 3052 2983 3062 3009
rect 3008 2971 3062 2983
rect 3108 3017 3162 3123
rect 3208 3157 3262 3169
rect 3208 3131 3218 3157
rect 3252 3131 3262 3157
rect 3208 3079 3209 3131
rect 3261 3079 3262 3131
rect 3208 3072 3262 3079
rect 3308 3157 3362 3263
rect 3408 3341 3462 3348
rect 3408 3289 3409 3341
rect 3461 3289 3462 3341
rect 3408 3263 3418 3289
rect 3452 3263 3462 3289
rect 3408 3251 3462 3263
rect 3508 3297 3562 3403
rect 3608 3437 3662 3449
rect 3608 3411 3618 3437
rect 3652 3411 3662 3437
rect 3608 3359 3609 3411
rect 3661 3359 3662 3411
rect 3608 3352 3662 3359
rect 3708 3437 3762 3543
rect 3808 3621 3862 3628
rect 3808 3569 3809 3621
rect 3861 3569 3862 3621
rect 3808 3543 3818 3569
rect 3852 3543 3862 3569
rect 3808 3531 3862 3543
rect 3908 3577 3962 3773
rect 4008 3807 4062 3819
rect 4008 3781 4018 3807
rect 4052 3781 4062 3807
rect 4008 3729 4009 3781
rect 4061 3729 4062 3781
rect 4008 3722 4062 3729
rect 4108 3807 4162 3913
rect 4208 3991 4262 3998
rect 4208 3939 4209 3991
rect 4261 3939 4262 3991
rect 4208 3913 4218 3939
rect 4252 3913 4262 3939
rect 4208 3901 4262 3913
rect 4308 3947 4362 4053
rect 4408 4087 4462 4099
rect 4408 4061 4418 4087
rect 4452 4061 4462 4087
rect 4408 4009 4409 4061
rect 4461 4009 4462 4061
rect 4408 4002 4462 4009
rect 4508 4087 4562 4193
rect 4608 4271 4662 4278
rect 4608 4219 4609 4271
rect 4661 4219 4662 4271
rect 4608 4193 4618 4219
rect 4652 4193 4662 4219
rect 4608 4181 4662 4193
rect 4708 4227 4762 4333
rect 4808 4367 4862 4379
rect 4808 4341 4818 4367
rect 4852 4341 4862 4367
rect 4808 4289 4809 4341
rect 4861 4289 4862 4341
rect 4808 4282 4862 4289
rect 4908 4367 4962 4473
rect 5008 4551 5062 4558
rect 5008 4499 5009 4551
rect 5061 4499 5062 4551
rect 5008 4473 5018 4499
rect 5052 4473 5062 4499
rect 5008 4461 5062 4473
rect 5108 4507 5162 4613
rect 5208 4647 5262 4659
rect 5208 4621 5218 4647
rect 5252 4621 5262 4647
rect 5208 4569 5209 4621
rect 5261 4569 5262 4621
rect 5208 4562 5262 4569
rect 5308 4647 5362 4753
rect 5408 4831 5462 4838
rect 5408 4779 5409 4831
rect 5461 4779 5462 4831
rect 5408 4753 5418 4779
rect 5452 4753 5462 4779
rect 5408 4741 5462 4753
rect 5508 4787 5562 4960
rect 5602 4903 5668 4904
rect 5602 4851 5609 4903
rect 5661 4851 5668 4903
rect 5602 4850 5668 4851
rect 5508 4753 5518 4787
rect 5552 4753 5562 4787
rect 5308 4613 5318 4647
rect 5352 4613 5362 4647
rect 5108 4473 5118 4507
rect 5152 4473 5162 4507
rect 4908 4333 4918 4367
rect 4952 4333 4962 4367
rect 4708 4193 4718 4227
rect 4752 4193 4762 4227
rect 4508 4053 4518 4087
rect 4552 4053 4562 4087
rect 4308 3913 4318 3947
rect 4352 3913 4362 3947
rect 4108 3773 4118 3807
rect 4152 3773 4162 3807
rect 4002 3693 4068 3694
rect 4002 3641 4009 3693
rect 4061 3641 4068 3693
rect 4002 3640 4068 3641
rect 3908 3543 3918 3577
rect 3952 3543 3962 3577
rect 3708 3403 3718 3437
rect 3752 3403 3762 3437
rect 3508 3263 3518 3297
rect 3552 3263 3562 3297
rect 3308 3123 3318 3157
rect 3352 3123 3362 3157
rect 3108 2983 3118 3017
rect 3152 2983 3162 3017
rect 2908 2843 2918 2877
rect 2952 2843 2962 2877
rect 2708 2703 2718 2737
rect 2752 2703 2762 2737
rect 2508 2563 2518 2597
rect 2552 2563 2562 2597
rect 2402 2483 2468 2484
rect 2402 2431 2409 2483
rect 2461 2431 2468 2483
rect 2402 2430 2468 2431
rect 2308 2333 2318 2367
rect 2352 2333 2362 2367
rect 2108 2193 2118 2227
rect 2152 2193 2162 2227
rect 1908 2053 1918 2087
rect 1952 2053 1962 2087
rect 1708 1913 1718 1947
rect 1752 1913 1762 1947
rect 1508 1773 1518 1807
rect 1552 1773 1562 1807
rect 1308 1633 1318 1667
rect 1352 1633 1362 1667
rect 1108 1493 1118 1527
rect 1152 1493 1162 1527
rect 908 1353 918 1387
rect 952 1353 962 1387
rect 802 1273 868 1274
rect 802 1221 809 1273
rect 861 1221 868 1273
rect 802 1220 868 1221
rect 708 1123 718 1157
rect 752 1123 762 1157
rect 508 983 518 1017
rect 552 983 562 1017
rect 308 843 318 877
rect 352 843 362 877
rect 108 703 118 737
rect 152 703 162 737
rect 8 597 62 609
rect 8 571 18 597
rect 52 571 62 597
rect 8 519 9 571
rect 61 519 62 571
rect 8 512 62 519
rect 108 597 162 703
rect 208 781 262 788
rect 208 729 209 781
rect 261 729 262 781
rect 208 703 218 729
rect 252 703 262 729
rect 208 691 262 703
rect 308 737 362 843
rect 408 877 462 889
rect 408 851 418 877
rect 452 851 462 877
rect 408 799 409 851
rect 461 799 462 851
rect 408 792 462 799
rect 508 877 562 983
rect 608 1061 662 1068
rect 608 1009 609 1061
rect 661 1009 662 1061
rect 608 983 618 1009
rect 652 983 662 1009
rect 608 971 662 983
rect 708 1017 762 1123
rect 808 1157 862 1169
rect 808 1131 818 1157
rect 852 1131 862 1157
rect 808 1079 809 1131
rect 861 1079 862 1131
rect 808 1072 862 1079
rect 908 1157 962 1353
rect 1008 1431 1062 1438
rect 1008 1379 1009 1431
rect 1061 1379 1062 1431
rect 1008 1353 1018 1379
rect 1052 1353 1062 1379
rect 1008 1341 1062 1353
rect 1108 1387 1162 1493
rect 1208 1527 1262 1539
rect 1208 1501 1218 1527
rect 1252 1501 1262 1527
rect 1208 1449 1209 1501
rect 1261 1449 1262 1501
rect 1208 1442 1262 1449
rect 1308 1527 1362 1633
rect 1408 1711 1462 1718
rect 1408 1659 1409 1711
rect 1461 1659 1462 1711
rect 1408 1633 1418 1659
rect 1452 1633 1462 1659
rect 1408 1621 1462 1633
rect 1508 1667 1562 1773
rect 1608 1807 1662 1819
rect 1608 1781 1618 1807
rect 1652 1781 1662 1807
rect 1608 1729 1609 1781
rect 1661 1729 1662 1781
rect 1608 1722 1662 1729
rect 1708 1807 1762 1913
rect 1808 1991 1862 1998
rect 1808 1939 1809 1991
rect 1861 1939 1862 1991
rect 1808 1913 1818 1939
rect 1852 1913 1862 1939
rect 1808 1901 1862 1913
rect 1908 1947 1962 2053
rect 2008 2087 2062 2099
rect 2008 2061 2018 2087
rect 2052 2061 2062 2087
rect 2008 2009 2009 2061
rect 2061 2009 2062 2061
rect 2008 2002 2062 2009
rect 2108 2087 2162 2193
rect 2208 2271 2262 2278
rect 2208 2219 2209 2271
rect 2261 2219 2262 2271
rect 2208 2193 2218 2219
rect 2252 2193 2262 2219
rect 2208 2181 2262 2193
rect 2308 2227 2362 2333
rect 2408 2367 2462 2379
rect 2408 2341 2418 2367
rect 2452 2341 2462 2367
rect 2408 2289 2409 2341
rect 2461 2289 2462 2341
rect 2408 2282 2462 2289
rect 2508 2367 2562 2563
rect 2608 2641 2662 2648
rect 2608 2589 2609 2641
rect 2661 2589 2662 2641
rect 2608 2563 2618 2589
rect 2652 2563 2662 2589
rect 2608 2551 2662 2563
rect 2708 2597 2762 2703
rect 2808 2737 2862 2749
rect 2808 2711 2818 2737
rect 2852 2711 2862 2737
rect 2808 2659 2809 2711
rect 2861 2659 2862 2711
rect 2808 2652 2862 2659
rect 2908 2737 2962 2843
rect 3008 2921 3062 2928
rect 3008 2869 3009 2921
rect 3061 2869 3062 2921
rect 3008 2843 3018 2869
rect 3052 2843 3062 2869
rect 3008 2831 3062 2843
rect 3108 2877 3162 2983
rect 3208 3017 3262 3029
rect 3208 2991 3218 3017
rect 3252 2991 3262 3017
rect 3208 2939 3209 2991
rect 3261 2939 3262 2991
rect 3208 2932 3262 2939
rect 3308 3017 3362 3123
rect 3408 3201 3462 3208
rect 3408 3149 3409 3201
rect 3461 3149 3462 3201
rect 3408 3123 3418 3149
rect 3452 3123 3462 3149
rect 3408 3111 3462 3123
rect 3508 3157 3562 3263
rect 3608 3297 3662 3309
rect 3608 3271 3618 3297
rect 3652 3271 3662 3297
rect 3608 3219 3609 3271
rect 3661 3219 3662 3271
rect 3608 3212 3662 3219
rect 3708 3297 3762 3403
rect 3808 3481 3862 3488
rect 3808 3429 3809 3481
rect 3861 3429 3862 3481
rect 3808 3403 3818 3429
rect 3852 3403 3862 3429
rect 3808 3391 3862 3403
rect 3908 3437 3962 3543
rect 4008 3577 4062 3589
rect 4008 3551 4018 3577
rect 4052 3551 4062 3577
rect 4008 3499 4009 3551
rect 4061 3499 4062 3551
rect 4008 3492 4062 3499
rect 4108 3577 4162 3773
rect 4208 3851 4262 3858
rect 4208 3799 4209 3851
rect 4261 3799 4262 3851
rect 4208 3773 4218 3799
rect 4252 3773 4262 3799
rect 4208 3761 4262 3773
rect 4308 3807 4362 3913
rect 4408 3947 4462 3959
rect 4408 3921 4418 3947
rect 4452 3921 4462 3947
rect 4408 3869 4409 3921
rect 4461 3869 4462 3921
rect 4408 3862 4462 3869
rect 4508 3947 4562 4053
rect 4608 4131 4662 4138
rect 4608 4079 4609 4131
rect 4661 4079 4662 4131
rect 4608 4053 4618 4079
rect 4652 4053 4662 4079
rect 4608 4041 4662 4053
rect 4708 4087 4762 4193
rect 4808 4227 4862 4239
rect 4808 4201 4818 4227
rect 4852 4201 4862 4227
rect 4808 4149 4809 4201
rect 4861 4149 4862 4201
rect 4808 4142 4862 4149
rect 4908 4227 4962 4333
rect 5008 4411 5062 4418
rect 5008 4359 5009 4411
rect 5061 4359 5062 4411
rect 5008 4333 5018 4359
rect 5052 4333 5062 4359
rect 5008 4321 5062 4333
rect 5108 4367 5162 4473
rect 5208 4507 5262 4519
rect 5208 4481 5218 4507
rect 5252 4481 5262 4507
rect 5208 4429 5209 4481
rect 5261 4429 5262 4481
rect 5208 4422 5262 4429
rect 5308 4507 5362 4613
rect 5408 4691 5462 4698
rect 5408 4639 5409 4691
rect 5461 4639 5462 4691
rect 5408 4613 5418 4639
rect 5452 4613 5462 4639
rect 5408 4601 5462 4613
rect 5508 4647 5562 4753
rect 5608 4787 5662 4799
rect 5608 4761 5618 4787
rect 5652 4761 5662 4787
rect 5608 4709 5609 4761
rect 5661 4709 5662 4761
rect 5608 4702 5662 4709
rect 5708 4787 5762 4960
rect 5802 4919 5868 4920
rect 5802 4867 5809 4919
rect 5861 4867 5868 4919
rect 5802 4866 5868 4867
rect 5708 4753 5718 4787
rect 5752 4753 5762 4787
rect 5508 4613 5518 4647
rect 5552 4613 5562 4647
rect 5308 4473 5318 4507
rect 5352 4473 5362 4507
rect 5108 4333 5118 4367
rect 5152 4333 5162 4367
rect 4908 4193 4918 4227
rect 4952 4193 4962 4227
rect 4708 4053 4718 4087
rect 4752 4053 4762 4087
rect 4508 3913 4518 3947
rect 4552 3913 4562 3947
rect 4308 3773 4318 3807
rect 4352 3773 4362 3807
rect 4202 3709 4268 3710
rect 4202 3657 4209 3709
rect 4261 3657 4268 3709
rect 4202 3656 4268 3657
rect 4108 3543 4118 3577
rect 4152 3543 4162 3577
rect 3908 3403 3918 3437
rect 3952 3403 3962 3437
rect 3708 3263 3718 3297
rect 3752 3263 3762 3297
rect 3508 3123 3518 3157
rect 3552 3123 3562 3157
rect 3308 2983 3318 3017
rect 3352 2983 3362 3017
rect 3108 2843 3118 2877
rect 3152 2843 3162 2877
rect 2908 2703 2918 2737
rect 2952 2703 2962 2737
rect 2708 2563 2718 2597
rect 2752 2563 2762 2597
rect 2602 2499 2668 2500
rect 2602 2447 2609 2499
rect 2661 2447 2668 2499
rect 2602 2446 2668 2447
rect 2508 2333 2518 2367
rect 2552 2333 2562 2367
rect 2308 2193 2318 2227
rect 2352 2193 2362 2227
rect 2108 2053 2118 2087
rect 2152 2053 2162 2087
rect 1908 1913 1918 1947
rect 1952 1913 1962 1947
rect 1708 1773 1718 1807
rect 1752 1773 1762 1807
rect 1508 1633 1518 1667
rect 1552 1633 1562 1667
rect 1308 1493 1318 1527
rect 1352 1493 1362 1527
rect 1108 1353 1118 1387
rect 1152 1353 1162 1387
rect 1002 1289 1068 1290
rect 1002 1237 1009 1289
rect 1061 1237 1068 1289
rect 1002 1236 1068 1237
rect 908 1123 918 1157
rect 952 1123 962 1157
rect 708 983 718 1017
rect 752 983 762 1017
rect 508 843 518 877
rect 552 843 562 877
rect 308 703 318 737
rect 352 703 362 737
rect 108 563 118 597
rect 152 563 162 597
rect 8 457 62 469
rect 8 431 18 457
rect 52 431 62 457
rect 8 379 9 431
rect 61 379 62 431
rect 8 372 62 379
rect 108 457 162 563
rect 208 641 262 648
rect 208 589 209 641
rect 261 589 262 641
rect 208 563 218 589
rect 252 563 262 589
rect 208 551 262 563
rect 308 597 362 703
rect 408 737 462 749
rect 408 711 418 737
rect 452 711 462 737
rect 408 659 409 711
rect 461 659 462 711
rect 408 652 462 659
rect 508 737 562 843
rect 608 921 662 928
rect 608 869 609 921
rect 661 869 662 921
rect 608 843 618 869
rect 652 843 662 869
rect 608 831 662 843
rect 708 877 762 983
rect 808 1017 862 1029
rect 808 991 818 1017
rect 852 991 862 1017
rect 808 939 809 991
rect 861 939 862 991
rect 808 932 862 939
rect 908 1017 962 1123
rect 1008 1201 1062 1208
rect 1008 1149 1009 1201
rect 1061 1149 1062 1201
rect 1008 1123 1018 1149
rect 1052 1123 1062 1149
rect 1008 1111 1062 1123
rect 1108 1157 1162 1353
rect 1208 1387 1262 1399
rect 1208 1361 1218 1387
rect 1252 1361 1262 1387
rect 1208 1309 1209 1361
rect 1261 1309 1262 1361
rect 1208 1302 1262 1309
rect 1308 1387 1362 1493
rect 1408 1571 1462 1578
rect 1408 1519 1409 1571
rect 1461 1519 1462 1571
rect 1408 1493 1418 1519
rect 1452 1493 1462 1519
rect 1408 1481 1462 1493
rect 1508 1527 1562 1633
rect 1608 1667 1662 1679
rect 1608 1641 1618 1667
rect 1652 1641 1662 1667
rect 1608 1589 1609 1641
rect 1661 1589 1662 1641
rect 1608 1582 1662 1589
rect 1708 1667 1762 1773
rect 1808 1851 1862 1858
rect 1808 1799 1809 1851
rect 1861 1799 1862 1851
rect 1808 1773 1818 1799
rect 1852 1773 1862 1799
rect 1808 1761 1862 1773
rect 1908 1807 1962 1913
rect 2008 1947 2062 1959
rect 2008 1921 2018 1947
rect 2052 1921 2062 1947
rect 2008 1869 2009 1921
rect 2061 1869 2062 1921
rect 2008 1862 2062 1869
rect 2108 1947 2162 2053
rect 2208 2131 2262 2138
rect 2208 2079 2209 2131
rect 2261 2079 2262 2131
rect 2208 2053 2218 2079
rect 2252 2053 2262 2079
rect 2208 2041 2262 2053
rect 2308 2087 2362 2193
rect 2408 2227 2462 2239
rect 2408 2201 2418 2227
rect 2452 2201 2462 2227
rect 2408 2149 2409 2201
rect 2461 2149 2462 2201
rect 2408 2142 2462 2149
rect 2508 2227 2562 2333
rect 2608 2411 2662 2418
rect 2608 2359 2609 2411
rect 2661 2359 2662 2411
rect 2608 2333 2618 2359
rect 2652 2333 2662 2359
rect 2608 2321 2662 2333
rect 2708 2367 2762 2563
rect 2808 2597 2862 2609
rect 2808 2571 2818 2597
rect 2852 2571 2862 2597
rect 2808 2519 2809 2571
rect 2861 2519 2862 2571
rect 2808 2512 2862 2519
rect 2908 2597 2962 2703
rect 3008 2781 3062 2788
rect 3008 2729 3009 2781
rect 3061 2729 3062 2781
rect 3008 2703 3018 2729
rect 3052 2703 3062 2729
rect 3008 2691 3062 2703
rect 3108 2737 3162 2843
rect 3208 2877 3262 2889
rect 3208 2851 3218 2877
rect 3252 2851 3262 2877
rect 3208 2799 3209 2851
rect 3261 2799 3262 2851
rect 3208 2792 3262 2799
rect 3308 2877 3362 2983
rect 3408 3061 3462 3068
rect 3408 3009 3409 3061
rect 3461 3009 3462 3061
rect 3408 2983 3418 3009
rect 3452 2983 3462 3009
rect 3408 2971 3462 2983
rect 3508 3017 3562 3123
rect 3608 3157 3662 3169
rect 3608 3131 3618 3157
rect 3652 3131 3662 3157
rect 3608 3079 3609 3131
rect 3661 3079 3662 3131
rect 3608 3072 3662 3079
rect 3708 3157 3762 3263
rect 3808 3341 3862 3348
rect 3808 3289 3809 3341
rect 3861 3289 3862 3341
rect 3808 3263 3818 3289
rect 3852 3263 3862 3289
rect 3808 3251 3862 3263
rect 3908 3297 3962 3403
rect 4008 3437 4062 3449
rect 4008 3411 4018 3437
rect 4052 3411 4062 3437
rect 4008 3359 4009 3411
rect 4061 3359 4062 3411
rect 4008 3352 4062 3359
rect 4108 3437 4162 3543
rect 4208 3621 4262 3628
rect 4208 3569 4209 3621
rect 4261 3569 4262 3621
rect 4208 3543 4218 3569
rect 4252 3543 4262 3569
rect 4208 3531 4262 3543
rect 4308 3577 4362 3773
rect 4408 3807 4462 3819
rect 4408 3781 4418 3807
rect 4452 3781 4462 3807
rect 4408 3729 4409 3781
rect 4461 3729 4462 3781
rect 4408 3722 4462 3729
rect 4508 3807 4562 3913
rect 4608 3991 4662 3998
rect 4608 3939 4609 3991
rect 4661 3939 4662 3991
rect 4608 3913 4618 3939
rect 4652 3913 4662 3939
rect 4608 3901 4662 3913
rect 4708 3947 4762 4053
rect 4808 4087 4862 4099
rect 4808 4061 4818 4087
rect 4852 4061 4862 4087
rect 4808 4009 4809 4061
rect 4861 4009 4862 4061
rect 4808 4002 4862 4009
rect 4908 4087 4962 4193
rect 5008 4271 5062 4278
rect 5008 4219 5009 4271
rect 5061 4219 5062 4271
rect 5008 4193 5018 4219
rect 5052 4193 5062 4219
rect 5008 4181 5062 4193
rect 5108 4227 5162 4333
rect 5208 4367 5262 4379
rect 5208 4341 5218 4367
rect 5252 4341 5262 4367
rect 5208 4289 5209 4341
rect 5261 4289 5262 4341
rect 5208 4282 5262 4289
rect 5308 4367 5362 4473
rect 5408 4551 5462 4558
rect 5408 4499 5409 4551
rect 5461 4499 5462 4551
rect 5408 4473 5418 4499
rect 5452 4473 5462 4499
rect 5408 4461 5462 4473
rect 5508 4507 5562 4613
rect 5608 4647 5662 4659
rect 5608 4621 5618 4647
rect 5652 4621 5662 4647
rect 5608 4569 5609 4621
rect 5661 4569 5662 4621
rect 5608 4562 5662 4569
rect 5708 4647 5762 4753
rect 5808 4831 5862 4838
rect 5808 4779 5809 4831
rect 5861 4779 5862 4831
rect 5808 4753 5818 4779
rect 5852 4753 5862 4779
rect 5808 4741 5862 4753
rect 5908 4787 5962 4960
rect 6002 4903 6068 4904
rect 6002 4851 6009 4903
rect 6061 4851 6068 4903
rect 6002 4850 6068 4851
rect 5908 4753 5918 4787
rect 5952 4753 5962 4787
rect 5708 4613 5718 4647
rect 5752 4613 5762 4647
rect 5508 4473 5518 4507
rect 5552 4473 5562 4507
rect 5308 4333 5318 4367
rect 5352 4333 5362 4367
rect 5108 4193 5118 4227
rect 5152 4193 5162 4227
rect 4908 4053 4918 4087
rect 4952 4053 4962 4087
rect 4708 3913 4718 3947
rect 4752 3913 4762 3947
rect 4508 3773 4518 3807
rect 4552 3773 4562 3807
rect 4402 3693 4468 3694
rect 4402 3641 4409 3693
rect 4461 3641 4468 3693
rect 4402 3640 4468 3641
rect 4308 3543 4318 3577
rect 4352 3543 4362 3577
rect 4108 3403 4118 3437
rect 4152 3403 4162 3437
rect 3908 3263 3918 3297
rect 3952 3263 3962 3297
rect 3708 3123 3718 3157
rect 3752 3123 3762 3157
rect 3508 2983 3518 3017
rect 3552 2983 3562 3017
rect 3308 2843 3318 2877
rect 3352 2843 3362 2877
rect 3108 2703 3118 2737
rect 3152 2703 3162 2737
rect 2908 2563 2918 2597
rect 2952 2563 2962 2597
rect 2802 2483 2868 2484
rect 2802 2431 2809 2483
rect 2861 2431 2868 2483
rect 2802 2430 2868 2431
rect 2708 2333 2718 2367
rect 2752 2333 2762 2367
rect 2508 2193 2518 2227
rect 2552 2193 2562 2227
rect 2308 2053 2318 2087
rect 2352 2053 2362 2087
rect 2108 1913 2118 1947
rect 2152 1913 2162 1947
rect 1908 1773 1918 1807
rect 1952 1773 1962 1807
rect 1708 1633 1718 1667
rect 1752 1633 1762 1667
rect 1508 1493 1518 1527
rect 1552 1493 1562 1527
rect 1308 1353 1318 1387
rect 1352 1353 1362 1387
rect 1202 1273 1268 1274
rect 1202 1221 1209 1273
rect 1261 1221 1268 1273
rect 1202 1220 1268 1221
rect 1108 1123 1118 1157
rect 1152 1123 1162 1157
rect 908 983 918 1017
rect 952 983 962 1017
rect 708 843 718 877
rect 752 843 762 877
rect 508 703 518 737
rect 552 703 562 737
rect 308 563 318 597
rect 352 563 362 597
rect 108 423 118 457
rect 152 423 162 457
rect 8 317 62 329
rect 8 291 18 317
rect 52 291 62 317
rect 8 239 9 291
rect 61 239 62 291
rect 8 232 62 239
rect 108 317 162 423
rect 208 501 262 508
rect 208 449 209 501
rect 261 449 262 501
rect 208 423 218 449
rect 252 423 262 449
rect 208 411 262 423
rect 308 457 362 563
rect 408 597 462 609
rect 408 571 418 597
rect 452 571 462 597
rect 408 519 409 571
rect 461 519 462 571
rect 408 512 462 519
rect 508 597 562 703
rect 608 781 662 788
rect 608 729 609 781
rect 661 729 662 781
rect 608 703 618 729
rect 652 703 662 729
rect 608 691 662 703
rect 708 737 762 843
rect 808 877 862 889
rect 808 851 818 877
rect 852 851 862 877
rect 808 799 809 851
rect 861 799 862 851
rect 808 792 862 799
rect 908 877 962 983
rect 1008 1061 1062 1068
rect 1008 1009 1009 1061
rect 1061 1009 1062 1061
rect 1008 983 1018 1009
rect 1052 983 1062 1009
rect 1008 971 1062 983
rect 1108 1017 1162 1123
rect 1208 1157 1262 1169
rect 1208 1131 1218 1157
rect 1252 1131 1262 1157
rect 1208 1079 1209 1131
rect 1261 1079 1262 1131
rect 1208 1072 1262 1079
rect 1308 1157 1362 1353
rect 1408 1431 1462 1438
rect 1408 1379 1409 1431
rect 1461 1379 1462 1431
rect 1408 1353 1418 1379
rect 1452 1353 1462 1379
rect 1408 1341 1462 1353
rect 1508 1387 1562 1493
rect 1608 1527 1662 1539
rect 1608 1501 1618 1527
rect 1652 1501 1662 1527
rect 1608 1449 1609 1501
rect 1661 1449 1662 1501
rect 1608 1442 1662 1449
rect 1708 1527 1762 1633
rect 1808 1711 1862 1718
rect 1808 1659 1809 1711
rect 1861 1659 1862 1711
rect 1808 1633 1818 1659
rect 1852 1633 1862 1659
rect 1808 1621 1862 1633
rect 1908 1667 1962 1773
rect 2008 1807 2062 1819
rect 2008 1781 2018 1807
rect 2052 1781 2062 1807
rect 2008 1729 2009 1781
rect 2061 1729 2062 1781
rect 2008 1722 2062 1729
rect 2108 1807 2162 1913
rect 2208 1991 2262 1998
rect 2208 1939 2209 1991
rect 2261 1939 2262 1991
rect 2208 1913 2218 1939
rect 2252 1913 2262 1939
rect 2208 1901 2262 1913
rect 2308 1947 2362 2053
rect 2408 2087 2462 2099
rect 2408 2061 2418 2087
rect 2452 2061 2462 2087
rect 2408 2009 2409 2061
rect 2461 2009 2462 2061
rect 2408 2002 2462 2009
rect 2508 2087 2562 2193
rect 2608 2271 2662 2278
rect 2608 2219 2609 2271
rect 2661 2219 2662 2271
rect 2608 2193 2618 2219
rect 2652 2193 2662 2219
rect 2608 2181 2662 2193
rect 2708 2227 2762 2333
rect 2808 2367 2862 2379
rect 2808 2341 2818 2367
rect 2852 2341 2862 2367
rect 2808 2289 2809 2341
rect 2861 2289 2862 2341
rect 2808 2282 2862 2289
rect 2908 2367 2962 2563
rect 3008 2641 3062 2648
rect 3008 2589 3009 2641
rect 3061 2589 3062 2641
rect 3008 2563 3018 2589
rect 3052 2563 3062 2589
rect 3008 2551 3062 2563
rect 3108 2597 3162 2703
rect 3208 2737 3262 2749
rect 3208 2711 3218 2737
rect 3252 2711 3262 2737
rect 3208 2659 3209 2711
rect 3261 2659 3262 2711
rect 3208 2652 3262 2659
rect 3308 2737 3362 2843
rect 3408 2921 3462 2928
rect 3408 2869 3409 2921
rect 3461 2869 3462 2921
rect 3408 2843 3418 2869
rect 3452 2843 3462 2869
rect 3408 2831 3462 2843
rect 3508 2877 3562 2983
rect 3608 3017 3662 3029
rect 3608 2991 3618 3017
rect 3652 2991 3662 3017
rect 3608 2939 3609 2991
rect 3661 2939 3662 2991
rect 3608 2932 3662 2939
rect 3708 3017 3762 3123
rect 3808 3201 3862 3208
rect 3808 3149 3809 3201
rect 3861 3149 3862 3201
rect 3808 3123 3818 3149
rect 3852 3123 3862 3149
rect 3808 3111 3862 3123
rect 3908 3157 3962 3263
rect 4008 3297 4062 3309
rect 4008 3271 4018 3297
rect 4052 3271 4062 3297
rect 4008 3219 4009 3271
rect 4061 3219 4062 3271
rect 4008 3212 4062 3219
rect 4108 3297 4162 3403
rect 4208 3481 4262 3488
rect 4208 3429 4209 3481
rect 4261 3429 4262 3481
rect 4208 3403 4218 3429
rect 4252 3403 4262 3429
rect 4208 3391 4262 3403
rect 4308 3437 4362 3543
rect 4408 3577 4462 3589
rect 4408 3551 4418 3577
rect 4452 3551 4462 3577
rect 4408 3499 4409 3551
rect 4461 3499 4462 3551
rect 4408 3492 4462 3499
rect 4508 3577 4562 3773
rect 4608 3851 4662 3858
rect 4608 3799 4609 3851
rect 4661 3799 4662 3851
rect 4608 3773 4618 3799
rect 4652 3773 4662 3799
rect 4608 3761 4662 3773
rect 4708 3807 4762 3913
rect 4808 3947 4862 3959
rect 4808 3921 4818 3947
rect 4852 3921 4862 3947
rect 4808 3869 4809 3921
rect 4861 3869 4862 3921
rect 4808 3862 4862 3869
rect 4908 3947 4962 4053
rect 5008 4131 5062 4138
rect 5008 4079 5009 4131
rect 5061 4079 5062 4131
rect 5008 4053 5018 4079
rect 5052 4053 5062 4079
rect 5008 4041 5062 4053
rect 5108 4087 5162 4193
rect 5208 4227 5262 4239
rect 5208 4201 5218 4227
rect 5252 4201 5262 4227
rect 5208 4149 5209 4201
rect 5261 4149 5262 4201
rect 5208 4142 5262 4149
rect 5308 4227 5362 4333
rect 5408 4411 5462 4418
rect 5408 4359 5409 4411
rect 5461 4359 5462 4411
rect 5408 4333 5418 4359
rect 5452 4333 5462 4359
rect 5408 4321 5462 4333
rect 5508 4367 5562 4473
rect 5608 4507 5662 4519
rect 5608 4481 5618 4507
rect 5652 4481 5662 4507
rect 5608 4429 5609 4481
rect 5661 4429 5662 4481
rect 5608 4422 5662 4429
rect 5708 4507 5762 4613
rect 5808 4691 5862 4698
rect 5808 4639 5809 4691
rect 5861 4639 5862 4691
rect 5808 4613 5818 4639
rect 5852 4613 5862 4639
rect 5808 4601 5862 4613
rect 5908 4647 5962 4753
rect 6008 4787 6062 4799
rect 6008 4761 6018 4787
rect 6052 4761 6062 4787
rect 6008 4709 6009 4761
rect 6061 4709 6062 4761
rect 6008 4702 6062 4709
rect 6108 4787 6162 4960
rect 6202 4919 6268 4920
rect 6202 4867 6209 4919
rect 6261 4867 6268 4919
rect 6202 4866 6268 4867
rect 6108 4753 6118 4787
rect 6152 4753 6162 4787
rect 5908 4613 5918 4647
rect 5952 4613 5962 4647
rect 5708 4473 5718 4507
rect 5752 4473 5762 4507
rect 5508 4333 5518 4367
rect 5552 4333 5562 4367
rect 5308 4193 5318 4227
rect 5352 4193 5362 4227
rect 5108 4053 5118 4087
rect 5152 4053 5162 4087
rect 4908 3913 4918 3947
rect 4952 3913 4962 3947
rect 4708 3773 4718 3807
rect 4752 3773 4762 3807
rect 4602 3709 4668 3710
rect 4602 3657 4609 3709
rect 4661 3657 4668 3709
rect 4602 3656 4668 3657
rect 4508 3543 4518 3577
rect 4552 3543 4562 3577
rect 4308 3403 4318 3437
rect 4352 3403 4362 3437
rect 4108 3263 4118 3297
rect 4152 3263 4162 3297
rect 3908 3123 3918 3157
rect 3952 3123 3962 3157
rect 3708 2983 3718 3017
rect 3752 2983 3762 3017
rect 3508 2843 3518 2877
rect 3552 2843 3562 2877
rect 3308 2703 3318 2737
rect 3352 2703 3362 2737
rect 3108 2563 3118 2597
rect 3152 2563 3162 2597
rect 3002 2499 3068 2500
rect 3002 2447 3009 2499
rect 3061 2447 3068 2499
rect 3002 2446 3068 2447
rect 2908 2333 2918 2367
rect 2952 2333 2962 2367
rect 2708 2193 2718 2227
rect 2752 2193 2762 2227
rect 2508 2053 2518 2087
rect 2552 2053 2562 2087
rect 2308 1913 2318 1947
rect 2352 1913 2362 1947
rect 2108 1773 2118 1807
rect 2152 1773 2162 1807
rect 1908 1633 1918 1667
rect 1952 1633 1962 1667
rect 1708 1493 1718 1527
rect 1752 1493 1762 1527
rect 1508 1353 1518 1387
rect 1552 1353 1562 1387
rect 1402 1289 1468 1290
rect 1402 1237 1409 1289
rect 1461 1237 1468 1289
rect 1402 1236 1468 1237
rect 1308 1123 1318 1157
rect 1352 1123 1362 1157
rect 1108 983 1118 1017
rect 1152 983 1162 1017
rect 908 843 918 877
rect 952 843 962 877
rect 708 703 718 737
rect 752 703 762 737
rect 508 563 518 597
rect 552 563 562 597
rect 308 423 318 457
rect 352 423 362 457
rect 108 283 118 317
rect 152 283 162 317
rect 8 177 62 189
rect 8 151 18 177
rect 52 151 62 177
rect 8 99 9 151
rect 61 99 62 151
rect 8 92 62 99
rect 108 177 162 283
rect 208 361 262 368
rect 208 309 209 361
rect 261 309 262 361
rect 208 283 218 309
rect 252 283 262 309
rect 208 271 262 283
rect 308 317 362 423
rect 408 457 462 469
rect 408 431 418 457
rect 452 431 462 457
rect 408 379 409 431
rect 461 379 462 431
rect 408 372 462 379
rect 508 457 562 563
rect 608 641 662 648
rect 608 589 609 641
rect 661 589 662 641
rect 608 563 618 589
rect 652 563 662 589
rect 608 551 662 563
rect 708 597 762 703
rect 808 737 862 749
rect 808 711 818 737
rect 852 711 862 737
rect 808 659 809 711
rect 861 659 862 711
rect 808 652 862 659
rect 908 737 962 843
rect 1008 921 1062 928
rect 1008 869 1009 921
rect 1061 869 1062 921
rect 1008 843 1018 869
rect 1052 843 1062 869
rect 1008 831 1062 843
rect 1108 877 1162 983
rect 1208 1017 1262 1029
rect 1208 991 1218 1017
rect 1252 991 1262 1017
rect 1208 939 1209 991
rect 1261 939 1262 991
rect 1208 932 1262 939
rect 1308 1017 1362 1123
rect 1408 1201 1462 1208
rect 1408 1149 1409 1201
rect 1461 1149 1462 1201
rect 1408 1123 1418 1149
rect 1452 1123 1462 1149
rect 1408 1111 1462 1123
rect 1508 1157 1562 1353
rect 1608 1387 1662 1399
rect 1608 1361 1618 1387
rect 1652 1361 1662 1387
rect 1608 1309 1609 1361
rect 1661 1309 1662 1361
rect 1608 1302 1662 1309
rect 1708 1387 1762 1493
rect 1808 1571 1862 1578
rect 1808 1519 1809 1571
rect 1861 1519 1862 1571
rect 1808 1493 1818 1519
rect 1852 1493 1862 1519
rect 1808 1481 1862 1493
rect 1908 1527 1962 1633
rect 2008 1667 2062 1679
rect 2008 1641 2018 1667
rect 2052 1641 2062 1667
rect 2008 1589 2009 1641
rect 2061 1589 2062 1641
rect 2008 1582 2062 1589
rect 2108 1667 2162 1773
rect 2208 1851 2262 1858
rect 2208 1799 2209 1851
rect 2261 1799 2262 1851
rect 2208 1773 2218 1799
rect 2252 1773 2262 1799
rect 2208 1761 2262 1773
rect 2308 1807 2362 1913
rect 2408 1947 2462 1959
rect 2408 1921 2418 1947
rect 2452 1921 2462 1947
rect 2408 1869 2409 1921
rect 2461 1869 2462 1921
rect 2408 1862 2462 1869
rect 2508 1947 2562 2053
rect 2608 2131 2662 2138
rect 2608 2079 2609 2131
rect 2661 2079 2662 2131
rect 2608 2053 2618 2079
rect 2652 2053 2662 2079
rect 2608 2041 2662 2053
rect 2708 2087 2762 2193
rect 2808 2227 2862 2239
rect 2808 2201 2818 2227
rect 2852 2201 2862 2227
rect 2808 2149 2809 2201
rect 2861 2149 2862 2201
rect 2808 2142 2862 2149
rect 2908 2227 2962 2333
rect 3008 2411 3062 2418
rect 3008 2359 3009 2411
rect 3061 2359 3062 2411
rect 3008 2333 3018 2359
rect 3052 2333 3062 2359
rect 3008 2321 3062 2333
rect 3108 2367 3162 2563
rect 3208 2597 3262 2609
rect 3208 2571 3218 2597
rect 3252 2571 3262 2597
rect 3208 2519 3209 2571
rect 3261 2519 3262 2571
rect 3208 2512 3262 2519
rect 3308 2597 3362 2703
rect 3408 2781 3462 2788
rect 3408 2729 3409 2781
rect 3461 2729 3462 2781
rect 3408 2703 3418 2729
rect 3452 2703 3462 2729
rect 3408 2691 3462 2703
rect 3508 2737 3562 2843
rect 3608 2877 3662 2889
rect 3608 2851 3618 2877
rect 3652 2851 3662 2877
rect 3608 2799 3609 2851
rect 3661 2799 3662 2851
rect 3608 2792 3662 2799
rect 3708 2877 3762 2983
rect 3808 3061 3862 3068
rect 3808 3009 3809 3061
rect 3861 3009 3862 3061
rect 3808 2983 3818 3009
rect 3852 2983 3862 3009
rect 3808 2971 3862 2983
rect 3908 3017 3962 3123
rect 4008 3157 4062 3169
rect 4008 3131 4018 3157
rect 4052 3131 4062 3157
rect 4008 3079 4009 3131
rect 4061 3079 4062 3131
rect 4008 3072 4062 3079
rect 4108 3157 4162 3263
rect 4208 3341 4262 3348
rect 4208 3289 4209 3341
rect 4261 3289 4262 3341
rect 4208 3263 4218 3289
rect 4252 3263 4262 3289
rect 4208 3251 4262 3263
rect 4308 3297 4362 3403
rect 4408 3437 4462 3449
rect 4408 3411 4418 3437
rect 4452 3411 4462 3437
rect 4408 3359 4409 3411
rect 4461 3359 4462 3411
rect 4408 3352 4462 3359
rect 4508 3437 4562 3543
rect 4608 3621 4662 3628
rect 4608 3569 4609 3621
rect 4661 3569 4662 3621
rect 4608 3543 4618 3569
rect 4652 3543 4662 3569
rect 4608 3531 4662 3543
rect 4708 3577 4762 3773
rect 4808 3807 4862 3819
rect 4808 3781 4818 3807
rect 4852 3781 4862 3807
rect 4808 3729 4809 3781
rect 4861 3729 4862 3781
rect 4808 3722 4862 3729
rect 4908 3807 4962 3913
rect 5008 3991 5062 3998
rect 5008 3939 5009 3991
rect 5061 3939 5062 3991
rect 5008 3913 5018 3939
rect 5052 3913 5062 3939
rect 5008 3901 5062 3913
rect 5108 3947 5162 4053
rect 5208 4087 5262 4099
rect 5208 4061 5218 4087
rect 5252 4061 5262 4087
rect 5208 4009 5209 4061
rect 5261 4009 5262 4061
rect 5208 4002 5262 4009
rect 5308 4087 5362 4193
rect 5408 4271 5462 4278
rect 5408 4219 5409 4271
rect 5461 4219 5462 4271
rect 5408 4193 5418 4219
rect 5452 4193 5462 4219
rect 5408 4181 5462 4193
rect 5508 4227 5562 4333
rect 5608 4367 5662 4379
rect 5608 4341 5618 4367
rect 5652 4341 5662 4367
rect 5608 4289 5609 4341
rect 5661 4289 5662 4341
rect 5608 4282 5662 4289
rect 5708 4367 5762 4473
rect 5808 4551 5862 4558
rect 5808 4499 5809 4551
rect 5861 4499 5862 4551
rect 5808 4473 5818 4499
rect 5852 4473 5862 4499
rect 5808 4461 5862 4473
rect 5908 4507 5962 4613
rect 6008 4647 6062 4659
rect 6008 4621 6018 4647
rect 6052 4621 6062 4647
rect 6008 4569 6009 4621
rect 6061 4569 6062 4621
rect 6008 4562 6062 4569
rect 6108 4647 6162 4753
rect 6208 4831 6262 4838
rect 6208 4779 6209 4831
rect 6261 4779 6262 4831
rect 6208 4753 6218 4779
rect 6252 4753 6262 4779
rect 6208 4741 6262 4753
rect 6308 4787 6362 4960
rect 6590 4897 6620 6201
rect 6504 4891 6620 4897
rect 6504 4857 6516 4891
rect 6550 4857 6620 4891
rect 6504 4851 6620 4857
rect 6506 4802 6560 4814
rect 6308 4753 6318 4787
rect 6352 4753 6362 4787
rect 6108 4613 6118 4647
rect 6152 4613 6162 4647
rect 5908 4473 5918 4507
rect 5952 4473 5962 4507
rect 5708 4333 5718 4367
rect 5752 4333 5762 4367
rect 5508 4193 5518 4227
rect 5552 4193 5562 4227
rect 5308 4053 5318 4087
rect 5352 4053 5362 4087
rect 5108 3913 5118 3947
rect 5152 3913 5162 3947
rect 4908 3773 4918 3807
rect 4952 3773 4962 3807
rect 4802 3693 4868 3694
rect 4802 3641 4809 3693
rect 4861 3641 4868 3693
rect 4802 3640 4868 3641
rect 4708 3543 4718 3577
rect 4752 3543 4762 3577
rect 4508 3403 4518 3437
rect 4552 3403 4562 3437
rect 4308 3263 4318 3297
rect 4352 3263 4362 3297
rect 4108 3123 4118 3157
rect 4152 3123 4162 3157
rect 3908 2983 3918 3017
rect 3952 2983 3962 3017
rect 3708 2843 3718 2877
rect 3752 2843 3762 2877
rect 3508 2703 3518 2737
rect 3552 2703 3562 2737
rect 3308 2563 3318 2597
rect 3352 2563 3362 2597
rect 3202 2483 3268 2484
rect 3202 2431 3209 2483
rect 3261 2431 3268 2483
rect 3202 2430 3268 2431
rect 3108 2333 3118 2367
rect 3152 2333 3162 2367
rect 2908 2193 2918 2227
rect 2952 2193 2962 2227
rect 2708 2053 2718 2087
rect 2752 2053 2762 2087
rect 2508 1913 2518 1947
rect 2552 1913 2562 1947
rect 2308 1773 2318 1807
rect 2352 1773 2362 1807
rect 2108 1633 2118 1667
rect 2152 1633 2162 1667
rect 1908 1493 1918 1527
rect 1952 1493 1962 1527
rect 1708 1353 1718 1387
rect 1752 1353 1762 1387
rect 1602 1273 1668 1274
rect 1602 1221 1609 1273
rect 1661 1221 1668 1273
rect 1602 1220 1668 1221
rect 1508 1123 1518 1157
rect 1552 1123 1562 1157
rect 1308 983 1318 1017
rect 1352 983 1362 1017
rect 1108 843 1118 877
rect 1152 843 1162 877
rect 908 703 918 737
rect 952 703 962 737
rect 708 563 718 597
rect 752 563 762 597
rect 508 423 518 457
rect 552 423 562 457
rect 308 283 318 317
rect 352 283 362 317
rect 108 143 118 177
rect 152 143 162 177
rect 2 63 68 64
rect 2 11 9 63
rect 61 11 68 63
rect 2 10 68 11
rect -92 -15 -38 0
rect -92 -67 -91 -15
rect -39 -67 -38 -15
rect -92 -79 -82 -67
rect -48 -79 -38 -67
rect -92 -131 -91 -79
rect -39 -131 -38 -79
rect 8 -22 62 10
rect 8 -74 9 -22
rect 61 -74 62 -22
rect 8 -81 62 -74
rect 108 -15 162 143
rect 208 221 262 228
rect 208 169 209 221
rect 261 169 262 221
rect 208 143 218 169
rect 252 143 262 169
rect 208 131 262 143
rect 308 177 362 283
rect 408 317 462 329
rect 408 291 418 317
rect 452 291 462 317
rect 408 239 409 291
rect 461 239 462 291
rect 408 232 462 239
rect 508 317 562 423
rect 608 501 662 508
rect 608 449 609 501
rect 661 449 662 501
rect 608 423 618 449
rect 652 423 662 449
rect 608 411 662 423
rect 708 457 762 563
rect 808 597 862 609
rect 808 571 818 597
rect 852 571 862 597
rect 808 519 809 571
rect 861 519 862 571
rect 808 512 862 519
rect 908 597 962 703
rect 1008 781 1062 788
rect 1008 729 1009 781
rect 1061 729 1062 781
rect 1008 703 1018 729
rect 1052 703 1062 729
rect 1008 691 1062 703
rect 1108 737 1162 843
rect 1208 877 1262 889
rect 1208 851 1218 877
rect 1252 851 1262 877
rect 1208 799 1209 851
rect 1261 799 1262 851
rect 1208 792 1262 799
rect 1308 877 1362 983
rect 1408 1061 1462 1068
rect 1408 1009 1409 1061
rect 1461 1009 1462 1061
rect 1408 983 1418 1009
rect 1452 983 1462 1009
rect 1408 971 1462 983
rect 1508 1017 1562 1123
rect 1608 1157 1662 1169
rect 1608 1131 1618 1157
rect 1652 1131 1662 1157
rect 1608 1079 1609 1131
rect 1661 1079 1662 1131
rect 1608 1072 1662 1079
rect 1708 1157 1762 1353
rect 1808 1431 1862 1438
rect 1808 1379 1809 1431
rect 1861 1379 1862 1431
rect 1808 1353 1818 1379
rect 1852 1353 1862 1379
rect 1808 1341 1862 1353
rect 1908 1387 1962 1493
rect 2008 1527 2062 1539
rect 2008 1501 2018 1527
rect 2052 1501 2062 1527
rect 2008 1449 2009 1501
rect 2061 1449 2062 1501
rect 2008 1442 2062 1449
rect 2108 1527 2162 1633
rect 2208 1711 2262 1718
rect 2208 1659 2209 1711
rect 2261 1659 2262 1711
rect 2208 1633 2218 1659
rect 2252 1633 2262 1659
rect 2208 1621 2262 1633
rect 2308 1667 2362 1773
rect 2408 1807 2462 1819
rect 2408 1781 2418 1807
rect 2452 1781 2462 1807
rect 2408 1729 2409 1781
rect 2461 1729 2462 1781
rect 2408 1722 2462 1729
rect 2508 1807 2562 1913
rect 2608 1991 2662 1998
rect 2608 1939 2609 1991
rect 2661 1939 2662 1991
rect 2608 1913 2618 1939
rect 2652 1913 2662 1939
rect 2608 1901 2662 1913
rect 2708 1947 2762 2053
rect 2808 2087 2862 2099
rect 2808 2061 2818 2087
rect 2852 2061 2862 2087
rect 2808 2009 2809 2061
rect 2861 2009 2862 2061
rect 2808 2002 2862 2009
rect 2908 2087 2962 2193
rect 3008 2271 3062 2278
rect 3008 2219 3009 2271
rect 3061 2219 3062 2271
rect 3008 2193 3018 2219
rect 3052 2193 3062 2219
rect 3008 2181 3062 2193
rect 3108 2227 3162 2333
rect 3208 2367 3262 2379
rect 3208 2341 3218 2367
rect 3252 2341 3262 2367
rect 3208 2289 3209 2341
rect 3261 2289 3262 2341
rect 3208 2282 3262 2289
rect 3308 2367 3362 2563
rect 3408 2641 3462 2648
rect 3408 2589 3409 2641
rect 3461 2589 3462 2641
rect 3408 2563 3418 2589
rect 3452 2563 3462 2589
rect 3408 2551 3462 2563
rect 3508 2597 3562 2703
rect 3608 2737 3662 2749
rect 3608 2711 3618 2737
rect 3652 2711 3662 2737
rect 3608 2659 3609 2711
rect 3661 2659 3662 2711
rect 3608 2652 3662 2659
rect 3708 2737 3762 2843
rect 3808 2921 3862 2928
rect 3808 2869 3809 2921
rect 3861 2869 3862 2921
rect 3808 2843 3818 2869
rect 3852 2843 3862 2869
rect 3808 2831 3862 2843
rect 3908 2877 3962 2983
rect 4008 3017 4062 3029
rect 4008 2991 4018 3017
rect 4052 2991 4062 3017
rect 4008 2939 4009 2991
rect 4061 2939 4062 2991
rect 4008 2932 4062 2939
rect 4108 3017 4162 3123
rect 4208 3201 4262 3208
rect 4208 3149 4209 3201
rect 4261 3149 4262 3201
rect 4208 3123 4218 3149
rect 4252 3123 4262 3149
rect 4208 3111 4262 3123
rect 4308 3157 4362 3263
rect 4408 3297 4462 3309
rect 4408 3271 4418 3297
rect 4452 3271 4462 3297
rect 4408 3219 4409 3271
rect 4461 3219 4462 3271
rect 4408 3212 4462 3219
rect 4508 3297 4562 3403
rect 4608 3481 4662 3488
rect 4608 3429 4609 3481
rect 4661 3429 4662 3481
rect 4608 3403 4618 3429
rect 4652 3403 4662 3429
rect 4608 3391 4662 3403
rect 4708 3437 4762 3543
rect 4808 3577 4862 3589
rect 4808 3551 4818 3577
rect 4852 3551 4862 3577
rect 4808 3499 4809 3551
rect 4861 3499 4862 3551
rect 4808 3492 4862 3499
rect 4908 3577 4962 3773
rect 5008 3851 5062 3858
rect 5008 3799 5009 3851
rect 5061 3799 5062 3851
rect 5008 3773 5018 3799
rect 5052 3773 5062 3799
rect 5008 3761 5062 3773
rect 5108 3807 5162 3913
rect 5208 3947 5262 3959
rect 5208 3921 5218 3947
rect 5252 3921 5262 3947
rect 5208 3869 5209 3921
rect 5261 3869 5262 3921
rect 5208 3862 5262 3869
rect 5308 3947 5362 4053
rect 5408 4131 5462 4138
rect 5408 4079 5409 4131
rect 5461 4079 5462 4131
rect 5408 4053 5418 4079
rect 5452 4053 5462 4079
rect 5408 4041 5462 4053
rect 5508 4087 5562 4193
rect 5608 4227 5662 4239
rect 5608 4201 5618 4227
rect 5652 4201 5662 4227
rect 5608 4149 5609 4201
rect 5661 4149 5662 4201
rect 5608 4142 5662 4149
rect 5708 4227 5762 4333
rect 5808 4411 5862 4418
rect 5808 4359 5809 4411
rect 5861 4359 5862 4411
rect 5808 4333 5818 4359
rect 5852 4333 5862 4359
rect 5808 4321 5862 4333
rect 5908 4367 5962 4473
rect 6008 4507 6062 4519
rect 6008 4481 6018 4507
rect 6052 4481 6062 4507
rect 6008 4429 6009 4481
rect 6061 4429 6062 4481
rect 6008 4422 6062 4429
rect 6108 4507 6162 4613
rect 6208 4691 6262 4698
rect 6208 4639 6209 4691
rect 6261 4639 6262 4691
rect 6208 4613 6218 4639
rect 6252 4613 6262 4639
rect 6208 4601 6262 4613
rect 6308 4647 6362 4753
rect 6408 4787 6462 4799
rect 6408 4761 6418 4787
rect 6452 4761 6462 4787
rect 6408 4709 6409 4761
rect 6461 4709 6462 4761
rect 6408 4702 6462 4709
rect 6506 4768 6516 4802
rect 6550 4768 6560 4802
rect 6506 4761 6560 4768
rect 6506 4709 6507 4761
rect 6559 4709 6560 4761
rect 6506 4702 6560 4709
rect 6506 4662 6560 4674
rect 6308 4613 6318 4647
rect 6352 4613 6362 4647
rect 6108 4473 6118 4507
rect 6152 4473 6162 4507
rect 5908 4333 5918 4367
rect 5952 4333 5962 4367
rect 5708 4193 5718 4227
rect 5752 4193 5762 4227
rect 5508 4053 5518 4087
rect 5552 4053 5562 4087
rect 5308 3913 5318 3947
rect 5352 3913 5362 3947
rect 5108 3773 5118 3807
rect 5152 3773 5162 3807
rect 5002 3709 5068 3710
rect 5002 3657 5009 3709
rect 5061 3657 5068 3709
rect 5002 3656 5068 3657
rect 4908 3543 4918 3577
rect 4952 3543 4962 3577
rect 4708 3403 4718 3437
rect 4752 3403 4762 3437
rect 4508 3263 4518 3297
rect 4552 3263 4562 3297
rect 4308 3123 4318 3157
rect 4352 3123 4362 3157
rect 4108 2983 4118 3017
rect 4152 2983 4162 3017
rect 3908 2843 3918 2877
rect 3952 2843 3962 2877
rect 3708 2703 3718 2737
rect 3752 2703 3762 2737
rect 3508 2563 3518 2597
rect 3552 2563 3562 2597
rect 3402 2499 3468 2500
rect 3402 2447 3409 2499
rect 3461 2447 3468 2499
rect 3402 2446 3468 2447
rect 3308 2333 3318 2367
rect 3352 2333 3362 2367
rect 3108 2193 3118 2227
rect 3152 2193 3162 2227
rect 2908 2053 2918 2087
rect 2952 2053 2962 2087
rect 2708 1913 2718 1947
rect 2752 1913 2762 1947
rect 2508 1773 2518 1807
rect 2552 1773 2562 1807
rect 2308 1633 2318 1667
rect 2352 1633 2362 1667
rect 2108 1493 2118 1527
rect 2152 1493 2162 1527
rect 1908 1353 1918 1387
rect 1952 1353 1962 1387
rect 1802 1289 1868 1290
rect 1802 1237 1809 1289
rect 1861 1237 1868 1289
rect 1802 1236 1868 1237
rect 1708 1123 1718 1157
rect 1752 1123 1762 1157
rect 1508 983 1518 1017
rect 1552 983 1562 1017
rect 1308 843 1318 877
rect 1352 843 1362 877
rect 1108 703 1118 737
rect 1152 703 1162 737
rect 908 563 918 597
rect 952 563 962 597
rect 708 423 718 457
rect 752 423 762 457
rect 508 283 518 317
rect 552 283 562 317
rect 308 143 318 177
rect 352 143 362 177
rect 202 79 268 80
rect 202 27 209 79
rect 261 27 268 79
rect 202 26 268 27
rect 108 -67 109 -15
rect 161 -67 162 -15
rect 108 -79 118 -67
rect 152 -79 162 -67
rect -92 -132 -38 -131
rect -92 -143 -82 -132
rect -48 -143 -38 -132
rect -92 -195 -91 -143
rect -39 -195 -38 -143
rect -92 -210 -38 -195
rect 12 -133 58 -81
rect 12 -167 18 -133
rect 52 -167 58 -133
rect -82 -291 -75 -239
rect -23 -291 -16 -239
rect -91 -326 -39 -320
rect -91 -390 -82 -378
rect -48 -390 -39 -378
rect -91 -454 -82 -442
rect -48 -454 -39 -442
rect -91 -555 -39 -506
rect 12 -363 58 -167
rect 108 -131 109 -79
rect 161 -131 162 -79
rect 208 -22 262 26
rect 208 -74 209 -22
rect 261 -74 262 -22
rect 208 -81 262 -74
rect 308 -15 362 143
rect 408 177 462 189
rect 408 151 418 177
rect 452 151 462 177
rect 408 99 409 151
rect 461 99 462 151
rect 408 92 462 99
rect 508 177 562 283
rect 608 361 662 368
rect 608 309 609 361
rect 661 309 662 361
rect 608 283 618 309
rect 652 283 662 309
rect 608 271 662 283
rect 708 317 762 423
rect 808 457 862 469
rect 808 431 818 457
rect 852 431 862 457
rect 808 379 809 431
rect 861 379 862 431
rect 808 372 862 379
rect 908 457 962 563
rect 1008 641 1062 648
rect 1008 589 1009 641
rect 1061 589 1062 641
rect 1008 563 1018 589
rect 1052 563 1062 589
rect 1008 551 1062 563
rect 1108 597 1162 703
rect 1208 737 1262 749
rect 1208 711 1218 737
rect 1252 711 1262 737
rect 1208 659 1209 711
rect 1261 659 1262 711
rect 1208 652 1262 659
rect 1308 737 1362 843
rect 1408 921 1462 928
rect 1408 869 1409 921
rect 1461 869 1462 921
rect 1408 843 1418 869
rect 1452 843 1462 869
rect 1408 831 1462 843
rect 1508 877 1562 983
rect 1608 1017 1662 1029
rect 1608 991 1618 1017
rect 1652 991 1662 1017
rect 1608 939 1609 991
rect 1661 939 1662 991
rect 1608 932 1662 939
rect 1708 1017 1762 1123
rect 1808 1201 1862 1208
rect 1808 1149 1809 1201
rect 1861 1149 1862 1201
rect 1808 1123 1818 1149
rect 1852 1123 1862 1149
rect 1808 1111 1862 1123
rect 1908 1157 1962 1353
rect 2008 1387 2062 1399
rect 2008 1361 2018 1387
rect 2052 1361 2062 1387
rect 2008 1309 2009 1361
rect 2061 1309 2062 1361
rect 2008 1302 2062 1309
rect 2108 1387 2162 1493
rect 2208 1571 2262 1578
rect 2208 1519 2209 1571
rect 2261 1519 2262 1571
rect 2208 1493 2218 1519
rect 2252 1493 2262 1519
rect 2208 1481 2262 1493
rect 2308 1527 2362 1633
rect 2408 1667 2462 1679
rect 2408 1641 2418 1667
rect 2452 1641 2462 1667
rect 2408 1589 2409 1641
rect 2461 1589 2462 1641
rect 2408 1582 2462 1589
rect 2508 1667 2562 1773
rect 2608 1851 2662 1858
rect 2608 1799 2609 1851
rect 2661 1799 2662 1851
rect 2608 1773 2618 1799
rect 2652 1773 2662 1799
rect 2608 1761 2662 1773
rect 2708 1807 2762 1913
rect 2808 1947 2862 1959
rect 2808 1921 2818 1947
rect 2852 1921 2862 1947
rect 2808 1869 2809 1921
rect 2861 1869 2862 1921
rect 2808 1862 2862 1869
rect 2908 1947 2962 2053
rect 3008 2131 3062 2138
rect 3008 2079 3009 2131
rect 3061 2079 3062 2131
rect 3008 2053 3018 2079
rect 3052 2053 3062 2079
rect 3008 2041 3062 2053
rect 3108 2087 3162 2193
rect 3208 2227 3262 2239
rect 3208 2201 3218 2227
rect 3252 2201 3262 2227
rect 3208 2149 3209 2201
rect 3261 2149 3262 2201
rect 3208 2142 3262 2149
rect 3308 2227 3362 2333
rect 3408 2411 3462 2418
rect 3408 2359 3409 2411
rect 3461 2359 3462 2411
rect 3408 2333 3418 2359
rect 3452 2333 3462 2359
rect 3408 2321 3462 2333
rect 3508 2367 3562 2563
rect 3608 2597 3662 2609
rect 3608 2571 3618 2597
rect 3652 2571 3662 2597
rect 3608 2519 3609 2571
rect 3661 2519 3662 2571
rect 3608 2512 3662 2519
rect 3708 2597 3762 2703
rect 3808 2781 3862 2788
rect 3808 2729 3809 2781
rect 3861 2729 3862 2781
rect 3808 2703 3818 2729
rect 3852 2703 3862 2729
rect 3808 2691 3862 2703
rect 3908 2737 3962 2843
rect 4008 2877 4062 2889
rect 4008 2851 4018 2877
rect 4052 2851 4062 2877
rect 4008 2799 4009 2851
rect 4061 2799 4062 2851
rect 4008 2792 4062 2799
rect 4108 2877 4162 2983
rect 4208 3061 4262 3068
rect 4208 3009 4209 3061
rect 4261 3009 4262 3061
rect 4208 2983 4218 3009
rect 4252 2983 4262 3009
rect 4208 2971 4262 2983
rect 4308 3017 4362 3123
rect 4408 3157 4462 3169
rect 4408 3131 4418 3157
rect 4452 3131 4462 3157
rect 4408 3079 4409 3131
rect 4461 3079 4462 3131
rect 4408 3072 4462 3079
rect 4508 3157 4562 3263
rect 4608 3341 4662 3348
rect 4608 3289 4609 3341
rect 4661 3289 4662 3341
rect 4608 3263 4618 3289
rect 4652 3263 4662 3289
rect 4608 3251 4662 3263
rect 4708 3297 4762 3403
rect 4808 3437 4862 3449
rect 4808 3411 4818 3437
rect 4852 3411 4862 3437
rect 4808 3359 4809 3411
rect 4861 3359 4862 3411
rect 4808 3352 4862 3359
rect 4908 3437 4962 3543
rect 5008 3621 5062 3628
rect 5008 3569 5009 3621
rect 5061 3569 5062 3621
rect 5008 3543 5018 3569
rect 5052 3543 5062 3569
rect 5008 3531 5062 3543
rect 5108 3577 5162 3773
rect 5208 3807 5262 3819
rect 5208 3781 5218 3807
rect 5252 3781 5262 3807
rect 5208 3729 5209 3781
rect 5261 3729 5262 3781
rect 5208 3722 5262 3729
rect 5308 3807 5362 3913
rect 5408 3991 5462 3998
rect 5408 3939 5409 3991
rect 5461 3939 5462 3991
rect 5408 3913 5418 3939
rect 5452 3913 5462 3939
rect 5408 3901 5462 3913
rect 5508 3947 5562 4053
rect 5608 4087 5662 4099
rect 5608 4061 5618 4087
rect 5652 4061 5662 4087
rect 5608 4009 5609 4061
rect 5661 4009 5662 4061
rect 5608 4002 5662 4009
rect 5708 4087 5762 4193
rect 5808 4271 5862 4278
rect 5808 4219 5809 4271
rect 5861 4219 5862 4271
rect 5808 4193 5818 4219
rect 5852 4193 5862 4219
rect 5808 4181 5862 4193
rect 5908 4227 5962 4333
rect 6008 4367 6062 4379
rect 6008 4341 6018 4367
rect 6052 4341 6062 4367
rect 6008 4289 6009 4341
rect 6061 4289 6062 4341
rect 6008 4282 6062 4289
rect 6108 4367 6162 4473
rect 6208 4551 6262 4558
rect 6208 4499 6209 4551
rect 6261 4499 6262 4551
rect 6208 4473 6218 4499
rect 6252 4473 6262 4499
rect 6208 4461 6262 4473
rect 6308 4507 6362 4613
rect 6408 4647 6462 4659
rect 6408 4621 6418 4647
rect 6452 4621 6462 4647
rect 6408 4569 6409 4621
rect 6461 4569 6462 4621
rect 6408 4562 6462 4569
rect 6506 4628 6516 4662
rect 6550 4628 6560 4662
rect 6506 4621 6560 4628
rect 6506 4569 6507 4621
rect 6559 4569 6560 4621
rect 6506 4562 6560 4569
rect 6506 4522 6560 4534
rect 6308 4473 6318 4507
rect 6352 4473 6362 4507
rect 6108 4333 6118 4367
rect 6152 4333 6162 4367
rect 5908 4193 5918 4227
rect 5952 4193 5962 4227
rect 5708 4053 5718 4087
rect 5752 4053 5762 4087
rect 5508 3913 5518 3947
rect 5552 3913 5562 3947
rect 5308 3773 5318 3807
rect 5352 3773 5362 3807
rect 5202 3693 5268 3694
rect 5202 3641 5209 3693
rect 5261 3641 5268 3693
rect 5202 3640 5268 3641
rect 5108 3543 5118 3577
rect 5152 3543 5162 3577
rect 4908 3403 4918 3437
rect 4952 3403 4962 3437
rect 4708 3263 4718 3297
rect 4752 3263 4762 3297
rect 4508 3123 4518 3157
rect 4552 3123 4562 3157
rect 4308 2983 4318 3017
rect 4352 2983 4362 3017
rect 4108 2843 4118 2877
rect 4152 2843 4162 2877
rect 3908 2703 3918 2737
rect 3952 2703 3962 2737
rect 3708 2563 3718 2597
rect 3752 2563 3762 2597
rect 3602 2483 3668 2484
rect 3602 2431 3609 2483
rect 3661 2431 3668 2483
rect 3602 2430 3668 2431
rect 3508 2333 3518 2367
rect 3552 2333 3562 2367
rect 3308 2193 3318 2227
rect 3352 2193 3362 2227
rect 3108 2053 3118 2087
rect 3152 2053 3162 2087
rect 2908 1913 2918 1947
rect 2952 1913 2962 1947
rect 2708 1773 2718 1807
rect 2752 1773 2762 1807
rect 2508 1633 2518 1667
rect 2552 1633 2562 1667
rect 2308 1493 2318 1527
rect 2352 1493 2362 1527
rect 2108 1353 2118 1387
rect 2152 1353 2162 1387
rect 2002 1273 2068 1274
rect 2002 1221 2009 1273
rect 2061 1221 2068 1273
rect 2002 1220 2068 1221
rect 1908 1123 1918 1157
rect 1952 1123 1962 1157
rect 1708 983 1718 1017
rect 1752 983 1762 1017
rect 1508 843 1518 877
rect 1552 843 1562 877
rect 1308 703 1318 737
rect 1352 703 1362 737
rect 1108 563 1118 597
rect 1152 563 1162 597
rect 908 423 918 457
rect 952 423 962 457
rect 708 283 718 317
rect 752 283 762 317
rect 508 143 518 177
rect 552 143 562 177
rect 402 63 468 64
rect 402 11 409 63
rect 461 11 468 63
rect 402 10 468 11
rect 308 -67 309 -15
rect 361 -67 362 -15
rect 308 -79 318 -67
rect 352 -79 362 -67
rect 108 -132 162 -131
rect 108 -143 118 -132
rect 152 -143 162 -132
rect 108 -195 109 -143
rect 161 -195 162 -143
rect 108 -210 162 -195
rect 212 -133 258 -81
rect 212 -167 218 -133
rect 252 -167 258 -133
rect 118 -291 125 -239
rect 177 -291 184 -239
rect 12 -397 18 -363
rect 52 -397 58 -363
rect 12 -435 58 -397
rect 12 -469 18 -435
rect 52 -469 58 -435
rect 12 -512 58 -469
rect 109 -326 161 -320
rect 109 -390 118 -378
rect 152 -390 161 -378
rect 109 -454 118 -442
rect 152 -454 161 -442
rect 109 -512 161 -506
rect 212 -363 258 -167
rect 308 -131 309 -79
rect 361 -131 362 -79
rect 408 -22 462 10
rect 408 -74 409 -22
rect 461 -74 462 -22
rect 408 -81 462 -74
rect 508 -15 562 143
rect 608 221 662 228
rect 608 169 609 221
rect 661 169 662 221
rect 608 143 618 169
rect 652 143 662 169
rect 608 131 662 143
rect 708 177 762 283
rect 808 317 862 329
rect 808 291 818 317
rect 852 291 862 317
rect 808 239 809 291
rect 861 239 862 291
rect 808 232 862 239
rect 908 317 962 423
rect 1008 501 1062 508
rect 1008 449 1009 501
rect 1061 449 1062 501
rect 1008 423 1018 449
rect 1052 423 1062 449
rect 1008 411 1062 423
rect 1108 457 1162 563
rect 1208 597 1262 609
rect 1208 571 1218 597
rect 1252 571 1262 597
rect 1208 519 1209 571
rect 1261 519 1262 571
rect 1208 512 1262 519
rect 1308 597 1362 703
rect 1408 781 1462 788
rect 1408 729 1409 781
rect 1461 729 1462 781
rect 1408 703 1418 729
rect 1452 703 1462 729
rect 1408 691 1462 703
rect 1508 737 1562 843
rect 1608 877 1662 889
rect 1608 851 1618 877
rect 1652 851 1662 877
rect 1608 799 1609 851
rect 1661 799 1662 851
rect 1608 792 1662 799
rect 1708 877 1762 983
rect 1808 1061 1862 1068
rect 1808 1009 1809 1061
rect 1861 1009 1862 1061
rect 1808 983 1818 1009
rect 1852 983 1862 1009
rect 1808 971 1862 983
rect 1908 1017 1962 1123
rect 2008 1157 2062 1169
rect 2008 1131 2018 1157
rect 2052 1131 2062 1157
rect 2008 1079 2009 1131
rect 2061 1079 2062 1131
rect 2008 1072 2062 1079
rect 2108 1157 2162 1353
rect 2208 1431 2262 1438
rect 2208 1379 2209 1431
rect 2261 1379 2262 1431
rect 2208 1353 2218 1379
rect 2252 1353 2262 1379
rect 2208 1341 2262 1353
rect 2308 1387 2362 1493
rect 2408 1527 2462 1539
rect 2408 1501 2418 1527
rect 2452 1501 2462 1527
rect 2408 1449 2409 1501
rect 2461 1449 2462 1501
rect 2408 1442 2462 1449
rect 2508 1527 2562 1633
rect 2608 1711 2662 1718
rect 2608 1659 2609 1711
rect 2661 1659 2662 1711
rect 2608 1633 2618 1659
rect 2652 1633 2662 1659
rect 2608 1621 2662 1633
rect 2708 1667 2762 1773
rect 2808 1807 2862 1819
rect 2808 1781 2818 1807
rect 2852 1781 2862 1807
rect 2808 1729 2809 1781
rect 2861 1729 2862 1781
rect 2808 1722 2862 1729
rect 2908 1807 2962 1913
rect 3008 1991 3062 1998
rect 3008 1939 3009 1991
rect 3061 1939 3062 1991
rect 3008 1913 3018 1939
rect 3052 1913 3062 1939
rect 3008 1901 3062 1913
rect 3108 1947 3162 2053
rect 3208 2087 3262 2099
rect 3208 2061 3218 2087
rect 3252 2061 3262 2087
rect 3208 2009 3209 2061
rect 3261 2009 3262 2061
rect 3208 2002 3262 2009
rect 3308 2087 3362 2193
rect 3408 2271 3462 2278
rect 3408 2219 3409 2271
rect 3461 2219 3462 2271
rect 3408 2193 3418 2219
rect 3452 2193 3462 2219
rect 3408 2181 3462 2193
rect 3508 2227 3562 2333
rect 3608 2367 3662 2379
rect 3608 2341 3618 2367
rect 3652 2341 3662 2367
rect 3608 2289 3609 2341
rect 3661 2289 3662 2341
rect 3608 2282 3662 2289
rect 3708 2367 3762 2563
rect 3808 2641 3862 2648
rect 3808 2589 3809 2641
rect 3861 2589 3862 2641
rect 3808 2563 3818 2589
rect 3852 2563 3862 2589
rect 3808 2551 3862 2563
rect 3908 2597 3962 2703
rect 4008 2737 4062 2749
rect 4008 2711 4018 2737
rect 4052 2711 4062 2737
rect 4008 2659 4009 2711
rect 4061 2659 4062 2711
rect 4008 2652 4062 2659
rect 4108 2737 4162 2843
rect 4208 2921 4262 2928
rect 4208 2869 4209 2921
rect 4261 2869 4262 2921
rect 4208 2843 4218 2869
rect 4252 2843 4262 2869
rect 4208 2831 4262 2843
rect 4308 2877 4362 2983
rect 4408 3017 4462 3029
rect 4408 2991 4418 3017
rect 4452 2991 4462 3017
rect 4408 2939 4409 2991
rect 4461 2939 4462 2991
rect 4408 2932 4462 2939
rect 4508 3017 4562 3123
rect 4608 3201 4662 3208
rect 4608 3149 4609 3201
rect 4661 3149 4662 3201
rect 4608 3123 4618 3149
rect 4652 3123 4662 3149
rect 4608 3111 4662 3123
rect 4708 3157 4762 3263
rect 4808 3297 4862 3309
rect 4808 3271 4818 3297
rect 4852 3271 4862 3297
rect 4808 3219 4809 3271
rect 4861 3219 4862 3271
rect 4808 3212 4862 3219
rect 4908 3297 4962 3403
rect 5008 3481 5062 3488
rect 5008 3429 5009 3481
rect 5061 3429 5062 3481
rect 5008 3403 5018 3429
rect 5052 3403 5062 3429
rect 5008 3391 5062 3403
rect 5108 3437 5162 3543
rect 5208 3577 5262 3589
rect 5208 3551 5218 3577
rect 5252 3551 5262 3577
rect 5208 3499 5209 3551
rect 5261 3499 5262 3551
rect 5208 3492 5262 3499
rect 5308 3577 5362 3773
rect 5408 3851 5462 3858
rect 5408 3799 5409 3851
rect 5461 3799 5462 3851
rect 5408 3773 5418 3799
rect 5452 3773 5462 3799
rect 5408 3761 5462 3773
rect 5508 3807 5562 3913
rect 5608 3947 5662 3959
rect 5608 3921 5618 3947
rect 5652 3921 5662 3947
rect 5608 3869 5609 3921
rect 5661 3869 5662 3921
rect 5608 3862 5662 3869
rect 5708 3947 5762 4053
rect 5808 4131 5862 4138
rect 5808 4079 5809 4131
rect 5861 4079 5862 4131
rect 5808 4053 5818 4079
rect 5852 4053 5862 4079
rect 5808 4041 5862 4053
rect 5908 4087 5962 4193
rect 6008 4227 6062 4239
rect 6008 4201 6018 4227
rect 6052 4201 6062 4227
rect 6008 4149 6009 4201
rect 6061 4149 6062 4201
rect 6008 4142 6062 4149
rect 6108 4227 6162 4333
rect 6208 4411 6262 4418
rect 6208 4359 6209 4411
rect 6261 4359 6262 4411
rect 6208 4333 6218 4359
rect 6252 4333 6262 4359
rect 6208 4321 6262 4333
rect 6308 4367 6362 4473
rect 6408 4507 6462 4519
rect 6408 4481 6418 4507
rect 6452 4481 6462 4507
rect 6408 4429 6409 4481
rect 6461 4429 6462 4481
rect 6408 4422 6462 4429
rect 6506 4488 6516 4522
rect 6550 4488 6560 4522
rect 6506 4481 6560 4488
rect 6506 4429 6507 4481
rect 6559 4429 6560 4481
rect 6506 4422 6560 4429
rect 6506 4382 6560 4394
rect 6308 4333 6318 4367
rect 6352 4333 6362 4367
rect 6108 4193 6118 4227
rect 6152 4193 6162 4227
rect 5908 4053 5918 4087
rect 5952 4053 5962 4087
rect 5708 3913 5718 3947
rect 5752 3913 5762 3947
rect 5508 3773 5518 3807
rect 5552 3773 5562 3807
rect 5402 3709 5468 3710
rect 5402 3657 5409 3709
rect 5461 3657 5468 3709
rect 5402 3656 5468 3657
rect 5308 3543 5318 3577
rect 5352 3543 5362 3577
rect 5108 3403 5118 3437
rect 5152 3403 5162 3437
rect 4908 3263 4918 3297
rect 4952 3263 4962 3297
rect 4708 3123 4718 3157
rect 4752 3123 4762 3157
rect 4508 2983 4518 3017
rect 4552 2983 4562 3017
rect 4308 2843 4318 2877
rect 4352 2843 4362 2877
rect 4108 2703 4118 2737
rect 4152 2703 4162 2737
rect 3908 2563 3918 2597
rect 3952 2563 3962 2597
rect 3802 2499 3868 2500
rect 3802 2447 3809 2499
rect 3861 2447 3868 2499
rect 3802 2446 3868 2447
rect 3708 2333 3718 2367
rect 3752 2333 3762 2367
rect 3508 2193 3518 2227
rect 3552 2193 3562 2227
rect 3308 2053 3318 2087
rect 3352 2053 3362 2087
rect 3108 1913 3118 1947
rect 3152 1913 3162 1947
rect 2908 1773 2918 1807
rect 2952 1773 2962 1807
rect 2708 1633 2718 1667
rect 2752 1633 2762 1667
rect 2508 1493 2518 1527
rect 2552 1493 2562 1527
rect 2308 1353 2318 1387
rect 2352 1353 2362 1387
rect 2202 1289 2268 1290
rect 2202 1237 2209 1289
rect 2261 1237 2268 1289
rect 2202 1236 2268 1237
rect 2108 1123 2118 1157
rect 2152 1123 2162 1157
rect 1908 983 1918 1017
rect 1952 983 1962 1017
rect 1708 843 1718 877
rect 1752 843 1762 877
rect 1508 703 1518 737
rect 1552 703 1562 737
rect 1308 563 1318 597
rect 1352 563 1362 597
rect 1108 423 1118 457
rect 1152 423 1162 457
rect 908 283 918 317
rect 952 283 962 317
rect 708 143 718 177
rect 752 143 762 177
rect 602 79 668 80
rect 602 27 609 79
rect 661 27 668 79
rect 602 26 668 27
rect 508 -67 509 -15
rect 561 -67 562 -15
rect 508 -79 518 -67
rect 552 -79 562 -67
rect 308 -132 362 -131
rect 308 -143 318 -132
rect 352 -143 362 -132
rect 308 -195 309 -143
rect 361 -195 362 -143
rect 308 -210 362 -195
rect 412 -133 458 -81
rect 412 -167 418 -133
rect 452 -167 458 -133
rect 318 -291 325 -239
rect 377 -291 384 -239
rect 212 -397 218 -363
rect 252 -397 258 -363
rect 212 -435 258 -397
rect 212 -469 218 -435
rect 252 -469 258 -435
rect 212 -512 258 -469
rect 309 -326 361 -320
rect 309 -390 318 -378
rect 352 -390 361 -378
rect 309 -454 318 -442
rect 352 -454 361 -442
rect 309 -555 361 -506
rect 412 -363 458 -167
rect 508 -131 509 -79
rect 561 -131 562 -79
rect 608 -22 662 26
rect 608 -74 609 -22
rect 661 -74 662 -22
rect 608 -81 662 -74
rect 708 -15 762 143
rect 808 177 862 189
rect 808 151 818 177
rect 852 151 862 177
rect 808 99 809 151
rect 861 99 862 151
rect 808 92 862 99
rect 908 177 962 283
rect 1008 361 1062 368
rect 1008 309 1009 361
rect 1061 309 1062 361
rect 1008 283 1018 309
rect 1052 283 1062 309
rect 1008 271 1062 283
rect 1108 317 1162 423
rect 1208 457 1262 469
rect 1208 431 1218 457
rect 1252 431 1262 457
rect 1208 379 1209 431
rect 1261 379 1262 431
rect 1208 372 1262 379
rect 1308 457 1362 563
rect 1408 641 1462 648
rect 1408 589 1409 641
rect 1461 589 1462 641
rect 1408 563 1418 589
rect 1452 563 1462 589
rect 1408 551 1462 563
rect 1508 597 1562 703
rect 1608 737 1662 749
rect 1608 711 1618 737
rect 1652 711 1662 737
rect 1608 659 1609 711
rect 1661 659 1662 711
rect 1608 652 1662 659
rect 1708 737 1762 843
rect 1808 921 1862 928
rect 1808 869 1809 921
rect 1861 869 1862 921
rect 1808 843 1818 869
rect 1852 843 1862 869
rect 1808 831 1862 843
rect 1908 877 1962 983
rect 2008 1017 2062 1029
rect 2008 991 2018 1017
rect 2052 991 2062 1017
rect 2008 939 2009 991
rect 2061 939 2062 991
rect 2008 932 2062 939
rect 2108 1017 2162 1123
rect 2208 1201 2262 1208
rect 2208 1149 2209 1201
rect 2261 1149 2262 1201
rect 2208 1123 2218 1149
rect 2252 1123 2262 1149
rect 2208 1111 2262 1123
rect 2308 1157 2362 1353
rect 2408 1387 2462 1399
rect 2408 1361 2418 1387
rect 2452 1361 2462 1387
rect 2408 1309 2409 1361
rect 2461 1309 2462 1361
rect 2408 1302 2462 1309
rect 2508 1387 2562 1493
rect 2608 1571 2662 1578
rect 2608 1519 2609 1571
rect 2661 1519 2662 1571
rect 2608 1493 2618 1519
rect 2652 1493 2662 1519
rect 2608 1481 2662 1493
rect 2708 1527 2762 1633
rect 2808 1667 2862 1679
rect 2808 1641 2818 1667
rect 2852 1641 2862 1667
rect 2808 1589 2809 1641
rect 2861 1589 2862 1641
rect 2808 1582 2862 1589
rect 2908 1667 2962 1773
rect 3008 1851 3062 1858
rect 3008 1799 3009 1851
rect 3061 1799 3062 1851
rect 3008 1773 3018 1799
rect 3052 1773 3062 1799
rect 3008 1761 3062 1773
rect 3108 1807 3162 1913
rect 3208 1947 3262 1959
rect 3208 1921 3218 1947
rect 3252 1921 3262 1947
rect 3208 1869 3209 1921
rect 3261 1869 3262 1921
rect 3208 1862 3262 1869
rect 3308 1947 3362 2053
rect 3408 2131 3462 2138
rect 3408 2079 3409 2131
rect 3461 2079 3462 2131
rect 3408 2053 3418 2079
rect 3452 2053 3462 2079
rect 3408 2041 3462 2053
rect 3508 2087 3562 2193
rect 3608 2227 3662 2239
rect 3608 2201 3618 2227
rect 3652 2201 3662 2227
rect 3608 2149 3609 2201
rect 3661 2149 3662 2201
rect 3608 2142 3662 2149
rect 3708 2227 3762 2333
rect 3808 2411 3862 2418
rect 3808 2359 3809 2411
rect 3861 2359 3862 2411
rect 3808 2333 3818 2359
rect 3852 2333 3862 2359
rect 3808 2321 3862 2333
rect 3908 2367 3962 2563
rect 4008 2597 4062 2609
rect 4008 2571 4018 2597
rect 4052 2571 4062 2597
rect 4008 2519 4009 2571
rect 4061 2519 4062 2571
rect 4008 2512 4062 2519
rect 4108 2597 4162 2703
rect 4208 2781 4262 2788
rect 4208 2729 4209 2781
rect 4261 2729 4262 2781
rect 4208 2703 4218 2729
rect 4252 2703 4262 2729
rect 4208 2691 4262 2703
rect 4308 2737 4362 2843
rect 4408 2877 4462 2889
rect 4408 2851 4418 2877
rect 4452 2851 4462 2877
rect 4408 2799 4409 2851
rect 4461 2799 4462 2851
rect 4408 2792 4462 2799
rect 4508 2877 4562 2983
rect 4608 3061 4662 3068
rect 4608 3009 4609 3061
rect 4661 3009 4662 3061
rect 4608 2983 4618 3009
rect 4652 2983 4662 3009
rect 4608 2971 4662 2983
rect 4708 3017 4762 3123
rect 4808 3157 4862 3169
rect 4808 3131 4818 3157
rect 4852 3131 4862 3157
rect 4808 3079 4809 3131
rect 4861 3079 4862 3131
rect 4808 3072 4862 3079
rect 4908 3157 4962 3263
rect 5008 3341 5062 3348
rect 5008 3289 5009 3341
rect 5061 3289 5062 3341
rect 5008 3263 5018 3289
rect 5052 3263 5062 3289
rect 5008 3251 5062 3263
rect 5108 3297 5162 3403
rect 5208 3437 5262 3449
rect 5208 3411 5218 3437
rect 5252 3411 5262 3437
rect 5208 3359 5209 3411
rect 5261 3359 5262 3411
rect 5208 3352 5262 3359
rect 5308 3437 5362 3543
rect 5408 3621 5462 3628
rect 5408 3569 5409 3621
rect 5461 3569 5462 3621
rect 5408 3543 5418 3569
rect 5452 3543 5462 3569
rect 5408 3531 5462 3543
rect 5508 3577 5562 3773
rect 5608 3807 5662 3819
rect 5608 3781 5618 3807
rect 5652 3781 5662 3807
rect 5608 3729 5609 3781
rect 5661 3729 5662 3781
rect 5608 3722 5662 3729
rect 5708 3807 5762 3913
rect 5808 3991 5862 3998
rect 5808 3939 5809 3991
rect 5861 3939 5862 3991
rect 5808 3913 5818 3939
rect 5852 3913 5862 3939
rect 5808 3901 5862 3913
rect 5908 3947 5962 4053
rect 6008 4087 6062 4099
rect 6008 4061 6018 4087
rect 6052 4061 6062 4087
rect 6008 4009 6009 4061
rect 6061 4009 6062 4061
rect 6008 4002 6062 4009
rect 6108 4087 6162 4193
rect 6208 4271 6262 4278
rect 6208 4219 6209 4271
rect 6261 4219 6262 4271
rect 6208 4193 6218 4219
rect 6252 4193 6262 4219
rect 6208 4181 6262 4193
rect 6308 4227 6362 4333
rect 6408 4367 6462 4379
rect 6408 4341 6418 4367
rect 6452 4341 6462 4367
rect 6408 4289 6409 4341
rect 6461 4289 6462 4341
rect 6408 4282 6462 4289
rect 6506 4348 6516 4382
rect 6550 4348 6560 4382
rect 6506 4341 6560 4348
rect 6506 4289 6507 4341
rect 6559 4289 6560 4341
rect 6506 4282 6560 4289
rect 6506 4242 6560 4254
rect 6308 4193 6318 4227
rect 6352 4193 6362 4227
rect 6108 4053 6118 4087
rect 6152 4053 6162 4087
rect 5908 3913 5918 3947
rect 5952 3913 5962 3947
rect 5708 3773 5718 3807
rect 5752 3773 5762 3807
rect 5602 3693 5668 3694
rect 5602 3641 5609 3693
rect 5661 3641 5668 3693
rect 5602 3640 5668 3641
rect 5508 3543 5518 3577
rect 5552 3543 5562 3577
rect 5308 3403 5318 3437
rect 5352 3403 5362 3437
rect 5108 3263 5118 3297
rect 5152 3263 5162 3297
rect 4908 3123 4918 3157
rect 4952 3123 4962 3157
rect 4708 2983 4718 3017
rect 4752 2983 4762 3017
rect 4508 2843 4518 2877
rect 4552 2843 4562 2877
rect 4308 2703 4318 2737
rect 4352 2703 4362 2737
rect 4108 2563 4118 2597
rect 4152 2563 4162 2597
rect 4002 2483 4068 2484
rect 4002 2431 4009 2483
rect 4061 2431 4068 2483
rect 4002 2430 4068 2431
rect 3908 2333 3918 2367
rect 3952 2333 3962 2367
rect 3708 2193 3718 2227
rect 3752 2193 3762 2227
rect 3508 2053 3518 2087
rect 3552 2053 3562 2087
rect 3308 1913 3318 1947
rect 3352 1913 3362 1947
rect 3108 1773 3118 1807
rect 3152 1773 3162 1807
rect 2908 1633 2918 1667
rect 2952 1633 2962 1667
rect 2708 1493 2718 1527
rect 2752 1493 2762 1527
rect 2508 1353 2518 1387
rect 2552 1353 2562 1387
rect 2402 1273 2468 1274
rect 2402 1221 2409 1273
rect 2461 1221 2468 1273
rect 2402 1220 2468 1221
rect 2308 1123 2318 1157
rect 2352 1123 2362 1157
rect 2108 983 2118 1017
rect 2152 983 2162 1017
rect 1908 843 1918 877
rect 1952 843 1962 877
rect 1708 703 1718 737
rect 1752 703 1762 737
rect 1508 563 1518 597
rect 1552 563 1562 597
rect 1308 423 1318 457
rect 1352 423 1362 457
rect 1108 283 1118 317
rect 1152 283 1162 317
rect 908 143 918 177
rect 952 143 962 177
rect 802 63 868 64
rect 802 11 809 63
rect 861 11 868 63
rect 802 10 868 11
rect 708 -67 709 -15
rect 761 -67 762 -15
rect 708 -79 718 -67
rect 752 -79 762 -67
rect 508 -132 562 -131
rect 508 -143 518 -132
rect 552 -143 562 -132
rect 508 -195 509 -143
rect 561 -195 562 -143
rect 508 -210 562 -195
rect 612 -133 658 -81
rect 612 -167 618 -133
rect 652 -167 658 -133
rect 518 -291 525 -239
rect 577 -291 584 -239
rect 412 -397 418 -363
rect 452 -397 458 -363
rect 412 -435 458 -397
rect 412 -469 418 -435
rect 452 -469 458 -435
rect 412 -512 458 -469
rect 509 -326 561 -320
rect 509 -390 518 -378
rect 552 -390 561 -378
rect 509 -454 518 -442
rect 552 -454 561 -442
rect 509 -512 561 -506
rect 612 -363 658 -167
rect 708 -131 709 -79
rect 761 -131 762 -79
rect 808 -22 862 10
rect 808 -74 809 -22
rect 861 -74 862 -22
rect 808 -81 862 -74
rect 908 -15 962 143
rect 1008 221 1062 228
rect 1008 169 1009 221
rect 1061 169 1062 221
rect 1008 143 1018 169
rect 1052 143 1062 169
rect 1008 131 1062 143
rect 1108 177 1162 283
rect 1208 317 1262 329
rect 1208 291 1218 317
rect 1252 291 1262 317
rect 1208 239 1209 291
rect 1261 239 1262 291
rect 1208 232 1262 239
rect 1308 317 1362 423
rect 1408 501 1462 508
rect 1408 449 1409 501
rect 1461 449 1462 501
rect 1408 423 1418 449
rect 1452 423 1462 449
rect 1408 411 1462 423
rect 1508 457 1562 563
rect 1608 597 1662 609
rect 1608 571 1618 597
rect 1652 571 1662 597
rect 1608 519 1609 571
rect 1661 519 1662 571
rect 1608 512 1662 519
rect 1708 597 1762 703
rect 1808 781 1862 788
rect 1808 729 1809 781
rect 1861 729 1862 781
rect 1808 703 1818 729
rect 1852 703 1862 729
rect 1808 691 1862 703
rect 1908 737 1962 843
rect 2008 877 2062 889
rect 2008 851 2018 877
rect 2052 851 2062 877
rect 2008 799 2009 851
rect 2061 799 2062 851
rect 2008 792 2062 799
rect 2108 877 2162 983
rect 2208 1061 2262 1068
rect 2208 1009 2209 1061
rect 2261 1009 2262 1061
rect 2208 983 2218 1009
rect 2252 983 2262 1009
rect 2208 971 2262 983
rect 2308 1017 2362 1123
rect 2408 1157 2462 1169
rect 2408 1131 2418 1157
rect 2452 1131 2462 1157
rect 2408 1079 2409 1131
rect 2461 1079 2462 1131
rect 2408 1072 2462 1079
rect 2508 1157 2562 1353
rect 2608 1431 2662 1438
rect 2608 1379 2609 1431
rect 2661 1379 2662 1431
rect 2608 1353 2618 1379
rect 2652 1353 2662 1379
rect 2608 1341 2662 1353
rect 2708 1387 2762 1493
rect 2808 1527 2862 1539
rect 2808 1501 2818 1527
rect 2852 1501 2862 1527
rect 2808 1449 2809 1501
rect 2861 1449 2862 1501
rect 2808 1442 2862 1449
rect 2908 1527 2962 1633
rect 3008 1711 3062 1718
rect 3008 1659 3009 1711
rect 3061 1659 3062 1711
rect 3008 1633 3018 1659
rect 3052 1633 3062 1659
rect 3008 1621 3062 1633
rect 3108 1667 3162 1773
rect 3208 1807 3262 1819
rect 3208 1781 3218 1807
rect 3252 1781 3262 1807
rect 3208 1729 3209 1781
rect 3261 1729 3262 1781
rect 3208 1722 3262 1729
rect 3308 1807 3362 1913
rect 3408 1991 3462 1998
rect 3408 1939 3409 1991
rect 3461 1939 3462 1991
rect 3408 1913 3418 1939
rect 3452 1913 3462 1939
rect 3408 1901 3462 1913
rect 3508 1947 3562 2053
rect 3608 2087 3662 2099
rect 3608 2061 3618 2087
rect 3652 2061 3662 2087
rect 3608 2009 3609 2061
rect 3661 2009 3662 2061
rect 3608 2002 3662 2009
rect 3708 2087 3762 2193
rect 3808 2271 3862 2278
rect 3808 2219 3809 2271
rect 3861 2219 3862 2271
rect 3808 2193 3818 2219
rect 3852 2193 3862 2219
rect 3808 2181 3862 2193
rect 3908 2227 3962 2333
rect 4008 2367 4062 2379
rect 4008 2341 4018 2367
rect 4052 2341 4062 2367
rect 4008 2289 4009 2341
rect 4061 2289 4062 2341
rect 4008 2282 4062 2289
rect 4108 2367 4162 2563
rect 4208 2641 4262 2648
rect 4208 2589 4209 2641
rect 4261 2589 4262 2641
rect 4208 2563 4218 2589
rect 4252 2563 4262 2589
rect 4208 2551 4262 2563
rect 4308 2597 4362 2703
rect 4408 2737 4462 2749
rect 4408 2711 4418 2737
rect 4452 2711 4462 2737
rect 4408 2659 4409 2711
rect 4461 2659 4462 2711
rect 4408 2652 4462 2659
rect 4508 2737 4562 2843
rect 4608 2921 4662 2928
rect 4608 2869 4609 2921
rect 4661 2869 4662 2921
rect 4608 2843 4618 2869
rect 4652 2843 4662 2869
rect 4608 2831 4662 2843
rect 4708 2877 4762 2983
rect 4808 3017 4862 3029
rect 4808 2991 4818 3017
rect 4852 2991 4862 3017
rect 4808 2939 4809 2991
rect 4861 2939 4862 2991
rect 4808 2932 4862 2939
rect 4908 3017 4962 3123
rect 5008 3201 5062 3208
rect 5008 3149 5009 3201
rect 5061 3149 5062 3201
rect 5008 3123 5018 3149
rect 5052 3123 5062 3149
rect 5008 3111 5062 3123
rect 5108 3157 5162 3263
rect 5208 3297 5262 3309
rect 5208 3271 5218 3297
rect 5252 3271 5262 3297
rect 5208 3219 5209 3271
rect 5261 3219 5262 3271
rect 5208 3212 5262 3219
rect 5308 3297 5362 3403
rect 5408 3481 5462 3488
rect 5408 3429 5409 3481
rect 5461 3429 5462 3481
rect 5408 3403 5418 3429
rect 5452 3403 5462 3429
rect 5408 3391 5462 3403
rect 5508 3437 5562 3543
rect 5608 3577 5662 3589
rect 5608 3551 5618 3577
rect 5652 3551 5662 3577
rect 5608 3499 5609 3551
rect 5661 3499 5662 3551
rect 5608 3492 5662 3499
rect 5708 3577 5762 3773
rect 5808 3851 5862 3858
rect 5808 3799 5809 3851
rect 5861 3799 5862 3851
rect 5808 3773 5818 3799
rect 5852 3773 5862 3799
rect 5808 3761 5862 3773
rect 5908 3807 5962 3913
rect 6008 3947 6062 3959
rect 6008 3921 6018 3947
rect 6052 3921 6062 3947
rect 6008 3869 6009 3921
rect 6061 3869 6062 3921
rect 6008 3862 6062 3869
rect 6108 3947 6162 4053
rect 6208 4131 6262 4138
rect 6208 4079 6209 4131
rect 6261 4079 6262 4131
rect 6208 4053 6218 4079
rect 6252 4053 6262 4079
rect 6208 4041 6262 4053
rect 6308 4087 6362 4193
rect 6408 4227 6462 4239
rect 6408 4201 6418 4227
rect 6452 4201 6462 4227
rect 6408 4149 6409 4201
rect 6461 4149 6462 4201
rect 6408 4142 6462 4149
rect 6506 4208 6516 4242
rect 6550 4208 6560 4242
rect 6506 4201 6560 4208
rect 6506 4149 6507 4201
rect 6559 4149 6560 4201
rect 6506 4142 6560 4149
rect 6506 4102 6560 4114
rect 6308 4053 6318 4087
rect 6352 4053 6362 4087
rect 6108 3913 6118 3947
rect 6152 3913 6162 3947
rect 5908 3773 5918 3807
rect 5952 3773 5962 3807
rect 5802 3709 5868 3710
rect 5802 3657 5809 3709
rect 5861 3657 5868 3709
rect 5802 3656 5868 3657
rect 5708 3543 5718 3577
rect 5752 3543 5762 3577
rect 5508 3403 5518 3437
rect 5552 3403 5562 3437
rect 5308 3263 5318 3297
rect 5352 3263 5362 3297
rect 5108 3123 5118 3157
rect 5152 3123 5162 3157
rect 4908 2983 4918 3017
rect 4952 2983 4962 3017
rect 4708 2843 4718 2877
rect 4752 2843 4762 2877
rect 4508 2703 4518 2737
rect 4552 2703 4562 2737
rect 4308 2563 4318 2597
rect 4352 2563 4362 2597
rect 4202 2499 4268 2500
rect 4202 2447 4209 2499
rect 4261 2447 4268 2499
rect 4202 2446 4268 2447
rect 4108 2333 4118 2367
rect 4152 2333 4162 2367
rect 3908 2193 3918 2227
rect 3952 2193 3962 2227
rect 3708 2053 3718 2087
rect 3752 2053 3762 2087
rect 3508 1913 3518 1947
rect 3552 1913 3562 1947
rect 3308 1773 3318 1807
rect 3352 1773 3362 1807
rect 3108 1633 3118 1667
rect 3152 1633 3162 1667
rect 2908 1493 2918 1527
rect 2952 1493 2962 1527
rect 2708 1353 2718 1387
rect 2752 1353 2762 1387
rect 2602 1289 2668 1290
rect 2602 1237 2609 1289
rect 2661 1237 2668 1289
rect 2602 1236 2668 1237
rect 2508 1123 2518 1157
rect 2552 1123 2562 1157
rect 2308 983 2318 1017
rect 2352 983 2362 1017
rect 2108 843 2118 877
rect 2152 843 2162 877
rect 1908 703 1918 737
rect 1952 703 1962 737
rect 1708 563 1718 597
rect 1752 563 1762 597
rect 1508 423 1518 457
rect 1552 423 1562 457
rect 1308 283 1318 317
rect 1352 283 1362 317
rect 1108 143 1118 177
rect 1152 143 1162 177
rect 1002 79 1068 80
rect 1002 27 1009 79
rect 1061 27 1068 79
rect 1002 26 1068 27
rect 908 -67 909 -15
rect 961 -67 962 -15
rect 908 -79 918 -67
rect 952 -79 962 -67
rect 708 -132 762 -131
rect 708 -143 718 -132
rect 752 -143 762 -132
rect 708 -195 709 -143
rect 761 -195 762 -143
rect 708 -210 762 -195
rect 812 -133 858 -81
rect 812 -167 818 -133
rect 852 -167 858 -133
rect 718 -291 725 -239
rect 777 -291 784 -239
rect 612 -397 618 -363
rect 652 -397 658 -363
rect 612 -435 658 -397
rect 612 -469 618 -435
rect 652 -469 658 -435
rect 612 -512 658 -469
rect 709 -326 761 -320
rect 709 -390 718 -378
rect 752 -390 761 -378
rect 709 -454 718 -442
rect 752 -454 761 -442
rect 709 -555 761 -506
rect 812 -363 858 -167
rect 908 -131 909 -79
rect 961 -131 962 -79
rect 1008 -22 1062 26
rect 1008 -74 1009 -22
rect 1061 -74 1062 -22
rect 1008 -81 1062 -74
rect 1108 -15 1162 143
rect 1208 177 1262 189
rect 1208 151 1218 177
rect 1252 151 1262 177
rect 1208 99 1209 151
rect 1261 99 1262 151
rect 1208 92 1262 99
rect 1308 177 1362 283
rect 1408 361 1462 368
rect 1408 309 1409 361
rect 1461 309 1462 361
rect 1408 283 1418 309
rect 1452 283 1462 309
rect 1408 271 1462 283
rect 1508 317 1562 423
rect 1608 457 1662 469
rect 1608 431 1618 457
rect 1652 431 1662 457
rect 1608 379 1609 431
rect 1661 379 1662 431
rect 1608 372 1662 379
rect 1708 457 1762 563
rect 1808 641 1862 648
rect 1808 589 1809 641
rect 1861 589 1862 641
rect 1808 563 1818 589
rect 1852 563 1862 589
rect 1808 551 1862 563
rect 1908 597 1962 703
rect 2008 737 2062 749
rect 2008 711 2018 737
rect 2052 711 2062 737
rect 2008 659 2009 711
rect 2061 659 2062 711
rect 2008 652 2062 659
rect 2108 737 2162 843
rect 2208 921 2262 928
rect 2208 869 2209 921
rect 2261 869 2262 921
rect 2208 843 2218 869
rect 2252 843 2262 869
rect 2208 831 2262 843
rect 2308 877 2362 983
rect 2408 1017 2462 1029
rect 2408 991 2418 1017
rect 2452 991 2462 1017
rect 2408 939 2409 991
rect 2461 939 2462 991
rect 2408 932 2462 939
rect 2508 1017 2562 1123
rect 2608 1201 2662 1208
rect 2608 1149 2609 1201
rect 2661 1149 2662 1201
rect 2608 1123 2618 1149
rect 2652 1123 2662 1149
rect 2608 1111 2662 1123
rect 2708 1157 2762 1353
rect 2808 1387 2862 1399
rect 2808 1361 2818 1387
rect 2852 1361 2862 1387
rect 2808 1309 2809 1361
rect 2861 1309 2862 1361
rect 2808 1302 2862 1309
rect 2908 1387 2962 1493
rect 3008 1571 3062 1578
rect 3008 1519 3009 1571
rect 3061 1519 3062 1571
rect 3008 1493 3018 1519
rect 3052 1493 3062 1519
rect 3008 1481 3062 1493
rect 3108 1527 3162 1633
rect 3208 1667 3262 1679
rect 3208 1641 3218 1667
rect 3252 1641 3262 1667
rect 3208 1589 3209 1641
rect 3261 1589 3262 1641
rect 3208 1582 3262 1589
rect 3308 1667 3362 1773
rect 3408 1851 3462 1858
rect 3408 1799 3409 1851
rect 3461 1799 3462 1851
rect 3408 1773 3418 1799
rect 3452 1773 3462 1799
rect 3408 1761 3462 1773
rect 3508 1807 3562 1913
rect 3608 1947 3662 1959
rect 3608 1921 3618 1947
rect 3652 1921 3662 1947
rect 3608 1869 3609 1921
rect 3661 1869 3662 1921
rect 3608 1862 3662 1869
rect 3708 1947 3762 2053
rect 3808 2131 3862 2138
rect 3808 2079 3809 2131
rect 3861 2079 3862 2131
rect 3808 2053 3818 2079
rect 3852 2053 3862 2079
rect 3808 2041 3862 2053
rect 3908 2087 3962 2193
rect 4008 2227 4062 2239
rect 4008 2201 4018 2227
rect 4052 2201 4062 2227
rect 4008 2149 4009 2201
rect 4061 2149 4062 2201
rect 4008 2142 4062 2149
rect 4108 2227 4162 2333
rect 4208 2411 4262 2418
rect 4208 2359 4209 2411
rect 4261 2359 4262 2411
rect 4208 2333 4218 2359
rect 4252 2333 4262 2359
rect 4208 2321 4262 2333
rect 4308 2367 4362 2563
rect 4408 2597 4462 2609
rect 4408 2571 4418 2597
rect 4452 2571 4462 2597
rect 4408 2519 4409 2571
rect 4461 2519 4462 2571
rect 4408 2512 4462 2519
rect 4508 2597 4562 2703
rect 4608 2781 4662 2788
rect 4608 2729 4609 2781
rect 4661 2729 4662 2781
rect 4608 2703 4618 2729
rect 4652 2703 4662 2729
rect 4608 2691 4662 2703
rect 4708 2737 4762 2843
rect 4808 2877 4862 2889
rect 4808 2851 4818 2877
rect 4852 2851 4862 2877
rect 4808 2799 4809 2851
rect 4861 2799 4862 2851
rect 4808 2792 4862 2799
rect 4908 2877 4962 2983
rect 5008 3061 5062 3068
rect 5008 3009 5009 3061
rect 5061 3009 5062 3061
rect 5008 2983 5018 3009
rect 5052 2983 5062 3009
rect 5008 2971 5062 2983
rect 5108 3017 5162 3123
rect 5208 3157 5262 3169
rect 5208 3131 5218 3157
rect 5252 3131 5262 3157
rect 5208 3079 5209 3131
rect 5261 3079 5262 3131
rect 5208 3072 5262 3079
rect 5308 3157 5362 3263
rect 5408 3341 5462 3348
rect 5408 3289 5409 3341
rect 5461 3289 5462 3341
rect 5408 3263 5418 3289
rect 5452 3263 5462 3289
rect 5408 3251 5462 3263
rect 5508 3297 5562 3403
rect 5608 3437 5662 3449
rect 5608 3411 5618 3437
rect 5652 3411 5662 3437
rect 5608 3359 5609 3411
rect 5661 3359 5662 3411
rect 5608 3352 5662 3359
rect 5708 3437 5762 3543
rect 5808 3621 5862 3628
rect 5808 3569 5809 3621
rect 5861 3569 5862 3621
rect 5808 3543 5818 3569
rect 5852 3543 5862 3569
rect 5808 3531 5862 3543
rect 5908 3577 5962 3773
rect 6008 3807 6062 3819
rect 6008 3781 6018 3807
rect 6052 3781 6062 3807
rect 6008 3729 6009 3781
rect 6061 3729 6062 3781
rect 6008 3722 6062 3729
rect 6108 3807 6162 3913
rect 6208 3991 6262 3998
rect 6208 3939 6209 3991
rect 6261 3939 6262 3991
rect 6208 3913 6218 3939
rect 6252 3913 6262 3939
rect 6208 3901 6262 3913
rect 6308 3947 6362 4053
rect 6408 4087 6462 4099
rect 6408 4061 6418 4087
rect 6452 4061 6462 4087
rect 6408 4009 6409 4061
rect 6461 4009 6462 4061
rect 6408 4002 6462 4009
rect 6506 4068 6516 4102
rect 6550 4068 6560 4102
rect 6506 4061 6560 4068
rect 6506 4009 6507 4061
rect 6559 4009 6560 4061
rect 6506 4002 6560 4009
rect 6506 3962 6560 3974
rect 6308 3913 6318 3947
rect 6352 3913 6362 3947
rect 6108 3773 6118 3807
rect 6152 3773 6162 3807
rect 6002 3693 6068 3694
rect 6002 3641 6009 3693
rect 6061 3641 6068 3693
rect 6002 3640 6068 3641
rect 5908 3543 5918 3577
rect 5952 3543 5962 3577
rect 5708 3403 5718 3437
rect 5752 3403 5762 3437
rect 5508 3263 5518 3297
rect 5552 3263 5562 3297
rect 5308 3123 5318 3157
rect 5352 3123 5362 3157
rect 5108 2983 5118 3017
rect 5152 2983 5162 3017
rect 4908 2843 4918 2877
rect 4952 2843 4962 2877
rect 4708 2703 4718 2737
rect 4752 2703 4762 2737
rect 4508 2563 4518 2597
rect 4552 2563 4562 2597
rect 4402 2483 4468 2484
rect 4402 2431 4409 2483
rect 4461 2431 4468 2483
rect 4402 2430 4468 2431
rect 4308 2333 4318 2367
rect 4352 2333 4362 2367
rect 4108 2193 4118 2227
rect 4152 2193 4162 2227
rect 3908 2053 3918 2087
rect 3952 2053 3962 2087
rect 3708 1913 3718 1947
rect 3752 1913 3762 1947
rect 3508 1773 3518 1807
rect 3552 1773 3562 1807
rect 3308 1633 3318 1667
rect 3352 1633 3362 1667
rect 3108 1493 3118 1527
rect 3152 1493 3162 1527
rect 2908 1353 2918 1387
rect 2952 1353 2962 1387
rect 2802 1273 2868 1274
rect 2802 1221 2809 1273
rect 2861 1221 2868 1273
rect 2802 1220 2868 1221
rect 2708 1123 2718 1157
rect 2752 1123 2762 1157
rect 2508 983 2518 1017
rect 2552 983 2562 1017
rect 2308 843 2318 877
rect 2352 843 2362 877
rect 2108 703 2118 737
rect 2152 703 2162 737
rect 1908 563 1918 597
rect 1952 563 1962 597
rect 1708 423 1718 457
rect 1752 423 1762 457
rect 1508 283 1518 317
rect 1552 283 1562 317
rect 1308 143 1318 177
rect 1352 143 1362 177
rect 1202 63 1268 64
rect 1202 11 1209 63
rect 1261 11 1268 63
rect 1202 10 1268 11
rect 1108 -67 1109 -15
rect 1161 -67 1162 -15
rect 1108 -79 1118 -67
rect 1152 -79 1162 -67
rect 908 -132 962 -131
rect 908 -143 918 -132
rect 952 -143 962 -132
rect 908 -195 909 -143
rect 961 -195 962 -143
rect 908 -210 962 -195
rect 1012 -133 1058 -81
rect 1012 -167 1018 -133
rect 1052 -167 1058 -133
rect 918 -291 925 -239
rect 977 -291 984 -239
rect 812 -397 818 -363
rect 852 -397 858 -363
rect 812 -435 858 -397
rect 812 -469 818 -435
rect 852 -469 858 -435
rect 812 -512 858 -469
rect 909 -326 961 -320
rect 909 -390 918 -378
rect 952 -390 961 -378
rect 909 -454 918 -442
rect 952 -454 961 -442
rect 909 -512 961 -506
rect 1012 -363 1058 -167
rect 1108 -131 1109 -79
rect 1161 -131 1162 -79
rect 1208 -22 1262 10
rect 1208 -74 1209 -22
rect 1261 -74 1262 -22
rect 1208 -81 1262 -74
rect 1308 -15 1362 143
rect 1408 221 1462 228
rect 1408 169 1409 221
rect 1461 169 1462 221
rect 1408 143 1418 169
rect 1452 143 1462 169
rect 1408 131 1462 143
rect 1508 177 1562 283
rect 1608 317 1662 329
rect 1608 291 1618 317
rect 1652 291 1662 317
rect 1608 239 1609 291
rect 1661 239 1662 291
rect 1608 232 1662 239
rect 1708 317 1762 423
rect 1808 501 1862 508
rect 1808 449 1809 501
rect 1861 449 1862 501
rect 1808 423 1818 449
rect 1852 423 1862 449
rect 1808 411 1862 423
rect 1908 457 1962 563
rect 2008 597 2062 609
rect 2008 571 2018 597
rect 2052 571 2062 597
rect 2008 519 2009 571
rect 2061 519 2062 571
rect 2008 512 2062 519
rect 2108 597 2162 703
rect 2208 781 2262 788
rect 2208 729 2209 781
rect 2261 729 2262 781
rect 2208 703 2218 729
rect 2252 703 2262 729
rect 2208 691 2262 703
rect 2308 737 2362 843
rect 2408 877 2462 889
rect 2408 851 2418 877
rect 2452 851 2462 877
rect 2408 799 2409 851
rect 2461 799 2462 851
rect 2408 792 2462 799
rect 2508 877 2562 983
rect 2608 1061 2662 1068
rect 2608 1009 2609 1061
rect 2661 1009 2662 1061
rect 2608 983 2618 1009
rect 2652 983 2662 1009
rect 2608 971 2662 983
rect 2708 1017 2762 1123
rect 2808 1157 2862 1169
rect 2808 1131 2818 1157
rect 2852 1131 2862 1157
rect 2808 1079 2809 1131
rect 2861 1079 2862 1131
rect 2808 1072 2862 1079
rect 2908 1157 2962 1353
rect 3008 1431 3062 1438
rect 3008 1379 3009 1431
rect 3061 1379 3062 1431
rect 3008 1353 3018 1379
rect 3052 1353 3062 1379
rect 3008 1341 3062 1353
rect 3108 1387 3162 1493
rect 3208 1527 3262 1539
rect 3208 1501 3218 1527
rect 3252 1501 3262 1527
rect 3208 1449 3209 1501
rect 3261 1449 3262 1501
rect 3208 1442 3262 1449
rect 3308 1527 3362 1633
rect 3408 1711 3462 1718
rect 3408 1659 3409 1711
rect 3461 1659 3462 1711
rect 3408 1633 3418 1659
rect 3452 1633 3462 1659
rect 3408 1621 3462 1633
rect 3508 1667 3562 1773
rect 3608 1807 3662 1819
rect 3608 1781 3618 1807
rect 3652 1781 3662 1807
rect 3608 1729 3609 1781
rect 3661 1729 3662 1781
rect 3608 1722 3662 1729
rect 3708 1807 3762 1913
rect 3808 1991 3862 1998
rect 3808 1939 3809 1991
rect 3861 1939 3862 1991
rect 3808 1913 3818 1939
rect 3852 1913 3862 1939
rect 3808 1901 3862 1913
rect 3908 1947 3962 2053
rect 4008 2087 4062 2099
rect 4008 2061 4018 2087
rect 4052 2061 4062 2087
rect 4008 2009 4009 2061
rect 4061 2009 4062 2061
rect 4008 2002 4062 2009
rect 4108 2087 4162 2193
rect 4208 2271 4262 2278
rect 4208 2219 4209 2271
rect 4261 2219 4262 2271
rect 4208 2193 4218 2219
rect 4252 2193 4262 2219
rect 4208 2181 4262 2193
rect 4308 2227 4362 2333
rect 4408 2367 4462 2379
rect 4408 2341 4418 2367
rect 4452 2341 4462 2367
rect 4408 2289 4409 2341
rect 4461 2289 4462 2341
rect 4408 2282 4462 2289
rect 4508 2367 4562 2563
rect 4608 2641 4662 2648
rect 4608 2589 4609 2641
rect 4661 2589 4662 2641
rect 4608 2563 4618 2589
rect 4652 2563 4662 2589
rect 4608 2551 4662 2563
rect 4708 2597 4762 2703
rect 4808 2737 4862 2749
rect 4808 2711 4818 2737
rect 4852 2711 4862 2737
rect 4808 2659 4809 2711
rect 4861 2659 4862 2711
rect 4808 2652 4862 2659
rect 4908 2737 4962 2843
rect 5008 2921 5062 2928
rect 5008 2869 5009 2921
rect 5061 2869 5062 2921
rect 5008 2843 5018 2869
rect 5052 2843 5062 2869
rect 5008 2831 5062 2843
rect 5108 2877 5162 2983
rect 5208 3017 5262 3029
rect 5208 2991 5218 3017
rect 5252 2991 5262 3017
rect 5208 2939 5209 2991
rect 5261 2939 5262 2991
rect 5208 2932 5262 2939
rect 5308 3017 5362 3123
rect 5408 3201 5462 3208
rect 5408 3149 5409 3201
rect 5461 3149 5462 3201
rect 5408 3123 5418 3149
rect 5452 3123 5462 3149
rect 5408 3111 5462 3123
rect 5508 3157 5562 3263
rect 5608 3297 5662 3309
rect 5608 3271 5618 3297
rect 5652 3271 5662 3297
rect 5608 3219 5609 3271
rect 5661 3219 5662 3271
rect 5608 3212 5662 3219
rect 5708 3297 5762 3403
rect 5808 3481 5862 3488
rect 5808 3429 5809 3481
rect 5861 3429 5862 3481
rect 5808 3403 5818 3429
rect 5852 3403 5862 3429
rect 5808 3391 5862 3403
rect 5908 3437 5962 3543
rect 6008 3577 6062 3589
rect 6008 3551 6018 3577
rect 6052 3551 6062 3577
rect 6008 3499 6009 3551
rect 6061 3499 6062 3551
rect 6008 3492 6062 3499
rect 6108 3577 6162 3773
rect 6208 3851 6262 3858
rect 6208 3799 6209 3851
rect 6261 3799 6262 3851
rect 6208 3773 6218 3799
rect 6252 3773 6262 3799
rect 6208 3761 6262 3773
rect 6308 3807 6362 3913
rect 6408 3947 6462 3959
rect 6408 3921 6418 3947
rect 6452 3921 6462 3947
rect 6408 3869 6409 3921
rect 6461 3869 6462 3921
rect 6408 3862 6462 3869
rect 6506 3928 6516 3962
rect 6550 3928 6560 3962
rect 6506 3921 6560 3928
rect 6506 3869 6507 3921
rect 6559 3869 6560 3921
rect 6506 3862 6560 3869
rect 6506 3822 6560 3834
rect 6308 3773 6318 3807
rect 6352 3773 6362 3807
rect 6202 3709 6268 3710
rect 6202 3657 6209 3709
rect 6261 3657 6268 3709
rect 6202 3656 6268 3657
rect 6108 3543 6118 3577
rect 6152 3543 6162 3577
rect 5908 3403 5918 3437
rect 5952 3403 5962 3437
rect 5708 3263 5718 3297
rect 5752 3263 5762 3297
rect 5508 3123 5518 3157
rect 5552 3123 5562 3157
rect 5308 2983 5318 3017
rect 5352 2983 5362 3017
rect 5108 2843 5118 2877
rect 5152 2843 5162 2877
rect 4908 2703 4918 2737
rect 4952 2703 4962 2737
rect 4708 2563 4718 2597
rect 4752 2563 4762 2597
rect 4602 2499 4668 2500
rect 4602 2447 4609 2499
rect 4661 2447 4668 2499
rect 4602 2446 4668 2447
rect 4508 2333 4518 2367
rect 4552 2333 4562 2367
rect 4308 2193 4318 2227
rect 4352 2193 4362 2227
rect 4108 2053 4118 2087
rect 4152 2053 4162 2087
rect 3908 1913 3918 1947
rect 3952 1913 3962 1947
rect 3708 1773 3718 1807
rect 3752 1773 3762 1807
rect 3508 1633 3518 1667
rect 3552 1633 3562 1667
rect 3308 1493 3318 1527
rect 3352 1493 3362 1527
rect 3108 1353 3118 1387
rect 3152 1353 3162 1387
rect 3002 1289 3068 1290
rect 3002 1237 3009 1289
rect 3061 1237 3068 1289
rect 3002 1236 3068 1237
rect 2908 1123 2918 1157
rect 2952 1123 2962 1157
rect 2708 983 2718 1017
rect 2752 983 2762 1017
rect 2508 843 2518 877
rect 2552 843 2562 877
rect 2308 703 2318 737
rect 2352 703 2362 737
rect 2108 563 2118 597
rect 2152 563 2162 597
rect 1908 423 1918 457
rect 1952 423 1962 457
rect 1708 283 1718 317
rect 1752 283 1762 317
rect 1508 143 1518 177
rect 1552 143 1562 177
rect 1402 79 1468 80
rect 1402 27 1409 79
rect 1461 27 1468 79
rect 1402 26 1468 27
rect 1308 -67 1309 -15
rect 1361 -67 1362 -15
rect 1308 -79 1318 -67
rect 1352 -79 1362 -67
rect 1108 -132 1162 -131
rect 1108 -143 1118 -132
rect 1152 -143 1162 -132
rect 1108 -195 1109 -143
rect 1161 -195 1162 -143
rect 1108 -210 1162 -195
rect 1212 -133 1258 -81
rect 1212 -167 1218 -133
rect 1252 -167 1258 -133
rect 1118 -291 1125 -239
rect 1177 -291 1184 -239
rect 1012 -397 1018 -363
rect 1052 -397 1058 -363
rect 1012 -435 1058 -397
rect 1012 -469 1018 -435
rect 1052 -469 1058 -435
rect 1012 -512 1058 -469
rect 1109 -326 1161 -320
rect 1109 -390 1118 -378
rect 1152 -390 1161 -378
rect 1109 -454 1118 -442
rect 1152 -454 1161 -442
rect 1109 -555 1161 -506
rect 1212 -363 1258 -167
rect 1308 -131 1309 -79
rect 1361 -131 1362 -79
rect 1408 -22 1462 26
rect 1408 -74 1409 -22
rect 1461 -74 1462 -22
rect 1408 -81 1462 -74
rect 1508 -15 1562 143
rect 1608 177 1662 189
rect 1608 151 1618 177
rect 1652 151 1662 177
rect 1608 99 1609 151
rect 1661 99 1662 151
rect 1608 92 1662 99
rect 1708 177 1762 283
rect 1808 361 1862 368
rect 1808 309 1809 361
rect 1861 309 1862 361
rect 1808 283 1818 309
rect 1852 283 1862 309
rect 1808 271 1862 283
rect 1908 317 1962 423
rect 2008 457 2062 469
rect 2008 431 2018 457
rect 2052 431 2062 457
rect 2008 379 2009 431
rect 2061 379 2062 431
rect 2008 372 2062 379
rect 2108 457 2162 563
rect 2208 641 2262 648
rect 2208 589 2209 641
rect 2261 589 2262 641
rect 2208 563 2218 589
rect 2252 563 2262 589
rect 2208 551 2262 563
rect 2308 597 2362 703
rect 2408 737 2462 749
rect 2408 711 2418 737
rect 2452 711 2462 737
rect 2408 659 2409 711
rect 2461 659 2462 711
rect 2408 652 2462 659
rect 2508 737 2562 843
rect 2608 921 2662 928
rect 2608 869 2609 921
rect 2661 869 2662 921
rect 2608 843 2618 869
rect 2652 843 2662 869
rect 2608 831 2662 843
rect 2708 877 2762 983
rect 2808 1017 2862 1029
rect 2808 991 2818 1017
rect 2852 991 2862 1017
rect 2808 939 2809 991
rect 2861 939 2862 991
rect 2808 932 2862 939
rect 2908 1017 2962 1123
rect 3008 1201 3062 1208
rect 3008 1149 3009 1201
rect 3061 1149 3062 1201
rect 3008 1123 3018 1149
rect 3052 1123 3062 1149
rect 3008 1111 3062 1123
rect 3108 1157 3162 1353
rect 3208 1387 3262 1399
rect 3208 1361 3218 1387
rect 3252 1361 3262 1387
rect 3208 1309 3209 1361
rect 3261 1309 3262 1361
rect 3208 1302 3262 1309
rect 3308 1387 3362 1493
rect 3408 1571 3462 1578
rect 3408 1519 3409 1571
rect 3461 1519 3462 1571
rect 3408 1493 3418 1519
rect 3452 1493 3462 1519
rect 3408 1481 3462 1493
rect 3508 1527 3562 1633
rect 3608 1667 3662 1679
rect 3608 1641 3618 1667
rect 3652 1641 3662 1667
rect 3608 1589 3609 1641
rect 3661 1589 3662 1641
rect 3608 1582 3662 1589
rect 3708 1667 3762 1773
rect 3808 1851 3862 1858
rect 3808 1799 3809 1851
rect 3861 1799 3862 1851
rect 3808 1773 3818 1799
rect 3852 1773 3862 1799
rect 3808 1761 3862 1773
rect 3908 1807 3962 1913
rect 4008 1947 4062 1959
rect 4008 1921 4018 1947
rect 4052 1921 4062 1947
rect 4008 1869 4009 1921
rect 4061 1869 4062 1921
rect 4008 1862 4062 1869
rect 4108 1947 4162 2053
rect 4208 2131 4262 2138
rect 4208 2079 4209 2131
rect 4261 2079 4262 2131
rect 4208 2053 4218 2079
rect 4252 2053 4262 2079
rect 4208 2041 4262 2053
rect 4308 2087 4362 2193
rect 4408 2227 4462 2239
rect 4408 2201 4418 2227
rect 4452 2201 4462 2227
rect 4408 2149 4409 2201
rect 4461 2149 4462 2201
rect 4408 2142 4462 2149
rect 4508 2227 4562 2333
rect 4608 2411 4662 2418
rect 4608 2359 4609 2411
rect 4661 2359 4662 2411
rect 4608 2333 4618 2359
rect 4652 2333 4662 2359
rect 4608 2321 4662 2333
rect 4708 2367 4762 2563
rect 4808 2597 4862 2609
rect 4808 2571 4818 2597
rect 4852 2571 4862 2597
rect 4808 2519 4809 2571
rect 4861 2519 4862 2571
rect 4808 2512 4862 2519
rect 4908 2597 4962 2703
rect 5008 2781 5062 2788
rect 5008 2729 5009 2781
rect 5061 2729 5062 2781
rect 5008 2703 5018 2729
rect 5052 2703 5062 2729
rect 5008 2691 5062 2703
rect 5108 2737 5162 2843
rect 5208 2877 5262 2889
rect 5208 2851 5218 2877
rect 5252 2851 5262 2877
rect 5208 2799 5209 2851
rect 5261 2799 5262 2851
rect 5208 2792 5262 2799
rect 5308 2877 5362 2983
rect 5408 3061 5462 3068
rect 5408 3009 5409 3061
rect 5461 3009 5462 3061
rect 5408 2983 5418 3009
rect 5452 2983 5462 3009
rect 5408 2971 5462 2983
rect 5508 3017 5562 3123
rect 5608 3157 5662 3169
rect 5608 3131 5618 3157
rect 5652 3131 5662 3157
rect 5608 3079 5609 3131
rect 5661 3079 5662 3131
rect 5608 3072 5662 3079
rect 5708 3157 5762 3263
rect 5808 3341 5862 3348
rect 5808 3289 5809 3341
rect 5861 3289 5862 3341
rect 5808 3263 5818 3289
rect 5852 3263 5862 3289
rect 5808 3251 5862 3263
rect 5908 3297 5962 3403
rect 6008 3437 6062 3449
rect 6008 3411 6018 3437
rect 6052 3411 6062 3437
rect 6008 3359 6009 3411
rect 6061 3359 6062 3411
rect 6008 3352 6062 3359
rect 6108 3437 6162 3543
rect 6208 3621 6262 3628
rect 6208 3569 6209 3621
rect 6261 3569 6262 3621
rect 6208 3543 6218 3569
rect 6252 3543 6262 3569
rect 6208 3531 6262 3543
rect 6308 3577 6362 3773
rect 6408 3807 6462 3819
rect 6408 3781 6418 3807
rect 6452 3781 6462 3807
rect 6408 3729 6409 3781
rect 6461 3729 6462 3781
rect 6408 3722 6462 3729
rect 6506 3788 6516 3822
rect 6550 3788 6560 3822
rect 6506 3781 6560 3788
rect 6506 3729 6507 3781
rect 6559 3729 6560 3781
rect 6506 3722 6560 3729
rect 6590 3687 6620 4851
rect 6504 3681 6620 3687
rect 6504 3647 6516 3681
rect 6550 3647 6620 3681
rect 6504 3641 6620 3647
rect 6506 3592 6560 3604
rect 6308 3543 6318 3577
rect 6352 3543 6362 3577
rect 6108 3403 6118 3437
rect 6152 3403 6162 3437
rect 5908 3263 5918 3297
rect 5952 3263 5962 3297
rect 5708 3123 5718 3157
rect 5752 3123 5762 3157
rect 5508 2983 5518 3017
rect 5552 2983 5562 3017
rect 5308 2843 5318 2877
rect 5352 2843 5362 2877
rect 5108 2703 5118 2737
rect 5152 2703 5162 2737
rect 4908 2563 4918 2597
rect 4952 2563 4962 2597
rect 4802 2483 4868 2484
rect 4802 2431 4809 2483
rect 4861 2431 4868 2483
rect 4802 2430 4868 2431
rect 4708 2333 4718 2367
rect 4752 2333 4762 2367
rect 4508 2193 4518 2227
rect 4552 2193 4562 2227
rect 4308 2053 4318 2087
rect 4352 2053 4362 2087
rect 4108 1913 4118 1947
rect 4152 1913 4162 1947
rect 3908 1773 3918 1807
rect 3952 1773 3962 1807
rect 3708 1633 3718 1667
rect 3752 1633 3762 1667
rect 3508 1493 3518 1527
rect 3552 1493 3562 1527
rect 3308 1353 3318 1387
rect 3352 1353 3362 1387
rect 3202 1273 3268 1274
rect 3202 1221 3209 1273
rect 3261 1221 3268 1273
rect 3202 1220 3268 1221
rect 3108 1123 3118 1157
rect 3152 1123 3162 1157
rect 2908 983 2918 1017
rect 2952 983 2962 1017
rect 2708 843 2718 877
rect 2752 843 2762 877
rect 2508 703 2518 737
rect 2552 703 2562 737
rect 2308 563 2318 597
rect 2352 563 2362 597
rect 2108 423 2118 457
rect 2152 423 2162 457
rect 1908 283 1918 317
rect 1952 283 1962 317
rect 1708 143 1718 177
rect 1752 143 1762 177
rect 1602 63 1668 64
rect 1602 11 1609 63
rect 1661 11 1668 63
rect 1602 10 1668 11
rect 1508 -67 1509 -15
rect 1561 -67 1562 -15
rect 1508 -79 1518 -67
rect 1552 -79 1562 -67
rect 1308 -132 1362 -131
rect 1308 -143 1318 -132
rect 1352 -143 1362 -132
rect 1308 -195 1309 -143
rect 1361 -195 1362 -143
rect 1308 -210 1362 -195
rect 1412 -133 1458 -81
rect 1412 -167 1418 -133
rect 1452 -167 1458 -133
rect 1318 -291 1325 -239
rect 1377 -291 1384 -239
rect 1212 -397 1218 -363
rect 1252 -397 1258 -363
rect 1212 -435 1258 -397
rect 1212 -469 1218 -435
rect 1252 -469 1258 -435
rect 1212 -512 1258 -469
rect 1309 -326 1361 -320
rect 1309 -390 1318 -378
rect 1352 -390 1361 -378
rect 1309 -454 1318 -442
rect 1352 -454 1361 -442
rect 1309 -512 1361 -506
rect 1412 -363 1458 -167
rect 1508 -131 1509 -79
rect 1561 -131 1562 -79
rect 1608 -22 1662 10
rect 1608 -74 1609 -22
rect 1661 -74 1662 -22
rect 1608 -81 1662 -74
rect 1708 -15 1762 143
rect 1808 221 1862 228
rect 1808 169 1809 221
rect 1861 169 1862 221
rect 1808 143 1818 169
rect 1852 143 1862 169
rect 1808 131 1862 143
rect 1908 177 1962 283
rect 2008 317 2062 329
rect 2008 291 2018 317
rect 2052 291 2062 317
rect 2008 239 2009 291
rect 2061 239 2062 291
rect 2008 232 2062 239
rect 2108 317 2162 423
rect 2208 501 2262 508
rect 2208 449 2209 501
rect 2261 449 2262 501
rect 2208 423 2218 449
rect 2252 423 2262 449
rect 2208 411 2262 423
rect 2308 457 2362 563
rect 2408 597 2462 609
rect 2408 571 2418 597
rect 2452 571 2462 597
rect 2408 519 2409 571
rect 2461 519 2462 571
rect 2408 512 2462 519
rect 2508 597 2562 703
rect 2608 781 2662 788
rect 2608 729 2609 781
rect 2661 729 2662 781
rect 2608 703 2618 729
rect 2652 703 2662 729
rect 2608 691 2662 703
rect 2708 737 2762 843
rect 2808 877 2862 889
rect 2808 851 2818 877
rect 2852 851 2862 877
rect 2808 799 2809 851
rect 2861 799 2862 851
rect 2808 792 2862 799
rect 2908 877 2962 983
rect 3008 1061 3062 1068
rect 3008 1009 3009 1061
rect 3061 1009 3062 1061
rect 3008 983 3018 1009
rect 3052 983 3062 1009
rect 3008 971 3062 983
rect 3108 1017 3162 1123
rect 3208 1157 3262 1169
rect 3208 1131 3218 1157
rect 3252 1131 3262 1157
rect 3208 1079 3209 1131
rect 3261 1079 3262 1131
rect 3208 1072 3262 1079
rect 3308 1157 3362 1353
rect 3408 1431 3462 1438
rect 3408 1379 3409 1431
rect 3461 1379 3462 1431
rect 3408 1353 3418 1379
rect 3452 1353 3462 1379
rect 3408 1341 3462 1353
rect 3508 1387 3562 1493
rect 3608 1527 3662 1539
rect 3608 1501 3618 1527
rect 3652 1501 3662 1527
rect 3608 1449 3609 1501
rect 3661 1449 3662 1501
rect 3608 1442 3662 1449
rect 3708 1527 3762 1633
rect 3808 1711 3862 1718
rect 3808 1659 3809 1711
rect 3861 1659 3862 1711
rect 3808 1633 3818 1659
rect 3852 1633 3862 1659
rect 3808 1621 3862 1633
rect 3908 1667 3962 1773
rect 4008 1807 4062 1819
rect 4008 1781 4018 1807
rect 4052 1781 4062 1807
rect 4008 1729 4009 1781
rect 4061 1729 4062 1781
rect 4008 1722 4062 1729
rect 4108 1807 4162 1913
rect 4208 1991 4262 1998
rect 4208 1939 4209 1991
rect 4261 1939 4262 1991
rect 4208 1913 4218 1939
rect 4252 1913 4262 1939
rect 4208 1901 4262 1913
rect 4308 1947 4362 2053
rect 4408 2087 4462 2099
rect 4408 2061 4418 2087
rect 4452 2061 4462 2087
rect 4408 2009 4409 2061
rect 4461 2009 4462 2061
rect 4408 2002 4462 2009
rect 4508 2087 4562 2193
rect 4608 2271 4662 2278
rect 4608 2219 4609 2271
rect 4661 2219 4662 2271
rect 4608 2193 4618 2219
rect 4652 2193 4662 2219
rect 4608 2181 4662 2193
rect 4708 2227 4762 2333
rect 4808 2367 4862 2379
rect 4808 2341 4818 2367
rect 4852 2341 4862 2367
rect 4808 2289 4809 2341
rect 4861 2289 4862 2341
rect 4808 2282 4862 2289
rect 4908 2367 4962 2563
rect 5008 2641 5062 2648
rect 5008 2589 5009 2641
rect 5061 2589 5062 2641
rect 5008 2563 5018 2589
rect 5052 2563 5062 2589
rect 5008 2551 5062 2563
rect 5108 2597 5162 2703
rect 5208 2737 5262 2749
rect 5208 2711 5218 2737
rect 5252 2711 5262 2737
rect 5208 2659 5209 2711
rect 5261 2659 5262 2711
rect 5208 2652 5262 2659
rect 5308 2737 5362 2843
rect 5408 2921 5462 2928
rect 5408 2869 5409 2921
rect 5461 2869 5462 2921
rect 5408 2843 5418 2869
rect 5452 2843 5462 2869
rect 5408 2831 5462 2843
rect 5508 2877 5562 2983
rect 5608 3017 5662 3029
rect 5608 2991 5618 3017
rect 5652 2991 5662 3017
rect 5608 2939 5609 2991
rect 5661 2939 5662 2991
rect 5608 2932 5662 2939
rect 5708 3017 5762 3123
rect 5808 3201 5862 3208
rect 5808 3149 5809 3201
rect 5861 3149 5862 3201
rect 5808 3123 5818 3149
rect 5852 3123 5862 3149
rect 5808 3111 5862 3123
rect 5908 3157 5962 3263
rect 6008 3297 6062 3309
rect 6008 3271 6018 3297
rect 6052 3271 6062 3297
rect 6008 3219 6009 3271
rect 6061 3219 6062 3271
rect 6008 3212 6062 3219
rect 6108 3297 6162 3403
rect 6208 3481 6262 3488
rect 6208 3429 6209 3481
rect 6261 3429 6262 3481
rect 6208 3403 6218 3429
rect 6252 3403 6262 3429
rect 6208 3391 6262 3403
rect 6308 3437 6362 3543
rect 6408 3577 6462 3589
rect 6408 3551 6418 3577
rect 6452 3551 6462 3577
rect 6408 3499 6409 3551
rect 6461 3499 6462 3551
rect 6408 3492 6462 3499
rect 6506 3558 6516 3592
rect 6550 3558 6560 3592
rect 6506 3551 6560 3558
rect 6506 3499 6507 3551
rect 6559 3499 6560 3551
rect 6506 3492 6560 3499
rect 6506 3452 6560 3464
rect 6308 3403 6318 3437
rect 6352 3403 6362 3437
rect 6108 3263 6118 3297
rect 6152 3263 6162 3297
rect 5908 3123 5918 3157
rect 5952 3123 5962 3157
rect 5708 2983 5718 3017
rect 5752 2983 5762 3017
rect 5508 2843 5518 2877
rect 5552 2843 5562 2877
rect 5308 2703 5318 2737
rect 5352 2703 5362 2737
rect 5108 2563 5118 2597
rect 5152 2563 5162 2597
rect 5002 2499 5068 2500
rect 5002 2447 5009 2499
rect 5061 2447 5068 2499
rect 5002 2446 5068 2447
rect 4908 2333 4918 2367
rect 4952 2333 4962 2367
rect 4708 2193 4718 2227
rect 4752 2193 4762 2227
rect 4508 2053 4518 2087
rect 4552 2053 4562 2087
rect 4308 1913 4318 1947
rect 4352 1913 4362 1947
rect 4108 1773 4118 1807
rect 4152 1773 4162 1807
rect 3908 1633 3918 1667
rect 3952 1633 3962 1667
rect 3708 1493 3718 1527
rect 3752 1493 3762 1527
rect 3508 1353 3518 1387
rect 3552 1353 3562 1387
rect 3402 1289 3468 1290
rect 3402 1237 3409 1289
rect 3461 1237 3468 1289
rect 3402 1236 3468 1237
rect 3308 1123 3318 1157
rect 3352 1123 3362 1157
rect 3108 983 3118 1017
rect 3152 983 3162 1017
rect 2908 843 2918 877
rect 2952 843 2962 877
rect 2708 703 2718 737
rect 2752 703 2762 737
rect 2508 563 2518 597
rect 2552 563 2562 597
rect 2308 423 2318 457
rect 2352 423 2362 457
rect 2108 283 2118 317
rect 2152 283 2162 317
rect 1908 143 1918 177
rect 1952 143 1962 177
rect 1802 79 1868 80
rect 1802 27 1809 79
rect 1861 27 1868 79
rect 1802 26 1868 27
rect 1708 -67 1709 -15
rect 1761 -67 1762 -15
rect 1708 -79 1718 -67
rect 1752 -79 1762 -67
rect 1508 -132 1562 -131
rect 1508 -143 1518 -132
rect 1552 -143 1562 -132
rect 1508 -195 1509 -143
rect 1561 -195 1562 -143
rect 1508 -210 1562 -195
rect 1612 -133 1658 -81
rect 1612 -167 1618 -133
rect 1652 -167 1658 -133
rect 1518 -291 1525 -239
rect 1577 -291 1584 -239
rect 1412 -397 1418 -363
rect 1452 -397 1458 -363
rect 1412 -435 1458 -397
rect 1412 -469 1418 -435
rect 1452 -469 1458 -435
rect 1412 -512 1458 -469
rect 1509 -326 1561 -320
rect 1509 -390 1518 -378
rect 1552 -390 1561 -378
rect 1509 -454 1518 -442
rect 1552 -454 1561 -442
rect 1509 -555 1561 -506
rect 1612 -363 1658 -167
rect 1708 -131 1709 -79
rect 1761 -131 1762 -79
rect 1808 -22 1862 26
rect 1808 -74 1809 -22
rect 1861 -74 1862 -22
rect 1808 -81 1862 -74
rect 1908 -15 1962 143
rect 2008 177 2062 189
rect 2008 151 2018 177
rect 2052 151 2062 177
rect 2008 99 2009 151
rect 2061 99 2062 151
rect 2008 92 2062 99
rect 2108 177 2162 283
rect 2208 361 2262 368
rect 2208 309 2209 361
rect 2261 309 2262 361
rect 2208 283 2218 309
rect 2252 283 2262 309
rect 2208 271 2262 283
rect 2308 317 2362 423
rect 2408 457 2462 469
rect 2408 431 2418 457
rect 2452 431 2462 457
rect 2408 379 2409 431
rect 2461 379 2462 431
rect 2408 372 2462 379
rect 2508 457 2562 563
rect 2608 641 2662 648
rect 2608 589 2609 641
rect 2661 589 2662 641
rect 2608 563 2618 589
rect 2652 563 2662 589
rect 2608 551 2662 563
rect 2708 597 2762 703
rect 2808 737 2862 749
rect 2808 711 2818 737
rect 2852 711 2862 737
rect 2808 659 2809 711
rect 2861 659 2862 711
rect 2808 652 2862 659
rect 2908 737 2962 843
rect 3008 921 3062 928
rect 3008 869 3009 921
rect 3061 869 3062 921
rect 3008 843 3018 869
rect 3052 843 3062 869
rect 3008 831 3062 843
rect 3108 877 3162 983
rect 3208 1017 3262 1029
rect 3208 991 3218 1017
rect 3252 991 3262 1017
rect 3208 939 3209 991
rect 3261 939 3262 991
rect 3208 932 3262 939
rect 3308 1017 3362 1123
rect 3408 1201 3462 1208
rect 3408 1149 3409 1201
rect 3461 1149 3462 1201
rect 3408 1123 3418 1149
rect 3452 1123 3462 1149
rect 3408 1111 3462 1123
rect 3508 1157 3562 1353
rect 3608 1387 3662 1399
rect 3608 1361 3618 1387
rect 3652 1361 3662 1387
rect 3608 1309 3609 1361
rect 3661 1309 3662 1361
rect 3608 1302 3662 1309
rect 3708 1387 3762 1493
rect 3808 1571 3862 1578
rect 3808 1519 3809 1571
rect 3861 1519 3862 1571
rect 3808 1493 3818 1519
rect 3852 1493 3862 1519
rect 3808 1481 3862 1493
rect 3908 1527 3962 1633
rect 4008 1667 4062 1679
rect 4008 1641 4018 1667
rect 4052 1641 4062 1667
rect 4008 1589 4009 1641
rect 4061 1589 4062 1641
rect 4008 1582 4062 1589
rect 4108 1667 4162 1773
rect 4208 1851 4262 1858
rect 4208 1799 4209 1851
rect 4261 1799 4262 1851
rect 4208 1773 4218 1799
rect 4252 1773 4262 1799
rect 4208 1761 4262 1773
rect 4308 1807 4362 1913
rect 4408 1947 4462 1959
rect 4408 1921 4418 1947
rect 4452 1921 4462 1947
rect 4408 1869 4409 1921
rect 4461 1869 4462 1921
rect 4408 1862 4462 1869
rect 4508 1947 4562 2053
rect 4608 2131 4662 2138
rect 4608 2079 4609 2131
rect 4661 2079 4662 2131
rect 4608 2053 4618 2079
rect 4652 2053 4662 2079
rect 4608 2041 4662 2053
rect 4708 2087 4762 2193
rect 4808 2227 4862 2239
rect 4808 2201 4818 2227
rect 4852 2201 4862 2227
rect 4808 2149 4809 2201
rect 4861 2149 4862 2201
rect 4808 2142 4862 2149
rect 4908 2227 4962 2333
rect 5008 2411 5062 2418
rect 5008 2359 5009 2411
rect 5061 2359 5062 2411
rect 5008 2333 5018 2359
rect 5052 2333 5062 2359
rect 5008 2321 5062 2333
rect 5108 2367 5162 2563
rect 5208 2597 5262 2609
rect 5208 2571 5218 2597
rect 5252 2571 5262 2597
rect 5208 2519 5209 2571
rect 5261 2519 5262 2571
rect 5208 2512 5262 2519
rect 5308 2597 5362 2703
rect 5408 2781 5462 2788
rect 5408 2729 5409 2781
rect 5461 2729 5462 2781
rect 5408 2703 5418 2729
rect 5452 2703 5462 2729
rect 5408 2691 5462 2703
rect 5508 2737 5562 2843
rect 5608 2877 5662 2889
rect 5608 2851 5618 2877
rect 5652 2851 5662 2877
rect 5608 2799 5609 2851
rect 5661 2799 5662 2851
rect 5608 2792 5662 2799
rect 5708 2877 5762 2983
rect 5808 3061 5862 3068
rect 5808 3009 5809 3061
rect 5861 3009 5862 3061
rect 5808 2983 5818 3009
rect 5852 2983 5862 3009
rect 5808 2971 5862 2983
rect 5908 3017 5962 3123
rect 6008 3157 6062 3169
rect 6008 3131 6018 3157
rect 6052 3131 6062 3157
rect 6008 3079 6009 3131
rect 6061 3079 6062 3131
rect 6008 3072 6062 3079
rect 6108 3157 6162 3263
rect 6208 3341 6262 3348
rect 6208 3289 6209 3341
rect 6261 3289 6262 3341
rect 6208 3263 6218 3289
rect 6252 3263 6262 3289
rect 6208 3251 6262 3263
rect 6308 3297 6362 3403
rect 6408 3437 6462 3449
rect 6408 3411 6418 3437
rect 6452 3411 6462 3437
rect 6408 3359 6409 3411
rect 6461 3359 6462 3411
rect 6408 3352 6462 3359
rect 6506 3418 6516 3452
rect 6550 3418 6560 3452
rect 6506 3411 6560 3418
rect 6506 3359 6507 3411
rect 6559 3359 6560 3411
rect 6506 3352 6560 3359
rect 6506 3312 6560 3324
rect 6308 3263 6318 3297
rect 6352 3263 6362 3297
rect 6108 3123 6118 3157
rect 6152 3123 6162 3157
rect 5908 2983 5918 3017
rect 5952 2983 5962 3017
rect 5708 2843 5718 2877
rect 5752 2843 5762 2877
rect 5508 2703 5518 2737
rect 5552 2703 5562 2737
rect 5308 2563 5318 2597
rect 5352 2563 5362 2597
rect 5202 2483 5268 2484
rect 5202 2431 5209 2483
rect 5261 2431 5268 2483
rect 5202 2430 5268 2431
rect 5108 2333 5118 2367
rect 5152 2333 5162 2367
rect 4908 2193 4918 2227
rect 4952 2193 4962 2227
rect 4708 2053 4718 2087
rect 4752 2053 4762 2087
rect 4508 1913 4518 1947
rect 4552 1913 4562 1947
rect 4308 1773 4318 1807
rect 4352 1773 4362 1807
rect 4108 1633 4118 1667
rect 4152 1633 4162 1667
rect 3908 1493 3918 1527
rect 3952 1493 3962 1527
rect 3708 1353 3718 1387
rect 3752 1353 3762 1387
rect 3602 1273 3668 1274
rect 3602 1221 3609 1273
rect 3661 1221 3668 1273
rect 3602 1220 3668 1221
rect 3508 1123 3518 1157
rect 3552 1123 3562 1157
rect 3308 983 3318 1017
rect 3352 983 3362 1017
rect 3108 843 3118 877
rect 3152 843 3162 877
rect 2908 703 2918 737
rect 2952 703 2962 737
rect 2708 563 2718 597
rect 2752 563 2762 597
rect 2508 423 2518 457
rect 2552 423 2562 457
rect 2308 283 2318 317
rect 2352 283 2362 317
rect 2108 143 2118 177
rect 2152 143 2162 177
rect 2002 63 2068 64
rect 2002 11 2009 63
rect 2061 11 2068 63
rect 2002 10 2068 11
rect 1908 -67 1909 -15
rect 1961 -67 1962 -15
rect 1908 -79 1918 -67
rect 1952 -79 1962 -67
rect 1708 -132 1762 -131
rect 1708 -143 1718 -132
rect 1752 -143 1762 -132
rect 1708 -195 1709 -143
rect 1761 -195 1762 -143
rect 1708 -210 1762 -195
rect 1812 -133 1858 -81
rect 1812 -167 1818 -133
rect 1852 -167 1858 -133
rect 1718 -291 1725 -239
rect 1777 -291 1784 -239
rect 1612 -397 1618 -363
rect 1652 -397 1658 -363
rect 1612 -435 1658 -397
rect 1612 -469 1618 -435
rect 1652 -469 1658 -435
rect 1612 -512 1658 -469
rect 1709 -326 1761 -320
rect 1709 -390 1718 -378
rect 1752 -390 1761 -378
rect 1709 -454 1718 -442
rect 1752 -454 1761 -442
rect 1709 -512 1761 -506
rect 1812 -363 1858 -167
rect 1908 -131 1909 -79
rect 1961 -131 1962 -79
rect 2008 -22 2062 10
rect 2008 -74 2009 -22
rect 2061 -74 2062 -22
rect 2008 -81 2062 -74
rect 2108 -15 2162 143
rect 2208 221 2262 228
rect 2208 169 2209 221
rect 2261 169 2262 221
rect 2208 143 2218 169
rect 2252 143 2262 169
rect 2208 131 2262 143
rect 2308 177 2362 283
rect 2408 317 2462 329
rect 2408 291 2418 317
rect 2452 291 2462 317
rect 2408 239 2409 291
rect 2461 239 2462 291
rect 2408 232 2462 239
rect 2508 317 2562 423
rect 2608 501 2662 508
rect 2608 449 2609 501
rect 2661 449 2662 501
rect 2608 423 2618 449
rect 2652 423 2662 449
rect 2608 411 2662 423
rect 2708 457 2762 563
rect 2808 597 2862 609
rect 2808 571 2818 597
rect 2852 571 2862 597
rect 2808 519 2809 571
rect 2861 519 2862 571
rect 2808 512 2862 519
rect 2908 597 2962 703
rect 3008 781 3062 788
rect 3008 729 3009 781
rect 3061 729 3062 781
rect 3008 703 3018 729
rect 3052 703 3062 729
rect 3008 691 3062 703
rect 3108 737 3162 843
rect 3208 877 3262 889
rect 3208 851 3218 877
rect 3252 851 3262 877
rect 3208 799 3209 851
rect 3261 799 3262 851
rect 3208 792 3262 799
rect 3308 877 3362 983
rect 3408 1061 3462 1068
rect 3408 1009 3409 1061
rect 3461 1009 3462 1061
rect 3408 983 3418 1009
rect 3452 983 3462 1009
rect 3408 971 3462 983
rect 3508 1017 3562 1123
rect 3608 1157 3662 1169
rect 3608 1131 3618 1157
rect 3652 1131 3662 1157
rect 3608 1079 3609 1131
rect 3661 1079 3662 1131
rect 3608 1072 3662 1079
rect 3708 1157 3762 1353
rect 3808 1431 3862 1438
rect 3808 1379 3809 1431
rect 3861 1379 3862 1431
rect 3808 1353 3818 1379
rect 3852 1353 3862 1379
rect 3808 1341 3862 1353
rect 3908 1387 3962 1493
rect 4008 1527 4062 1539
rect 4008 1501 4018 1527
rect 4052 1501 4062 1527
rect 4008 1449 4009 1501
rect 4061 1449 4062 1501
rect 4008 1442 4062 1449
rect 4108 1527 4162 1633
rect 4208 1711 4262 1718
rect 4208 1659 4209 1711
rect 4261 1659 4262 1711
rect 4208 1633 4218 1659
rect 4252 1633 4262 1659
rect 4208 1621 4262 1633
rect 4308 1667 4362 1773
rect 4408 1807 4462 1819
rect 4408 1781 4418 1807
rect 4452 1781 4462 1807
rect 4408 1729 4409 1781
rect 4461 1729 4462 1781
rect 4408 1722 4462 1729
rect 4508 1807 4562 1913
rect 4608 1991 4662 1998
rect 4608 1939 4609 1991
rect 4661 1939 4662 1991
rect 4608 1913 4618 1939
rect 4652 1913 4662 1939
rect 4608 1901 4662 1913
rect 4708 1947 4762 2053
rect 4808 2087 4862 2099
rect 4808 2061 4818 2087
rect 4852 2061 4862 2087
rect 4808 2009 4809 2061
rect 4861 2009 4862 2061
rect 4808 2002 4862 2009
rect 4908 2087 4962 2193
rect 5008 2271 5062 2278
rect 5008 2219 5009 2271
rect 5061 2219 5062 2271
rect 5008 2193 5018 2219
rect 5052 2193 5062 2219
rect 5008 2181 5062 2193
rect 5108 2227 5162 2333
rect 5208 2367 5262 2379
rect 5208 2341 5218 2367
rect 5252 2341 5262 2367
rect 5208 2289 5209 2341
rect 5261 2289 5262 2341
rect 5208 2282 5262 2289
rect 5308 2367 5362 2563
rect 5408 2641 5462 2648
rect 5408 2589 5409 2641
rect 5461 2589 5462 2641
rect 5408 2563 5418 2589
rect 5452 2563 5462 2589
rect 5408 2551 5462 2563
rect 5508 2597 5562 2703
rect 5608 2737 5662 2749
rect 5608 2711 5618 2737
rect 5652 2711 5662 2737
rect 5608 2659 5609 2711
rect 5661 2659 5662 2711
rect 5608 2652 5662 2659
rect 5708 2737 5762 2843
rect 5808 2921 5862 2928
rect 5808 2869 5809 2921
rect 5861 2869 5862 2921
rect 5808 2843 5818 2869
rect 5852 2843 5862 2869
rect 5808 2831 5862 2843
rect 5908 2877 5962 2983
rect 6008 3017 6062 3029
rect 6008 2991 6018 3017
rect 6052 2991 6062 3017
rect 6008 2939 6009 2991
rect 6061 2939 6062 2991
rect 6008 2932 6062 2939
rect 6108 3017 6162 3123
rect 6208 3201 6262 3208
rect 6208 3149 6209 3201
rect 6261 3149 6262 3201
rect 6208 3123 6218 3149
rect 6252 3123 6262 3149
rect 6208 3111 6262 3123
rect 6308 3157 6362 3263
rect 6408 3297 6462 3309
rect 6408 3271 6418 3297
rect 6452 3271 6462 3297
rect 6408 3219 6409 3271
rect 6461 3219 6462 3271
rect 6408 3212 6462 3219
rect 6506 3278 6516 3312
rect 6550 3278 6560 3312
rect 6506 3271 6560 3278
rect 6506 3219 6507 3271
rect 6559 3219 6560 3271
rect 6506 3212 6560 3219
rect 6506 3172 6560 3184
rect 6308 3123 6318 3157
rect 6352 3123 6362 3157
rect 6108 2983 6118 3017
rect 6152 2983 6162 3017
rect 5908 2843 5918 2877
rect 5952 2843 5962 2877
rect 5708 2703 5718 2737
rect 5752 2703 5762 2737
rect 5508 2563 5518 2597
rect 5552 2563 5562 2597
rect 5402 2499 5468 2500
rect 5402 2447 5409 2499
rect 5461 2447 5468 2499
rect 5402 2446 5468 2447
rect 5308 2333 5318 2367
rect 5352 2333 5362 2367
rect 5108 2193 5118 2227
rect 5152 2193 5162 2227
rect 4908 2053 4918 2087
rect 4952 2053 4962 2087
rect 4708 1913 4718 1947
rect 4752 1913 4762 1947
rect 4508 1773 4518 1807
rect 4552 1773 4562 1807
rect 4308 1633 4318 1667
rect 4352 1633 4362 1667
rect 4108 1493 4118 1527
rect 4152 1493 4162 1527
rect 3908 1353 3918 1387
rect 3952 1353 3962 1387
rect 3802 1289 3868 1290
rect 3802 1237 3809 1289
rect 3861 1237 3868 1289
rect 3802 1236 3868 1237
rect 3708 1123 3718 1157
rect 3752 1123 3762 1157
rect 3508 983 3518 1017
rect 3552 983 3562 1017
rect 3308 843 3318 877
rect 3352 843 3362 877
rect 3108 703 3118 737
rect 3152 703 3162 737
rect 2908 563 2918 597
rect 2952 563 2962 597
rect 2708 423 2718 457
rect 2752 423 2762 457
rect 2508 283 2518 317
rect 2552 283 2562 317
rect 2308 143 2318 177
rect 2352 143 2362 177
rect 2202 79 2268 80
rect 2202 27 2209 79
rect 2261 27 2268 79
rect 2202 26 2268 27
rect 2108 -67 2109 -15
rect 2161 -67 2162 -15
rect 2108 -79 2118 -67
rect 2152 -79 2162 -67
rect 1908 -132 1962 -131
rect 1908 -143 1918 -132
rect 1952 -143 1962 -132
rect 1908 -195 1909 -143
rect 1961 -195 1962 -143
rect 1908 -210 1962 -195
rect 2012 -133 2058 -81
rect 2012 -167 2018 -133
rect 2052 -167 2058 -133
rect 1918 -291 1925 -239
rect 1977 -291 1984 -239
rect 1812 -397 1818 -363
rect 1852 -397 1858 -363
rect 1812 -435 1858 -397
rect 1812 -469 1818 -435
rect 1852 -469 1858 -435
rect 1812 -512 1858 -469
rect 1909 -326 1961 -320
rect 1909 -390 1918 -378
rect 1952 -390 1961 -378
rect 1909 -454 1918 -442
rect 1952 -454 1961 -442
rect 1909 -555 1961 -506
rect 2012 -363 2058 -167
rect 2108 -131 2109 -79
rect 2161 -131 2162 -79
rect 2208 -22 2262 26
rect 2208 -74 2209 -22
rect 2261 -74 2262 -22
rect 2208 -81 2262 -74
rect 2308 -15 2362 143
rect 2408 177 2462 189
rect 2408 151 2418 177
rect 2452 151 2462 177
rect 2408 99 2409 151
rect 2461 99 2462 151
rect 2408 92 2462 99
rect 2508 177 2562 283
rect 2608 361 2662 368
rect 2608 309 2609 361
rect 2661 309 2662 361
rect 2608 283 2618 309
rect 2652 283 2662 309
rect 2608 271 2662 283
rect 2708 317 2762 423
rect 2808 457 2862 469
rect 2808 431 2818 457
rect 2852 431 2862 457
rect 2808 379 2809 431
rect 2861 379 2862 431
rect 2808 372 2862 379
rect 2908 457 2962 563
rect 3008 641 3062 648
rect 3008 589 3009 641
rect 3061 589 3062 641
rect 3008 563 3018 589
rect 3052 563 3062 589
rect 3008 551 3062 563
rect 3108 597 3162 703
rect 3208 737 3262 749
rect 3208 711 3218 737
rect 3252 711 3262 737
rect 3208 659 3209 711
rect 3261 659 3262 711
rect 3208 652 3262 659
rect 3308 737 3362 843
rect 3408 921 3462 928
rect 3408 869 3409 921
rect 3461 869 3462 921
rect 3408 843 3418 869
rect 3452 843 3462 869
rect 3408 831 3462 843
rect 3508 877 3562 983
rect 3608 1017 3662 1029
rect 3608 991 3618 1017
rect 3652 991 3662 1017
rect 3608 939 3609 991
rect 3661 939 3662 991
rect 3608 932 3662 939
rect 3708 1017 3762 1123
rect 3808 1201 3862 1208
rect 3808 1149 3809 1201
rect 3861 1149 3862 1201
rect 3808 1123 3818 1149
rect 3852 1123 3862 1149
rect 3808 1111 3862 1123
rect 3908 1157 3962 1353
rect 4008 1387 4062 1399
rect 4008 1361 4018 1387
rect 4052 1361 4062 1387
rect 4008 1309 4009 1361
rect 4061 1309 4062 1361
rect 4008 1302 4062 1309
rect 4108 1387 4162 1493
rect 4208 1571 4262 1578
rect 4208 1519 4209 1571
rect 4261 1519 4262 1571
rect 4208 1493 4218 1519
rect 4252 1493 4262 1519
rect 4208 1481 4262 1493
rect 4308 1527 4362 1633
rect 4408 1667 4462 1679
rect 4408 1641 4418 1667
rect 4452 1641 4462 1667
rect 4408 1589 4409 1641
rect 4461 1589 4462 1641
rect 4408 1582 4462 1589
rect 4508 1667 4562 1773
rect 4608 1851 4662 1858
rect 4608 1799 4609 1851
rect 4661 1799 4662 1851
rect 4608 1773 4618 1799
rect 4652 1773 4662 1799
rect 4608 1761 4662 1773
rect 4708 1807 4762 1913
rect 4808 1947 4862 1959
rect 4808 1921 4818 1947
rect 4852 1921 4862 1947
rect 4808 1869 4809 1921
rect 4861 1869 4862 1921
rect 4808 1862 4862 1869
rect 4908 1947 4962 2053
rect 5008 2131 5062 2138
rect 5008 2079 5009 2131
rect 5061 2079 5062 2131
rect 5008 2053 5018 2079
rect 5052 2053 5062 2079
rect 5008 2041 5062 2053
rect 5108 2087 5162 2193
rect 5208 2227 5262 2239
rect 5208 2201 5218 2227
rect 5252 2201 5262 2227
rect 5208 2149 5209 2201
rect 5261 2149 5262 2201
rect 5208 2142 5262 2149
rect 5308 2227 5362 2333
rect 5408 2411 5462 2418
rect 5408 2359 5409 2411
rect 5461 2359 5462 2411
rect 5408 2333 5418 2359
rect 5452 2333 5462 2359
rect 5408 2321 5462 2333
rect 5508 2367 5562 2563
rect 5608 2597 5662 2609
rect 5608 2571 5618 2597
rect 5652 2571 5662 2597
rect 5608 2519 5609 2571
rect 5661 2519 5662 2571
rect 5608 2512 5662 2519
rect 5708 2597 5762 2703
rect 5808 2781 5862 2788
rect 5808 2729 5809 2781
rect 5861 2729 5862 2781
rect 5808 2703 5818 2729
rect 5852 2703 5862 2729
rect 5808 2691 5862 2703
rect 5908 2737 5962 2843
rect 6008 2877 6062 2889
rect 6008 2851 6018 2877
rect 6052 2851 6062 2877
rect 6008 2799 6009 2851
rect 6061 2799 6062 2851
rect 6008 2792 6062 2799
rect 6108 2877 6162 2983
rect 6208 3061 6262 3068
rect 6208 3009 6209 3061
rect 6261 3009 6262 3061
rect 6208 2983 6218 3009
rect 6252 2983 6262 3009
rect 6208 2971 6262 2983
rect 6308 3017 6362 3123
rect 6408 3157 6462 3169
rect 6408 3131 6418 3157
rect 6452 3131 6462 3157
rect 6408 3079 6409 3131
rect 6461 3079 6462 3131
rect 6408 3072 6462 3079
rect 6506 3138 6516 3172
rect 6550 3138 6560 3172
rect 6506 3131 6560 3138
rect 6506 3079 6507 3131
rect 6559 3079 6560 3131
rect 6506 3072 6560 3079
rect 6506 3032 6560 3044
rect 6308 2983 6318 3017
rect 6352 2983 6362 3017
rect 6108 2843 6118 2877
rect 6152 2843 6162 2877
rect 5908 2703 5918 2737
rect 5952 2703 5962 2737
rect 5708 2563 5718 2597
rect 5752 2563 5762 2597
rect 5602 2483 5668 2484
rect 5602 2431 5609 2483
rect 5661 2431 5668 2483
rect 5602 2430 5668 2431
rect 5508 2333 5518 2367
rect 5552 2333 5562 2367
rect 5308 2193 5318 2227
rect 5352 2193 5362 2227
rect 5108 2053 5118 2087
rect 5152 2053 5162 2087
rect 4908 1913 4918 1947
rect 4952 1913 4962 1947
rect 4708 1773 4718 1807
rect 4752 1773 4762 1807
rect 4508 1633 4518 1667
rect 4552 1633 4562 1667
rect 4308 1493 4318 1527
rect 4352 1493 4362 1527
rect 4108 1353 4118 1387
rect 4152 1353 4162 1387
rect 4002 1273 4068 1274
rect 4002 1221 4009 1273
rect 4061 1221 4068 1273
rect 4002 1220 4068 1221
rect 3908 1123 3918 1157
rect 3952 1123 3962 1157
rect 3708 983 3718 1017
rect 3752 983 3762 1017
rect 3508 843 3518 877
rect 3552 843 3562 877
rect 3308 703 3318 737
rect 3352 703 3362 737
rect 3108 563 3118 597
rect 3152 563 3162 597
rect 2908 423 2918 457
rect 2952 423 2962 457
rect 2708 283 2718 317
rect 2752 283 2762 317
rect 2508 143 2518 177
rect 2552 143 2562 177
rect 2402 63 2468 64
rect 2402 11 2409 63
rect 2461 11 2468 63
rect 2402 10 2468 11
rect 2308 -67 2309 -15
rect 2361 -67 2362 -15
rect 2308 -79 2318 -67
rect 2352 -79 2362 -67
rect 2108 -132 2162 -131
rect 2108 -143 2118 -132
rect 2152 -143 2162 -132
rect 2108 -195 2109 -143
rect 2161 -195 2162 -143
rect 2108 -210 2162 -195
rect 2212 -133 2258 -81
rect 2212 -167 2218 -133
rect 2252 -167 2258 -133
rect 2118 -291 2125 -239
rect 2177 -291 2184 -239
rect 2012 -397 2018 -363
rect 2052 -397 2058 -363
rect 2012 -435 2058 -397
rect 2012 -469 2018 -435
rect 2052 -469 2058 -435
rect 2012 -512 2058 -469
rect 2109 -326 2161 -320
rect 2109 -390 2118 -378
rect 2152 -390 2161 -378
rect 2109 -454 2118 -442
rect 2152 -454 2161 -442
rect 2109 -512 2161 -506
rect 2212 -363 2258 -167
rect 2308 -131 2309 -79
rect 2361 -131 2362 -79
rect 2408 -22 2462 10
rect 2408 -74 2409 -22
rect 2461 -74 2462 -22
rect 2408 -81 2462 -74
rect 2508 -15 2562 143
rect 2608 221 2662 228
rect 2608 169 2609 221
rect 2661 169 2662 221
rect 2608 143 2618 169
rect 2652 143 2662 169
rect 2608 131 2662 143
rect 2708 177 2762 283
rect 2808 317 2862 329
rect 2808 291 2818 317
rect 2852 291 2862 317
rect 2808 239 2809 291
rect 2861 239 2862 291
rect 2808 232 2862 239
rect 2908 317 2962 423
rect 3008 501 3062 508
rect 3008 449 3009 501
rect 3061 449 3062 501
rect 3008 423 3018 449
rect 3052 423 3062 449
rect 3008 411 3062 423
rect 3108 457 3162 563
rect 3208 597 3262 609
rect 3208 571 3218 597
rect 3252 571 3262 597
rect 3208 519 3209 571
rect 3261 519 3262 571
rect 3208 512 3262 519
rect 3308 597 3362 703
rect 3408 781 3462 788
rect 3408 729 3409 781
rect 3461 729 3462 781
rect 3408 703 3418 729
rect 3452 703 3462 729
rect 3408 691 3462 703
rect 3508 737 3562 843
rect 3608 877 3662 889
rect 3608 851 3618 877
rect 3652 851 3662 877
rect 3608 799 3609 851
rect 3661 799 3662 851
rect 3608 792 3662 799
rect 3708 877 3762 983
rect 3808 1061 3862 1068
rect 3808 1009 3809 1061
rect 3861 1009 3862 1061
rect 3808 983 3818 1009
rect 3852 983 3862 1009
rect 3808 971 3862 983
rect 3908 1017 3962 1123
rect 4008 1157 4062 1169
rect 4008 1131 4018 1157
rect 4052 1131 4062 1157
rect 4008 1079 4009 1131
rect 4061 1079 4062 1131
rect 4008 1072 4062 1079
rect 4108 1157 4162 1353
rect 4208 1431 4262 1438
rect 4208 1379 4209 1431
rect 4261 1379 4262 1431
rect 4208 1353 4218 1379
rect 4252 1353 4262 1379
rect 4208 1341 4262 1353
rect 4308 1387 4362 1493
rect 4408 1527 4462 1539
rect 4408 1501 4418 1527
rect 4452 1501 4462 1527
rect 4408 1449 4409 1501
rect 4461 1449 4462 1501
rect 4408 1442 4462 1449
rect 4508 1527 4562 1633
rect 4608 1711 4662 1718
rect 4608 1659 4609 1711
rect 4661 1659 4662 1711
rect 4608 1633 4618 1659
rect 4652 1633 4662 1659
rect 4608 1621 4662 1633
rect 4708 1667 4762 1773
rect 4808 1807 4862 1819
rect 4808 1781 4818 1807
rect 4852 1781 4862 1807
rect 4808 1729 4809 1781
rect 4861 1729 4862 1781
rect 4808 1722 4862 1729
rect 4908 1807 4962 1913
rect 5008 1991 5062 1998
rect 5008 1939 5009 1991
rect 5061 1939 5062 1991
rect 5008 1913 5018 1939
rect 5052 1913 5062 1939
rect 5008 1901 5062 1913
rect 5108 1947 5162 2053
rect 5208 2087 5262 2099
rect 5208 2061 5218 2087
rect 5252 2061 5262 2087
rect 5208 2009 5209 2061
rect 5261 2009 5262 2061
rect 5208 2002 5262 2009
rect 5308 2087 5362 2193
rect 5408 2271 5462 2278
rect 5408 2219 5409 2271
rect 5461 2219 5462 2271
rect 5408 2193 5418 2219
rect 5452 2193 5462 2219
rect 5408 2181 5462 2193
rect 5508 2227 5562 2333
rect 5608 2367 5662 2379
rect 5608 2341 5618 2367
rect 5652 2341 5662 2367
rect 5608 2289 5609 2341
rect 5661 2289 5662 2341
rect 5608 2282 5662 2289
rect 5708 2367 5762 2563
rect 5808 2641 5862 2648
rect 5808 2589 5809 2641
rect 5861 2589 5862 2641
rect 5808 2563 5818 2589
rect 5852 2563 5862 2589
rect 5808 2551 5862 2563
rect 5908 2597 5962 2703
rect 6008 2737 6062 2749
rect 6008 2711 6018 2737
rect 6052 2711 6062 2737
rect 6008 2659 6009 2711
rect 6061 2659 6062 2711
rect 6008 2652 6062 2659
rect 6108 2737 6162 2843
rect 6208 2921 6262 2928
rect 6208 2869 6209 2921
rect 6261 2869 6262 2921
rect 6208 2843 6218 2869
rect 6252 2843 6262 2869
rect 6208 2831 6262 2843
rect 6308 2877 6362 2983
rect 6408 3017 6462 3029
rect 6408 2991 6418 3017
rect 6452 2991 6462 3017
rect 6408 2939 6409 2991
rect 6461 2939 6462 2991
rect 6408 2932 6462 2939
rect 6506 2998 6516 3032
rect 6550 2998 6560 3032
rect 6506 2991 6560 2998
rect 6506 2939 6507 2991
rect 6559 2939 6560 2991
rect 6506 2932 6560 2939
rect 6506 2892 6560 2904
rect 6308 2843 6318 2877
rect 6352 2843 6362 2877
rect 6108 2703 6118 2737
rect 6152 2703 6162 2737
rect 5908 2563 5918 2597
rect 5952 2563 5962 2597
rect 5802 2499 5868 2500
rect 5802 2447 5809 2499
rect 5861 2447 5868 2499
rect 5802 2446 5868 2447
rect 5708 2333 5718 2367
rect 5752 2333 5762 2367
rect 5508 2193 5518 2227
rect 5552 2193 5562 2227
rect 5308 2053 5318 2087
rect 5352 2053 5362 2087
rect 5108 1913 5118 1947
rect 5152 1913 5162 1947
rect 4908 1773 4918 1807
rect 4952 1773 4962 1807
rect 4708 1633 4718 1667
rect 4752 1633 4762 1667
rect 4508 1493 4518 1527
rect 4552 1493 4562 1527
rect 4308 1353 4318 1387
rect 4352 1353 4362 1387
rect 4202 1289 4268 1290
rect 4202 1237 4209 1289
rect 4261 1237 4268 1289
rect 4202 1236 4268 1237
rect 4108 1123 4118 1157
rect 4152 1123 4162 1157
rect 3908 983 3918 1017
rect 3952 983 3962 1017
rect 3708 843 3718 877
rect 3752 843 3762 877
rect 3508 703 3518 737
rect 3552 703 3562 737
rect 3308 563 3318 597
rect 3352 563 3362 597
rect 3108 423 3118 457
rect 3152 423 3162 457
rect 2908 283 2918 317
rect 2952 283 2962 317
rect 2708 143 2718 177
rect 2752 143 2762 177
rect 2602 79 2668 80
rect 2602 27 2609 79
rect 2661 27 2668 79
rect 2602 26 2668 27
rect 2508 -67 2509 -15
rect 2561 -67 2562 -15
rect 2508 -79 2518 -67
rect 2552 -79 2562 -67
rect 2308 -132 2362 -131
rect 2308 -143 2318 -132
rect 2352 -143 2362 -132
rect 2308 -195 2309 -143
rect 2361 -195 2362 -143
rect 2308 -210 2362 -195
rect 2412 -133 2458 -81
rect 2412 -167 2418 -133
rect 2452 -167 2458 -133
rect 2318 -291 2325 -239
rect 2377 -291 2384 -239
rect 2212 -397 2218 -363
rect 2252 -397 2258 -363
rect 2212 -435 2258 -397
rect 2212 -469 2218 -435
rect 2252 -469 2258 -435
rect 2212 -512 2258 -469
rect 2309 -326 2361 -320
rect 2309 -390 2318 -378
rect 2352 -390 2361 -378
rect 2309 -454 2318 -442
rect 2352 -454 2361 -442
rect 2309 -555 2361 -506
rect 2412 -363 2458 -167
rect 2508 -131 2509 -79
rect 2561 -131 2562 -79
rect 2608 -22 2662 26
rect 2608 -74 2609 -22
rect 2661 -74 2662 -22
rect 2608 -81 2662 -74
rect 2708 -15 2762 143
rect 2808 177 2862 189
rect 2808 151 2818 177
rect 2852 151 2862 177
rect 2808 99 2809 151
rect 2861 99 2862 151
rect 2808 92 2862 99
rect 2908 177 2962 283
rect 3008 361 3062 368
rect 3008 309 3009 361
rect 3061 309 3062 361
rect 3008 283 3018 309
rect 3052 283 3062 309
rect 3008 271 3062 283
rect 3108 317 3162 423
rect 3208 457 3262 469
rect 3208 431 3218 457
rect 3252 431 3262 457
rect 3208 379 3209 431
rect 3261 379 3262 431
rect 3208 372 3262 379
rect 3308 457 3362 563
rect 3408 641 3462 648
rect 3408 589 3409 641
rect 3461 589 3462 641
rect 3408 563 3418 589
rect 3452 563 3462 589
rect 3408 551 3462 563
rect 3508 597 3562 703
rect 3608 737 3662 749
rect 3608 711 3618 737
rect 3652 711 3662 737
rect 3608 659 3609 711
rect 3661 659 3662 711
rect 3608 652 3662 659
rect 3708 737 3762 843
rect 3808 921 3862 928
rect 3808 869 3809 921
rect 3861 869 3862 921
rect 3808 843 3818 869
rect 3852 843 3862 869
rect 3808 831 3862 843
rect 3908 877 3962 983
rect 4008 1017 4062 1029
rect 4008 991 4018 1017
rect 4052 991 4062 1017
rect 4008 939 4009 991
rect 4061 939 4062 991
rect 4008 932 4062 939
rect 4108 1017 4162 1123
rect 4208 1201 4262 1208
rect 4208 1149 4209 1201
rect 4261 1149 4262 1201
rect 4208 1123 4218 1149
rect 4252 1123 4262 1149
rect 4208 1111 4262 1123
rect 4308 1157 4362 1353
rect 4408 1387 4462 1399
rect 4408 1361 4418 1387
rect 4452 1361 4462 1387
rect 4408 1309 4409 1361
rect 4461 1309 4462 1361
rect 4408 1302 4462 1309
rect 4508 1387 4562 1493
rect 4608 1571 4662 1578
rect 4608 1519 4609 1571
rect 4661 1519 4662 1571
rect 4608 1493 4618 1519
rect 4652 1493 4662 1519
rect 4608 1481 4662 1493
rect 4708 1527 4762 1633
rect 4808 1667 4862 1679
rect 4808 1641 4818 1667
rect 4852 1641 4862 1667
rect 4808 1589 4809 1641
rect 4861 1589 4862 1641
rect 4808 1582 4862 1589
rect 4908 1667 4962 1773
rect 5008 1851 5062 1858
rect 5008 1799 5009 1851
rect 5061 1799 5062 1851
rect 5008 1773 5018 1799
rect 5052 1773 5062 1799
rect 5008 1761 5062 1773
rect 5108 1807 5162 1913
rect 5208 1947 5262 1959
rect 5208 1921 5218 1947
rect 5252 1921 5262 1947
rect 5208 1869 5209 1921
rect 5261 1869 5262 1921
rect 5208 1862 5262 1869
rect 5308 1947 5362 2053
rect 5408 2131 5462 2138
rect 5408 2079 5409 2131
rect 5461 2079 5462 2131
rect 5408 2053 5418 2079
rect 5452 2053 5462 2079
rect 5408 2041 5462 2053
rect 5508 2087 5562 2193
rect 5608 2227 5662 2239
rect 5608 2201 5618 2227
rect 5652 2201 5662 2227
rect 5608 2149 5609 2201
rect 5661 2149 5662 2201
rect 5608 2142 5662 2149
rect 5708 2227 5762 2333
rect 5808 2411 5862 2418
rect 5808 2359 5809 2411
rect 5861 2359 5862 2411
rect 5808 2333 5818 2359
rect 5852 2333 5862 2359
rect 5808 2321 5862 2333
rect 5908 2367 5962 2563
rect 6008 2597 6062 2609
rect 6008 2571 6018 2597
rect 6052 2571 6062 2597
rect 6008 2519 6009 2571
rect 6061 2519 6062 2571
rect 6008 2512 6062 2519
rect 6108 2597 6162 2703
rect 6208 2781 6262 2788
rect 6208 2729 6209 2781
rect 6261 2729 6262 2781
rect 6208 2703 6218 2729
rect 6252 2703 6262 2729
rect 6208 2691 6262 2703
rect 6308 2737 6362 2843
rect 6408 2877 6462 2889
rect 6408 2851 6418 2877
rect 6452 2851 6462 2877
rect 6408 2799 6409 2851
rect 6461 2799 6462 2851
rect 6408 2792 6462 2799
rect 6506 2858 6516 2892
rect 6550 2858 6560 2892
rect 6506 2851 6560 2858
rect 6506 2799 6507 2851
rect 6559 2799 6560 2851
rect 6506 2792 6560 2799
rect 6506 2752 6560 2764
rect 6308 2703 6318 2737
rect 6352 2703 6362 2737
rect 6108 2563 6118 2597
rect 6152 2563 6162 2597
rect 6002 2483 6068 2484
rect 6002 2431 6009 2483
rect 6061 2431 6068 2483
rect 6002 2430 6068 2431
rect 5908 2333 5918 2367
rect 5952 2333 5962 2367
rect 5708 2193 5718 2227
rect 5752 2193 5762 2227
rect 5508 2053 5518 2087
rect 5552 2053 5562 2087
rect 5308 1913 5318 1947
rect 5352 1913 5362 1947
rect 5108 1773 5118 1807
rect 5152 1773 5162 1807
rect 4908 1633 4918 1667
rect 4952 1633 4962 1667
rect 4708 1493 4718 1527
rect 4752 1493 4762 1527
rect 4508 1353 4518 1387
rect 4552 1353 4562 1387
rect 4402 1273 4468 1274
rect 4402 1221 4409 1273
rect 4461 1221 4468 1273
rect 4402 1220 4468 1221
rect 4308 1123 4318 1157
rect 4352 1123 4362 1157
rect 4108 983 4118 1017
rect 4152 983 4162 1017
rect 3908 843 3918 877
rect 3952 843 3962 877
rect 3708 703 3718 737
rect 3752 703 3762 737
rect 3508 563 3518 597
rect 3552 563 3562 597
rect 3308 423 3318 457
rect 3352 423 3362 457
rect 3108 283 3118 317
rect 3152 283 3162 317
rect 2908 143 2918 177
rect 2952 143 2962 177
rect 2802 63 2868 64
rect 2802 11 2809 63
rect 2861 11 2868 63
rect 2802 10 2868 11
rect 2708 -67 2709 -15
rect 2761 -67 2762 -15
rect 2708 -79 2718 -67
rect 2752 -79 2762 -67
rect 2508 -132 2562 -131
rect 2508 -143 2518 -132
rect 2552 -143 2562 -132
rect 2508 -195 2509 -143
rect 2561 -195 2562 -143
rect 2508 -210 2562 -195
rect 2612 -133 2658 -81
rect 2612 -167 2618 -133
rect 2652 -167 2658 -133
rect 2518 -291 2525 -239
rect 2577 -291 2584 -239
rect 2412 -397 2418 -363
rect 2452 -397 2458 -363
rect 2412 -435 2458 -397
rect 2412 -469 2418 -435
rect 2452 -469 2458 -435
rect 2412 -512 2458 -469
rect 2509 -326 2561 -320
rect 2509 -390 2518 -378
rect 2552 -390 2561 -378
rect 2509 -454 2518 -442
rect 2552 -454 2561 -442
rect 2509 -512 2561 -506
rect 2612 -363 2658 -167
rect 2708 -131 2709 -79
rect 2761 -131 2762 -79
rect 2808 -22 2862 10
rect 2808 -74 2809 -22
rect 2861 -74 2862 -22
rect 2808 -81 2862 -74
rect 2908 -15 2962 143
rect 3008 221 3062 228
rect 3008 169 3009 221
rect 3061 169 3062 221
rect 3008 143 3018 169
rect 3052 143 3062 169
rect 3008 131 3062 143
rect 3108 177 3162 283
rect 3208 317 3262 329
rect 3208 291 3218 317
rect 3252 291 3262 317
rect 3208 239 3209 291
rect 3261 239 3262 291
rect 3208 232 3262 239
rect 3308 317 3362 423
rect 3408 501 3462 508
rect 3408 449 3409 501
rect 3461 449 3462 501
rect 3408 423 3418 449
rect 3452 423 3462 449
rect 3408 411 3462 423
rect 3508 457 3562 563
rect 3608 597 3662 609
rect 3608 571 3618 597
rect 3652 571 3662 597
rect 3608 519 3609 571
rect 3661 519 3662 571
rect 3608 512 3662 519
rect 3708 597 3762 703
rect 3808 781 3862 788
rect 3808 729 3809 781
rect 3861 729 3862 781
rect 3808 703 3818 729
rect 3852 703 3862 729
rect 3808 691 3862 703
rect 3908 737 3962 843
rect 4008 877 4062 889
rect 4008 851 4018 877
rect 4052 851 4062 877
rect 4008 799 4009 851
rect 4061 799 4062 851
rect 4008 792 4062 799
rect 4108 877 4162 983
rect 4208 1061 4262 1068
rect 4208 1009 4209 1061
rect 4261 1009 4262 1061
rect 4208 983 4218 1009
rect 4252 983 4262 1009
rect 4208 971 4262 983
rect 4308 1017 4362 1123
rect 4408 1157 4462 1169
rect 4408 1131 4418 1157
rect 4452 1131 4462 1157
rect 4408 1079 4409 1131
rect 4461 1079 4462 1131
rect 4408 1072 4462 1079
rect 4508 1157 4562 1353
rect 4608 1431 4662 1438
rect 4608 1379 4609 1431
rect 4661 1379 4662 1431
rect 4608 1353 4618 1379
rect 4652 1353 4662 1379
rect 4608 1341 4662 1353
rect 4708 1387 4762 1493
rect 4808 1527 4862 1539
rect 4808 1501 4818 1527
rect 4852 1501 4862 1527
rect 4808 1449 4809 1501
rect 4861 1449 4862 1501
rect 4808 1442 4862 1449
rect 4908 1527 4962 1633
rect 5008 1711 5062 1718
rect 5008 1659 5009 1711
rect 5061 1659 5062 1711
rect 5008 1633 5018 1659
rect 5052 1633 5062 1659
rect 5008 1621 5062 1633
rect 5108 1667 5162 1773
rect 5208 1807 5262 1819
rect 5208 1781 5218 1807
rect 5252 1781 5262 1807
rect 5208 1729 5209 1781
rect 5261 1729 5262 1781
rect 5208 1722 5262 1729
rect 5308 1807 5362 1913
rect 5408 1991 5462 1998
rect 5408 1939 5409 1991
rect 5461 1939 5462 1991
rect 5408 1913 5418 1939
rect 5452 1913 5462 1939
rect 5408 1901 5462 1913
rect 5508 1947 5562 2053
rect 5608 2087 5662 2099
rect 5608 2061 5618 2087
rect 5652 2061 5662 2087
rect 5608 2009 5609 2061
rect 5661 2009 5662 2061
rect 5608 2002 5662 2009
rect 5708 2087 5762 2193
rect 5808 2271 5862 2278
rect 5808 2219 5809 2271
rect 5861 2219 5862 2271
rect 5808 2193 5818 2219
rect 5852 2193 5862 2219
rect 5808 2181 5862 2193
rect 5908 2227 5962 2333
rect 6008 2367 6062 2379
rect 6008 2341 6018 2367
rect 6052 2341 6062 2367
rect 6008 2289 6009 2341
rect 6061 2289 6062 2341
rect 6008 2282 6062 2289
rect 6108 2367 6162 2563
rect 6208 2641 6262 2648
rect 6208 2589 6209 2641
rect 6261 2589 6262 2641
rect 6208 2563 6218 2589
rect 6252 2563 6262 2589
rect 6208 2551 6262 2563
rect 6308 2597 6362 2703
rect 6408 2737 6462 2749
rect 6408 2711 6418 2737
rect 6452 2711 6462 2737
rect 6408 2659 6409 2711
rect 6461 2659 6462 2711
rect 6408 2652 6462 2659
rect 6506 2718 6516 2752
rect 6550 2718 6560 2752
rect 6506 2711 6560 2718
rect 6506 2659 6507 2711
rect 6559 2659 6560 2711
rect 6506 2652 6560 2659
rect 6506 2612 6560 2624
rect 6308 2563 6318 2597
rect 6352 2563 6362 2597
rect 6202 2499 6268 2500
rect 6202 2447 6209 2499
rect 6261 2447 6268 2499
rect 6202 2446 6268 2447
rect 6108 2333 6118 2367
rect 6152 2333 6162 2367
rect 5908 2193 5918 2227
rect 5952 2193 5962 2227
rect 5708 2053 5718 2087
rect 5752 2053 5762 2087
rect 5508 1913 5518 1947
rect 5552 1913 5562 1947
rect 5308 1773 5318 1807
rect 5352 1773 5362 1807
rect 5108 1633 5118 1667
rect 5152 1633 5162 1667
rect 4908 1493 4918 1527
rect 4952 1493 4962 1527
rect 4708 1353 4718 1387
rect 4752 1353 4762 1387
rect 4602 1289 4668 1290
rect 4602 1237 4609 1289
rect 4661 1237 4668 1289
rect 4602 1236 4668 1237
rect 4508 1123 4518 1157
rect 4552 1123 4562 1157
rect 4308 983 4318 1017
rect 4352 983 4362 1017
rect 4108 843 4118 877
rect 4152 843 4162 877
rect 3908 703 3918 737
rect 3952 703 3962 737
rect 3708 563 3718 597
rect 3752 563 3762 597
rect 3508 423 3518 457
rect 3552 423 3562 457
rect 3308 283 3318 317
rect 3352 283 3362 317
rect 3108 143 3118 177
rect 3152 143 3162 177
rect 3002 79 3068 80
rect 3002 27 3009 79
rect 3061 27 3068 79
rect 3002 26 3068 27
rect 2908 -67 2909 -15
rect 2961 -67 2962 -15
rect 2908 -79 2918 -67
rect 2952 -79 2962 -67
rect 2708 -132 2762 -131
rect 2708 -143 2718 -132
rect 2752 -143 2762 -132
rect 2708 -195 2709 -143
rect 2761 -195 2762 -143
rect 2708 -210 2762 -195
rect 2812 -133 2858 -81
rect 2812 -167 2818 -133
rect 2852 -167 2858 -133
rect 2718 -291 2725 -239
rect 2777 -291 2784 -239
rect 2612 -397 2618 -363
rect 2652 -397 2658 -363
rect 2612 -435 2658 -397
rect 2612 -469 2618 -435
rect 2652 -469 2658 -435
rect 2612 -512 2658 -469
rect 2709 -326 2761 -320
rect 2709 -390 2718 -378
rect 2752 -390 2761 -378
rect 2709 -454 2718 -442
rect 2752 -454 2761 -442
rect 2709 -555 2761 -506
rect 2812 -363 2858 -167
rect 2908 -131 2909 -79
rect 2961 -131 2962 -79
rect 3008 -22 3062 26
rect 3008 -74 3009 -22
rect 3061 -74 3062 -22
rect 3008 -81 3062 -74
rect 3108 -15 3162 143
rect 3208 177 3262 189
rect 3208 151 3218 177
rect 3252 151 3262 177
rect 3208 99 3209 151
rect 3261 99 3262 151
rect 3208 92 3262 99
rect 3308 177 3362 283
rect 3408 361 3462 368
rect 3408 309 3409 361
rect 3461 309 3462 361
rect 3408 283 3418 309
rect 3452 283 3462 309
rect 3408 271 3462 283
rect 3508 317 3562 423
rect 3608 457 3662 469
rect 3608 431 3618 457
rect 3652 431 3662 457
rect 3608 379 3609 431
rect 3661 379 3662 431
rect 3608 372 3662 379
rect 3708 457 3762 563
rect 3808 641 3862 648
rect 3808 589 3809 641
rect 3861 589 3862 641
rect 3808 563 3818 589
rect 3852 563 3862 589
rect 3808 551 3862 563
rect 3908 597 3962 703
rect 4008 737 4062 749
rect 4008 711 4018 737
rect 4052 711 4062 737
rect 4008 659 4009 711
rect 4061 659 4062 711
rect 4008 652 4062 659
rect 4108 737 4162 843
rect 4208 921 4262 928
rect 4208 869 4209 921
rect 4261 869 4262 921
rect 4208 843 4218 869
rect 4252 843 4262 869
rect 4208 831 4262 843
rect 4308 877 4362 983
rect 4408 1017 4462 1029
rect 4408 991 4418 1017
rect 4452 991 4462 1017
rect 4408 939 4409 991
rect 4461 939 4462 991
rect 4408 932 4462 939
rect 4508 1017 4562 1123
rect 4608 1201 4662 1208
rect 4608 1149 4609 1201
rect 4661 1149 4662 1201
rect 4608 1123 4618 1149
rect 4652 1123 4662 1149
rect 4608 1111 4662 1123
rect 4708 1157 4762 1353
rect 4808 1387 4862 1399
rect 4808 1361 4818 1387
rect 4852 1361 4862 1387
rect 4808 1309 4809 1361
rect 4861 1309 4862 1361
rect 4808 1302 4862 1309
rect 4908 1387 4962 1493
rect 5008 1571 5062 1578
rect 5008 1519 5009 1571
rect 5061 1519 5062 1571
rect 5008 1493 5018 1519
rect 5052 1493 5062 1519
rect 5008 1481 5062 1493
rect 5108 1527 5162 1633
rect 5208 1667 5262 1679
rect 5208 1641 5218 1667
rect 5252 1641 5262 1667
rect 5208 1589 5209 1641
rect 5261 1589 5262 1641
rect 5208 1582 5262 1589
rect 5308 1667 5362 1773
rect 5408 1851 5462 1858
rect 5408 1799 5409 1851
rect 5461 1799 5462 1851
rect 5408 1773 5418 1799
rect 5452 1773 5462 1799
rect 5408 1761 5462 1773
rect 5508 1807 5562 1913
rect 5608 1947 5662 1959
rect 5608 1921 5618 1947
rect 5652 1921 5662 1947
rect 5608 1869 5609 1921
rect 5661 1869 5662 1921
rect 5608 1862 5662 1869
rect 5708 1947 5762 2053
rect 5808 2131 5862 2138
rect 5808 2079 5809 2131
rect 5861 2079 5862 2131
rect 5808 2053 5818 2079
rect 5852 2053 5862 2079
rect 5808 2041 5862 2053
rect 5908 2087 5962 2193
rect 6008 2227 6062 2239
rect 6008 2201 6018 2227
rect 6052 2201 6062 2227
rect 6008 2149 6009 2201
rect 6061 2149 6062 2201
rect 6008 2142 6062 2149
rect 6108 2227 6162 2333
rect 6208 2411 6262 2418
rect 6208 2359 6209 2411
rect 6261 2359 6262 2411
rect 6208 2333 6218 2359
rect 6252 2333 6262 2359
rect 6208 2321 6262 2333
rect 6308 2367 6362 2563
rect 6408 2597 6462 2609
rect 6408 2571 6418 2597
rect 6452 2571 6462 2597
rect 6408 2519 6409 2571
rect 6461 2519 6462 2571
rect 6408 2512 6462 2519
rect 6506 2578 6516 2612
rect 6550 2578 6560 2612
rect 6506 2571 6560 2578
rect 6506 2519 6507 2571
rect 6559 2519 6560 2571
rect 6506 2512 6560 2519
rect 6590 2477 6620 3641
rect 6504 2471 6620 2477
rect 6504 2437 6516 2471
rect 6550 2437 6620 2471
rect 6504 2431 6620 2437
rect 6506 2382 6560 2394
rect 6308 2333 6318 2367
rect 6352 2333 6362 2367
rect 6108 2193 6118 2227
rect 6152 2193 6162 2227
rect 5908 2053 5918 2087
rect 5952 2053 5962 2087
rect 5708 1913 5718 1947
rect 5752 1913 5762 1947
rect 5508 1773 5518 1807
rect 5552 1773 5562 1807
rect 5308 1633 5318 1667
rect 5352 1633 5362 1667
rect 5108 1493 5118 1527
rect 5152 1493 5162 1527
rect 4908 1353 4918 1387
rect 4952 1353 4962 1387
rect 4802 1273 4868 1274
rect 4802 1221 4809 1273
rect 4861 1221 4868 1273
rect 4802 1220 4868 1221
rect 4708 1123 4718 1157
rect 4752 1123 4762 1157
rect 4508 983 4518 1017
rect 4552 983 4562 1017
rect 4308 843 4318 877
rect 4352 843 4362 877
rect 4108 703 4118 737
rect 4152 703 4162 737
rect 3908 563 3918 597
rect 3952 563 3962 597
rect 3708 423 3718 457
rect 3752 423 3762 457
rect 3508 283 3518 317
rect 3552 283 3562 317
rect 3308 143 3318 177
rect 3352 143 3362 177
rect 3202 63 3268 64
rect 3202 11 3209 63
rect 3261 11 3268 63
rect 3202 10 3268 11
rect 3108 -67 3109 -15
rect 3161 -67 3162 -15
rect 3108 -79 3118 -67
rect 3152 -79 3162 -67
rect 2908 -132 2962 -131
rect 2908 -143 2918 -132
rect 2952 -143 2962 -132
rect 2908 -195 2909 -143
rect 2961 -195 2962 -143
rect 2908 -210 2962 -195
rect 3012 -133 3058 -81
rect 3012 -167 3018 -133
rect 3052 -167 3058 -133
rect 2918 -291 2925 -239
rect 2977 -291 2984 -239
rect 2812 -397 2818 -363
rect 2852 -397 2858 -363
rect 2812 -435 2858 -397
rect 2812 -469 2818 -435
rect 2852 -469 2858 -435
rect 2812 -512 2858 -469
rect 2909 -326 2961 -320
rect 2909 -390 2918 -378
rect 2952 -390 2961 -378
rect 2909 -454 2918 -442
rect 2952 -454 2961 -442
rect 2909 -512 2961 -506
rect 3012 -363 3058 -167
rect 3108 -131 3109 -79
rect 3161 -131 3162 -79
rect 3208 -22 3262 10
rect 3208 -74 3209 -22
rect 3261 -74 3262 -22
rect 3208 -81 3262 -74
rect 3308 -15 3362 143
rect 3408 221 3462 228
rect 3408 169 3409 221
rect 3461 169 3462 221
rect 3408 143 3418 169
rect 3452 143 3462 169
rect 3408 131 3462 143
rect 3508 177 3562 283
rect 3608 317 3662 329
rect 3608 291 3618 317
rect 3652 291 3662 317
rect 3608 239 3609 291
rect 3661 239 3662 291
rect 3608 232 3662 239
rect 3708 317 3762 423
rect 3808 501 3862 508
rect 3808 449 3809 501
rect 3861 449 3862 501
rect 3808 423 3818 449
rect 3852 423 3862 449
rect 3808 411 3862 423
rect 3908 457 3962 563
rect 4008 597 4062 609
rect 4008 571 4018 597
rect 4052 571 4062 597
rect 4008 519 4009 571
rect 4061 519 4062 571
rect 4008 512 4062 519
rect 4108 597 4162 703
rect 4208 781 4262 788
rect 4208 729 4209 781
rect 4261 729 4262 781
rect 4208 703 4218 729
rect 4252 703 4262 729
rect 4208 691 4262 703
rect 4308 737 4362 843
rect 4408 877 4462 889
rect 4408 851 4418 877
rect 4452 851 4462 877
rect 4408 799 4409 851
rect 4461 799 4462 851
rect 4408 792 4462 799
rect 4508 877 4562 983
rect 4608 1061 4662 1068
rect 4608 1009 4609 1061
rect 4661 1009 4662 1061
rect 4608 983 4618 1009
rect 4652 983 4662 1009
rect 4608 971 4662 983
rect 4708 1017 4762 1123
rect 4808 1157 4862 1169
rect 4808 1131 4818 1157
rect 4852 1131 4862 1157
rect 4808 1079 4809 1131
rect 4861 1079 4862 1131
rect 4808 1072 4862 1079
rect 4908 1157 4962 1353
rect 5008 1431 5062 1438
rect 5008 1379 5009 1431
rect 5061 1379 5062 1431
rect 5008 1353 5018 1379
rect 5052 1353 5062 1379
rect 5008 1341 5062 1353
rect 5108 1387 5162 1493
rect 5208 1527 5262 1539
rect 5208 1501 5218 1527
rect 5252 1501 5262 1527
rect 5208 1449 5209 1501
rect 5261 1449 5262 1501
rect 5208 1442 5262 1449
rect 5308 1527 5362 1633
rect 5408 1711 5462 1718
rect 5408 1659 5409 1711
rect 5461 1659 5462 1711
rect 5408 1633 5418 1659
rect 5452 1633 5462 1659
rect 5408 1621 5462 1633
rect 5508 1667 5562 1773
rect 5608 1807 5662 1819
rect 5608 1781 5618 1807
rect 5652 1781 5662 1807
rect 5608 1729 5609 1781
rect 5661 1729 5662 1781
rect 5608 1722 5662 1729
rect 5708 1807 5762 1913
rect 5808 1991 5862 1998
rect 5808 1939 5809 1991
rect 5861 1939 5862 1991
rect 5808 1913 5818 1939
rect 5852 1913 5862 1939
rect 5808 1901 5862 1913
rect 5908 1947 5962 2053
rect 6008 2087 6062 2099
rect 6008 2061 6018 2087
rect 6052 2061 6062 2087
rect 6008 2009 6009 2061
rect 6061 2009 6062 2061
rect 6008 2002 6062 2009
rect 6108 2087 6162 2193
rect 6208 2271 6262 2278
rect 6208 2219 6209 2271
rect 6261 2219 6262 2271
rect 6208 2193 6218 2219
rect 6252 2193 6262 2219
rect 6208 2181 6262 2193
rect 6308 2227 6362 2333
rect 6408 2367 6462 2379
rect 6408 2341 6418 2367
rect 6452 2341 6462 2367
rect 6408 2289 6409 2341
rect 6461 2289 6462 2341
rect 6408 2282 6462 2289
rect 6506 2348 6516 2382
rect 6550 2348 6560 2382
rect 6506 2341 6560 2348
rect 6506 2289 6507 2341
rect 6559 2289 6560 2341
rect 6506 2282 6560 2289
rect 6506 2242 6560 2254
rect 6308 2193 6318 2227
rect 6352 2193 6362 2227
rect 6108 2053 6118 2087
rect 6152 2053 6162 2087
rect 5908 1913 5918 1947
rect 5952 1913 5962 1947
rect 5708 1773 5718 1807
rect 5752 1773 5762 1807
rect 5508 1633 5518 1667
rect 5552 1633 5562 1667
rect 5308 1493 5318 1527
rect 5352 1493 5362 1527
rect 5108 1353 5118 1387
rect 5152 1353 5162 1387
rect 5002 1289 5068 1290
rect 5002 1237 5009 1289
rect 5061 1237 5068 1289
rect 5002 1236 5068 1237
rect 4908 1123 4918 1157
rect 4952 1123 4962 1157
rect 4708 983 4718 1017
rect 4752 983 4762 1017
rect 4508 843 4518 877
rect 4552 843 4562 877
rect 4308 703 4318 737
rect 4352 703 4362 737
rect 4108 563 4118 597
rect 4152 563 4162 597
rect 3908 423 3918 457
rect 3952 423 3962 457
rect 3708 283 3718 317
rect 3752 283 3762 317
rect 3508 143 3518 177
rect 3552 143 3562 177
rect 3402 79 3468 80
rect 3402 27 3409 79
rect 3461 27 3468 79
rect 3402 26 3468 27
rect 3308 -67 3309 -15
rect 3361 -67 3362 -15
rect 3308 -79 3318 -67
rect 3352 -79 3362 -67
rect 3108 -132 3162 -131
rect 3108 -143 3118 -132
rect 3152 -143 3162 -132
rect 3108 -195 3109 -143
rect 3161 -195 3162 -143
rect 3108 -210 3162 -195
rect 3212 -133 3258 -81
rect 3212 -167 3218 -133
rect 3252 -167 3258 -133
rect 3118 -291 3125 -239
rect 3177 -291 3184 -239
rect 3012 -397 3018 -363
rect 3052 -397 3058 -363
rect 3012 -435 3058 -397
rect 3012 -469 3018 -435
rect 3052 -469 3058 -435
rect 3012 -512 3058 -469
rect 3109 -326 3161 -320
rect 3109 -390 3118 -378
rect 3152 -390 3161 -378
rect 3109 -454 3118 -442
rect 3152 -454 3161 -442
rect 3109 -555 3161 -506
rect 3212 -363 3258 -167
rect 3308 -131 3309 -79
rect 3361 -131 3362 -79
rect 3408 -22 3462 26
rect 3408 -74 3409 -22
rect 3461 -74 3462 -22
rect 3408 -81 3462 -74
rect 3508 -15 3562 143
rect 3608 177 3662 189
rect 3608 151 3618 177
rect 3652 151 3662 177
rect 3608 99 3609 151
rect 3661 99 3662 151
rect 3608 92 3662 99
rect 3708 177 3762 283
rect 3808 361 3862 368
rect 3808 309 3809 361
rect 3861 309 3862 361
rect 3808 283 3818 309
rect 3852 283 3862 309
rect 3808 271 3862 283
rect 3908 317 3962 423
rect 4008 457 4062 469
rect 4008 431 4018 457
rect 4052 431 4062 457
rect 4008 379 4009 431
rect 4061 379 4062 431
rect 4008 372 4062 379
rect 4108 457 4162 563
rect 4208 641 4262 648
rect 4208 589 4209 641
rect 4261 589 4262 641
rect 4208 563 4218 589
rect 4252 563 4262 589
rect 4208 551 4262 563
rect 4308 597 4362 703
rect 4408 737 4462 749
rect 4408 711 4418 737
rect 4452 711 4462 737
rect 4408 659 4409 711
rect 4461 659 4462 711
rect 4408 652 4462 659
rect 4508 737 4562 843
rect 4608 921 4662 928
rect 4608 869 4609 921
rect 4661 869 4662 921
rect 4608 843 4618 869
rect 4652 843 4662 869
rect 4608 831 4662 843
rect 4708 877 4762 983
rect 4808 1017 4862 1029
rect 4808 991 4818 1017
rect 4852 991 4862 1017
rect 4808 939 4809 991
rect 4861 939 4862 991
rect 4808 932 4862 939
rect 4908 1017 4962 1123
rect 5008 1201 5062 1208
rect 5008 1149 5009 1201
rect 5061 1149 5062 1201
rect 5008 1123 5018 1149
rect 5052 1123 5062 1149
rect 5008 1111 5062 1123
rect 5108 1157 5162 1353
rect 5208 1387 5262 1399
rect 5208 1361 5218 1387
rect 5252 1361 5262 1387
rect 5208 1309 5209 1361
rect 5261 1309 5262 1361
rect 5208 1302 5262 1309
rect 5308 1387 5362 1493
rect 5408 1571 5462 1578
rect 5408 1519 5409 1571
rect 5461 1519 5462 1571
rect 5408 1493 5418 1519
rect 5452 1493 5462 1519
rect 5408 1481 5462 1493
rect 5508 1527 5562 1633
rect 5608 1667 5662 1679
rect 5608 1641 5618 1667
rect 5652 1641 5662 1667
rect 5608 1589 5609 1641
rect 5661 1589 5662 1641
rect 5608 1582 5662 1589
rect 5708 1667 5762 1773
rect 5808 1851 5862 1858
rect 5808 1799 5809 1851
rect 5861 1799 5862 1851
rect 5808 1773 5818 1799
rect 5852 1773 5862 1799
rect 5808 1761 5862 1773
rect 5908 1807 5962 1913
rect 6008 1947 6062 1959
rect 6008 1921 6018 1947
rect 6052 1921 6062 1947
rect 6008 1869 6009 1921
rect 6061 1869 6062 1921
rect 6008 1862 6062 1869
rect 6108 1947 6162 2053
rect 6208 2131 6262 2138
rect 6208 2079 6209 2131
rect 6261 2079 6262 2131
rect 6208 2053 6218 2079
rect 6252 2053 6262 2079
rect 6208 2041 6262 2053
rect 6308 2087 6362 2193
rect 6408 2227 6462 2239
rect 6408 2201 6418 2227
rect 6452 2201 6462 2227
rect 6408 2149 6409 2201
rect 6461 2149 6462 2201
rect 6408 2142 6462 2149
rect 6506 2208 6516 2242
rect 6550 2208 6560 2242
rect 6506 2201 6560 2208
rect 6506 2149 6507 2201
rect 6559 2149 6560 2201
rect 6506 2142 6560 2149
rect 6506 2102 6560 2114
rect 6308 2053 6318 2087
rect 6352 2053 6362 2087
rect 6108 1913 6118 1947
rect 6152 1913 6162 1947
rect 5908 1773 5918 1807
rect 5952 1773 5962 1807
rect 5708 1633 5718 1667
rect 5752 1633 5762 1667
rect 5508 1493 5518 1527
rect 5552 1493 5562 1527
rect 5308 1353 5318 1387
rect 5352 1353 5362 1387
rect 5202 1273 5268 1274
rect 5202 1221 5209 1273
rect 5261 1221 5268 1273
rect 5202 1220 5268 1221
rect 5108 1123 5118 1157
rect 5152 1123 5162 1157
rect 4908 983 4918 1017
rect 4952 983 4962 1017
rect 4708 843 4718 877
rect 4752 843 4762 877
rect 4508 703 4518 737
rect 4552 703 4562 737
rect 4308 563 4318 597
rect 4352 563 4362 597
rect 4108 423 4118 457
rect 4152 423 4162 457
rect 3908 283 3918 317
rect 3952 283 3962 317
rect 3708 143 3718 177
rect 3752 143 3762 177
rect 3602 63 3668 64
rect 3602 11 3609 63
rect 3661 11 3668 63
rect 3602 10 3668 11
rect 3508 -67 3509 -15
rect 3561 -67 3562 -15
rect 3508 -79 3518 -67
rect 3552 -79 3562 -67
rect 3308 -132 3362 -131
rect 3308 -143 3318 -132
rect 3352 -143 3362 -132
rect 3308 -195 3309 -143
rect 3361 -195 3362 -143
rect 3308 -210 3362 -195
rect 3412 -133 3458 -81
rect 3412 -167 3418 -133
rect 3452 -167 3458 -133
rect 3318 -291 3325 -239
rect 3377 -291 3384 -239
rect 3212 -397 3218 -363
rect 3252 -397 3258 -363
rect 3212 -435 3258 -397
rect 3212 -469 3218 -435
rect 3252 -469 3258 -435
rect 3212 -512 3258 -469
rect 3309 -326 3361 -320
rect 3309 -390 3318 -378
rect 3352 -390 3361 -378
rect 3309 -454 3318 -442
rect 3352 -454 3361 -442
rect 3309 -512 3361 -506
rect 3412 -363 3458 -167
rect 3508 -131 3509 -79
rect 3561 -131 3562 -79
rect 3608 -22 3662 10
rect 3608 -74 3609 -22
rect 3661 -74 3662 -22
rect 3608 -81 3662 -74
rect 3708 -15 3762 143
rect 3808 221 3862 228
rect 3808 169 3809 221
rect 3861 169 3862 221
rect 3808 143 3818 169
rect 3852 143 3862 169
rect 3808 131 3862 143
rect 3908 177 3962 283
rect 4008 317 4062 329
rect 4008 291 4018 317
rect 4052 291 4062 317
rect 4008 239 4009 291
rect 4061 239 4062 291
rect 4008 232 4062 239
rect 4108 317 4162 423
rect 4208 501 4262 508
rect 4208 449 4209 501
rect 4261 449 4262 501
rect 4208 423 4218 449
rect 4252 423 4262 449
rect 4208 411 4262 423
rect 4308 457 4362 563
rect 4408 597 4462 609
rect 4408 571 4418 597
rect 4452 571 4462 597
rect 4408 519 4409 571
rect 4461 519 4462 571
rect 4408 512 4462 519
rect 4508 597 4562 703
rect 4608 781 4662 788
rect 4608 729 4609 781
rect 4661 729 4662 781
rect 4608 703 4618 729
rect 4652 703 4662 729
rect 4608 691 4662 703
rect 4708 737 4762 843
rect 4808 877 4862 889
rect 4808 851 4818 877
rect 4852 851 4862 877
rect 4808 799 4809 851
rect 4861 799 4862 851
rect 4808 792 4862 799
rect 4908 877 4962 983
rect 5008 1061 5062 1068
rect 5008 1009 5009 1061
rect 5061 1009 5062 1061
rect 5008 983 5018 1009
rect 5052 983 5062 1009
rect 5008 971 5062 983
rect 5108 1017 5162 1123
rect 5208 1157 5262 1169
rect 5208 1131 5218 1157
rect 5252 1131 5262 1157
rect 5208 1079 5209 1131
rect 5261 1079 5262 1131
rect 5208 1072 5262 1079
rect 5308 1157 5362 1353
rect 5408 1431 5462 1438
rect 5408 1379 5409 1431
rect 5461 1379 5462 1431
rect 5408 1353 5418 1379
rect 5452 1353 5462 1379
rect 5408 1341 5462 1353
rect 5508 1387 5562 1493
rect 5608 1527 5662 1539
rect 5608 1501 5618 1527
rect 5652 1501 5662 1527
rect 5608 1449 5609 1501
rect 5661 1449 5662 1501
rect 5608 1442 5662 1449
rect 5708 1527 5762 1633
rect 5808 1711 5862 1718
rect 5808 1659 5809 1711
rect 5861 1659 5862 1711
rect 5808 1633 5818 1659
rect 5852 1633 5862 1659
rect 5808 1621 5862 1633
rect 5908 1667 5962 1773
rect 6008 1807 6062 1819
rect 6008 1781 6018 1807
rect 6052 1781 6062 1807
rect 6008 1729 6009 1781
rect 6061 1729 6062 1781
rect 6008 1722 6062 1729
rect 6108 1807 6162 1913
rect 6208 1991 6262 1998
rect 6208 1939 6209 1991
rect 6261 1939 6262 1991
rect 6208 1913 6218 1939
rect 6252 1913 6262 1939
rect 6208 1901 6262 1913
rect 6308 1947 6362 2053
rect 6408 2087 6462 2099
rect 6408 2061 6418 2087
rect 6452 2061 6462 2087
rect 6408 2009 6409 2061
rect 6461 2009 6462 2061
rect 6408 2002 6462 2009
rect 6506 2068 6516 2102
rect 6550 2068 6560 2102
rect 6506 2061 6560 2068
rect 6506 2009 6507 2061
rect 6559 2009 6560 2061
rect 6506 2002 6560 2009
rect 6506 1962 6560 1974
rect 6308 1913 6318 1947
rect 6352 1913 6362 1947
rect 6108 1773 6118 1807
rect 6152 1773 6162 1807
rect 5908 1633 5918 1667
rect 5952 1633 5962 1667
rect 5708 1493 5718 1527
rect 5752 1493 5762 1527
rect 5508 1353 5518 1387
rect 5552 1353 5562 1387
rect 5402 1289 5468 1290
rect 5402 1237 5409 1289
rect 5461 1237 5468 1289
rect 5402 1236 5468 1237
rect 5308 1123 5318 1157
rect 5352 1123 5362 1157
rect 5108 983 5118 1017
rect 5152 983 5162 1017
rect 4908 843 4918 877
rect 4952 843 4962 877
rect 4708 703 4718 737
rect 4752 703 4762 737
rect 4508 563 4518 597
rect 4552 563 4562 597
rect 4308 423 4318 457
rect 4352 423 4362 457
rect 4108 283 4118 317
rect 4152 283 4162 317
rect 3908 143 3918 177
rect 3952 143 3962 177
rect 3802 79 3868 80
rect 3802 27 3809 79
rect 3861 27 3868 79
rect 3802 26 3868 27
rect 3708 -67 3709 -15
rect 3761 -67 3762 -15
rect 3708 -79 3718 -67
rect 3752 -79 3762 -67
rect 3508 -132 3562 -131
rect 3508 -143 3518 -132
rect 3552 -143 3562 -132
rect 3508 -195 3509 -143
rect 3561 -195 3562 -143
rect 3508 -210 3562 -195
rect 3612 -133 3658 -81
rect 3612 -167 3618 -133
rect 3652 -167 3658 -133
rect 3518 -291 3525 -239
rect 3577 -291 3584 -239
rect 3412 -397 3418 -363
rect 3452 -397 3458 -363
rect 3412 -435 3458 -397
rect 3412 -469 3418 -435
rect 3452 -469 3458 -435
rect 3412 -512 3458 -469
rect 3509 -326 3561 -320
rect 3509 -390 3518 -378
rect 3552 -390 3561 -378
rect 3509 -454 3518 -442
rect 3552 -454 3561 -442
rect 3509 -555 3561 -506
rect 3612 -363 3658 -167
rect 3708 -131 3709 -79
rect 3761 -131 3762 -79
rect 3808 -22 3862 26
rect 3808 -74 3809 -22
rect 3861 -74 3862 -22
rect 3808 -81 3862 -74
rect 3908 -15 3962 143
rect 4008 177 4062 189
rect 4008 151 4018 177
rect 4052 151 4062 177
rect 4008 99 4009 151
rect 4061 99 4062 151
rect 4008 92 4062 99
rect 4108 177 4162 283
rect 4208 361 4262 368
rect 4208 309 4209 361
rect 4261 309 4262 361
rect 4208 283 4218 309
rect 4252 283 4262 309
rect 4208 271 4262 283
rect 4308 317 4362 423
rect 4408 457 4462 469
rect 4408 431 4418 457
rect 4452 431 4462 457
rect 4408 379 4409 431
rect 4461 379 4462 431
rect 4408 372 4462 379
rect 4508 457 4562 563
rect 4608 641 4662 648
rect 4608 589 4609 641
rect 4661 589 4662 641
rect 4608 563 4618 589
rect 4652 563 4662 589
rect 4608 551 4662 563
rect 4708 597 4762 703
rect 4808 737 4862 749
rect 4808 711 4818 737
rect 4852 711 4862 737
rect 4808 659 4809 711
rect 4861 659 4862 711
rect 4808 652 4862 659
rect 4908 737 4962 843
rect 5008 921 5062 928
rect 5008 869 5009 921
rect 5061 869 5062 921
rect 5008 843 5018 869
rect 5052 843 5062 869
rect 5008 831 5062 843
rect 5108 877 5162 983
rect 5208 1017 5262 1029
rect 5208 991 5218 1017
rect 5252 991 5262 1017
rect 5208 939 5209 991
rect 5261 939 5262 991
rect 5208 932 5262 939
rect 5308 1017 5362 1123
rect 5408 1201 5462 1208
rect 5408 1149 5409 1201
rect 5461 1149 5462 1201
rect 5408 1123 5418 1149
rect 5452 1123 5462 1149
rect 5408 1111 5462 1123
rect 5508 1157 5562 1353
rect 5608 1387 5662 1399
rect 5608 1361 5618 1387
rect 5652 1361 5662 1387
rect 5608 1309 5609 1361
rect 5661 1309 5662 1361
rect 5608 1302 5662 1309
rect 5708 1387 5762 1493
rect 5808 1571 5862 1578
rect 5808 1519 5809 1571
rect 5861 1519 5862 1571
rect 5808 1493 5818 1519
rect 5852 1493 5862 1519
rect 5808 1481 5862 1493
rect 5908 1527 5962 1633
rect 6008 1667 6062 1679
rect 6008 1641 6018 1667
rect 6052 1641 6062 1667
rect 6008 1589 6009 1641
rect 6061 1589 6062 1641
rect 6008 1582 6062 1589
rect 6108 1667 6162 1773
rect 6208 1851 6262 1858
rect 6208 1799 6209 1851
rect 6261 1799 6262 1851
rect 6208 1773 6218 1799
rect 6252 1773 6262 1799
rect 6208 1761 6262 1773
rect 6308 1807 6362 1913
rect 6408 1947 6462 1959
rect 6408 1921 6418 1947
rect 6452 1921 6462 1947
rect 6408 1869 6409 1921
rect 6461 1869 6462 1921
rect 6408 1862 6462 1869
rect 6506 1928 6516 1962
rect 6550 1928 6560 1962
rect 6506 1921 6560 1928
rect 6506 1869 6507 1921
rect 6559 1869 6560 1921
rect 6506 1862 6560 1869
rect 6506 1822 6560 1834
rect 6308 1773 6318 1807
rect 6352 1773 6362 1807
rect 6108 1633 6118 1667
rect 6152 1633 6162 1667
rect 5908 1493 5918 1527
rect 5952 1493 5962 1527
rect 5708 1353 5718 1387
rect 5752 1353 5762 1387
rect 5602 1273 5668 1274
rect 5602 1221 5609 1273
rect 5661 1221 5668 1273
rect 5602 1220 5668 1221
rect 5508 1123 5518 1157
rect 5552 1123 5562 1157
rect 5308 983 5318 1017
rect 5352 983 5362 1017
rect 5108 843 5118 877
rect 5152 843 5162 877
rect 4908 703 4918 737
rect 4952 703 4962 737
rect 4708 563 4718 597
rect 4752 563 4762 597
rect 4508 423 4518 457
rect 4552 423 4562 457
rect 4308 283 4318 317
rect 4352 283 4362 317
rect 4108 143 4118 177
rect 4152 143 4162 177
rect 4002 63 4068 64
rect 4002 11 4009 63
rect 4061 11 4068 63
rect 4002 10 4068 11
rect 3908 -67 3909 -15
rect 3961 -67 3962 -15
rect 3908 -79 3918 -67
rect 3952 -79 3962 -67
rect 3708 -132 3762 -131
rect 3708 -143 3718 -132
rect 3752 -143 3762 -132
rect 3708 -195 3709 -143
rect 3761 -195 3762 -143
rect 3708 -210 3762 -195
rect 3812 -133 3858 -81
rect 3812 -167 3818 -133
rect 3852 -167 3858 -133
rect 3718 -291 3725 -239
rect 3777 -291 3784 -239
rect 3612 -397 3618 -363
rect 3652 -397 3658 -363
rect 3612 -435 3658 -397
rect 3612 -469 3618 -435
rect 3652 -469 3658 -435
rect 3612 -512 3658 -469
rect 3709 -326 3761 -320
rect 3709 -390 3718 -378
rect 3752 -390 3761 -378
rect 3709 -454 3718 -442
rect 3752 -454 3761 -442
rect 3709 -512 3761 -506
rect 3812 -363 3858 -167
rect 3908 -131 3909 -79
rect 3961 -131 3962 -79
rect 4008 -22 4062 10
rect 4008 -74 4009 -22
rect 4061 -74 4062 -22
rect 4008 -81 4062 -74
rect 4108 -15 4162 143
rect 4208 221 4262 228
rect 4208 169 4209 221
rect 4261 169 4262 221
rect 4208 143 4218 169
rect 4252 143 4262 169
rect 4208 131 4262 143
rect 4308 177 4362 283
rect 4408 317 4462 329
rect 4408 291 4418 317
rect 4452 291 4462 317
rect 4408 239 4409 291
rect 4461 239 4462 291
rect 4408 232 4462 239
rect 4508 317 4562 423
rect 4608 501 4662 508
rect 4608 449 4609 501
rect 4661 449 4662 501
rect 4608 423 4618 449
rect 4652 423 4662 449
rect 4608 411 4662 423
rect 4708 457 4762 563
rect 4808 597 4862 609
rect 4808 571 4818 597
rect 4852 571 4862 597
rect 4808 519 4809 571
rect 4861 519 4862 571
rect 4808 512 4862 519
rect 4908 597 4962 703
rect 5008 781 5062 788
rect 5008 729 5009 781
rect 5061 729 5062 781
rect 5008 703 5018 729
rect 5052 703 5062 729
rect 5008 691 5062 703
rect 5108 737 5162 843
rect 5208 877 5262 889
rect 5208 851 5218 877
rect 5252 851 5262 877
rect 5208 799 5209 851
rect 5261 799 5262 851
rect 5208 792 5262 799
rect 5308 877 5362 983
rect 5408 1061 5462 1068
rect 5408 1009 5409 1061
rect 5461 1009 5462 1061
rect 5408 983 5418 1009
rect 5452 983 5462 1009
rect 5408 971 5462 983
rect 5508 1017 5562 1123
rect 5608 1157 5662 1169
rect 5608 1131 5618 1157
rect 5652 1131 5662 1157
rect 5608 1079 5609 1131
rect 5661 1079 5662 1131
rect 5608 1072 5662 1079
rect 5708 1157 5762 1353
rect 5808 1431 5862 1438
rect 5808 1379 5809 1431
rect 5861 1379 5862 1431
rect 5808 1353 5818 1379
rect 5852 1353 5862 1379
rect 5808 1341 5862 1353
rect 5908 1387 5962 1493
rect 6008 1527 6062 1539
rect 6008 1501 6018 1527
rect 6052 1501 6062 1527
rect 6008 1449 6009 1501
rect 6061 1449 6062 1501
rect 6008 1442 6062 1449
rect 6108 1527 6162 1633
rect 6208 1711 6262 1718
rect 6208 1659 6209 1711
rect 6261 1659 6262 1711
rect 6208 1633 6218 1659
rect 6252 1633 6262 1659
rect 6208 1621 6262 1633
rect 6308 1667 6362 1773
rect 6408 1807 6462 1819
rect 6408 1781 6418 1807
rect 6452 1781 6462 1807
rect 6408 1729 6409 1781
rect 6461 1729 6462 1781
rect 6408 1722 6462 1729
rect 6506 1788 6516 1822
rect 6550 1788 6560 1822
rect 6506 1781 6560 1788
rect 6506 1729 6507 1781
rect 6559 1729 6560 1781
rect 6506 1722 6560 1729
rect 6506 1682 6560 1694
rect 6308 1633 6318 1667
rect 6352 1633 6362 1667
rect 6108 1493 6118 1527
rect 6152 1493 6162 1527
rect 5908 1353 5918 1387
rect 5952 1353 5962 1387
rect 5802 1289 5868 1290
rect 5802 1237 5809 1289
rect 5861 1237 5868 1289
rect 5802 1236 5868 1237
rect 5708 1123 5718 1157
rect 5752 1123 5762 1157
rect 5508 983 5518 1017
rect 5552 983 5562 1017
rect 5308 843 5318 877
rect 5352 843 5362 877
rect 5108 703 5118 737
rect 5152 703 5162 737
rect 4908 563 4918 597
rect 4952 563 4962 597
rect 4708 423 4718 457
rect 4752 423 4762 457
rect 4508 283 4518 317
rect 4552 283 4562 317
rect 4308 143 4318 177
rect 4352 143 4362 177
rect 4202 79 4268 80
rect 4202 27 4209 79
rect 4261 27 4268 79
rect 4202 26 4268 27
rect 4108 -67 4109 -15
rect 4161 -67 4162 -15
rect 4108 -79 4118 -67
rect 4152 -79 4162 -67
rect 3908 -132 3962 -131
rect 3908 -143 3918 -132
rect 3952 -143 3962 -132
rect 3908 -195 3909 -143
rect 3961 -195 3962 -143
rect 3908 -210 3962 -195
rect 4012 -133 4058 -81
rect 4012 -167 4018 -133
rect 4052 -167 4058 -133
rect 3918 -291 3925 -239
rect 3977 -291 3984 -239
rect 3812 -397 3818 -363
rect 3852 -397 3858 -363
rect 3812 -435 3858 -397
rect 3812 -469 3818 -435
rect 3852 -469 3858 -435
rect 3812 -512 3858 -469
rect 3909 -326 3961 -320
rect 3909 -390 3918 -378
rect 3952 -390 3961 -378
rect 3909 -454 3918 -442
rect 3952 -454 3961 -442
rect 3909 -555 3961 -506
rect 4012 -363 4058 -167
rect 4108 -131 4109 -79
rect 4161 -131 4162 -79
rect 4208 -22 4262 26
rect 4208 -74 4209 -22
rect 4261 -74 4262 -22
rect 4208 -81 4262 -74
rect 4308 -15 4362 143
rect 4408 177 4462 189
rect 4408 151 4418 177
rect 4452 151 4462 177
rect 4408 99 4409 151
rect 4461 99 4462 151
rect 4408 92 4462 99
rect 4508 177 4562 283
rect 4608 361 4662 368
rect 4608 309 4609 361
rect 4661 309 4662 361
rect 4608 283 4618 309
rect 4652 283 4662 309
rect 4608 271 4662 283
rect 4708 317 4762 423
rect 4808 457 4862 469
rect 4808 431 4818 457
rect 4852 431 4862 457
rect 4808 379 4809 431
rect 4861 379 4862 431
rect 4808 372 4862 379
rect 4908 457 4962 563
rect 5008 641 5062 648
rect 5008 589 5009 641
rect 5061 589 5062 641
rect 5008 563 5018 589
rect 5052 563 5062 589
rect 5008 551 5062 563
rect 5108 597 5162 703
rect 5208 737 5262 749
rect 5208 711 5218 737
rect 5252 711 5262 737
rect 5208 659 5209 711
rect 5261 659 5262 711
rect 5208 652 5262 659
rect 5308 737 5362 843
rect 5408 921 5462 928
rect 5408 869 5409 921
rect 5461 869 5462 921
rect 5408 843 5418 869
rect 5452 843 5462 869
rect 5408 831 5462 843
rect 5508 877 5562 983
rect 5608 1017 5662 1029
rect 5608 991 5618 1017
rect 5652 991 5662 1017
rect 5608 939 5609 991
rect 5661 939 5662 991
rect 5608 932 5662 939
rect 5708 1017 5762 1123
rect 5808 1201 5862 1208
rect 5808 1149 5809 1201
rect 5861 1149 5862 1201
rect 5808 1123 5818 1149
rect 5852 1123 5862 1149
rect 5808 1111 5862 1123
rect 5908 1157 5962 1353
rect 6008 1387 6062 1399
rect 6008 1361 6018 1387
rect 6052 1361 6062 1387
rect 6008 1309 6009 1361
rect 6061 1309 6062 1361
rect 6008 1302 6062 1309
rect 6108 1387 6162 1493
rect 6208 1571 6262 1578
rect 6208 1519 6209 1571
rect 6261 1519 6262 1571
rect 6208 1493 6218 1519
rect 6252 1493 6262 1519
rect 6208 1481 6262 1493
rect 6308 1527 6362 1633
rect 6408 1667 6462 1679
rect 6408 1641 6418 1667
rect 6452 1641 6462 1667
rect 6408 1589 6409 1641
rect 6461 1589 6462 1641
rect 6408 1582 6462 1589
rect 6506 1648 6516 1682
rect 6550 1648 6560 1682
rect 6506 1641 6560 1648
rect 6506 1589 6507 1641
rect 6559 1589 6560 1641
rect 6506 1582 6560 1589
rect 6506 1542 6560 1554
rect 6308 1493 6318 1527
rect 6352 1493 6362 1527
rect 6108 1353 6118 1387
rect 6152 1353 6162 1387
rect 6002 1273 6068 1274
rect 6002 1221 6009 1273
rect 6061 1221 6068 1273
rect 6002 1220 6068 1221
rect 5908 1123 5918 1157
rect 5952 1123 5962 1157
rect 5708 983 5718 1017
rect 5752 983 5762 1017
rect 5508 843 5518 877
rect 5552 843 5562 877
rect 5308 703 5318 737
rect 5352 703 5362 737
rect 5108 563 5118 597
rect 5152 563 5162 597
rect 4908 423 4918 457
rect 4952 423 4962 457
rect 4708 283 4718 317
rect 4752 283 4762 317
rect 4508 143 4518 177
rect 4552 143 4562 177
rect 4402 63 4468 64
rect 4402 11 4409 63
rect 4461 11 4468 63
rect 4402 10 4468 11
rect 4308 -67 4309 -15
rect 4361 -67 4362 -15
rect 4308 -79 4318 -67
rect 4352 -79 4362 -67
rect 4108 -132 4162 -131
rect 4108 -143 4118 -132
rect 4152 -143 4162 -132
rect 4108 -195 4109 -143
rect 4161 -195 4162 -143
rect 4108 -210 4162 -195
rect 4212 -133 4258 -81
rect 4212 -167 4218 -133
rect 4252 -167 4258 -133
rect 4118 -291 4125 -239
rect 4177 -291 4184 -239
rect 4012 -397 4018 -363
rect 4052 -397 4058 -363
rect 4012 -435 4058 -397
rect 4012 -469 4018 -435
rect 4052 -469 4058 -435
rect 4012 -512 4058 -469
rect 4109 -326 4161 -320
rect 4109 -390 4118 -378
rect 4152 -390 4161 -378
rect 4109 -454 4118 -442
rect 4152 -454 4161 -442
rect 4109 -512 4161 -506
rect 4212 -363 4258 -167
rect 4308 -131 4309 -79
rect 4361 -131 4362 -79
rect 4408 -22 4462 10
rect 4408 -74 4409 -22
rect 4461 -74 4462 -22
rect 4408 -81 4462 -74
rect 4508 -15 4562 143
rect 4608 221 4662 228
rect 4608 169 4609 221
rect 4661 169 4662 221
rect 4608 143 4618 169
rect 4652 143 4662 169
rect 4608 131 4662 143
rect 4708 177 4762 283
rect 4808 317 4862 329
rect 4808 291 4818 317
rect 4852 291 4862 317
rect 4808 239 4809 291
rect 4861 239 4862 291
rect 4808 232 4862 239
rect 4908 317 4962 423
rect 5008 501 5062 508
rect 5008 449 5009 501
rect 5061 449 5062 501
rect 5008 423 5018 449
rect 5052 423 5062 449
rect 5008 411 5062 423
rect 5108 457 5162 563
rect 5208 597 5262 609
rect 5208 571 5218 597
rect 5252 571 5262 597
rect 5208 519 5209 571
rect 5261 519 5262 571
rect 5208 512 5262 519
rect 5308 597 5362 703
rect 5408 781 5462 788
rect 5408 729 5409 781
rect 5461 729 5462 781
rect 5408 703 5418 729
rect 5452 703 5462 729
rect 5408 691 5462 703
rect 5508 737 5562 843
rect 5608 877 5662 889
rect 5608 851 5618 877
rect 5652 851 5662 877
rect 5608 799 5609 851
rect 5661 799 5662 851
rect 5608 792 5662 799
rect 5708 877 5762 983
rect 5808 1061 5862 1068
rect 5808 1009 5809 1061
rect 5861 1009 5862 1061
rect 5808 983 5818 1009
rect 5852 983 5862 1009
rect 5808 971 5862 983
rect 5908 1017 5962 1123
rect 6008 1157 6062 1169
rect 6008 1131 6018 1157
rect 6052 1131 6062 1157
rect 6008 1079 6009 1131
rect 6061 1079 6062 1131
rect 6008 1072 6062 1079
rect 6108 1157 6162 1353
rect 6208 1431 6262 1438
rect 6208 1379 6209 1431
rect 6261 1379 6262 1431
rect 6208 1353 6218 1379
rect 6252 1353 6262 1379
rect 6208 1341 6262 1353
rect 6308 1387 6362 1493
rect 6408 1527 6462 1539
rect 6408 1501 6418 1527
rect 6452 1501 6462 1527
rect 6408 1449 6409 1501
rect 6461 1449 6462 1501
rect 6408 1442 6462 1449
rect 6506 1508 6516 1542
rect 6550 1508 6560 1542
rect 6506 1501 6560 1508
rect 6506 1449 6507 1501
rect 6559 1449 6560 1501
rect 6506 1442 6560 1449
rect 6506 1402 6560 1414
rect 6308 1353 6318 1387
rect 6352 1353 6362 1387
rect 6202 1289 6268 1290
rect 6202 1237 6209 1289
rect 6261 1237 6268 1289
rect 6202 1236 6268 1237
rect 6108 1123 6118 1157
rect 6152 1123 6162 1157
rect 5908 983 5918 1017
rect 5952 983 5962 1017
rect 5708 843 5718 877
rect 5752 843 5762 877
rect 5508 703 5518 737
rect 5552 703 5562 737
rect 5308 563 5318 597
rect 5352 563 5362 597
rect 5108 423 5118 457
rect 5152 423 5162 457
rect 4908 283 4918 317
rect 4952 283 4962 317
rect 4708 143 4718 177
rect 4752 143 4762 177
rect 4602 79 4668 80
rect 4602 27 4609 79
rect 4661 27 4668 79
rect 4602 26 4668 27
rect 4508 -67 4509 -15
rect 4561 -67 4562 -15
rect 4508 -79 4518 -67
rect 4552 -79 4562 -67
rect 4308 -132 4362 -131
rect 4308 -143 4318 -132
rect 4352 -143 4362 -132
rect 4308 -195 4309 -143
rect 4361 -195 4362 -143
rect 4308 -210 4362 -195
rect 4412 -133 4458 -81
rect 4412 -167 4418 -133
rect 4452 -167 4458 -133
rect 4318 -291 4325 -239
rect 4377 -291 4384 -239
rect 4212 -397 4218 -363
rect 4252 -397 4258 -363
rect 4212 -435 4258 -397
rect 4212 -469 4218 -435
rect 4252 -469 4258 -435
rect 4212 -512 4258 -469
rect 4309 -326 4361 -320
rect 4309 -390 4318 -378
rect 4352 -390 4361 -378
rect 4309 -454 4318 -442
rect 4352 -454 4361 -442
rect 4309 -555 4361 -506
rect 4412 -363 4458 -167
rect 4508 -131 4509 -79
rect 4561 -131 4562 -79
rect 4608 -22 4662 26
rect 4608 -74 4609 -22
rect 4661 -74 4662 -22
rect 4608 -81 4662 -74
rect 4708 -15 4762 143
rect 4808 177 4862 189
rect 4808 151 4818 177
rect 4852 151 4862 177
rect 4808 99 4809 151
rect 4861 99 4862 151
rect 4808 92 4862 99
rect 4908 177 4962 283
rect 5008 361 5062 368
rect 5008 309 5009 361
rect 5061 309 5062 361
rect 5008 283 5018 309
rect 5052 283 5062 309
rect 5008 271 5062 283
rect 5108 317 5162 423
rect 5208 457 5262 469
rect 5208 431 5218 457
rect 5252 431 5262 457
rect 5208 379 5209 431
rect 5261 379 5262 431
rect 5208 372 5262 379
rect 5308 457 5362 563
rect 5408 641 5462 648
rect 5408 589 5409 641
rect 5461 589 5462 641
rect 5408 563 5418 589
rect 5452 563 5462 589
rect 5408 551 5462 563
rect 5508 597 5562 703
rect 5608 737 5662 749
rect 5608 711 5618 737
rect 5652 711 5662 737
rect 5608 659 5609 711
rect 5661 659 5662 711
rect 5608 652 5662 659
rect 5708 737 5762 843
rect 5808 921 5862 928
rect 5808 869 5809 921
rect 5861 869 5862 921
rect 5808 843 5818 869
rect 5852 843 5862 869
rect 5808 831 5862 843
rect 5908 877 5962 983
rect 6008 1017 6062 1029
rect 6008 991 6018 1017
rect 6052 991 6062 1017
rect 6008 939 6009 991
rect 6061 939 6062 991
rect 6008 932 6062 939
rect 6108 1017 6162 1123
rect 6208 1201 6262 1208
rect 6208 1149 6209 1201
rect 6261 1149 6262 1201
rect 6208 1123 6218 1149
rect 6252 1123 6262 1149
rect 6208 1111 6262 1123
rect 6308 1157 6362 1353
rect 6408 1387 6462 1399
rect 6408 1361 6418 1387
rect 6452 1361 6462 1387
rect 6408 1309 6409 1361
rect 6461 1309 6462 1361
rect 6408 1302 6462 1309
rect 6506 1368 6516 1402
rect 6550 1368 6560 1402
rect 6506 1361 6560 1368
rect 6506 1309 6507 1361
rect 6559 1309 6560 1361
rect 6506 1302 6560 1309
rect 6590 1267 6620 2431
rect 6504 1261 6620 1267
rect 6504 1227 6516 1261
rect 6550 1227 6620 1261
rect 6504 1221 6620 1227
rect 6506 1172 6560 1184
rect 6308 1123 6318 1157
rect 6352 1123 6362 1157
rect 6108 983 6118 1017
rect 6152 983 6162 1017
rect 5908 843 5918 877
rect 5952 843 5962 877
rect 5708 703 5718 737
rect 5752 703 5762 737
rect 5508 563 5518 597
rect 5552 563 5562 597
rect 5308 423 5318 457
rect 5352 423 5362 457
rect 5108 283 5118 317
rect 5152 283 5162 317
rect 4908 143 4918 177
rect 4952 143 4962 177
rect 4802 63 4868 64
rect 4802 11 4809 63
rect 4861 11 4868 63
rect 4802 10 4868 11
rect 4708 -67 4709 -15
rect 4761 -67 4762 -15
rect 4708 -79 4718 -67
rect 4752 -79 4762 -67
rect 4508 -132 4562 -131
rect 4508 -143 4518 -132
rect 4552 -143 4562 -132
rect 4508 -195 4509 -143
rect 4561 -195 4562 -143
rect 4508 -210 4562 -195
rect 4612 -133 4658 -81
rect 4612 -167 4618 -133
rect 4652 -167 4658 -133
rect 4518 -291 4525 -239
rect 4577 -291 4584 -239
rect 4412 -397 4418 -363
rect 4452 -397 4458 -363
rect 4412 -435 4458 -397
rect 4412 -469 4418 -435
rect 4452 -469 4458 -435
rect 4412 -512 4458 -469
rect 4509 -326 4561 -320
rect 4509 -390 4518 -378
rect 4552 -390 4561 -378
rect 4509 -454 4518 -442
rect 4552 -454 4561 -442
rect 4509 -512 4561 -506
rect 4612 -363 4658 -167
rect 4708 -131 4709 -79
rect 4761 -131 4762 -79
rect 4808 -22 4862 10
rect 4808 -74 4809 -22
rect 4861 -74 4862 -22
rect 4808 -81 4862 -74
rect 4908 -15 4962 143
rect 5008 221 5062 228
rect 5008 169 5009 221
rect 5061 169 5062 221
rect 5008 143 5018 169
rect 5052 143 5062 169
rect 5008 131 5062 143
rect 5108 177 5162 283
rect 5208 317 5262 329
rect 5208 291 5218 317
rect 5252 291 5262 317
rect 5208 239 5209 291
rect 5261 239 5262 291
rect 5208 232 5262 239
rect 5308 317 5362 423
rect 5408 501 5462 508
rect 5408 449 5409 501
rect 5461 449 5462 501
rect 5408 423 5418 449
rect 5452 423 5462 449
rect 5408 411 5462 423
rect 5508 457 5562 563
rect 5608 597 5662 609
rect 5608 571 5618 597
rect 5652 571 5662 597
rect 5608 519 5609 571
rect 5661 519 5662 571
rect 5608 512 5662 519
rect 5708 597 5762 703
rect 5808 781 5862 788
rect 5808 729 5809 781
rect 5861 729 5862 781
rect 5808 703 5818 729
rect 5852 703 5862 729
rect 5808 691 5862 703
rect 5908 737 5962 843
rect 6008 877 6062 889
rect 6008 851 6018 877
rect 6052 851 6062 877
rect 6008 799 6009 851
rect 6061 799 6062 851
rect 6008 792 6062 799
rect 6108 877 6162 983
rect 6208 1061 6262 1068
rect 6208 1009 6209 1061
rect 6261 1009 6262 1061
rect 6208 983 6218 1009
rect 6252 983 6262 1009
rect 6208 971 6262 983
rect 6308 1017 6362 1123
rect 6408 1157 6462 1169
rect 6408 1131 6418 1157
rect 6452 1131 6462 1157
rect 6408 1079 6409 1131
rect 6461 1079 6462 1131
rect 6408 1072 6462 1079
rect 6506 1138 6516 1172
rect 6550 1138 6560 1172
rect 6506 1131 6560 1138
rect 6506 1079 6507 1131
rect 6559 1079 6560 1131
rect 6506 1072 6560 1079
rect 6506 1032 6560 1044
rect 6308 983 6318 1017
rect 6352 983 6362 1017
rect 6108 843 6118 877
rect 6152 843 6162 877
rect 5908 703 5918 737
rect 5952 703 5962 737
rect 5708 563 5718 597
rect 5752 563 5762 597
rect 5508 423 5518 457
rect 5552 423 5562 457
rect 5308 283 5318 317
rect 5352 283 5362 317
rect 5108 143 5118 177
rect 5152 143 5162 177
rect 5002 79 5068 80
rect 5002 27 5009 79
rect 5061 27 5068 79
rect 5002 26 5068 27
rect 4908 -67 4909 -15
rect 4961 -67 4962 -15
rect 4908 -79 4918 -67
rect 4952 -79 4962 -67
rect 4708 -132 4762 -131
rect 4708 -143 4718 -132
rect 4752 -143 4762 -132
rect 4708 -195 4709 -143
rect 4761 -195 4762 -143
rect 4708 -210 4762 -195
rect 4812 -133 4858 -81
rect 4812 -167 4818 -133
rect 4852 -167 4858 -133
rect 4718 -291 4725 -239
rect 4777 -291 4784 -239
rect 4612 -397 4618 -363
rect 4652 -397 4658 -363
rect 4612 -435 4658 -397
rect 4612 -469 4618 -435
rect 4652 -469 4658 -435
rect 4612 -512 4658 -469
rect 4709 -326 4761 -320
rect 4709 -390 4718 -378
rect 4752 -390 4761 -378
rect 4709 -454 4718 -442
rect 4752 -454 4761 -442
rect 4709 -555 4761 -506
rect 4812 -363 4858 -167
rect 4908 -131 4909 -79
rect 4961 -131 4962 -79
rect 5008 -22 5062 26
rect 5008 -74 5009 -22
rect 5061 -74 5062 -22
rect 5008 -81 5062 -74
rect 5108 -15 5162 143
rect 5208 177 5262 189
rect 5208 151 5218 177
rect 5252 151 5262 177
rect 5208 99 5209 151
rect 5261 99 5262 151
rect 5208 92 5262 99
rect 5308 177 5362 283
rect 5408 361 5462 368
rect 5408 309 5409 361
rect 5461 309 5462 361
rect 5408 283 5418 309
rect 5452 283 5462 309
rect 5408 271 5462 283
rect 5508 317 5562 423
rect 5608 457 5662 469
rect 5608 431 5618 457
rect 5652 431 5662 457
rect 5608 379 5609 431
rect 5661 379 5662 431
rect 5608 372 5662 379
rect 5708 457 5762 563
rect 5808 641 5862 648
rect 5808 589 5809 641
rect 5861 589 5862 641
rect 5808 563 5818 589
rect 5852 563 5862 589
rect 5808 551 5862 563
rect 5908 597 5962 703
rect 6008 737 6062 749
rect 6008 711 6018 737
rect 6052 711 6062 737
rect 6008 659 6009 711
rect 6061 659 6062 711
rect 6008 652 6062 659
rect 6108 737 6162 843
rect 6208 921 6262 928
rect 6208 869 6209 921
rect 6261 869 6262 921
rect 6208 843 6218 869
rect 6252 843 6262 869
rect 6208 831 6262 843
rect 6308 877 6362 983
rect 6408 1017 6462 1029
rect 6408 991 6418 1017
rect 6452 991 6462 1017
rect 6408 939 6409 991
rect 6461 939 6462 991
rect 6408 932 6462 939
rect 6506 998 6516 1032
rect 6550 998 6560 1032
rect 6506 991 6560 998
rect 6506 939 6507 991
rect 6559 939 6560 991
rect 6506 932 6560 939
rect 6506 892 6560 904
rect 6308 843 6318 877
rect 6352 843 6362 877
rect 6108 703 6118 737
rect 6152 703 6162 737
rect 5908 563 5918 597
rect 5952 563 5962 597
rect 5708 423 5718 457
rect 5752 423 5762 457
rect 5508 283 5518 317
rect 5552 283 5562 317
rect 5308 143 5318 177
rect 5352 143 5362 177
rect 5202 63 5268 64
rect 5202 11 5209 63
rect 5261 11 5268 63
rect 5202 10 5268 11
rect 5108 -67 5109 -15
rect 5161 -67 5162 -15
rect 5108 -79 5118 -67
rect 5152 -79 5162 -67
rect 4908 -132 4962 -131
rect 4908 -143 4918 -132
rect 4952 -143 4962 -132
rect 4908 -195 4909 -143
rect 4961 -195 4962 -143
rect 4908 -210 4962 -195
rect 5012 -133 5058 -81
rect 5012 -167 5018 -133
rect 5052 -167 5058 -133
rect 4918 -291 4925 -239
rect 4977 -291 4984 -239
rect 4812 -397 4818 -363
rect 4852 -397 4858 -363
rect 4812 -435 4858 -397
rect 4812 -469 4818 -435
rect 4852 -469 4858 -435
rect 4812 -512 4858 -469
rect 4909 -326 4961 -320
rect 4909 -390 4918 -378
rect 4952 -390 4961 -378
rect 4909 -454 4918 -442
rect 4952 -454 4961 -442
rect 4909 -512 4961 -506
rect 5012 -363 5058 -167
rect 5108 -131 5109 -79
rect 5161 -131 5162 -79
rect 5208 -22 5262 10
rect 5208 -74 5209 -22
rect 5261 -74 5262 -22
rect 5208 -81 5262 -74
rect 5308 -15 5362 143
rect 5408 221 5462 228
rect 5408 169 5409 221
rect 5461 169 5462 221
rect 5408 143 5418 169
rect 5452 143 5462 169
rect 5408 131 5462 143
rect 5508 177 5562 283
rect 5608 317 5662 329
rect 5608 291 5618 317
rect 5652 291 5662 317
rect 5608 239 5609 291
rect 5661 239 5662 291
rect 5608 232 5662 239
rect 5708 317 5762 423
rect 5808 501 5862 508
rect 5808 449 5809 501
rect 5861 449 5862 501
rect 5808 423 5818 449
rect 5852 423 5862 449
rect 5808 411 5862 423
rect 5908 457 5962 563
rect 6008 597 6062 609
rect 6008 571 6018 597
rect 6052 571 6062 597
rect 6008 519 6009 571
rect 6061 519 6062 571
rect 6008 512 6062 519
rect 6108 597 6162 703
rect 6208 781 6262 788
rect 6208 729 6209 781
rect 6261 729 6262 781
rect 6208 703 6218 729
rect 6252 703 6262 729
rect 6208 691 6262 703
rect 6308 737 6362 843
rect 6408 877 6462 889
rect 6408 851 6418 877
rect 6452 851 6462 877
rect 6408 799 6409 851
rect 6461 799 6462 851
rect 6408 792 6462 799
rect 6506 858 6516 892
rect 6550 858 6560 892
rect 6506 851 6560 858
rect 6506 799 6507 851
rect 6559 799 6560 851
rect 6506 792 6560 799
rect 6506 752 6560 764
rect 6308 703 6318 737
rect 6352 703 6362 737
rect 6108 563 6118 597
rect 6152 563 6162 597
rect 5908 423 5918 457
rect 5952 423 5962 457
rect 5708 283 5718 317
rect 5752 283 5762 317
rect 5508 143 5518 177
rect 5552 143 5562 177
rect 5402 79 5468 80
rect 5402 27 5409 79
rect 5461 27 5468 79
rect 5402 26 5468 27
rect 5308 -67 5309 -15
rect 5361 -67 5362 -15
rect 5308 -79 5318 -67
rect 5352 -79 5362 -67
rect 5108 -132 5162 -131
rect 5108 -143 5118 -132
rect 5152 -143 5162 -132
rect 5108 -195 5109 -143
rect 5161 -195 5162 -143
rect 5108 -210 5162 -195
rect 5212 -133 5258 -81
rect 5212 -167 5218 -133
rect 5252 -167 5258 -133
rect 5118 -291 5125 -239
rect 5177 -291 5184 -239
rect 5012 -397 5018 -363
rect 5052 -397 5058 -363
rect 5012 -435 5058 -397
rect 5012 -469 5018 -435
rect 5052 -469 5058 -435
rect 5012 -512 5058 -469
rect 5109 -326 5161 -320
rect 5109 -390 5118 -378
rect 5152 -390 5161 -378
rect 5109 -454 5118 -442
rect 5152 -454 5161 -442
rect 5109 -555 5161 -506
rect 5212 -363 5258 -167
rect 5308 -131 5309 -79
rect 5361 -131 5362 -79
rect 5408 -22 5462 26
rect 5408 -74 5409 -22
rect 5461 -74 5462 -22
rect 5408 -81 5462 -74
rect 5508 -15 5562 143
rect 5608 177 5662 189
rect 5608 151 5618 177
rect 5652 151 5662 177
rect 5608 99 5609 151
rect 5661 99 5662 151
rect 5608 92 5662 99
rect 5708 177 5762 283
rect 5808 361 5862 368
rect 5808 309 5809 361
rect 5861 309 5862 361
rect 5808 283 5818 309
rect 5852 283 5862 309
rect 5808 271 5862 283
rect 5908 317 5962 423
rect 6008 457 6062 469
rect 6008 431 6018 457
rect 6052 431 6062 457
rect 6008 379 6009 431
rect 6061 379 6062 431
rect 6008 372 6062 379
rect 6108 457 6162 563
rect 6208 641 6262 648
rect 6208 589 6209 641
rect 6261 589 6262 641
rect 6208 563 6218 589
rect 6252 563 6262 589
rect 6208 551 6262 563
rect 6308 597 6362 703
rect 6408 737 6462 749
rect 6408 711 6418 737
rect 6452 711 6462 737
rect 6408 659 6409 711
rect 6461 659 6462 711
rect 6408 652 6462 659
rect 6506 718 6516 752
rect 6550 718 6560 752
rect 6506 711 6560 718
rect 6506 659 6507 711
rect 6559 659 6560 711
rect 6506 652 6560 659
rect 6506 612 6560 624
rect 6308 563 6318 597
rect 6352 563 6362 597
rect 6108 423 6118 457
rect 6152 423 6162 457
rect 5908 283 5918 317
rect 5952 283 5962 317
rect 5708 143 5718 177
rect 5752 143 5762 177
rect 5602 63 5668 64
rect 5602 11 5609 63
rect 5661 11 5668 63
rect 5602 10 5668 11
rect 5508 -67 5509 -15
rect 5561 -67 5562 -15
rect 5508 -79 5518 -67
rect 5552 -79 5562 -67
rect 5308 -132 5362 -131
rect 5308 -143 5318 -132
rect 5352 -143 5362 -132
rect 5308 -195 5309 -143
rect 5361 -195 5362 -143
rect 5308 -210 5362 -195
rect 5412 -133 5458 -81
rect 5412 -167 5418 -133
rect 5452 -167 5458 -133
rect 5318 -291 5325 -239
rect 5377 -291 5384 -239
rect 5212 -397 5218 -363
rect 5252 -397 5258 -363
rect 5212 -435 5258 -397
rect 5212 -469 5218 -435
rect 5252 -469 5258 -435
rect 5212 -512 5258 -469
rect 5309 -326 5361 -320
rect 5309 -390 5318 -378
rect 5352 -390 5361 -378
rect 5309 -454 5318 -442
rect 5352 -454 5361 -442
rect 5309 -512 5361 -506
rect 5412 -363 5458 -167
rect 5508 -131 5509 -79
rect 5561 -131 5562 -79
rect 5608 -22 5662 10
rect 5608 -74 5609 -22
rect 5661 -74 5662 -22
rect 5608 -81 5662 -74
rect 5708 -15 5762 143
rect 5808 221 5862 228
rect 5808 169 5809 221
rect 5861 169 5862 221
rect 5808 143 5818 169
rect 5852 143 5862 169
rect 5808 131 5862 143
rect 5908 177 5962 283
rect 6008 317 6062 329
rect 6008 291 6018 317
rect 6052 291 6062 317
rect 6008 239 6009 291
rect 6061 239 6062 291
rect 6008 232 6062 239
rect 6108 317 6162 423
rect 6208 501 6262 508
rect 6208 449 6209 501
rect 6261 449 6262 501
rect 6208 423 6218 449
rect 6252 423 6262 449
rect 6208 411 6262 423
rect 6308 457 6362 563
rect 6408 597 6462 609
rect 6408 571 6418 597
rect 6452 571 6462 597
rect 6408 519 6409 571
rect 6461 519 6462 571
rect 6408 512 6462 519
rect 6506 578 6516 612
rect 6550 578 6560 612
rect 6506 571 6560 578
rect 6506 519 6507 571
rect 6559 519 6560 571
rect 6506 512 6560 519
rect 6506 472 6560 484
rect 6308 423 6318 457
rect 6352 423 6362 457
rect 6108 283 6118 317
rect 6152 283 6162 317
rect 5908 143 5918 177
rect 5952 143 5962 177
rect 5802 79 5868 80
rect 5802 27 5809 79
rect 5861 27 5868 79
rect 5802 26 5868 27
rect 5708 -67 5709 -15
rect 5761 -67 5762 -15
rect 5708 -79 5718 -67
rect 5752 -79 5762 -67
rect 5508 -132 5562 -131
rect 5508 -143 5518 -132
rect 5552 -143 5562 -132
rect 5508 -195 5509 -143
rect 5561 -195 5562 -143
rect 5508 -210 5562 -195
rect 5612 -133 5658 -81
rect 5612 -167 5618 -133
rect 5652 -167 5658 -133
rect 5518 -291 5525 -239
rect 5577 -291 5584 -239
rect 5412 -397 5418 -363
rect 5452 -397 5458 -363
rect 5412 -435 5458 -397
rect 5412 -469 5418 -435
rect 5452 -469 5458 -435
rect 5412 -512 5458 -469
rect 5509 -326 5561 -320
rect 5509 -390 5518 -378
rect 5552 -390 5561 -378
rect 5509 -454 5518 -442
rect 5552 -454 5561 -442
rect 5509 -555 5561 -506
rect 5612 -363 5658 -167
rect 5708 -131 5709 -79
rect 5761 -131 5762 -79
rect 5808 -22 5862 26
rect 5808 -74 5809 -22
rect 5861 -74 5862 -22
rect 5808 -81 5862 -74
rect 5908 -15 5962 143
rect 6008 177 6062 189
rect 6008 151 6018 177
rect 6052 151 6062 177
rect 6008 99 6009 151
rect 6061 99 6062 151
rect 6008 92 6062 99
rect 6108 177 6162 283
rect 6208 361 6262 368
rect 6208 309 6209 361
rect 6261 309 6262 361
rect 6208 283 6218 309
rect 6252 283 6262 309
rect 6208 271 6262 283
rect 6308 317 6362 423
rect 6408 457 6462 469
rect 6408 431 6418 457
rect 6452 431 6462 457
rect 6408 379 6409 431
rect 6461 379 6462 431
rect 6408 372 6462 379
rect 6506 438 6516 472
rect 6550 438 6560 472
rect 6506 431 6560 438
rect 6506 379 6507 431
rect 6559 379 6560 431
rect 6506 372 6560 379
rect 6506 332 6560 344
rect 6308 283 6318 317
rect 6352 283 6362 317
rect 6108 143 6118 177
rect 6152 143 6162 177
rect 6002 63 6068 64
rect 6002 11 6009 63
rect 6061 11 6068 63
rect 6002 10 6068 11
rect 5908 -67 5909 -15
rect 5961 -67 5962 -15
rect 5908 -79 5918 -67
rect 5952 -79 5962 -67
rect 5708 -132 5762 -131
rect 5708 -143 5718 -132
rect 5752 -143 5762 -132
rect 5708 -195 5709 -143
rect 5761 -195 5762 -143
rect 5708 -210 5762 -195
rect 5812 -133 5858 -81
rect 5812 -167 5818 -133
rect 5852 -167 5858 -133
rect 5718 -291 5725 -239
rect 5777 -291 5784 -239
rect 5612 -397 5618 -363
rect 5652 -397 5658 -363
rect 5612 -435 5658 -397
rect 5612 -469 5618 -435
rect 5652 -469 5658 -435
rect 5612 -512 5658 -469
rect 5709 -326 5761 -320
rect 5709 -390 5718 -378
rect 5752 -390 5761 -378
rect 5709 -454 5718 -442
rect 5752 -454 5761 -442
rect 5709 -512 5761 -506
rect 5812 -363 5858 -167
rect 5908 -131 5909 -79
rect 5961 -131 5962 -79
rect 6008 -22 6062 10
rect 6008 -74 6009 -22
rect 6061 -74 6062 -22
rect 6008 -81 6062 -74
rect 6108 -15 6162 143
rect 6208 221 6262 228
rect 6208 169 6209 221
rect 6261 169 6262 221
rect 6208 143 6218 169
rect 6252 143 6262 169
rect 6208 131 6262 143
rect 6308 177 6362 283
rect 6408 317 6462 329
rect 6408 291 6418 317
rect 6452 291 6462 317
rect 6408 239 6409 291
rect 6461 239 6462 291
rect 6408 232 6462 239
rect 6506 298 6516 332
rect 6550 298 6560 332
rect 6506 291 6560 298
rect 6506 239 6507 291
rect 6559 239 6560 291
rect 6506 232 6560 239
rect 6506 192 6560 204
rect 6308 143 6318 177
rect 6352 143 6362 177
rect 6202 79 6268 80
rect 6202 27 6209 79
rect 6261 27 6268 79
rect 6202 26 6268 27
rect 6108 -67 6109 -15
rect 6161 -67 6162 -15
rect 6108 -79 6118 -67
rect 6152 -79 6162 -67
rect 5908 -132 5962 -131
rect 5908 -143 5918 -132
rect 5952 -143 5962 -132
rect 5908 -195 5909 -143
rect 5961 -195 5962 -143
rect 5908 -210 5962 -195
rect 6012 -133 6058 -81
rect 6012 -167 6018 -133
rect 6052 -167 6058 -133
rect 5918 -291 5925 -239
rect 5977 -291 5984 -239
rect 5812 -397 5818 -363
rect 5852 -397 5858 -363
rect 5812 -435 5858 -397
rect 5812 -469 5818 -435
rect 5852 -469 5858 -435
rect 5812 -512 5858 -469
rect 5909 -326 5961 -320
rect 5909 -390 5918 -378
rect 5952 -390 5961 -378
rect 5909 -454 5918 -442
rect 5952 -454 5961 -442
rect 5909 -555 5961 -506
rect 6012 -363 6058 -167
rect 6108 -131 6109 -79
rect 6161 -131 6162 -79
rect 6208 -22 6262 26
rect 6208 -74 6209 -22
rect 6261 -74 6262 -22
rect 6208 -81 6262 -74
rect 6308 -15 6362 143
rect 6408 177 6462 189
rect 6408 151 6418 177
rect 6452 151 6462 177
rect 6408 99 6409 151
rect 6461 99 6462 151
rect 6408 92 6462 99
rect 6506 158 6516 192
rect 6550 158 6560 192
rect 6506 151 6560 158
rect 6506 99 6507 151
rect 6559 99 6560 151
rect 6506 92 6560 99
rect 6590 57 6620 1221
rect 6504 51 6620 57
rect 6504 17 6516 51
rect 6550 17 6620 51
rect 6504 11 6620 17
rect 6590 0 6620 11
rect 6650 9899 6680 10050
rect 6880 9900 6910 10050
rect 6980 9900 7010 10050
rect 7080 9900 7110 10050
rect 7180 9900 7210 10050
rect 7280 9900 7310 10050
rect 7380 9900 7410 10050
rect 6650 9893 6766 9899
rect 6650 9859 6720 9893
rect 6754 9859 6766 9893
rect 6650 9853 6766 9859
rect 6872 9888 6918 9900
rect 6872 9854 6878 9888
rect 6912 9854 6918 9888
rect 6650 8689 6680 9853
rect 6872 9842 6918 9854
rect 6972 9888 7018 9900
rect 6972 9854 6978 9888
rect 7012 9854 7018 9888
rect 6972 9842 7018 9854
rect 7072 9888 7118 9900
rect 7072 9854 7078 9888
rect 7112 9854 7118 9888
rect 7072 9842 7118 9854
rect 7172 9888 7218 9900
rect 7172 9854 7178 9888
rect 7212 9854 7218 9888
rect 7172 9842 7218 9854
rect 7272 9888 7318 9900
rect 7272 9854 7278 9888
rect 7312 9854 7318 9888
rect 7272 9842 7318 9854
rect 7372 9888 7418 9900
rect 7372 9854 7378 9888
rect 7412 9854 7418 9888
rect 7372 9842 7418 9854
rect 6710 9811 6764 9818
rect 6710 9759 6711 9811
rect 6763 9759 6764 9811
rect 6710 9752 6764 9759
rect 6710 9718 6720 9752
rect 6754 9718 6764 9752
rect 6710 9706 6764 9718
rect 6710 9671 6764 9678
rect 6710 9619 6711 9671
rect 6763 9619 6764 9671
rect 6710 9612 6764 9619
rect 6710 9578 6720 9612
rect 6754 9578 6764 9612
rect 6710 9566 6764 9578
rect 6710 9531 6764 9538
rect 6710 9479 6711 9531
rect 6763 9479 6764 9531
rect 6710 9472 6764 9479
rect 6710 9438 6720 9472
rect 6754 9438 6764 9472
rect 6710 9426 6764 9438
rect 6710 9391 6764 9398
rect 6710 9339 6711 9391
rect 6763 9339 6764 9391
rect 6710 9332 6764 9339
rect 6710 9298 6720 9332
rect 6754 9298 6764 9332
rect 6710 9286 6764 9298
rect 6710 9251 6764 9258
rect 6710 9199 6711 9251
rect 6763 9199 6764 9251
rect 6710 9192 6764 9199
rect 6710 9158 6720 9192
rect 6754 9158 6764 9192
rect 6710 9146 6764 9158
rect 6710 9111 6764 9118
rect 6710 9059 6711 9111
rect 6763 9059 6764 9111
rect 6710 9052 6764 9059
rect 6710 9018 6720 9052
rect 6754 9018 6764 9052
rect 6710 9006 6764 9018
rect 6710 8971 6764 8978
rect 6710 8919 6711 8971
rect 6763 8919 6764 8971
rect 6710 8912 6764 8919
rect 6710 8878 6720 8912
rect 6754 8878 6764 8912
rect 6710 8866 6764 8878
rect 6710 8831 6764 8838
rect 6710 8779 6711 8831
rect 6763 8779 6764 8831
rect 6710 8772 6764 8779
rect 6710 8738 6720 8772
rect 6754 8738 6764 8772
rect 6710 8726 6764 8738
rect 6880 8690 6910 9842
rect 6980 8690 7010 9842
rect 7080 8690 7110 9842
rect 7180 8690 7210 9842
rect 7280 8690 7310 9842
rect 7380 8690 7410 9842
rect 6650 8683 6766 8689
rect 6650 8649 6720 8683
rect 6754 8649 6766 8683
rect 6650 8643 6766 8649
rect 6872 8678 6918 8690
rect 6872 8644 6878 8678
rect 6912 8644 6918 8678
rect 6650 7479 6680 8643
rect 6872 8632 6918 8644
rect 6972 8678 7018 8690
rect 6972 8644 6978 8678
rect 7012 8644 7018 8678
rect 6972 8632 7018 8644
rect 7072 8678 7118 8690
rect 7072 8644 7078 8678
rect 7112 8644 7118 8678
rect 7072 8632 7118 8644
rect 7172 8678 7218 8690
rect 7172 8644 7178 8678
rect 7212 8644 7218 8678
rect 7172 8632 7218 8644
rect 7272 8678 7318 8690
rect 7272 8644 7278 8678
rect 7312 8644 7318 8678
rect 7272 8632 7318 8644
rect 7372 8678 7418 8690
rect 7372 8644 7378 8678
rect 7412 8644 7418 8678
rect 7372 8632 7418 8644
rect 6710 8601 6764 8608
rect 6710 8549 6711 8601
rect 6763 8549 6764 8601
rect 6710 8542 6764 8549
rect 6710 8508 6720 8542
rect 6754 8508 6764 8542
rect 6710 8496 6764 8508
rect 6710 8461 6764 8468
rect 6710 8409 6711 8461
rect 6763 8409 6764 8461
rect 6710 8402 6764 8409
rect 6710 8368 6720 8402
rect 6754 8368 6764 8402
rect 6710 8356 6764 8368
rect 6710 8321 6764 8328
rect 6710 8269 6711 8321
rect 6763 8269 6764 8321
rect 6710 8262 6764 8269
rect 6710 8228 6720 8262
rect 6754 8228 6764 8262
rect 6710 8216 6764 8228
rect 6710 8181 6764 8188
rect 6710 8129 6711 8181
rect 6763 8129 6764 8181
rect 6710 8122 6764 8129
rect 6710 8088 6720 8122
rect 6754 8088 6764 8122
rect 6710 8076 6764 8088
rect 6710 8041 6764 8048
rect 6710 7989 6711 8041
rect 6763 7989 6764 8041
rect 6710 7982 6764 7989
rect 6710 7948 6720 7982
rect 6754 7948 6764 7982
rect 6710 7936 6764 7948
rect 6710 7901 6764 7908
rect 6710 7849 6711 7901
rect 6763 7849 6764 7901
rect 6710 7842 6764 7849
rect 6710 7808 6720 7842
rect 6754 7808 6764 7842
rect 6710 7796 6764 7808
rect 6710 7761 6764 7768
rect 6710 7709 6711 7761
rect 6763 7709 6764 7761
rect 6710 7702 6764 7709
rect 6710 7668 6720 7702
rect 6754 7668 6764 7702
rect 6710 7656 6764 7668
rect 6710 7621 6764 7628
rect 6710 7569 6711 7621
rect 6763 7569 6764 7621
rect 6710 7562 6764 7569
rect 6710 7528 6720 7562
rect 6754 7528 6764 7562
rect 6710 7516 6764 7528
rect 6880 7480 6910 8632
rect 6980 7480 7010 8632
rect 7080 7480 7110 8632
rect 7180 7480 7210 8632
rect 7280 7480 7310 8632
rect 7380 7480 7410 8632
rect 6650 7473 6766 7479
rect 6650 7439 6720 7473
rect 6754 7439 6766 7473
rect 6650 7433 6766 7439
rect 6872 7468 6918 7480
rect 6872 7434 6878 7468
rect 6912 7434 6918 7468
rect 6650 6269 6680 7433
rect 6872 7422 6918 7434
rect 6972 7468 7018 7480
rect 6972 7434 6978 7468
rect 7012 7434 7018 7468
rect 6972 7422 7018 7434
rect 7072 7468 7118 7480
rect 7072 7434 7078 7468
rect 7112 7434 7118 7468
rect 7072 7422 7118 7434
rect 7172 7468 7218 7480
rect 7172 7434 7178 7468
rect 7212 7434 7218 7468
rect 7172 7422 7218 7434
rect 7272 7468 7318 7480
rect 7272 7434 7278 7468
rect 7312 7434 7318 7468
rect 7272 7422 7318 7434
rect 7372 7468 7418 7480
rect 7372 7434 7378 7468
rect 7412 7434 7418 7468
rect 7372 7422 7418 7434
rect 6710 7391 6764 7398
rect 6710 7339 6711 7391
rect 6763 7339 6764 7391
rect 6710 7332 6764 7339
rect 6710 7298 6720 7332
rect 6754 7298 6764 7332
rect 6710 7286 6764 7298
rect 6710 7251 6764 7258
rect 6710 7199 6711 7251
rect 6763 7199 6764 7251
rect 6710 7192 6764 7199
rect 6710 7158 6720 7192
rect 6754 7158 6764 7192
rect 6710 7146 6764 7158
rect 6710 7111 6764 7118
rect 6710 7059 6711 7111
rect 6763 7059 6764 7111
rect 6710 7052 6764 7059
rect 6710 7018 6720 7052
rect 6754 7018 6764 7052
rect 6710 7006 6764 7018
rect 6710 6971 6764 6978
rect 6710 6919 6711 6971
rect 6763 6919 6764 6971
rect 6710 6912 6764 6919
rect 6710 6878 6720 6912
rect 6754 6878 6764 6912
rect 6710 6866 6764 6878
rect 6710 6831 6764 6838
rect 6710 6779 6711 6831
rect 6763 6779 6764 6831
rect 6710 6772 6764 6779
rect 6710 6738 6720 6772
rect 6754 6738 6764 6772
rect 6710 6726 6764 6738
rect 6710 6691 6764 6698
rect 6710 6639 6711 6691
rect 6763 6639 6764 6691
rect 6710 6632 6764 6639
rect 6710 6598 6720 6632
rect 6754 6598 6764 6632
rect 6710 6586 6764 6598
rect 6710 6551 6764 6558
rect 6710 6499 6711 6551
rect 6763 6499 6764 6551
rect 6710 6492 6764 6499
rect 6710 6458 6720 6492
rect 6754 6458 6764 6492
rect 6710 6446 6764 6458
rect 6710 6411 6764 6418
rect 6710 6359 6711 6411
rect 6763 6359 6764 6411
rect 6710 6352 6764 6359
rect 6710 6318 6720 6352
rect 6754 6318 6764 6352
rect 6710 6306 6764 6318
rect 6880 6270 6910 7422
rect 6980 6270 7010 7422
rect 7080 6270 7110 7422
rect 7180 6270 7210 7422
rect 7280 6270 7310 7422
rect 7380 6270 7410 7422
rect 6650 6263 6766 6269
rect 6650 6229 6720 6263
rect 6754 6229 6766 6263
rect 6650 6223 6766 6229
rect 6872 6258 6918 6270
rect 6872 6224 6878 6258
rect 6912 6224 6918 6258
rect 6650 4919 6680 6223
rect 6872 6212 6918 6224
rect 6972 6258 7018 6270
rect 6972 6224 6978 6258
rect 7012 6224 7018 6258
rect 6972 6212 7018 6224
rect 7072 6258 7118 6270
rect 7072 6224 7078 6258
rect 7112 6224 7118 6258
rect 7072 6212 7118 6224
rect 7172 6258 7218 6270
rect 7172 6224 7178 6258
rect 7212 6224 7218 6258
rect 7172 6212 7218 6224
rect 7272 6258 7318 6270
rect 7272 6224 7278 6258
rect 7312 6224 7318 6258
rect 7272 6212 7318 6224
rect 7372 6258 7418 6270
rect 7372 6224 7378 6258
rect 7412 6224 7418 6258
rect 7372 6212 7418 6224
rect 6710 6181 6764 6188
rect 6710 6129 6711 6181
rect 6763 6129 6764 6181
rect 6710 6122 6764 6129
rect 6710 6088 6720 6122
rect 6754 6088 6764 6122
rect 6710 6076 6764 6088
rect 6710 6041 6764 6048
rect 6710 5989 6711 6041
rect 6763 5989 6764 6041
rect 6710 5982 6764 5989
rect 6710 5948 6720 5982
rect 6754 5948 6764 5982
rect 6710 5936 6764 5948
rect 6710 5901 6764 5908
rect 6710 5849 6711 5901
rect 6763 5849 6764 5901
rect 6710 5842 6764 5849
rect 6710 5808 6720 5842
rect 6754 5808 6764 5842
rect 6710 5796 6764 5808
rect 6710 5761 6764 5768
rect 6710 5709 6711 5761
rect 6763 5709 6764 5761
rect 6710 5702 6764 5709
rect 6710 5668 6720 5702
rect 6754 5668 6764 5702
rect 6710 5656 6764 5668
rect 6710 5621 6764 5628
rect 6710 5569 6711 5621
rect 6763 5569 6764 5621
rect 6710 5562 6764 5569
rect 6710 5528 6720 5562
rect 6754 5528 6764 5562
rect 6710 5516 6764 5528
rect 6710 5481 6764 5488
rect 6710 5429 6711 5481
rect 6763 5429 6764 5481
rect 6710 5422 6764 5429
rect 6710 5388 6720 5422
rect 6754 5388 6764 5422
rect 6710 5376 6764 5388
rect 6710 5341 6764 5348
rect 6710 5289 6711 5341
rect 6763 5289 6764 5341
rect 6710 5282 6764 5289
rect 6710 5248 6720 5282
rect 6754 5248 6764 5282
rect 6710 5236 6764 5248
rect 6710 5201 6764 5208
rect 6710 5149 6711 5201
rect 6763 5149 6764 5201
rect 6710 5142 6764 5149
rect 6710 5108 6720 5142
rect 6754 5108 6764 5142
rect 6710 5096 6764 5108
rect 6880 4920 6910 6212
rect 6980 4920 7010 6212
rect 7080 4920 7110 6212
rect 7180 4920 7210 6212
rect 7280 4920 7310 6212
rect 7380 4920 7410 6212
rect 6650 4913 6766 4919
rect 6650 4879 6720 4913
rect 6754 4879 6766 4913
rect 6650 4873 6766 4879
rect 6872 4908 6918 4920
rect 6872 4874 6878 4908
rect 6912 4874 6918 4908
rect 6650 3709 6680 4873
rect 6872 4862 6918 4874
rect 6972 4908 7018 4920
rect 6972 4874 6978 4908
rect 7012 4874 7018 4908
rect 6972 4862 7018 4874
rect 7072 4908 7118 4920
rect 7072 4874 7078 4908
rect 7112 4874 7118 4908
rect 7072 4862 7118 4874
rect 7172 4908 7218 4920
rect 7172 4874 7178 4908
rect 7212 4874 7218 4908
rect 7172 4862 7218 4874
rect 7272 4908 7318 4920
rect 7272 4874 7278 4908
rect 7312 4874 7318 4908
rect 7272 4862 7318 4874
rect 7372 4908 7418 4920
rect 7372 4874 7378 4908
rect 7412 4874 7418 4908
rect 7372 4862 7418 4874
rect 6710 4831 6764 4838
rect 6710 4779 6711 4831
rect 6763 4779 6764 4831
rect 6710 4772 6764 4779
rect 6710 4738 6720 4772
rect 6754 4738 6764 4772
rect 6710 4726 6764 4738
rect 6710 4691 6764 4698
rect 6710 4639 6711 4691
rect 6763 4639 6764 4691
rect 6710 4632 6764 4639
rect 6710 4598 6720 4632
rect 6754 4598 6764 4632
rect 6710 4586 6764 4598
rect 6710 4551 6764 4558
rect 6710 4499 6711 4551
rect 6763 4499 6764 4551
rect 6710 4492 6764 4499
rect 6710 4458 6720 4492
rect 6754 4458 6764 4492
rect 6710 4446 6764 4458
rect 6710 4411 6764 4418
rect 6710 4359 6711 4411
rect 6763 4359 6764 4411
rect 6710 4352 6764 4359
rect 6710 4318 6720 4352
rect 6754 4318 6764 4352
rect 6710 4306 6764 4318
rect 6710 4271 6764 4278
rect 6710 4219 6711 4271
rect 6763 4219 6764 4271
rect 6710 4212 6764 4219
rect 6710 4178 6720 4212
rect 6754 4178 6764 4212
rect 6710 4166 6764 4178
rect 6710 4131 6764 4138
rect 6710 4079 6711 4131
rect 6763 4079 6764 4131
rect 6710 4072 6764 4079
rect 6710 4038 6720 4072
rect 6754 4038 6764 4072
rect 6710 4026 6764 4038
rect 6710 3991 6764 3998
rect 6710 3939 6711 3991
rect 6763 3939 6764 3991
rect 6710 3932 6764 3939
rect 6710 3898 6720 3932
rect 6754 3898 6764 3932
rect 6710 3886 6764 3898
rect 6710 3851 6764 3858
rect 6710 3799 6711 3851
rect 6763 3799 6764 3851
rect 6710 3792 6764 3799
rect 6710 3758 6720 3792
rect 6754 3758 6764 3792
rect 6710 3746 6764 3758
rect 6880 3710 6910 4862
rect 6980 3710 7010 4862
rect 7080 3710 7110 4862
rect 7180 3710 7210 4862
rect 7280 3710 7310 4862
rect 7380 3710 7410 4862
rect 6650 3703 6766 3709
rect 6650 3669 6720 3703
rect 6754 3669 6766 3703
rect 6650 3663 6766 3669
rect 6872 3698 6918 3710
rect 6872 3664 6878 3698
rect 6912 3664 6918 3698
rect 6650 2499 6680 3663
rect 6872 3652 6918 3664
rect 6972 3698 7018 3710
rect 6972 3664 6978 3698
rect 7012 3664 7018 3698
rect 6972 3652 7018 3664
rect 7072 3698 7118 3710
rect 7072 3664 7078 3698
rect 7112 3664 7118 3698
rect 7072 3652 7118 3664
rect 7172 3698 7218 3710
rect 7172 3664 7178 3698
rect 7212 3664 7218 3698
rect 7172 3652 7218 3664
rect 7272 3698 7318 3710
rect 7272 3664 7278 3698
rect 7312 3664 7318 3698
rect 7272 3652 7318 3664
rect 7372 3698 7418 3710
rect 7372 3664 7378 3698
rect 7412 3664 7418 3698
rect 7372 3652 7418 3664
rect 6710 3621 6764 3628
rect 6710 3569 6711 3621
rect 6763 3569 6764 3621
rect 6710 3562 6764 3569
rect 6710 3528 6720 3562
rect 6754 3528 6764 3562
rect 6710 3516 6764 3528
rect 6710 3481 6764 3488
rect 6710 3429 6711 3481
rect 6763 3429 6764 3481
rect 6710 3422 6764 3429
rect 6710 3388 6720 3422
rect 6754 3388 6764 3422
rect 6710 3376 6764 3388
rect 6710 3341 6764 3348
rect 6710 3289 6711 3341
rect 6763 3289 6764 3341
rect 6710 3282 6764 3289
rect 6710 3248 6720 3282
rect 6754 3248 6764 3282
rect 6710 3236 6764 3248
rect 6710 3201 6764 3208
rect 6710 3149 6711 3201
rect 6763 3149 6764 3201
rect 6710 3142 6764 3149
rect 6710 3108 6720 3142
rect 6754 3108 6764 3142
rect 6710 3096 6764 3108
rect 6710 3061 6764 3068
rect 6710 3009 6711 3061
rect 6763 3009 6764 3061
rect 6710 3002 6764 3009
rect 6710 2968 6720 3002
rect 6754 2968 6764 3002
rect 6710 2956 6764 2968
rect 6710 2921 6764 2928
rect 6710 2869 6711 2921
rect 6763 2869 6764 2921
rect 6710 2862 6764 2869
rect 6710 2828 6720 2862
rect 6754 2828 6764 2862
rect 6710 2816 6764 2828
rect 6710 2781 6764 2788
rect 6710 2729 6711 2781
rect 6763 2729 6764 2781
rect 6710 2722 6764 2729
rect 6710 2688 6720 2722
rect 6754 2688 6764 2722
rect 6710 2676 6764 2688
rect 6710 2641 6764 2648
rect 6710 2589 6711 2641
rect 6763 2589 6764 2641
rect 6710 2582 6764 2589
rect 6710 2548 6720 2582
rect 6754 2548 6764 2582
rect 6710 2536 6764 2548
rect 6880 2500 6910 3652
rect 6980 2500 7010 3652
rect 7080 2500 7110 3652
rect 7180 2500 7210 3652
rect 7280 2500 7310 3652
rect 7380 2500 7410 3652
rect 6650 2493 6766 2499
rect 6650 2459 6720 2493
rect 6754 2459 6766 2493
rect 6650 2453 6766 2459
rect 6872 2488 6918 2500
rect 6872 2454 6878 2488
rect 6912 2454 6918 2488
rect 6650 1289 6680 2453
rect 6872 2442 6918 2454
rect 6972 2488 7018 2500
rect 6972 2454 6978 2488
rect 7012 2454 7018 2488
rect 6972 2442 7018 2454
rect 7072 2488 7118 2500
rect 7072 2454 7078 2488
rect 7112 2454 7118 2488
rect 7072 2442 7118 2454
rect 7172 2488 7218 2500
rect 7172 2454 7178 2488
rect 7212 2454 7218 2488
rect 7172 2442 7218 2454
rect 7272 2488 7318 2500
rect 7272 2454 7278 2488
rect 7312 2454 7318 2488
rect 7272 2442 7318 2454
rect 7372 2488 7418 2500
rect 7372 2454 7378 2488
rect 7412 2454 7418 2488
rect 7372 2442 7418 2454
rect 6710 2411 6764 2418
rect 6710 2359 6711 2411
rect 6763 2359 6764 2411
rect 6710 2352 6764 2359
rect 6710 2318 6720 2352
rect 6754 2318 6764 2352
rect 6710 2306 6764 2318
rect 6710 2271 6764 2278
rect 6710 2219 6711 2271
rect 6763 2219 6764 2271
rect 6710 2212 6764 2219
rect 6710 2178 6720 2212
rect 6754 2178 6764 2212
rect 6710 2166 6764 2178
rect 6710 2131 6764 2138
rect 6710 2079 6711 2131
rect 6763 2079 6764 2131
rect 6710 2072 6764 2079
rect 6710 2038 6720 2072
rect 6754 2038 6764 2072
rect 6710 2026 6764 2038
rect 6710 1991 6764 1998
rect 6710 1939 6711 1991
rect 6763 1939 6764 1991
rect 6710 1932 6764 1939
rect 6710 1898 6720 1932
rect 6754 1898 6764 1932
rect 6710 1886 6764 1898
rect 6710 1851 6764 1858
rect 6710 1799 6711 1851
rect 6763 1799 6764 1851
rect 6710 1792 6764 1799
rect 6710 1758 6720 1792
rect 6754 1758 6764 1792
rect 6710 1746 6764 1758
rect 6710 1711 6764 1718
rect 6710 1659 6711 1711
rect 6763 1659 6764 1711
rect 6710 1652 6764 1659
rect 6710 1618 6720 1652
rect 6754 1618 6764 1652
rect 6710 1606 6764 1618
rect 6710 1571 6764 1578
rect 6710 1519 6711 1571
rect 6763 1519 6764 1571
rect 6710 1512 6764 1519
rect 6710 1478 6720 1512
rect 6754 1478 6764 1512
rect 6710 1466 6764 1478
rect 6710 1431 6764 1438
rect 6710 1379 6711 1431
rect 6763 1379 6764 1431
rect 6710 1372 6764 1379
rect 6710 1338 6720 1372
rect 6754 1338 6764 1372
rect 6710 1326 6764 1338
rect 6880 1290 6910 2442
rect 6980 1290 7010 2442
rect 7080 1290 7110 2442
rect 7180 1290 7210 2442
rect 7280 1290 7310 2442
rect 7380 1290 7410 2442
rect 6650 1283 6766 1289
rect 6650 1249 6720 1283
rect 6754 1249 6766 1283
rect 6650 1243 6766 1249
rect 6872 1278 6918 1290
rect 6872 1244 6878 1278
rect 6912 1244 6918 1278
rect 6650 79 6680 1243
rect 6872 1232 6918 1244
rect 6972 1278 7018 1290
rect 6972 1244 6978 1278
rect 7012 1244 7018 1278
rect 6972 1232 7018 1244
rect 7072 1278 7118 1290
rect 7072 1244 7078 1278
rect 7112 1244 7118 1278
rect 7072 1232 7118 1244
rect 7172 1278 7218 1290
rect 7172 1244 7178 1278
rect 7212 1244 7218 1278
rect 7172 1232 7218 1244
rect 7272 1278 7318 1290
rect 7272 1244 7278 1278
rect 7312 1244 7318 1278
rect 7272 1232 7318 1244
rect 7372 1278 7418 1290
rect 7372 1244 7378 1278
rect 7412 1244 7418 1278
rect 7372 1232 7418 1244
rect 6710 1201 6764 1208
rect 6710 1149 6711 1201
rect 6763 1149 6764 1201
rect 6710 1142 6764 1149
rect 6710 1108 6720 1142
rect 6754 1108 6764 1142
rect 6710 1096 6764 1108
rect 6710 1061 6764 1068
rect 6710 1009 6711 1061
rect 6763 1009 6764 1061
rect 6710 1002 6764 1009
rect 6710 968 6720 1002
rect 6754 968 6764 1002
rect 6710 956 6764 968
rect 6710 921 6764 928
rect 6710 869 6711 921
rect 6763 869 6764 921
rect 6710 862 6764 869
rect 6710 828 6720 862
rect 6754 828 6764 862
rect 6710 816 6764 828
rect 6710 781 6764 788
rect 6710 729 6711 781
rect 6763 729 6764 781
rect 6710 722 6764 729
rect 6710 688 6720 722
rect 6754 688 6764 722
rect 6710 676 6764 688
rect 6710 641 6764 648
rect 6710 589 6711 641
rect 6763 589 6764 641
rect 6710 582 6764 589
rect 6710 548 6720 582
rect 6754 548 6764 582
rect 6710 536 6764 548
rect 6710 501 6764 508
rect 6710 449 6711 501
rect 6763 449 6764 501
rect 6710 442 6764 449
rect 6710 408 6720 442
rect 6754 408 6764 442
rect 6710 396 6764 408
rect 6710 361 6764 368
rect 6710 309 6711 361
rect 6763 309 6764 361
rect 6710 302 6764 309
rect 6710 268 6720 302
rect 6754 268 6764 302
rect 6710 256 6764 268
rect 6710 221 6764 228
rect 6710 169 6711 221
rect 6763 169 6764 221
rect 6710 162 6764 169
rect 6710 128 6720 162
rect 6754 128 6764 162
rect 6710 116 6764 128
rect 6880 80 6910 1232
rect 6980 80 7010 1232
rect 7080 80 7110 1232
rect 7180 80 7210 1232
rect 7280 80 7310 1232
rect 7380 80 7410 1232
rect 6650 73 6766 79
rect 6650 39 6720 73
rect 6754 39 6766 73
rect 6650 33 6766 39
rect 6872 68 6918 80
rect 6872 34 6878 68
rect 6912 34 6918 68
rect 6650 0 6680 33
rect 6872 22 6918 34
rect 6972 68 7018 80
rect 6972 34 6978 68
rect 7012 34 7018 68
rect 6972 22 7018 34
rect 7072 68 7118 80
rect 7072 34 7078 68
rect 7112 34 7118 68
rect 7072 22 7118 34
rect 7172 68 7218 80
rect 7172 34 7178 68
rect 7212 34 7218 68
rect 7172 22 7218 34
rect 7272 68 7318 80
rect 7272 34 7278 68
rect 7312 34 7318 68
rect 7272 22 7318 34
rect 7372 68 7418 80
rect 7372 34 7378 68
rect 7412 34 7418 68
rect 7372 22 7418 34
rect 6880 0 6910 22
rect 6980 0 7010 22
rect 7080 0 7110 22
rect 7180 0 7210 22
rect 7280 0 7310 22
rect 7380 0 7410 22
rect 8126 1 8297 7
rect 6308 -67 6309 -15
rect 6361 -67 6362 -15
rect 8126 -51 8153 1
rect 8205 -51 8217 1
rect 8269 -51 8297 1
rect 8126 -57 8297 -51
rect 8405 1 8736 7
rect 8405 -51 8416 1
rect 8468 -8 8480 1
rect 8532 -8 8544 1
rect 8596 -8 8608 1
rect 8660 -8 8672 1
rect 8476 -42 8480 -8
rect 8468 -51 8480 -42
rect 8532 -51 8544 -42
rect 8596 -51 8608 -42
rect 8660 -51 8672 -42
rect 8724 -51 8736 1
rect 8405 -57 8736 -51
rect 8806 1 9137 7
rect 8806 -51 8817 1
rect 8869 -8 8881 1
rect 8933 -8 8945 1
rect 8997 -8 9009 1
rect 9061 -8 9073 1
rect 9061 -42 9065 -8
rect 8869 -51 8881 -42
rect 8933 -51 8945 -42
rect 8997 -51 9009 -42
rect 9061 -51 9073 -42
rect 9125 -51 9137 1
rect 8806 -57 9137 -51
rect 9245 1 9416 7
rect 9245 -51 9272 1
rect 9324 -51 9336 1
rect 9388 -51 9416 1
rect 9245 -57 9416 -51
rect 6308 -79 6318 -67
rect 6352 -79 6362 -67
rect 6108 -132 6162 -131
rect 6108 -143 6118 -132
rect 6152 -143 6162 -132
rect 6108 -195 6109 -143
rect 6161 -195 6162 -143
rect 6108 -210 6162 -195
rect 6212 -133 6258 -81
rect 6212 -167 6218 -133
rect 6252 -167 6258 -133
rect 6118 -291 6125 -239
rect 6177 -291 6184 -239
rect 6012 -397 6018 -363
rect 6052 -397 6058 -363
rect 6012 -435 6058 -397
rect 6012 -469 6018 -435
rect 6052 -469 6058 -435
rect 6012 -512 6058 -469
rect 6109 -326 6161 -320
rect 6109 -390 6118 -378
rect 6152 -390 6161 -378
rect 6109 -454 6118 -442
rect 6152 -454 6161 -442
rect 6109 -512 6161 -506
rect 6212 -363 6258 -167
rect 6308 -131 6309 -79
rect 6361 -131 6362 -79
rect 8120 -108 8736 -102
rect 8120 -110 8160 -108
rect 6308 -132 6362 -131
rect 6308 -143 6318 -132
rect 6352 -143 6362 -132
rect 8000 -140 8160 -110
rect 6308 -195 6309 -143
rect 6361 -195 6362 -143
rect 8120 -142 8160 -140
rect 8194 -142 8232 -108
rect 8266 -142 8441 -108
rect 8475 -142 8513 -108
rect 8547 -142 8585 -108
rect 8619 -142 8657 -108
rect 8691 -142 8736 -108
rect 8120 -148 8736 -142
rect 8806 -151 8812 -99
rect 8864 -102 8870 -99
rect 8864 -108 9422 -102
rect 8885 -142 8923 -108
rect 8957 -142 8995 -108
rect 9029 -142 9067 -108
rect 9101 -142 9276 -108
rect 9310 -142 9348 -108
rect 9382 -142 9422 -108
rect 8864 -148 9422 -142
rect 8864 -151 8870 -148
rect 6308 -210 6362 -195
rect 8126 -199 8297 -193
rect 8034 -210 8040 -199
rect 8000 -240 8040 -210
rect 8034 -251 8040 -240
rect 8092 -251 8098 -199
rect 8126 -251 8153 -199
rect 8205 -251 8217 -199
rect 8269 -251 8297 -199
rect 8126 -257 8297 -251
rect 8325 -199 8377 -193
rect 8325 -257 8377 -251
rect 8405 -199 8736 -193
rect 8405 -251 8416 -199
rect 8468 -208 8480 -199
rect 8532 -208 8544 -199
rect 8596 -208 8608 -199
rect 8660 -208 8672 -199
rect 8476 -242 8480 -208
rect 8468 -251 8480 -242
rect 8532 -251 8544 -242
rect 8596 -251 8608 -242
rect 8660 -251 8672 -242
rect 8724 -251 8736 -199
rect 8405 -257 8736 -251
rect 8806 -199 9137 -193
rect 8806 -251 8817 -199
rect 8869 -208 8881 -199
rect 8933 -208 8945 -199
rect 8997 -208 9009 -199
rect 9061 -208 9073 -199
rect 9061 -242 9065 -208
rect 8869 -251 8881 -242
rect 8933 -251 8945 -242
rect 8997 -251 9009 -242
rect 9061 -251 9073 -242
rect 9125 -251 9137 -199
rect 8806 -257 9137 -251
rect 9165 -199 9217 -193
rect 9165 -257 9217 -251
rect 9245 -199 9416 -193
rect 9245 -251 9272 -199
rect 9324 -251 9336 -199
rect 9388 -251 9416 -199
rect 9245 -257 9416 -251
rect 8120 -308 8736 -302
rect 8120 -310 8160 -308
rect 6212 -397 6218 -363
rect 6252 -397 6258 -363
rect 6212 -435 6258 -397
rect 6212 -469 6218 -435
rect 6252 -469 6258 -435
rect 6212 -512 6258 -469
rect 6309 -326 6361 -320
rect 8000 -340 8160 -310
rect 8120 -342 8160 -340
rect 8194 -342 8232 -308
rect 8266 -342 8441 -308
rect 8475 -342 8513 -308
rect 8547 -342 8585 -308
rect 8619 -342 8657 -308
rect 8691 -342 8736 -308
rect 8120 -348 8736 -342
rect 8806 -351 8812 -299
rect 8864 -302 8870 -299
rect 8864 -308 9422 -302
rect 8885 -342 8923 -308
rect 8957 -342 8995 -308
rect 9029 -342 9067 -308
rect 9101 -342 9276 -308
rect 9310 -342 9348 -308
rect 9382 -342 9422 -308
rect 8864 -348 9422 -342
rect 8864 -351 8870 -348
rect 6309 -390 6318 -378
rect 6352 -390 6361 -378
rect 8126 -399 8297 -393
rect 8034 -410 8040 -399
rect 8000 -440 8040 -410
rect 6309 -454 6318 -442
rect 6352 -454 6361 -442
rect 8034 -451 8040 -440
rect 8092 -451 8098 -399
rect 8126 -451 8153 -399
rect 8205 -451 8217 -399
rect 8269 -451 8297 -399
rect 8126 -457 8297 -451
rect 8325 -399 8377 -393
rect 8325 -457 8377 -451
rect 8405 -399 8736 -393
rect 8405 -451 8416 -399
rect 8468 -408 8480 -399
rect 8532 -408 8544 -399
rect 8596 -408 8608 -399
rect 8660 -408 8672 -399
rect 8476 -442 8480 -408
rect 8468 -451 8480 -442
rect 8532 -451 8544 -442
rect 8596 -451 8608 -442
rect 8660 -451 8672 -442
rect 8724 -451 8736 -399
rect 8405 -457 8736 -451
rect 8806 -399 9137 -393
rect 8806 -451 8817 -399
rect 8869 -408 8881 -399
rect 8933 -408 8945 -399
rect 8997 -408 9009 -399
rect 9061 -408 9073 -399
rect 9061 -442 9065 -408
rect 8869 -451 8881 -442
rect 8933 -451 8945 -442
rect 8997 -451 9009 -442
rect 9061 -451 9073 -442
rect 9125 -451 9137 -399
rect 8806 -457 9137 -451
rect 9165 -399 9217 -393
rect 9165 -457 9217 -451
rect 9245 -399 9416 -393
rect 9245 -451 9272 -399
rect 9324 -451 9336 -399
rect 9388 -451 9416 -399
rect 9245 -457 9416 -451
rect 6309 -555 6361 -506
rect 8120 -508 8736 -502
rect 8120 -510 8160 -508
rect 8000 -540 8160 -510
rect 8120 -542 8160 -540
rect 8194 -542 8232 -508
rect 8266 -542 8441 -508
rect 8475 -542 8513 -508
rect 8547 -542 8585 -508
rect 8619 -542 8657 -508
rect 8691 -542 8736 -508
rect 8120 -548 8736 -542
rect 8806 -551 8812 -499
rect 8864 -502 8870 -499
rect 8864 -508 9422 -502
rect 8885 -542 8923 -508
rect 8957 -542 8995 -508
rect 9029 -542 9067 -508
rect 9101 -542 9276 -508
rect 9310 -542 9348 -508
rect 9382 -542 9422 -508
rect 8864 -548 9422 -542
rect 8864 -551 8870 -548
rect -137 -561 7 -555
rect -137 -595 -118 -561
rect -84 -595 -46 -561
rect -12 -595 7 -561
rect -137 -601 7 -595
rect 263 -561 407 -555
rect 263 -595 282 -561
rect 316 -595 354 -561
rect 388 -595 407 -561
rect 263 -601 407 -595
rect 663 -561 807 -555
rect 663 -595 682 -561
rect 716 -595 754 -561
rect 788 -595 807 -561
rect 663 -601 807 -595
rect 1063 -561 1207 -555
rect 1063 -595 1082 -561
rect 1116 -595 1154 -561
rect 1188 -595 1207 -561
rect 1063 -601 1207 -595
rect 1463 -561 1607 -555
rect 1463 -595 1482 -561
rect 1516 -595 1554 -561
rect 1588 -595 1607 -561
rect 1463 -601 1607 -595
rect 1863 -561 2007 -555
rect 1863 -595 1882 -561
rect 1916 -595 1954 -561
rect 1988 -595 2007 -561
rect 1863 -601 2007 -595
rect 2263 -561 2407 -555
rect 2263 -595 2282 -561
rect 2316 -595 2354 -561
rect 2388 -595 2407 -561
rect 2263 -601 2407 -595
rect 2663 -561 2807 -555
rect 2663 -595 2682 -561
rect 2716 -595 2754 -561
rect 2788 -595 2807 -561
rect 2663 -601 2807 -595
rect 3063 -561 3207 -555
rect 3063 -595 3082 -561
rect 3116 -595 3154 -561
rect 3188 -595 3207 -561
rect 3063 -601 3207 -595
rect 3463 -561 3607 -555
rect 3463 -595 3482 -561
rect 3516 -595 3554 -561
rect 3588 -595 3607 -561
rect 3463 -601 3607 -595
rect 3863 -561 4007 -555
rect 3863 -595 3882 -561
rect 3916 -595 3954 -561
rect 3988 -595 4007 -561
rect 3863 -601 4007 -595
rect 4263 -561 4407 -555
rect 4263 -595 4282 -561
rect 4316 -595 4354 -561
rect 4388 -595 4407 -561
rect 4263 -601 4407 -595
rect 4663 -561 4807 -555
rect 4663 -595 4682 -561
rect 4716 -595 4754 -561
rect 4788 -595 4807 -561
rect 4663 -601 4807 -595
rect 5063 -561 5207 -555
rect 5063 -595 5082 -561
rect 5116 -595 5154 -561
rect 5188 -595 5207 -561
rect 5063 -601 5207 -595
rect 5463 -561 5607 -555
rect 5463 -595 5482 -561
rect 5516 -595 5554 -561
rect 5588 -595 5607 -561
rect 5463 -601 5607 -595
rect 5863 -561 6007 -555
rect 5863 -595 5882 -561
rect 5916 -595 5954 -561
rect 5988 -595 6007 -561
rect 5863 -601 6007 -595
rect 6263 -561 6407 -555
rect 6263 -595 6282 -561
rect 6316 -595 6354 -561
rect 6388 -595 6407 -561
rect 6263 -601 6407 -595
rect 8126 -599 8297 -593
rect 8034 -610 8040 -599
rect 32 -630 90 -624
rect 32 -632 44 -630
rect -148 -662 44 -632
rect 32 -664 44 -662
rect 78 -632 90 -630
rect 180 -630 238 -624
rect 180 -632 192 -630
rect 78 -662 192 -632
rect 78 -664 90 -662
rect 32 -670 90 -664
rect 180 -664 192 -662
rect 226 -632 238 -630
rect 432 -630 490 -624
rect 432 -632 444 -630
rect 226 -662 444 -632
rect 226 -664 238 -662
rect 180 -670 238 -664
rect 432 -664 444 -662
rect 478 -632 490 -630
rect 580 -630 638 -624
rect 580 -632 592 -630
rect 478 -662 592 -632
rect 478 -664 490 -662
rect 432 -670 490 -664
rect 580 -664 592 -662
rect 626 -632 638 -630
rect 832 -630 890 -624
rect 832 -632 844 -630
rect 626 -662 844 -632
rect 626 -664 638 -662
rect 580 -670 638 -664
rect 832 -664 844 -662
rect 878 -632 890 -630
rect 980 -630 1038 -624
rect 980 -632 992 -630
rect 878 -662 992 -632
rect 878 -664 890 -662
rect 832 -670 890 -664
rect 980 -664 992 -662
rect 1026 -632 1038 -630
rect 1232 -630 1290 -624
rect 1232 -632 1244 -630
rect 1026 -662 1244 -632
rect 1026 -664 1038 -662
rect 980 -670 1038 -664
rect 1232 -664 1244 -662
rect 1278 -632 1290 -630
rect 1380 -630 1438 -624
rect 1380 -632 1392 -630
rect 1278 -662 1392 -632
rect 1278 -664 1290 -662
rect 1232 -670 1290 -664
rect 1380 -664 1392 -662
rect 1426 -632 1438 -630
rect 1632 -630 1690 -624
rect 1632 -632 1644 -630
rect 1426 -662 1644 -632
rect 1426 -664 1438 -662
rect 1380 -670 1438 -664
rect 1632 -664 1644 -662
rect 1678 -632 1690 -630
rect 1780 -630 1838 -624
rect 1780 -632 1792 -630
rect 1678 -662 1792 -632
rect 1678 -664 1690 -662
rect 1632 -670 1690 -664
rect 1780 -664 1792 -662
rect 1826 -632 1838 -630
rect 2032 -630 2090 -624
rect 2032 -632 2044 -630
rect 1826 -662 2044 -632
rect 1826 -664 1838 -662
rect 1780 -670 1838 -664
rect 2032 -664 2044 -662
rect 2078 -632 2090 -630
rect 2180 -630 2238 -624
rect 2180 -632 2192 -630
rect 2078 -662 2192 -632
rect 2078 -664 2090 -662
rect 2032 -670 2090 -664
rect 2180 -664 2192 -662
rect 2226 -632 2238 -630
rect 2432 -630 2490 -624
rect 2432 -632 2444 -630
rect 2226 -662 2444 -632
rect 2226 -664 2238 -662
rect 2180 -670 2238 -664
rect 2432 -664 2444 -662
rect 2478 -632 2490 -630
rect 2580 -630 2638 -624
rect 2580 -632 2592 -630
rect 2478 -662 2592 -632
rect 2478 -664 2490 -662
rect 2432 -670 2490 -664
rect 2580 -664 2592 -662
rect 2626 -632 2638 -630
rect 2832 -630 2890 -624
rect 2832 -632 2844 -630
rect 2626 -662 2844 -632
rect 2626 -664 2638 -662
rect 2580 -670 2638 -664
rect 2832 -664 2844 -662
rect 2878 -632 2890 -630
rect 2980 -630 3038 -624
rect 2980 -632 2992 -630
rect 2878 -662 2992 -632
rect 2878 -664 2890 -662
rect 2832 -670 2890 -664
rect 2980 -664 2992 -662
rect 3026 -632 3038 -630
rect 3232 -630 3290 -624
rect 3232 -632 3244 -630
rect 3026 -662 3244 -632
rect 3026 -664 3038 -662
rect 2980 -670 3038 -664
rect 3232 -664 3244 -662
rect 3278 -632 3290 -630
rect 3380 -630 3438 -624
rect 3380 -632 3392 -630
rect 3278 -662 3392 -632
rect 3278 -664 3290 -662
rect 3232 -670 3290 -664
rect 3380 -664 3392 -662
rect 3426 -632 3438 -630
rect 3632 -630 3690 -624
rect 3632 -632 3644 -630
rect 3426 -662 3644 -632
rect 3426 -664 3438 -662
rect 3380 -670 3438 -664
rect 3632 -664 3644 -662
rect 3678 -632 3690 -630
rect 3780 -630 3838 -624
rect 3780 -632 3792 -630
rect 3678 -662 3792 -632
rect 3678 -664 3690 -662
rect 3632 -670 3690 -664
rect 3780 -664 3792 -662
rect 3826 -632 3838 -630
rect 4032 -630 4090 -624
rect 4032 -632 4044 -630
rect 3826 -662 4044 -632
rect 3826 -664 3838 -662
rect 3780 -670 3838 -664
rect 4032 -664 4044 -662
rect 4078 -632 4090 -630
rect 4180 -630 4238 -624
rect 4180 -632 4192 -630
rect 4078 -662 4192 -632
rect 4078 -664 4090 -662
rect 4032 -670 4090 -664
rect 4180 -664 4192 -662
rect 4226 -632 4238 -630
rect 4432 -630 4490 -624
rect 4432 -632 4444 -630
rect 4226 -662 4444 -632
rect 4226 -664 4238 -662
rect 4180 -670 4238 -664
rect 4432 -664 4444 -662
rect 4478 -632 4490 -630
rect 4580 -630 4638 -624
rect 4580 -632 4592 -630
rect 4478 -662 4592 -632
rect 4478 -664 4490 -662
rect 4432 -670 4490 -664
rect 4580 -664 4592 -662
rect 4626 -632 4638 -630
rect 4832 -630 4890 -624
rect 4832 -632 4844 -630
rect 4626 -662 4844 -632
rect 4626 -664 4638 -662
rect 4580 -670 4638 -664
rect 4832 -664 4844 -662
rect 4878 -632 4890 -630
rect 4980 -630 5038 -624
rect 4980 -632 4992 -630
rect 4878 -662 4992 -632
rect 4878 -664 4890 -662
rect 4832 -670 4890 -664
rect 4980 -664 4992 -662
rect 5026 -632 5038 -630
rect 5232 -630 5290 -624
rect 5232 -632 5244 -630
rect 5026 -662 5244 -632
rect 5026 -664 5038 -662
rect 4980 -670 5038 -664
rect 5232 -664 5244 -662
rect 5278 -632 5290 -630
rect 5380 -630 5438 -624
rect 5380 -632 5392 -630
rect 5278 -662 5392 -632
rect 5278 -664 5290 -662
rect 5232 -670 5290 -664
rect 5380 -664 5392 -662
rect 5426 -632 5438 -630
rect 5632 -630 5690 -624
rect 5632 -632 5644 -630
rect 5426 -662 5644 -632
rect 5426 -664 5438 -662
rect 5380 -670 5438 -664
rect 5632 -664 5644 -662
rect 5678 -632 5690 -630
rect 5780 -630 5838 -624
rect 5780 -632 5792 -630
rect 5678 -662 5792 -632
rect 5678 -664 5690 -662
rect 5632 -670 5690 -664
rect 5780 -664 5792 -662
rect 5826 -632 5838 -630
rect 6032 -630 6090 -624
rect 6032 -632 6044 -630
rect 5826 -662 6044 -632
rect 5826 -664 5838 -662
rect 5780 -670 5838 -664
rect 6032 -664 6044 -662
rect 6078 -632 6090 -630
rect 6180 -630 6238 -624
rect 6180 -632 6192 -630
rect 6078 -662 6192 -632
rect 6078 -664 6090 -662
rect 6032 -670 6090 -664
rect 6180 -664 6192 -662
rect 6226 -632 6238 -630
rect 6226 -662 6418 -632
rect 8000 -640 8040 -610
rect 8034 -651 8040 -640
rect 8092 -651 8098 -599
rect 8126 -651 8153 -599
rect 8205 -651 8217 -599
rect 8269 -651 8297 -599
rect 8126 -657 8297 -651
rect 8325 -599 8377 -593
rect 8325 -657 8377 -651
rect 8405 -599 8736 -593
rect 8405 -651 8416 -599
rect 8468 -608 8480 -599
rect 8532 -608 8544 -599
rect 8596 -608 8608 -599
rect 8660 -608 8672 -599
rect 8476 -642 8480 -608
rect 8468 -651 8480 -642
rect 8532 -651 8544 -642
rect 8596 -651 8608 -642
rect 8660 -651 8672 -642
rect 8724 -651 8736 -599
rect 8405 -657 8736 -651
rect 8806 -599 9137 -593
rect 8806 -651 8817 -599
rect 8869 -608 8881 -599
rect 8933 -608 8945 -599
rect 8997 -608 9009 -599
rect 9061 -608 9073 -599
rect 9061 -642 9065 -608
rect 8869 -651 8881 -642
rect 8933 -651 8945 -642
rect 8997 -651 9009 -642
rect 9061 -651 9073 -642
rect 9125 -651 9137 -599
rect 8806 -657 9137 -651
rect 9165 -599 9217 -593
rect 9165 -657 9217 -651
rect 9245 -599 9416 -593
rect 9245 -651 9272 -599
rect 9324 -651 9336 -599
rect 9388 -651 9416 -599
rect 9245 -657 9416 -651
rect 6226 -664 6238 -662
rect 6180 -670 6238 -664
rect 8120 -708 8736 -702
rect 8120 -710 8160 -708
rect 8000 -740 8160 -710
rect 8120 -742 8160 -740
rect 8194 -742 8232 -708
rect 8266 -742 8441 -708
rect 8475 -742 8513 -708
rect 8547 -742 8585 -708
rect 8619 -742 8657 -708
rect 8691 -742 8736 -708
rect 8120 -748 8736 -742
rect 8806 -751 8812 -699
rect 8864 -702 8870 -699
rect 8864 -708 9422 -702
rect 8885 -742 8923 -708
rect 8957 -742 8995 -708
rect 9029 -742 9067 -708
rect 9101 -742 9276 -708
rect 9310 -742 9348 -708
rect 9382 -742 9422 -708
rect 8864 -748 9422 -742
rect 8864 -751 8870 -748
rect 8126 -799 8297 -793
rect 8034 -810 8040 -799
rect -18 -880 -9 -828
rect 43 -880 55 -828
rect 107 -880 116 -828
rect 154 -880 163 -828
rect 215 -880 227 -828
rect 279 -880 288 -828
rect 382 -880 391 -828
rect 443 -880 455 -828
rect 507 -880 516 -828
rect 554 -880 563 -828
rect 615 -880 627 -828
rect 679 -880 688 -828
rect 782 -880 791 -828
rect 843 -880 855 -828
rect 907 -880 916 -828
rect 954 -880 963 -828
rect 1015 -880 1027 -828
rect 1079 -880 1088 -828
rect 1182 -880 1191 -828
rect 1243 -880 1255 -828
rect 1307 -880 1316 -828
rect 1354 -880 1363 -828
rect 1415 -880 1427 -828
rect 1479 -880 1488 -828
rect 1582 -880 1591 -828
rect 1643 -880 1655 -828
rect 1707 -880 1716 -828
rect 1754 -880 1763 -828
rect 1815 -880 1827 -828
rect 1879 -880 1888 -828
rect 1982 -880 1991 -828
rect 2043 -880 2055 -828
rect 2107 -880 2116 -828
rect 2154 -880 2163 -828
rect 2215 -880 2227 -828
rect 2279 -880 2288 -828
rect 2382 -880 2391 -828
rect 2443 -880 2455 -828
rect 2507 -880 2516 -828
rect 2554 -880 2563 -828
rect 2615 -880 2627 -828
rect 2679 -880 2688 -828
rect 2782 -880 2791 -828
rect 2843 -880 2855 -828
rect 2907 -880 2916 -828
rect 2954 -880 2963 -828
rect 3015 -880 3027 -828
rect 3079 -880 3088 -828
rect 3182 -880 3191 -828
rect 3243 -880 3255 -828
rect 3307 -880 3316 -828
rect 3354 -880 3363 -828
rect 3415 -880 3427 -828
rect 3479 -880 3488 -828
rect 3582 -880 3591 -828
rect 3643 -880 3655 -828
rect 3707 -880 3716 -828
rect 3754 -880 3763 -828
rect 3815 -880 3827 -828
rect 3879 -880 3888 -828
rect 3982 -880 3991 -828
rect 4043 -880 4055 -828
rect 4107 -880 4116 -828
rect 4154 -880 4163 -828
rect 4215 -880 4227 -828
rect 4279 -880 4288 -828
rect 4382 -880 4391 -828
rect 4443 -880 4455 -828
rect 4507 -880 4516 -828
rect 4554 -880 4563 -828
rect 4615 -880 4627 -828
rect 4679 -880 4688 -828
rect 4782 -880 4791 -828
rect 4843 -880 4855 -828
rect 4907 -880 4916 -828
rect 4954 -880 4963 -828
rect 5015 -880 5027 -828
rect 5079 -880 5088 -828
rect 5182 -880 5191 -828
rect 5243 -880 5255 -828
rect 5307 -880 5316 -828
rect 5354 -880 5363 -828
rect 5415 -880 5427 -828
rect 5479 -880 5488 -828
rect 5582 -880 5591 -828
rect 5643 -880 5655 -828
rect 5707 -880 5716 -828
rect 5754 -880 5763 -828
rect 5815 -880 5827 -828
rect 5879 -880 5888 -828
rect 5982 -880 5991 -828
rect 6043 -880 6055 -828
rect 6107 -880 6116 -828
rect 6154 -880 6163 -828
rect 6215 -880 6227 -828
rect 6279 -880 6288 -828
rect 8000 -840 8040 -810
rect 8034 -851 8040 -840
rect 8092 -851 8098 -799
rect 8126 -851 8153 -799
rect 8205 -851 8217 -799
rect 8269 -851 8297 -799
rect 8126 -857 8297 -851
rect 8325 -799 8377 -793
rect 8325 -857 8377 -851
rect 8405 -799 8736 -793
rect 8405 -851 8416 -799
rect 8468 -808 8480 -799
rect 8532 -808 8544 -799
rect 8596 -808 8608 -799
rect 8660 -808 8672 -799
rect 8476 -842 8480 -808
rect 8468 -851 8480 -842
rect 8532 -851 8544 -842
rect 8596 -851 8608 -842
rect 8660 -851 8672 -842
rect 8724 -851 8736 -799
rect 8405 -857 8736 -851
rect 8806 -799 9137 -793
rect 8806 -851 8817 -799
rect 8869 -808 8881 -799
rect 8933 -808 8945 -799
rect 8997 -808 9009 -799
rect 9061 -808 9073 -799
rect 9061 -842 9065 -808
rect 8869 -851 8881 -842
rect 8933 -851 8945 -842
rect 8997 -851 9009 -842
rect 9061 -851 9073 -842
rect 9125 -851 9137 -799
rect 8806 -857 9137 -851
rect 9165 -799 9217 -793
rect 9165 -857 9217 -851
rect 9245 -799 9416 -793
rect 9245 -851 9272 -799
rect 9324 -851 9336 -799
rect 9388 -851 9416 -799
rect 9245 -857 9416 -851
rect -94 -908 -36 -902
rect -94 -910 -82 -908
rect -106 -940 -82 -910
rect -94 -942 -82 -940
rect -48 -910 -36 -908
rect 706 -908 764 -902
rect 706 -910 718 -908
rect -48 -940 718 -910
rect -48 -942 -36 -940
rect -94 -948 -36 -942
rect 706 -942 718 -940
rect 752 -910 764 -908
rect 1506 -908 1564 -902
rect 1506 -910 1518 -908
rect 752 -940 1518 -910
rect 752 -942 764 -940
rect 706 -948 764 -942
rect 1506 -942 1518 -940
rect 1552 -910 1564 -908
rect 2306 -908 2364 -902
rect 2306 -910 2318 -908
rect 1552 -940 2318 -910
rect 1552 -942 1564 -940
rect 1506 -948 1564 -942
rect 2306 -942 2318 -940
rect 2352 -910 2364 -908
rect 3106 -908 3164 -902
rect 3106 -910 3118 -908
rect 2352 -940 3118 -910
rect 2352 -942 2364 -940
rect 2306 -948 2364 -942
rect 3106 -942 3118 -940
rect 3152 -910 3164 -908
rect 3906 -908 3964 -902
rect 3906 -910 3918 -908
rect 3152 -940 3918 -910
rect 3152 -942 3164 -940
rect 3106 -948 3164 -942
rect 3906 -942 3918 -940
rect 3952 -910 3964 -908
rect 4706 -908 4764 -902
rect 4706 -910 4718 -908
rect 3952 -940 4718 -910
rect 3952 -942 3964 -940
rect 3906 -948 3964 -942
rect 4706 -942 4718 -940
rect 4752 -910 4764 -908
rect 5506 -908 5564 -902
rect 5506 -910 5518 -908
rect 4752 -940 5518 -910
rect 4752 -942 4764 -940
rect 4706 -948 4764 -942
rect 5506 -942 5518 -940
rect 5552 -910 5564 -908
rect 6306 -908 6364 -902
rect 6306 -910 6318 -908
rect 5552 -940 6318 -910
rect 5552 -942 5564 -940
rect 5506 -948 5564 -942
rect 6306 -942 6318 -940
rect 6352 -910 6364 -908
rect 8120 -908 8736 -902
rect 8120 -910 8160 -908
rect 6352 -940 6376 -910
rect 8000 -940 8160 -910
rect 6352 -942 6364 -940
rect 6306 -948 6364 -942
rect 8120 -942 8160 -940
rect 8194 -942 8232 -908
rect 8266 -942 8441 -908
rect 8475 -942 8513 -908
rect 8547 -942 8585 -908
rect 8619 -942 8657 -908
rect 8691 -942 8736 -908
rect 8120 -948 8736 -942
rect 8806 -951 8812 -899
rect 8864 -902 8870 -899
rect 8864 -908 9422 -902
rect 8885 -942 8923 -908
rect 8957 -942 8995 -908
rect 9029 -942 9067 -908
rect 9101 -942 9276 -908
rect 9310 -942 9348 -908
rect 9382 -942 9422 -908
rect 8864 -948 9422 -942
rect 8864 -951 8870 -948
rect 8126 -999 8297 -993
rect -94 -1008 -36 -1002
rect -94 -1010 -82 -1008
rect -106 -1040 -82 -1010
rect -94 -1042 -82 -1040
rect -48 -1010 -36 -1008
rect 706 -1008 764 -1002
rect 706 -1010 718 -1008
rect -48 -1040 718 -1010
rect -48 -1042 -36 -1040
rect -94 -1048 -36 -1042
rect 706 -1042 718 -1040
rect 752 -1010 764 -1008
rect 1506 -1008 1564 -1002
rect 1506 -1010 1518 -1008
rect 752 -1040 1518 -1010
rect 752 -1042 764 -1040
rect 706 -1048 764 -1042
rect 1506 -1042 1518 -1040
rect 1552 -1010 1564 -1008
rect 2306 -1008 2364 -1002
rect 2306 -1010 2318 -1008
rect 1552 -1040 2318 -1010
rect 1552 -1042 1564 -1040
rect 1506 -1048 1564 -1042
rect 2306 -1042 2318 -1040
rect 2352 -1010 2364 -1008
rect 3106 -1008 3164 -1002
rect 3106 -1010 3118 -1008
rect 2352 -1040 3118 -1010
rect 2352 -1042 2364 -1040
rect 2306 -1048 2364 -1042
rect 3106 -1042 3118 -1040
rect 3152 -1010 3164 -1008
rect 3906 -1008 3964 -1002
rect 3906 -1010 3918 -1008
rect 3152 -1040 3918 -1010
rect 3152 -1042 3164 -1040
rect 3106 -1048 3164 -1042
rect 3906 -1042 3918 -1040
rect 3952 -1010 3964 -1008
rect 4706 -1008 4764 -1002
rect 4706 -1010 4718 -1008
rect 3952 -1040 4718 -1010
rect 3952 -1042 3964 -1040
rect 3906 -1048 3964 -1042
rect 4706 -1042 4718 -1040
rect 4752 -1010 4764 -1008
rect 5506 -1008 5564 -1002
rect 5506 -1010 5518 -1008
rect 4752 -1040 5518 -1010
rect 4752 -1042 4764 -1040
rect 4706 -1048 4764 -1042
rect 5506 -1042 5518 -1040
rect 5552 -1010 5564 -1008
rect 6306 -1008 6364 -1002
rect 6306 -1010 6318 -1008
rect 5552 -1040 6318 -1010
rect 5552 -1042 5564 -1040
rect 5506 -1048 5564 -1042
rect 6306 -1042 6318 -1040
rect 6352 -1010 6364 -1008
rect 8034 -1010 8040 -999
rect 6352 -1040 6376 -1010
rect 8000 -1040 8040 -1010
rect 6352 -1042 6364 -1040
rect 6306 -1048 6364 -1042
rect 8034 -1051 8040 -1040
rect 8092 -1051 8098 -999
rect 8126 -1051 8153 -999
rect 8205 -1051 8217 -999
rect 8269 -1051 8297 -999
rect 8126 -1057 8297 -1051
rect 8325 -999 8377 -993
rect 8325 -1057 8377 -1051
rect 8405 -999 8736 -993
rect 8405 -1051 8416 -999
rect 8468 -1008 8480 -999
rect 8532 -1008 8544 -999
rect 8596 -1008 8608 -999
rect 8660 -1008 8672 -999
rect 8476 -1042 8480 -1008
rect 8468 -1051 8480 -1042
rect 8532 -1051 8544 -1042
rect 8596 -1051 8608 -1042
rect 8660 -1051 8672 -1042
rect 8724 -1051 8736 -999
rect 8405 -1057 8736 -1051
rect 8806 -999 9137 -993
rect 8806 -1051 8817 -999
rect 8869 -1008 8881 -999
rect 8933 -1008 8945 -999
rect 8997 -1008 9009 -999
rect 9061 -1008 9073 -999
rect 9061 -1042 9065 -1008
rect 8869 -1051 8881 -1042
rect 8933 -1051 8945 -1042
rect 8997 -1051 9009 -1042
rect 9061 -1051 9073 -1042
rect 9125 -1051 9137 -999
rect 8806 -1057 9137 -1051
rect 9165 -999 9217 -993
rect 9165 -1057 9217 -1051
rect 9245 -999 9416 -993
rect 9245 -1051 9272 -999
rect 9324 -1051 9336 -999
rect 9388 -1051 9416 -999
rect 9245 -1057 9416 -1051
rect -94 -1108 -36 -1102
rect -94 -1110 -82 -1108
rect -106 -1140 -82 -1110
rect -94 -1142 -82 -1140
rect -48 -1110 -36 -1108
rect 706 -1108 764 -1102
rect 706 -1110 718 -1108
rect -48 -1140 718 -1110
rect -48 -1142 -36 -1140
rect -94 -1148 -36 -1142
rect 706 -1142 718 -1140
rect 752 -1110 764 -1108
rect 1506 -1108 1564 -1102
rect 1506 -1110 1518 -1108
rect 752 -1140 1518 -1110
rect 752 -1142 764 -1140
rect 706 -1148 764 -1142
rect 1506 -1142 1518 -1140
rect 1552 -1110 1564 -1108
rect 2306 -1108 2364 -1102
rect 2306 -1110 2318 -1108
rect 1552 -1140 2318 -1110
rect 1552 -1142 1564 -1140
rect 1506 -1148 1564 -1142
rect 2306 -1142 2318 -1140
rect 2352 -1110 2364 -1108
rect 3106 -1108 3164 -1102
rect 3106 -1110 3118 -1108
rect 2352 -1140 3118 -1110
rect 2352 -1142 2364 -1140
rect 2306 -1148 2364 -1142
rect 3106 -1142 3118 -1140
rect 3152 -1110 3164 -1108
rect 3906 -1108 3964 -1102
rect 3906 -1110 3918 -1108
rect 3152 -1140 3918 -1110
rect 3152 -1142 3164 -1140
rect 3106 -1148 3164 -1142
rect 3906 -1142 3918 -1140
rect 3952 -1110 3964 -1108
rect 4706 -1108 4764 -1102
rect 4706 -1110 4718 -1108
rect 3952 -1140 4718 -1110
rect 3952 -1142 3964 -1140
rect 3906 -1148 3964 -1142
rect 4706 -1142 4718 -1140
rect 4752 -1110 4764 -1108
rect 5506 -1108 5564 -1102
rect 5506 -1110 5518 -1108
rect 4752 -1140 5518 -1110
rect 4752 -1142 4764 -1140
rect 4706 -1148 4764 -1142
rect 5506 -1142 5518 -1140
rect 5552 -1110 5564 -1108
rect 6306 -1108 6364 -1102
rect 6306 -1110 6318 -1108
rect 5552 -1140 6318 -1110
rect 5552 -1142 5564 -1140
rect 5506 -1148 5564 -1142
rect 6306 -1142 6318 -1140
rect 6352 -1110 6364 -1108
rect 8120 -1108 8736 -1102
rect 8120 -1110 8160 -1108
rect 6352 -1140 6376 -1110
rect 8000 -1140 8160 -1110
rect 6352 -1142 6364 -1140
rect 6306 -1148 6364 -1142
rect 8120 -1142 8160 -1140
rect 8194 -1142 8232 -1108
rect 8266 -1142 8441 -1108
rect 8475 -1142 8513 -1108
rect 8547 -1142 8585 -1108
rect 8619 -1142 8657 -1108
rect 8691 -1142 8736 -1108
rect 8120 -1148 8736 -1142
rect 8806 -1151 8812 -1099
rect 8864 -1102 8870 -1099
rect 8864 -1108 9422 -1102
rect 8885 -1142 8923 -1108
rect 8957 -1142 8995 -1108
rect 9029 -1142 9067 -1108
rect 9101 -1142 9276 -1108
rect 9310 -1142 9348 -1108
rect 9382 -1142 9422 -1108
rect 8864 -1148 9422 -1142
rect 8864 -1151 8870 -1148
rect 8126 -1199 8297 -1193
rect -94 -1208 -36 -1202
rect -94 -1210 -82 -1208
rect -106 -1240 -82 -1210
rect -94 -1242 -82 -1240
rect -48 -1210 -36 -1208
rect 706 -1208 764 -1202
rect 706 -1210 718 -1208
rect -48 -1240 718 -1210
rect -48 -1242 -36 -1240
rect -94 -1248 -36 -1242
rect 706 -1242 718 -1240
rect 752 -1210 764 -1208
rect 1506 -1208 1564 -1202
rect 1506 -1210 1518 -1208
rect 752 -1240 1518 -1210
rect 752 -1242 764 -1240
rect 706 -1248 764 -1242
rect 1506 -1242 1518 -1240
rect 1552 -1210 1564 -1208
rect 2306 -1208 2364 -1202
rect 2306 -1210 2318 -1208
rect 1552 -1240 2318 -1210
rect 1552 -1242 1564 -1240
rect 1506 -1248 1564 -1242
rect 2306 -1242 2318 -1240
rect 2352 -1210 2364 -1208
rect 3106 -1208 3164 -1202
rect 3106 -1210 3118 -1208
rect 2352 -1240 3118 -1210
rect 2352 -1242 2364 -1240
rect 2306 -1248 2364 -1242
rect 3106 -1242 3118 -1240
rect 3152 -1210 3164 -1208
rect 3906 -1208 3964 -1202
rect 3906 -1210 3918 -1208
rect 3152 -1240 3918 -1210
rect 3152 -1242 3164 -1240
rect 3106 -1248 3164 -1242
rect 3906 -1242 3918 -1240
rect 3952 -1210 3964 -1208
rect 4706 -1208 4764 -1202
rect 4706 -1210 4718 -1208
rect 3952 -1240 4718 -1210
rect 3952 -1242 3964 -1240
rect 3906 -1248 3964 -1242
rect 4706 -1242 4718 -1240
rect 4752 -1210 4764 -1208
rect 5506 -1208 5564 -1202
rect 5506 -1210 5518 -1208
rect 4752 -1240 5518 -1210
rect 4752 -1242 4764 -1240
rect 4706 -1248 4764 -1242
rect 5506 -1242 5518 -1240
rect 5552 -1210 5564 -1208
rect 6306 -1208 6364 -1202
rect 6306 -1210 6318 -1208
rect 5552 -1240 6318 -1210
rect 5552 -1242 5564 -1240
rect 5506 -1248 5564 -1242
rect 6306 -1242 6318 -1240
rect 6352 -1210 6364 -1208
rect 8034 -1210 8040 -1199
rect 6352 -1240 6376 -1210
rect 8000 -1240 8040 -1210
rect 6352 -1242 6364 -1240
rect 6306 -1248 6364 -1242
rect 8034 -1251 8040 -1240
rect 8092 -1251 8098 -1199
rect 8126 -1251 8153 -1199
rect 8205 -1251 8217 -1199
rect 8269 -1251 8297 -1199
rect 8126 -1257 8297 -1251
rect 8325 -1199 8377 -1193
rect 8325 -1257 8377 -1251
rect 8405 -1199 8736 -1193
rect 8405 -1251 8416 -1199
rect 8468 -1208 8480 -1199
rect 8532 -1208 8544 -1199
rect 8596 -1208 8608 -1199
rect 8660 -1208 8672 -1199
rect 8476 -1242 8480 -1208
rect 8468 -1251 8480 -1242
rect 8532 -1251 8544 -1242
rect 8596 -1251 8608 -1242
rect 8660 -1251 8672 -1242
rect 8724 -1251 8736 -1199
rect 8405 -1257 8736 -1251
rect 8806 -1199 9137 -1193
rect 8806 -1251 8817 -1199
rect 8869 -1208 8881 -1199
rect 8933 -1208 8945 -1199
rect 8997 -1208 9009 -1199
rect 9061 -1208 9073 -1199
rect 9061 -1242 9065 -1208
rect 8869 -1251 8881 -1242
rect 8933 -1251 8945 -1242
rect 8997 -1251 9009 -1242
rect 9061 -1251 9073 -1242
rect 9125 -1251 9137 -1199
rect 8806 -1257 9137 -1251
rect 9165 -1199 9217 -1193
rect 9165 -1257 9217 -1251
rect 9245 -1199 9416 -1193
rect 9245 -1251 9272 -1199
rect 9324 -1251 9336 -1199
rect 9388 -1251 9416 -1199
rect 9245 -1257 9416 -1251
rect -94 -1308 -36 -1302
rect -94 -1310 -82 -1308
rect -106 -1340 -82 -1310
rect -94 -1342 -82 -1340
rect -48 -1310 -36 -1308
rect 706 -1308 764 -1302
rect 706 -1310 718 -1308
rect -48 -1340 718 -1310
rect -48 -1342 -36 -1340
rect -94 -1348 -36 -1342
rect 706 -1342 718 -1340
rect 752 -1310 764 -1308
rect 1506 -1308 1564 -1302
rect 1506 -1310 1518 -1308
rect 752 -1340 1518 -1310
rect 752 -1342 764 -1340
rect 706 -1348 764 -1342
rect 1506 -1342 1518 -1340
rect 1552 -1310 1564 -1308
rect 2306 -1308 2364 -1302
rect 2306 -1310 2318 -1308
rect 1552 -1340 2318 -1310
rect 1552 -1342 1564 -1340
rect 1506 -1348 1564 -1342
rect 2306 -1342 2318 -1340
rect 2352 -1310 2364 -1308
rect 3106 -1308 3164 -1302
rect 3106 -1310 3118 -1308
rect 2352 -1340 3118 -1310
rect 2352 -1342 2364 -1340
rect 2306 -1348 2364 -1342
rect 3106 -1342 3118 -1340
rect 3152 -1310 3164 -1308
rect 3906 -1308 3964 -1302
rect 3906 -1310 3918 -1308
rect 3152 -1340 3918 -1310
rect 3152 -1342 3164 -1340
rect 3106 -1348 3164 -1342
rect 3906 -1342 3918 -1340
rect 3952 -1310 3964 -1308
rect 4706 -1308 4764 -1302
rect 4706 -1310 4718 -1308
rect 3952 -1340 4718 -1310
rect 3952 -1342 3964 -1340
rect 3906 -1348 3964 -1342
rect 4706 -1342 4718 -1340
rect 4752 -1310 4764 -1308
rect 5506 -1308 5564 -1302
rect 5506 -1310 5518 -1308
rect 4752 -1340 5518 -1310
rect 4752 -1342 4764 -1340
rect 4706 -1348 4764 -1342
rect 5506 -1342 5518 -1340
rect 5552 -1310 5564 -1308
rect 6306 -1308 6364 -1302
rect 6306 -1310 6318 -1308
rect 5552 -1340 6318 -1310
rect 5552 -1342 5564 -1340
rect 5506 -1348 5564 -1342
rect 6306 -1342 6318 -1340
rect 6352 -1310 6364 -1308
rect 8120 -1308 8736 -1302
rect 8120 -1310 8160 -1308
rect 6352 -1340 6376 -1310
rect 8000 -1340 8160 -1310
rect 6352 -1342 6364 -1340
rect 6306 -1348 6364 -1342
rect 8120 -1342 8160 -1340
rect 8194 -1342 8232 -1308
rect 8266 -1342 8441 -1308
rect 8475 -1342 8513 -1308
rect 8547 -1342 8585 -1308
rect 8619 -1342 8657 -1308
rect 8691 -1342 8736 -1308
rect 8120 -1348 8736 -1342
rect 8806 -1351 8812 -1299
rect 8864 -1302 8870 -1299
rect 8864 -1308 9422 -1302
rect 8885 -1342 8923 -1308
rect 8957 -1342 8995 -1308
rect 9029 -1342 9067 -1308
rect 9101 -1342 9276 -1308
rect 9310 -1342 9348 -1308
rect 9382 -1342 9422 -1308
rect 8864 -1348 9422 -1342
rect 8864 -1351 8870 -1348
rect 8126 -1399 8297 -1393
rect -94 -1408 -36 -1402
rect -94 -1410 -82 -1408
rect -106 -1440 -82 -1410
rect -94 -1442 -82 -1440
rect -48 -1410 -36 -1408
rect 706 -1408 764 -1402
rect 706 -1410 718 -1408
rect -48 -1440 718 -1410
rect -48 -1442 -36 -1440
rect -94 -1448 -36 -1442
rect 706 -1442 718 -1440
rect 752 -1410 764 -1408
rect 1506 -1408 1564 -1402
rect 1506 -1410 1518 -1408
rect 752 -1440 1518 -1410
rect 752 -1442 764 -1440
rect 706 -1448 764 -1442
rect 1506 -1442 1518 -1440
rect 1552 -1410 1564 -1408
rect 2306 -1408 2364 -1402
rect 2306 -1410 2318 -1408
rect 1552 -1440 2318 -1410
rect 1552 -1442 1564 -1440
rect 1506 -1448 1564 -1442
rect 2306 -1442 2318 -1440
rect 2352 -1410 2364 -1408
rect 3106 -1408 3164 -1402
rect 3106 -1410 3118 -1408
rect 2352 -1440 3118 -1410
rect 2352 -1442 2364 -1440
rect 2306 -1448 2364 -1442
rect 3106 -1442 3118 -1440
rect 3152 -1410 3164 -1408
rect 3906 -1408 3964 -1402
rect 3906 -1410 3918 -1408
rect 3152 -1440 3918 -1410
rect 3152 -1442 3164 -1440
rect 3106 -1448 3164 -1442
rect 3906 -1442 3918 -1440
rect 3952 -1410 3964 -1408
rect 4706 -1408 4764 -1402
rect 4706 -1410 4718 -1408
rect 3952 -1440 4718 -1410
rect 3952 -1442 3964 -1440
rect 3906 -1448 3964 -1442
rect 4706 -1442 4718 -1440
rect 4752 -1410 4764 -1408
rect 5506 -1408 5564 -1402
rect 5506 -1410 5518 -1408
rect 4752 -1440 5518 -1410
rect 4752 -1442 4764 -1440
rect 4706 -1448 4764 -1442
rect 5506 -1442 5518 -1440
rect 5552 -1410 5564 -1408
rect 6306 -1408 6364 -1402
rect 6306 -1410 6318 -1408
rect 5552 -1440 6318 -1410
rect 5552 -1442 5564 -1440
rect 5506 -1448 5564 -1442
rect 6306 -1442 6318 -1440
rect 6352 -1410 6364 -1408
rect 8034 -1410 8040 -1399
rect 6352 -1440 6376 -1410
rect 8000 -1440 8040 -1410
rect 6352 -1442 6364 -1440
rect 6306 -1448 6364 -1442
rect 8034 -1451 8040 -1440
rect 8092 -1451 8098 -1399
rect 8126 -1451 8153 -1399
rect 8205 -1451 8217 -1399
rect 8269 -1451 8297 -1399
rect 8126 -1457 8297 -1451
rect 8325 -1399 8377 -1393
rect 8325 -1457 8377 -1451
rect 8405 -1399 8736 -1393
rect 8405 -1451 8416 -1399
rect 8468 -1408 8480 -1399
rect 8532 -1408 8544 -1399
rect 8596 -1408 8608 -1399
rect 8660 -1408 8672 -1399
rect 8476 -1442 8480 -1408
rect 8468 -1451 8480 -1442
rect 8532 -1451 8544 -1442
rect 8596 -1451 8608 -1442
rect 8660 -1451 8672 -1442
rect 8724 -1451 8736 -1399
rect 8405 -1457 8736 -1451
rect 8806 -1399 9137 -1393
rect 8806 -1451 8817 -1399
rect 8869 -1408 8881 -1399
rect 8933 -1408 8945 -1399
rect 8997 -1408 9009 -1399
rect 9061 -1408 9073 -1399
rect 9061 -1442 9065 -1408
rect 8869 -1451 8881 -1442
rect 8933 -1451 8945 -1442
rect 8997 -1451 9009 -1442
rect 9061 -1451 9073 -1442
rect 9125 -1451 9137 -1399
rect 8806 -1457 9137 -1451
rect 9165 -1399 9217 -1393
rect 9165 -1457 9217 -1451
rect 9245 -1399 9416 -1393
rect 9245 -1451 9272 -1399
rect 9324 -1451 9336 -1399
rect 9388 -1451 9416 -1399
rect 9245 -1457 9416 -1451
rect -94 -1508 -36 -1502
rect -94 -1510 -82 -1508
rect -106 -1540 -82 -1510
rect -94 -1542 -82 -1540
rect -48 -1510 -36 -1508
rect 706 -1508 764 -1502
rect 706 -1510 718 -1508
rect -48 -1540 718 -1510
rect -48 -1542 -36 -1540
rect -94 -1548 -36 -1542
rect 706 -1542 718 -1540
rect 752 -1510 764 -1508
rect 1506 -1508 1564 -1502
rect 1506 -1510 1518 -1508
rect 752 -1540 1518 -1510
rect 752 -1542 764 -1540
rect 706 -1548 764 -1542
rect 1506 -1542 1518 -1540
rect 1552 -1510 1564 -1508
rect 2306 -1508 2364 -1502
rect 2306 -1510 2318 -1508
rect 1552 -1540 2318 -1510
rect 1552 -1542 1564 -1540
rect 1506 -1548 1564 -1542
rect 2306 -1542 2318 -1540
rect 2352 -1510 2364 -1508
rect 3106 -1508 3164 -1502
rect 3106 -1510 3118 -1508
rect 2352 -1540 3118 -1510
rect 2352 -1542 2364 -1540
rect 2306 -1548 2364 -1542
rect 3106 -1542 3118 -1540
rect 3152 -1510 3164 -1508
rect 3906 -1508 3964 -1502
rect 3906 -1510 3918 -1508
rect 3152 -1540 3918 -1510
rect 3152 -1542 3164 -1540
rect 3106 -1548 3164 -1542
rect 3906 -1542 3918 -1540
rect 3952 -1510 3964 -1508
rect 4706 -1508 4764 -1502
rect 4706 -1510 4718 -1508
rect 3952 -1540 4718 -1510
rect 3952 -1542 3964 -1540
rect 3906 -1548 3964 -1542
rect 4706 -1542 4718 -1540
rect 4752 -1510 4764 -1508
rect 5506 -1508 5564 -1502
rect 5506 -1510 5518 -1508
rect 4752 -1540 5518 -1510
rect 4752 -1542 4764 -1540
rect 4706 -1548 4764 -1542
rect 5506 -1542 5518 -1540
rect 5552 -1510 5564 -1508
rect 6306 -1508 6364 -1502
rect 6306 -1510 6318 -1508
rect 5552 -1540 6318 -1510
rect 5552 -1542 5564 -1540
rect 5506 -1548 5564 -1542
rect 6306 -1542 6318 -1540
rect 6352 -1510 6364 -1508
rect 8120 -1508 8736 -1502
rect 8120 -1510 8160 -1508
rect 6352 -1540 6376 -1510
rect 8000 -1540 8160 -1510
rect 6352 -1542 6364 -1540
rect 6306 -1548 6364 -1542
rect 8120 -1542 8160 -1540
rect 8194 -1542 8232 -1508
rect 8266 -1542 8441 -1508
rect 8475 -1542 8513 -1508
rect 8547 -1542 8585 -1508
rect 8619 -1542 8657 -1508
rect 8691 -1542 8736 -1508
rect 8120 -1548 8736 -1542
rect 8806 -1551 8812 -1499
rect 8864 -1502 8870 -1499
rect 8864 -1508 9422 -1502
rect 8885 -1542 8923 -1508
rect 8957 -1542 8995 -1508
rect 9029 -1542 9067 -1508
rect 9101 -1542 9276 -1508
rect 9310 -1542 9348 -1508
rect 9382 -1542 9422 -1508
rect 8864 -1548 9422 -1542
rect 8864 -1551 8870 -1548
rect 8126 -1599 8297 -1593
rect -94 -1608 -36 -1602
rect -94 -1610 -82 -1608
rect -106 -1640 -82 -1610
rect -94 -1642 -82 -1640
rect -48 -1610 -36 -1608
rect 706 -1608 764 -1602
rect 706 -1610 718 -1608
rect -48 -1640 718 -1610
rect -48 -1642 -36 -1640
rect -94 -1648 -36 -1642
rect 706 -1642 718 -1640
rect 752 -1610 764 -1608
rect 1506 -1608 1564 -1602
rect 1506 -1610 1518 -1608
rect 752 -1640 1518 -1610
rect 752 -1642 764 -1640
rect 706 -1648 764 -1642
rect 1506 -1642 1518 -1640
rect 1552 -1610 1564 -1608
rect 2306 -1608 2364 -1602
rect 2306 -1610 2318 -1608
rect 1552 -1640 2318 -1610
rect 1552 -1642 1564 -1640
rect 1506 -1648 1564 -1642
rect 2306 -1642 2318 -1640
rect 2352 -1610 2364 -1608
rect 3106 -1608 3164 -1602
rect 3106 -1610 3118 -1608
rect 2352 -1640 3118 -1610
rect 2352 -1642 2364 -1640
rect 2306 -1648 2364 -1642
rect 3106 -1642 3118 -1640
rect 3152 -1610 3164 -1608
rect 3906 -1608 3964 -1602
rect 3906 -1610 3918 -1608
rect 3152 -1640 3918 -1610
rect 3152 -1642 3164 -1640
rect 3106 -1648 3164 -1642
rect 3906 -1642 3918 -1640
rect 3952 -1610 3964 -1608
rect 4706 -1608 4764 -1602
rect 4706 -1610 4718 -1608
rect 3952 -1640 4718 -1610
rect 3952 -1642 3964 -1640
rect 3906 -1648 3964 -1642
rect 4706 -1642 4718 -1640
rect 4752 -1610 4764 -1608
rect 5506 -1608 5564 -1602
rect 5506 -1610 5518 -1608
rect 4752 -1640 5518 -1610
rect 4752 -1642 4764 -1640
rect 4706 -1648 4764 -1642
rect 5506 -1642 5518 -1640
rect 5552 -1610 5564 -1608
rect 6306 -1608 6364 -1602
rect 6306 -1610 6318 -1608
rect 5552 -1640 6318 -1610
rect 5552 -1642 5564 -1640
rect 5506 -1648 5564 -1642
rect 6306 -1642 6318 -1640
rect 6352 -1610 6364 -1608
rect 8034 -1610 8040 -1599
rect 6352 -1640 6376 -1610
rect 8000 -1640 8040 -1610
rect 6352 -1642 6364 -1640
rect 6306 -1648 6364 -1642
rect 8034 -1651 8040 -1640
rect 8092 -1651 8098 -1599
rect 8126 -1651 8153 -1599
rect 8205 -1651 8217 -1599
rect 8269 -1651 8297 -1599
rect 8126 -1657 8297 -1651
rect 8325 -1599 8377 -1593
rect 8325 -1657 8377 -1651
rect 8405 -1599 8736 -1593
rect 8405 -1651 8416 -1599
rect 8468 -1608 8480 -1599
rect 8532 -1608 8544 -1599
rect 8596 -1608 8608 -1599
rect 8660 -1608 8672 -1599
rect 8476 -1642 8480 -1608
rect 8468 -1651 8480 -1642
rect 8532 -1651 8544 -1642
rect 8596 -1651 8608 -1642
rect 8660 -1651 8672 -1642
rect 8724 -1651 8736 -1599
rect 8405 -1657 8736 -1651
rect 8806 -1599 9137 -1593
rect 8806 -1651 8817 -1599
rect 8869 -1608 8881 -1599
rect 8933 -1608 8945 -1599
rect 8997 -1608 9009 -1599
rect 9061 -1608 9073 -1599
rect 9061 -1642 9065 -1608
rect 8869 -1651 8881 -1642
rect 8933 -1651 8945 -1642
rect 8997 -1651 9009 -1642
rect 9061 -1651 9073 -1642
rect 9125 -1651 9137 -1599
rect 8806 -1657 9137 -1651
rect 9165 -1599 9217 -1593
rect 9165 -1657 9217 -1651
rect 9245 -1599 9416 -1593
rect 9245 -1651 9272 -1599
rect 9324 -1651 9336 -1599
rect 9388 -1651 9416 -1599
rect 9245 -1657 9416 -1651
rect -94 -1708 -36 -1702
rect -94 -1710 -82 -1708
rect -106 -1740 -82 -1710
rect -94 -1742 -82 -1740
rect -48 -1710 -36 -1708
rect 706 -1708 764 -1702
rect 706 -1710 718 -1708
rect -48 -1740 718 -1710
rect -48 -1742 -36 -1740
rect -94 -1748 -36 -1742
rect 706 -1742 718 -1740
rect 752 -1710 764 -1708
rect 1506 -1708 1564 -1702
rect 1506 -1710 1518 -1708
rect 752 -1740 1518 -1710
rect 752 -1742 764 -1740
rect 706 -1748 764 -1742
rect 1506 -1742 1518 -1740
rect 1552 -1710 1564 -1708
rect 2306 -1708 2364 -1702
rect 2306 -1710 2318 -1708
rect 1552 -1740 2318 -1710
rect 1552 -1742 1564 -1740
rect 1506 -1748 1564 -1742
rect 2306 -1742 2318 -1740
rect 2352 -1710 2364 -1708
rect 3106 -1708 3164 -1702
rect 3106 -1710 3118 -1708
rect 2352 -1740 3118 -1710
rect 2352 -1742 2364 -1740
rect 2306 -1748 2364 -1742
rect 3106 -1742 3118 -1740
rect 3152 -1710 3164 -1708
rect 3906 -1708 3964 -1702
rect 3906 -1710 3918 -1708
rect 3152 -1740 3918 -1710
rect 3152 -1742 3164 -1740
rect 3106 -1748 3164 -1742
rect 3906 -1742 3918 -1740
rect 3952 -1710 3964 -1708
rect 4706 -1708 4764 -1702
rect 4706 -1710 4718 -1708
rect 3952 -1740 4718 -1710
rect 3952 -1742 3964 -1740
rect 3906 -1748 3964 -1742
rect 4706 -1742 4718 -1740
rect 4752 -1710 4764 -1708
rect 5506 -1708 5564 -1702
rect 5506 -1710 5518 -1708
rect 4752 -1740 5518 -1710
rect 4752 -1742 4764 -1740
rect 4706 -1748 4764 -1742
rect 5506 -1742 5518 -1740
rect 5552 -1710 5564 -1708
rect 6306 -1708 6364 -1702
rect 6306 -1710 6318 -1708
rect 5552 -1740 6318 -1710
rect 5552 -1742 5564 -1740
rect 5506 -1748 5564 -1742
rect 6306 -1742 6318 -1740
rect 6352 -1710 6364 -1708
rect 8120 -1708 8736 -1702
rect 8120 -1710 8160 -1708
rect 6352 -1740 6376 -1710
rect 8000 -1740 8160 -1710
rect 6352 -1742 6364 -1740
rect 6306 -1748 6364 -1742
rect 8120 -1742 8160 -1740
rect 8194 -1742 8232 -1708
rect 8266 -1742 8441 -1708
rect 8475 -1742 8513 -1708
rect 8547 -1742 8585 -1708
rect 8619 -1742 8657 -1708
rect 8691 -1742 8736 -1708
rect 8120 -1748 8736 -1742
rect 8806 -1751 8812 -1699
rect 8864 -1702 8870 -1699
rect 8864 -1708 9422 -1702
rect 8885 -1742 8923 -1708
rect 8957 -1742 8995 -1708
rect 9029 -1742 9067 -1708
rect 9101 -1742 9276 -1708
rect 9310 -1742 9348 -1708
rect 9382 -1742 9422 -1708
rect 8864 -1748 9422 -1742
rect 8864 -1751 8870 -1748
rect 8126 -1799 8297 -1793
rect -94 -1808 -36 -1802
rect -94 -1810 -82 -1808
rect -106 -1840 -82 -1810
rect -94 -1842 -82 -1840
rect -48 -1810 -36 -1808
rect 706 -1808 764 -1802
rect 706 -1810 718 -1808
rect -48 -1840 718 -1810
rect -48 -1842 -36 -1840
rect -94 -1848 -36 -1842
rect 706 -1842 718 -1840
rect 752 -1810 764 -1808
rect 1506 -1808 1564 -1802
rect 1506 -1810 1518 -1808
rect 752 -1840 1518 -1810
rect 752 -1842 764 -1840
rect 706 -1848 764 -1842
rect 1506 -1842 1518 -1840
rect 1552 -1810 1564 -1808
rect 2306 -1808 2364 -1802
rect 2306 -1810 2318 -1808
rect 1552 -1840 2318 -1810
rect 1552 -1842 1564 -1840
rect 1506 -1848 1564 -1842
rect 2306 -1842 2318 -1840
rect 2352 -1810 2364 -1808
rect 3106 -1808 3164 -1802
rect 3106 -1810 3118 -1808
rect 2352 -1840 3118 -1810
rect 2352 -1842 2364 -1840
rect 2306 -1848 2364 -1842
rect 3106 -1842 3118 -1840
rect 3152 -1810 3164 -1808
rect 3906 -1808 3964 -1802
rect 3906 -1810 3918 -1808
rect 3152 -1840 3918 -1810
rect 3152 -1842 3164 -1840
rect 3106 -1848 3164 -1842
rect 3906 -1842 3918 -1840
rect 3952 -1810 3964 -1808
rect 4706 -1808 4764 -1802
rect 4706 -1810 4718 -1808
rect 3952 -1840 4718 -1810
rect 3952 -1842 3964 -1840
rect 3906 -1848 3964 -1842
rect 4706 -1842 4718 -1840
rect 4752 -1810 4764 -1808
rect 5506 -1808 5564 -1802
rect 5506 -1810 5518 -1808
rect 4752 -1840 5518 -1810
rect 4752 -1842 4764 -1840
rect 4706 -1848 4764 -1842
rect 5506 -1842 5518 -1840
rect 5552 -1810 5564 -1808
rect 6306 -1808 6364 -1802
rect 6306 -1810 6318 -1808
rect 5552 -1840 6318 -1810
rect 5552 -1842 5564 -1840
rect 5506 -1848 5564 -1842
rect 6306 -1842 6318 -1840
rect 6352 -1810 6364 -1808
rect 8034 -1810 8040 -1799
rect 6352 -1840 6376 -1810
rect 8000 -1840 8040 -1810
rect 6352 -1842 6364 -1840
rect 6306 -1848 6364 -1842
rect 8034 -1851 8040 -1840
rect 8092 -1851 8098 -1799
rect 8126 -1851 8153 -1799
rect 8205 -1851 8217 -1799
rect 8269 -1851 8297 -1799
rect 8126 -1857 8297 -1851
rect 8325 -1799 8377 -1793
rect 8325 -1857 8377 -1851
rect 8405 -1799 8736 -1793
rect 8405 -1851 8416 -1799
rect 8468 -1808 8480 -1799
rect 8532 -1808 8544 -1799
rect 8596 -1808 8608 -1799
rect 8660 -1808 8672 -1799
rect 8476 -1842 8480 -1808
rect 8468 -1851 8480 -1842
rect 8532 -1851 8544 -1842
rect 8596 -1851 8608 -1842
rect 8660 -1851 8672 -1842
rect 8724 -1851 8736 -1799
rect 8405 -1857 8736 -1851
rect 8806 -1799 9137 -1793
rect 8806 -1851 8817 -1799
rect 8869 -1808 8881 -1799
rect 8933 -1808 8945 -1799
rect 8997 -1808 9009 -1799
rect 9061 -1808 9073 -1799
rect 9061 -1842 9065 -1808
rect 8869 -1851 8881 -1842
rect 8933 -1851 8945 -1842
rect 8997 -1851 9009 -1842
rect 9061 -1851 9073 -1842
rect 9125 -1851 9137 -1799
rect 8806 -1857 9137 -1851
rect 9165 -1799 9217 -1793
rect 9165 -1857 9217 -1851
rect 9245 -1799 9416 -1793
rect 9245 -1851 9272 -1799
rect 9324 -1851 9336 -1799
rect 9388 -1851 9416 -1799
rect 9245 -1857 9416 -1851
rect -65 -1935 6335 -1917
rect -65 -1969 -4 -1935
rect 30 -1969 68 -1935
rect 102 -1969 168 -1935
rect 202 -1969 240 -1935
rect 274 -1969 396 -1935
rect 430 -1969 468 -1935
rect 502 -1969 568 -1935
rect 602 -1969 640 -1935
rect 674 -1969 796 -1935
rect 830 -1969 868 -1935
rect 902 -1969 968 -1935
rect 1002 -1969 1040 -1935
rect 1074 -1969 1196 -1935
rect 1230 -1969 1268 -1935
rect 1302 -1969 1368 -1935
rect 1402 -1969 1440 -1935
rect 1474 -1969 1596 -1935
rect 1630 -1969 1668 -1935
rect 1702 -1969 1768 -1935
rect 1802 -1969 1840 -1935
rect 1874 -1969 1996 -1935
rect 2030 -1969 2068 -1935
rect 2102 -1969 2168 -1935
rect 2202 -1969 2240 -1935
rect 2274 -1969 2396 -1935
rect 2430 -1969 2468 -1935
rect 2502 -1969 2568 -1935
rect 2602 -1969 2640 -1935
rect 2674 -1969 2796 -1935
rect 2830 -1969 2868 -1935
rect 2902 -1969 2968 -1935
rect 3002 -1969 3040 -1935
rect 3074 -1969 3196 -1935
rect 3230 -1969 3268 -1935
rect 3302 -1969 3368 -1935
rect 3402 -1969 3440 -1935
rect 3474 -1969 3596 -1935
rect 3630 -1969 3668 -1935
rect 3702 -1969 3768 -1935
rect 3802 -1969 3840 -1935
rect 3874 -1969 3996 -1935
rect 4030 -1969 4068 -1935
rect 4102 -1969 4168 -1935
rect 4202 -1969 4240 -1935
rect 4274 -1969 4396 -1935
rect 4430 -1969 4468 -1935
rect 4502 -1969 4568 -1935
rect 4602 -1969 4640 -1935
rect 4674 -1969 4796 -1935
rect 4830 -1969 4868 -1935
rect 4902 -1969 4968 -1935
rect 5002 -1969 5040 -1935
rect 5074 -1969 5196 -1935
rect 5230 -1969 5268 -1935
rect 5302 -1969 5368 -1935
rect 5402 -1969 5440 -1935
rect 5474 -1969 5596 -1935
rect 5630 -1969 5668 -1935
rect 5702 -1969 5768 -1935
rect 5802 -1969 5840 -1935
rect 5874 -1969 5996 -1935
rect 6030 -1969 6068 -1935
rect 6102 -1969 6168 -1935
rect 6202 -1969 6240 -1935
rect 6274 -1969 6335 -1935
rect -65 -1987 6335 -1969
<< via1 >>
rect 9 9874 61 9883
rect 9 9840 18 9874
rect 18 9840 52 9874
rect 52 9840 61 9874
rect 9 9831 61 9840
rect 9 9733 18 9741
rect 18 9733 52 9741
rect 52 9733 61 9741
rect 9 9689 61 9733
rect 209 9890 261 9899
rect 209 9856 218 9890
rect 218 9856 252 9890
rect 252 9856 261 9890
rect 209 9847 261 9856
rect 9 9593 18 9601
rect 18 9593 52 9601
rect 52 9593 61 9601
rect 9 9549 61 9593
rect 209 9767 261 9811
rect 209 9759 218 9767
rect 218 9759 252 9767
rect 252 9759 261 9767
rect 409 9874 461 9883
rect 409 9840 418 9874
rect 418 9840 452 9874
rect 452 9840 461 9874
rect 409 9831 461 9840
rect 9 9453 18 9461
rect 18 9453 52 9461
rect 52 9453 61 9461
rect 9 9409 61 9453
rect 209 9627 261 9671
rect 209 9619 218 9627
rect 218 9619 252 9627
rect 252 9619 261 9627
rect 409 9733 418 9741
rect 418 9733 452 9741
rect 452 9733 461 9741
rect 409 9689 461 9733
rect 609 9890 661 9899
rect 609 9856 618 9890
rect 618 9856 652 9890
rect 652 9856 661 9890
rect 609 9847 661 9856
rect 9 9313 18 9321
rect 18 9313 52 9321
rect 52 9313 61 9321
rect 9 9269 61 9313
rect 209 9487 261 9531
rect 209 9479 218 9487
rect 218 9479 252 9487
rect 252 9479 261 9487
rect 409 9593 418 9601
rect 418 9593 452 9601
rect 452 9593 461 9601
rect 409 9549 461 9593
rect 609 9767 661 9811
rect 609 9759 618 9767
rect 618 9759 652 9767
rect 652 9759 661 9767
rect 809 9874 861 9883
rect 809 9840 818 9874
rect 818 9840 852 9874
rect 852 9840 861 9874
rect 809 9831 861 9840
rect 9 9173 18 9181
rect 18 9173 52 9181
rect 52 9173 61 9181
rect 9 9129 61 9173
rect 209 9347 261 9391
rect 209 9339 218 9347
rect 218 9339 252 9347
rect 252 9339 261 9347
rect 409 9453 418 9461
rect 418 9453 452 9461
rect 452 9453 461 9461
rect 409 9409 461 9453
rect 609 9627 661 9671
rect 609 9619 618 9627
rect 618 9619 652 9627
rect 652 9619 661 9627
rect 809 9733 818 9741
rect 818 9733 852 9741
rect 852 9733 861 9741
rect 809 9689 861 9733
rect 1009 9890 1061 9899
rect 1009 9856 1018 9890
rect 1018 9856 1052 9890
rect 1052 9856 1061 9890
rect 1009 9847 1061 9856
rect 9 9033 18 9041
rect 18 9033 52 9041
rect 52 9033 61 9041
rect 9 8989 61 9033
rect 209 9207 261 9251
rect 209 9199 218 9207
rect 218 9199 252 9207
rect 252 9199 261 9207
rect 409 9313 418 9321
rect 418 9313 452 9321
rect 452 9313 461 9321
rect 409 9269 461 9313
rect 609 9487 661 9531
rect 609 9479 618 9487
rect 618 9479 652 9487
rect 652 9479 661 9487
rect 809 9593 818 9601
rect 818 9593 852 9601
rect 852 9593 861 9601
rect 809 9549 861 9593
rect 1009 9767 1061 9811
rect 1009 9759 1018 9767
rect 1018 9759 1052 9767
rect 1052 9759 1061 9767
rect 1209 9874 1261 9883
rect 1209 9840 1218 9874
rect 1218 9840 1252 9874
rect 1252 9840 1261 9874
rect 1209 9831 1261 9840
rect 9 8893 18 8901
rect 18 8893 52 8901
rect 52 8893 61 8901
rect 9 8849 61 8893
rect 209 9067 261 9111
rect 209 9059 218 9067
rect 218 9059 252 9067
rect 252 9059 261 9067
rect 409 9173 418 9181
rect 418 9173 452 9181
rect 452 9173 461 9181
rect 409 9129 461 9173
rect 609 9347 661 9391
rect 609 9339 618 9347
rect 618 9339 652 9347
rect 652 9339 661 9347
rect 809 9453 818 9461
rect 818 9453 852 9461
rect 852 9453 861 9461
rect 809 9409 861 9453
rect 1009 9627 1061 9671
rect 1009 9619 1018 9627
rect 1018 9619 1052 9627
rect 1052 9619 1061 9627
rect 1209 9733 1218 9741
rect 1218 9733 1252 9741
rect 1252 9733 1261 9741
rect 1209 9689 1261 9733
rect 1409 9890 1461 9899
rect 1409 9856 1418 9890
rect 1418 9856 1452 9890
rect 1452 9856 1461 9890
rect 1409 9847 1461 9856
rect 9 8753 18 8761
rect 18 8753 52 8761
rect 52 8753 61 8761
rect 9 8709 61 8753
rect 209 8927 261 8971
rect 209 8919 218 8927
rect 218 8919 252 8927
rect 252 8919 261 8927
rect 409 9033 418 9041
rect 418 9033 452 9041
rect 452 9033 461 9041
rect 409 8989 461 9033
rect 609 9207 661 9251
rect 609 9199 618 9207
rect 618 9199 652 9207
rect 652 9199 661 9207
rect 809 9313 818 9321
rect 818 9313 852 9321
rect 852 9313 861 9321
rect 809 9269 861 9313
rect 1009 9487 1061 9531
rect 1009 9479 1018 9487
rect 1018 9479 1052 9487
rect 1052 9479 1061 9487
rect 1209 9593 1218 9601
rect 1218 9593 1252 9601
rect 1252 9593 1261 9601
rect 1209 9549 1261 9593
rect 1409 9767 1461 9811
rect 1409 9759 1418 9767
rect 1418 9759 1452 9767
rect 1452 9759 1461 9767
rect 1609 9874 1661 9883
rect 1609 9840 1618 9874
rect 1618 9840 1652 9874
rect 1652 9840 1661 9874
rect 1609 9831 1661 9840
rect 9 8664 61 8673
rect 9 8630 18 8664
rect 18 8630 52 8664
rect 52 8630 61 8664
rect 9 8621 61 8630
rect 9 8523 18 8531
rect 18 8523 52 8531
rect 52 8523 61 8531
rect 9 8479 61 8523
rect 209 8787 261 8831
rect 209 8779 218 8787
rect 218 8779 252 8787
rect 252 8779 261 8787
rect 409 8893 418 8901
rect 418 8893 452 8901
rect 452 8893 461 8901
rect 409 8849 461 8893
rect 609 9067 661 9111
rect 609 9059 618 9067
rect 618 9059 652 9067
rect 652 9059 661 9067
rect 809 9173 818 9181
rect 818 9173 852 9181
rect 852 9173 861 9181
rect 809 9129 861 9173
rect 1009 9347 1061 9391
rect 1009 9339 1018 9347
rect 1018 9339 1052 9347
rect 1052 9339 1061 9347
rect 1209 9453 1218 9461
rect 1218 9453 1252 9461
rect 1252 9453 1261 9461
rect 1209 9409 1261 9453
rect 1409 9627 1461 9671
rect 1409 9619 1418 9627
rect 1418 9619 1452 9627
rect 1452 9619 1461 9627
rect 1609 9733 1618 9741
rect 1618 9733 1652 9741
rect 1652 9733 1661 9741
rect 1609 9689 1661 9733
rect 1809 9890 1861 9899
rect 1809 9856 1818 9890
rect 1818 9856 1852 9890
rect 1852 9856 1861 9890
rect 1809 9847 1861 9856
rect 209 8680 261 8689
rect 209 8646 218 8680
rect 218 8646 252 8680
rect 252 8646 261 8680
rect 209 8637 261 8646
rect 9 8383 18 8391
rect 18 8383 52 8391
rect 52 8383 61 8391
rect 9 8339 61 8383
rect 209 8557 261 8601
rect 209 8549 218 8557
rect 218 8549 252 8557
rect 252 8549 261 8557
rect 409 8753 418 8761
rect 418 8753 452 8761
rect 452 8753 461 8761
rect 409 8709 461 8753
rect 609 8927 661 8971
rect 609 8919 618 8927
rect 618 8919 652 8927
rect 652 8919 661 8927
rect 809 9033 818 9041
rect 818 9033 852 9041
rect 852 9033 861 9041
rect 809 8989 861 9033
rect 1009 9207 1061 9251
rect 1009 9199 1018 9207
rect 1018 9199 1052 9207
rect 1052 9199 1061 9207
rect 1209 9313 1218 9321
rect 1218 9313 1252 9321
rect 1252 9313 1261 9321
rect 1209 9269 1261 9313
rect 1409 9487 1461 9531
rect 1409 9479 1418 9487
rect 1418 9479 1452 9487
rect 1452 9479 1461 9487
rect 1609 9593 1618 9601
rect 1618 9593 1652 9601
rect 1652 9593 1661 9601
rect 1609 9549 1661 9593
rect 1809 9767 1861 9811
rect 1809 9759 1818 9767
rect 1818 9759 1852 9767
rect 1852 9759 1861 9767
rect 2009 9874 2061 9883
rect 2009 9840 2018 9874
rect 2018 9840 2052 9874
rect 2052 9840 2061 9874
rect 2009 9831 2061 9840
rect 409 8664 461 8673
rect 409 8630 418 8664
rect 418 8630 452 8664
rect 452 8630 461 8664
rect 409 8621 461 8630
rect 9 8243 18 8251
rect 18 8243 52 8251
rect 52 8243 61 8251
rect 9 8199 61 8243
rect 209 8417 261 8461
rect 209 8409 218 8417
rect 218 8409 252 8417
rect 252 8409 261 8417
rect 409 8523 418 8531
rect 418 8523 452 8531
rect 452 8523 461 8531
rect 409 8479 461 8523
rect 609 8787 661 8831
rect 609 8779 618 8787
rect 618 8779 652 8787
rect 652 8779 661 8787
rect 809 8893 818 8901
rect 818 8893 852 8901
rect 852 8893 861 8901
rect 809 8849 861 8893
rect 1009 9067 1061 9111
rect 1009 9059 1018 9067
rect 1018 9059 1052 9067
rect 1052 9059 1061 9067
rect 1209 9173 1218 9181
rect 1218 9173 1252 9181
rect 1252 9173 1261 9181
rect 1209 9129 1261 9173
rect 1409 9347 1461 9391
rect 1409 9339 1418 9347
rect 1418 9339 1452 9347
rect 1452 9339 1461 9347
rect 1609 9453 1618 9461
rect 1618 9453 1652 9461
rect 1652 9453 1661 9461
rect 1609 9409 1661 9453
rect 1809 9627 1861 9671
rect 1809 9619 1818 9627
rect 1818 9619 1852 9627
rect 1852 9619 1861 9627
rect 2009 9733 2018 9741
rect 2018 9733 2052 9741
rect 2052 9733 2061 9741
rect 2009 9689 2061 9733
rect 2209 9890 2261 9899
rect 2209 9856 2218 9890
rect 2218 9856 2252 9890
rect 2252 9856 2261 9890
rect 2209 9847 2261 9856
rect 609 8680 661 8689
rect 609 8646 618 8680
rect 618 8646 652 8680
rect 652 8646 661 8680
rect 609 8637 661 8646
rect 9 8103 18 8111
rect 18 8103 52 8111
rect 52 8103 61 8111
rect 9 8059 61 8103
rect 209 8277 261 8321
rect 209 8269 218 8277
rect 218 8269 252 8277
rect 252 8269 261 8277
rect 409 8383 418 8391
rect 418 8383 452 8391
rect 452 8383 461 8391
rect 409 8339 461 8383
rect 609 8557 661 8601
rect 609 8549 618 8557
rect 618 8549 652 8557
rect 652 8549 661 8557
rect 809 8753 818 8761
rect 818 8753 852 8761
rect 852 8753 861 8761
rect 809 8709 861 8753
rect 1009 8927 1061 8971
rect 1009 8919 1018 8927
rect 1018 8919 1052 8927
rect 1052 8919 1061 8927
rect 1209 9033 1218 9041
rect 1218 9033 1252 9041
rect 1252 9033 1261 9041
rect 1209 8989 1261 9033
rect 1409 9207 1461 9251
rect 1409 9199 1418 9207
rect 1418 9199 1452 9207
rect 1452 9199 1461 9207
rect 1609 9313 1618 9321
rect 1618 9313 1652 9321
rect 1652 9313 1661 9321
rect 1609 9269 1661 9313
rect 1809 9487 1861 9531
rect 1809 9479 1818 9487
rect 1818 9479 1852 9487
rect 1852 9479 1861 9487
rect 2009 9593 2018 9601
rect 2018 9593 2052 9601
rect 2052 9593 2061 9601
rect 2009 9549 2061 9593
rect 2209 9767 2261 9811
rect 2209 9759 2218 9767
rect 2218 9759 2252 9767
rect 2252 9759 2261 9767
rect 2409 9874 2461 9883
rect 2409 9840 2418 9874
rect 2418 9840 2452 9874
rect 2452 9840 2461 9874
rect 2409 9831 2461 9840
rect 809 8664 861 8673
rect 809 8630 818 8664
rect 818 8630 852 8664
rect 852 8630 861 8664
rect 809 8621 861 8630
rect 9 7963 18 7971
rect 18 7963 52 7971
rect 52 7963 61 7971
rect 9 7919 61 7963
rect 209 8137 261 8181
rect 209 8129 218 8137
rect 218 8129 252 8137
rect 252 8129 261 8137
rect 409 8243 418 8251
rect 418 8243 452 8251
rect 452 8243 461 8251
rect 409 8199 461 8243
rect 609 8417 661 8461
rect 609 8409 618 8417
rect 618 8409 652 8417
rect 652 8409 661 8417
rect 809 8523 818 8531
rect 818 8523 852 8531
rect 852 8523 861 8531
rect 809 8479 861 8523
rect 1009 8787 1061 8831
rect 1009 8779 1018 8787
rect 1018 8779 1052 8787
rect 1052 8779 1061 8787
rect 1209 8893 1218 8901
rect 1218 8893 1252 8901
rect 1252 8893 1261 8901
rect 1209 8849 1261 8893
rect 1409 9067 1461 9111
rect 1409 9059 1418 9067
rect 1418 9059 1452 9067
rect 1452 9059 1461 9067
rect 1609 9173 1618 9181
rect 1618 9173 1652 9181
rect 1652 9173 1661 9181
rect 1609 9129 1661 9173
rect 1809 9347 1861 9391
rect 1809 9339 1818 9347
rect 1818 9339 1852 9347
rect 1852 9339 1861 9347
rect 2009 9453 2018 9461
rect 2018 9453 2052 9461
rect 2052 9453 2061 9461
rect 2009 9409 2061 9453
rect 2209 9627 2261 9671
rect 2209 9619 2218 9627
rect 2218 9619 2252 9627
rect 2252 9619 2261 9627
rect 2409 9733 2418 9741
rect 2418 9733 2452 9741
rect 2452 9733 2461 9741
rect 2409 9689 2461 9733
rect 2609 9890 2661 9899
rect 2609 9856 2618 9890
rect 2618 9856 2652 9890
rect 2652 9856 2661 9890
rect 2609 9847 2661 9856
rect 1009 8680 1061 8689
rect 1009 8646 1018 8680
rect 1018 8646 1052 8680
rect 1052 8646 1061 8680
rect 1009 8637 1061 8646
rect 9 7823 18 7831
rect 18 7823 52 7831
rect 52 7823 61 7831
rect 9 7779 61 7823
rect 209 7997 261 8041
rect 209 7989 218 7997
rect 218 7989 252 7997
rect 252 7989 261 7997
rect 409 8103 418 8111
rect 418 8103 452 8111
rect 452 8103 461 8111
rect 409 8059 461 8103
rect 609 8277 661 8321
rect 609 8269 618 8277
rect 618 8269 652 8277
rect 652 8269 661 8277
rect 809 8383 818 8391
rect 818 8383 852 8391
rect 852 8383 861 8391
rect 809 8339 861 8383
rect 1009 8557 1061 8601
rect 1009 8549 1018 8557
rect 1018 8549 1052 8557
rect 1052 8549 1061 8557
rect 1209 8753 1218 8761
rect 1218 8753 1252 8761
rect 1252 8753 1261 8761
rect 1209 8709 1261 8753
rect 1409 8927 1461 8971
rect 1409 8919 1418 8927
rect 1418 8919 1452 8927
rect 1452 8919 1461 8927
rect 1609 9033 1618 9041
rect 1618 9033 1652 9041
rect 1652 9033 1661 9041
rect 1609 8989 1661 9033
rect 1809 9207 1861 9251
rect 1809 9199 1818 9207
rect 1818 9199 1852 9207
rect 1852 9199 1861 9207
rect 2009 9313 2018 9321
rect 2018 9313 2052 9321
rect 2052 9313 2061 9321
rect 2009 9269 2061 9313
rect 2209 9487 2261 9531
rect 2209 9479 2218 9487
rect 2218 9479 2252 9487
rect 2252 9479 2261 9487
rect 2409 9593 2418 9601
rect 2418 9593 2452 9601
rect 2452 9593 2461 9601
rect 2409 9549 2461 9593
rect 2609 9767 2661 9811
rect 2609 9759 2618 9767
rect 2618 9759 2652 9767
rect 2652 9759 2661 9767
rect 2809 9874 2861 9883
rect 2809 9840 2818 9874
rect 2818 9840 2852 9874
rect 2852 9840 2861 9874
rect 2809 9831 2861 9840
rect 1209 8664 1261 8673
rect 1209 8630 1218 8664
rect 1218 8630 1252 8664
rect 1252 8630 1261 8664
rect 1209 8621 1261 8630
rect 9 7683 18 7691
rect 18 7683 52 7691
rect 52 7683 61 7691
rect 9 7639 61 7683
rect 209 7857 261 7901
rect 209 7849 218 7857
rect 218 7849 252 7857
rect 252 7849 261 7857
rect 409 7963 418 7971
rect 418 7963 452 7971
rect 452 7963 461 7971
rect 409 7919 461 7963
rect 609 8137 661 8181
rect 609 8129 618 8137
rect 618 8129 652 8137
rect 652 8129 661 8137
rect 809 8243 818 8251
rect 818 8243 852 8251
rect 852 8243 861 8251
rect 809 8199 861 8243
rect 1009 8417 1061 8461
rect 1009 8409 1018 8417
rect 1018 8409 1052 8417
rect 1052 8409 1061 8417
rect 1209 8523 1218 8531
rect 1218 8523 1252 8531
rect 1252 8523 1261 8531
rect 1209 8479 1261 8523
rect 1409 8787 1461 8831
rect 1409 8779 1418 8787
rect 1418 8779 1452 8787
rect 1452 8779 1461 8787
rect 1609 8893 1618 8901
rect 1618 8893 1652 8901
rect 1652 8893 1661 8901
rect 1609 8849 1661 8893
rect 1809 9067 1861 9111
rect 1809 9059 1818 9067
rect 1818 9059 1852 9067
rect 1852 9059 1861 9067
rect 2009 9173 2018 9181
rect 2018 9173 2052 9181
rect 2052 9173 2061 9181
rect 2009 9129 2061 9173
rect 2209 9347 2261 9391
rect 2209 9339 2218 9347
rect 2218 9339 2252 9347
rect 2252 9339 2261 9347
rect 2409 9453 2418 9461
rect 2418 9453 2452 9461
rect 2452 9453 2461 9461
rect 2409 9409 2461 9453
rect 2609 9627 2661 9671
rect 2609 9619 2618 9627
rect 2618 9619 2652 9627
rect 2652 9619 2661 9627
rect 2809 9733 2818 9741
rect 2818 9733 2852 9741
rect 2852 9733 2861 9741
rect 2809 9689 2861 9733
rect 3009 9890 3061 9899
rect 3009 9856 3018 9890
rect 3018 9856 3052 9890
rect 3052 9856 3061 9890
rect 3009 9847 3061 9856
rect 1409 8680 1461 8689
rect 1409 8646 1418 8680
rect 1418 8646 1452 8680
rect 1452 8646 1461 8680
rect 1409 8637 1461 8646
rect 9 7543 18 7551
rect 18 7543 52 7551
rect 52 7543 61 7551
rect 9 7499 61 7543
rect 209 7717 261 7761
rect 209 7709 218 7717
rect 218 7709 252 7717
rect 252 7709 261 7717
rect 409 7823 418 7831
rect 418 7823 452 7831
rect 452 7823 461 7831
rect 409 7779 461 7823
rect 609 7997 661 8041
rect 609 7989 618 7997
rect 618 7989 652 7997
rect 652 7989 661 7997
rect 809 8103 818 8111
rect 818 8103 852 8111
rect 852 8103 861 8111
rect 809 8059 861 8103
rect 1009 8277 1061 8321
rect 1009 8269 1018 8277
rect 1018 8269 1052 8277
rect 1052 8269 1061 8277
rect 1209 8383 1218 8391
rect 1218 8383 1252 8391
rect 1252 8383 1261 8391
rect 1209 8339 1261 8383
rect 1409 8557 1461 8601
rect 1409 8549 1418 8557
rect 1418 8549 1452 8557
rect 1452 8549 1461 8557
rect 1609 8753 1618 8761
rect 1618 8753 1652 8761
rect 1652 8753 1661 8761
rect 1609 8709 1661 8753
rect 1809 8927 1861 8971
rect 1809 8919 1818 8927
rect 1818 8919 1852 8927
rect 1852 8919 1861 8927
rect 2009 9033 2018 9041
rect 2018 9033 2052 9041
rect 2052 9033 2061 9041
rect 2009 8989 2061 9033
rect 2209 9207 2261 9251
rect 2209 9199 2218 9207
rect 2218 9199 2252 9207
rect 2252 9199 2261 9207
rect 2409 9313 2418 9321
rect 2418 9313 2452 9321
rect 2452 9313 2461 9321
rect 2409 9269 2461 9313
rect 2609 9487 2661 9531
rect 2609 9479 2618 9487
rect 2618 9479 2652 9487
rect 2652 9479 2661 9487
rect 2809 9593 2818 9601
rect 2818 9593 2852 9601
rect 2852 9593 2861 9601
rect 2809 9549 2861 9593
rect 3009 9767 3061 9811
rect 3009 9759 3018 9767
rect 3018 9759 3052 9767
rect 3052 9759 3061 9767
rect 3209 9874 3261 9883
rect 3209 9840 3218 9874
rect 3218 9840 3252 9874
rect 3252 9840 3261 9874
rect 3209 9831 3261 9840
rect 1609 8664 1661 8673
rect 1609 8630 1618 8664
rect 1618 8630 1652 8664
rect 1652 8630 1661 8664
rect 1609 8621 1661 8630
rect 9 7454 61 7463
rect 9 7420 18 7454
rect 18 7420 52 7454
rect 52 7420 61 7454
rect 9 7411 61 7420
rect 9 7313 18 7321
rect 18 7313 52 7321
rect 52 7313 61 7321
rect 9 7269 61 7313
rect 209 7577 261 7621
rect 209 7569 218 7577
rect 218 7569 252 7577
rect 252 7569 261 7577
rect 409 7683 418 7691
rect 418 7683 452 7691
rect 452 7683 461 7691
rect 409 7639 461 7683
rect 609 7857 661 7901
rect 609 7849 618 7857
rect 618 7849 652 7857
rect 652 7849 661 7857
rect 809 7963 818 7971
rect 818 7963 852 7971
rect 852 7963 861 7971
rect 809 7919 861 7963
rect 1009 8137 1061 8181
rect 1009 8129 1018 8137
rect 1018 8129 1052 8137
rect 1052 8129 1061 8137
rect 1209 8243 1218 8251
rect 1218 8243 1252 8251
rect 1252 8243 1261 8251
rect 1209 8199 1261 8243
rect 1409 8417 1461 8461
rect 1409 8409 1418 8417
rect 1418 8409 1452 8417
rect 1452 8409 1461 8417
rect 1609 8523 1618 8531
rect 1618 8523 1652 8531
rect 1652 8523 1661 8531
rect 1609 8479 1661 8523
rect 1809 8787 1861 8831
rect 1809 8779 1818 8787
rect 1818 8779 1852 8787
rect 1852 8779 1861 8787
rect 2009 8893 2018 8901
rect 2018 8893 2052 8901
rect 2052 8893 2061 8901
rect 2009 8849 2061 8893
rect 2209 9067 2261 9111
rect 2209 9059 2218 9067
rect 2218 9059 2252 9067
rect 2252 9059 2261 9067
rect 2409 9173 2418 9181
rect 2418 9173 2452 9181
rect 2452 9173 2461 9181
rect 2409 9129 2461 9173
rect 2609 9347 2661 9391
rect 2609 9339 2618 9347
rect 2618 9339 2652 9347
rect 2652 9339 2661 9347
rect 2809 9453 2818 9461
rect 2818 9453 2852 9461
rect 2852 9453 2861 9461
rect 2809 9409 2861 9453
rect 3009 9627 3061 9671
rect 3009 9619 3018 9627
rect 3018 9619 3052 9627
rect 3052 9619 3061 9627
rect 3209 9733 3218 9741
rect 3218 9733 3252 9741
rect 3252 9733 3261 9741
rect 3209 9689 3261 9733
rect 3409 9890 3461 9899
rect 3409 9856 3418 9890
rect 3418 9856 3452 9890
rect 3452 9856 3461 9890
rect 3409 9847 3461 9856
rect 1809 8680 1861 8689
rect 1809 8646 1818 8680
rect 1818 8646 1852 8680
rect 1852 8646 1861 8680
rect 1809 8637 1861 8646
rect 209 7470 261 7479
rect 209 7436 218 7470
rect 218 7436 252 7470
rect 252 7436 261 7470
rect 209 7427 261 7436
rect 9 7173 18 7181
rect 18 7173 52 7181
rect 52 7173 61 7181
rect 9 7129 61 7173
rect 209 7347 261 7391
rect 209 7339 218 7347
rect 218 7339 252 7347
rect 252 7339 261 7347
rect 409 7543 418 7551
rect 418 7543 452 7551
rect 452 7543 461 7551
rect 409 7499 461 7543
rect 609 7717 661 7761
rect 609 7709 618 7717
rect 618 7709 652 7717
rect 652 7709 661 7717
rect 809 7823 818 7831
rect 818 7823 852 7831
rect 852 7823 861 7831
rect 809 7779 861 7823
rect 1009 7997 1061 8041
rect 1009 7989 1018 7997
rect 1018 7989 1052 7997
rect 1052 7989 1061 7997
rect 1209 8103 1218 8111
rect 1218 8103 1252 8111
rect 1252 8103 1261 8111
rect 1209 8059 1261 8103
rect 1409 8277 1461 8321
rect 1409 8269 1418 8277
rect 1418 8269 1452 8277
rect 1452 8269 1461 8277
rect 1609 8383 1618 8391
rect 1618 8383 1652 8391
rect 1652 8383 1661 8391
rect 1609 8339 1661 8383
rect 1809 8557 1861 8601
rect 1809 8549 1818 8557
rect 1818 8549 1852 8557
rect 1852 8549 1861 8557
rect 2009 8753 2018 8761
rect 2018 8753 2052 8761
rect 2052 8753 2061 8761
rect 2009 8709 2061 8753
rect 2209 8927 2261 8971
rect 2209 8919 2218 8927
rect 2218 8919 2252 8927
rect 2252 8919 2261 8927
rect 2409 9033 2418 9041
rect 2418 9033 2452 9041
rect 2452 9033 2461 9041
rect 2409 8989 2461 9033
rect 2609 9207 2661 9251
rect 2609 9199 2618 9207
rect 2618 9199 2652 9207
rect 2652 9199 2661 9207
rect 2809 9313 2818 9321
rect 2818 9313 2852 9321
rect 2852 9313 2861 9321
rect 2809 9269 2861 9313
rect 3009 9487 3061 9531
rect 3009 9479 3018 9487
rect 3018 9479 3052 9487
rect 3052 9479 3061 9487
rect 3209 9593 3218 9601
rect 3218 9593 3252 9601
rect 3252 9593 3261 9601
rect 3209 9549 3261 9593
rect 3409 9767 3461 9811
rect 3409 9759 3418 9767
rect 3418 9759 3452 9767
rect 3452 9759 3461 9767
rect 3609 9874 3661 9883
rect 3609 9840 3618 9874
rect 3618 9840 3652 9874
rect 3652 9840 3661 9874
rect 3609 9831 3661 9840
rect 2009 8664 2061 8673
rect 2009 8630 2018 8664
rect 2018 8630 2052 8664
rect 2052 8630 2061 8664
rect 2009 8621 2061 8630
rect 409 7454 461 7463
rect 409 7420 418 7454
rect 418 7420 452 7454
rect 452 7420 461 7454
rect 409 7411 461 7420
rect 9 7033 18 7041
rect 18 7033 52 7041
rect 52 7033 61 7041
rect 9 6989 61 7033
rect 209 7207 261 7251
rect 209 7199 218 7207
rect 218 7199 252 7207
rect 252 7199 261 7207
rect 409 7313 418 7321
rect 418 7313 452 7321
rect 452 7313 461 7321
rect 409 7269 461 7313
rect 609 7577 661 7621
rect 609 7569 618 7577
rect 618 7569 652 7577
rect 652 7569 661 7577
rect 809 7683 818 7691
rect 818 7683 852 7691
rect 852 7683 861 7691
rect 809 7639 861 7683
rect 1009 7857 1061 7901
rect 1009 7849 1018 7857
rect 1018 7849 1052 7857
rect 1052 7849 1061 7857
rect 1209 7963 1218 7971
rect 1218 7963 1252 7971
rect 1252 7963 1261 7971
rect 1209 7919 1261 7963
rect 1409 8137 1461 8181
rect 1409 8129 1418 8137
rect 1418 8129 1452 8137
rect 1452 8129 1461 8137
rect 1609 8243 1618 8251
rect 1618 8243 1652 8251
rect 1652 8243 1661 8251
rect 1609 8199 1661 8243
rect 1809 8417 1861 8461
rect 1809 8409 1818 8417
rect 1818 8409 1852 8417
rect 1852 8409 1861 8417
rect 2009 8523 2018 8531
rect 2018 8523 2052 8531
rect 2052 8523 2061 8531
rect 2009 8479 2061 8523
rect 2209 8787 2261 8831
rect 2209 8779 2218 8787
rect 2218 8779 2252 8787
rect 2252 8779 2261 8787
rect 2409 8893 2418 8901
rect 2418 8893 2452 8901
rect 2452 8893 2461 8901
rect 2409 8849 2461 8893
rect 2609 9067 2661 9111
rect 2609 9059 2618 9067
rect 2618 9059 2652 9067
rect 2652 9059 2661 9067
rect 2809 9173 2818 9181
rect 2818 9173 2852 9181
rect 2852 9173 2861 9181
rect 2809 9129 2861 9173
rect 3009 9347 3061 9391
rect 3009 9339 3018 9347
rect 3018 9339 3052 9347
rect 3052 9339 3061 9347
rect 3209 9453 3218 9461
rect 3218 9453 3252 9461
rect 3252 9453 3261 9461
rect 3209 9409 3261 9453
rect 3409 9627 3461 9671
rect 3409 9619 3418 9627
rect 3418 9619 3452 9627
rect 3452 9619 3461 9627
rect 3609 9733 3618 9741
rect 3618 9733 3652 9741
rect 3652 9733 3661 9741
rect 3609 9689 3661 9733
rect 3809 9890 3861 9899
rect 3809 9856 3818 9890
rect 3818 9856 3852 9890
rect 3852 9856 3861 9890
rect 3809 9847 3861 9856
rect 2209 8680 2261 8689
rect 2209 8646 2218 8680
rect 2218 8646 2252 8680
rect 2252 8646 2261 8680
rect 2209 8637 2261 8646
rect 609 7470 661 7479
rect 609 7436 618 7470
rect 618 7436 652 7470
rect 652 7436 661 7470
rect 609 7427 661 7436
rect 9 6893 18 6901
rect 18 6893 52 6901
rect 52 6893 61 6901
rect 9 6849 61 6893
rect 209 7067 261 7111
rect 209 7059 218 7067
rect 218 7059 252 7067
rect 252 7059 261 7067
rect 409 7173 418 7181
rect 418 7173 452 7181
rect 452 7173 461 7181
rect 409 7129 461 7173
rect 609 7347 661 7391
rect 609 7339 618 7347
rect 618 7339 652 7347
rect 652 7339 661 7347
rect 809 7543 818 7551
rect 818 7543 852 7551
rect 852 7543 861 7551
rect 809 7499 861 7543
rect 1009 7717 1061 7761
rect 1009 7709 1018 7717
rect 1018 7709 1052 7717
rect 1052 7709 1061 7717
rect 1209 7823 1218 7831
rect 1218 7823 1252 7831
rect 1252 7823 1261 7831
rect 1209 7779 1261 7823
rect 1409 7997 1461 8041
rect 1409 7989 1418 7997
rect 1418 7989 1452 7997
rect 1452 7989 1461 7997
rect 1609 8103 1618 8111
rect 1618 8103 1652 8111
rect 1652 8103 1661 8111
rect 1609 8059 1661 8103
rect 1809 8277 1861 8321
rect 1809 8269 1818 8277
rect 1818 8269 1852 8277
rect 1852 8269 1861 8277
rect 2009 8383 2018 8391
rect 2018 8383 2052 8391
rect 2052 8383 2061 8391
rect 2009 8339 2061 8383
rect 2209 8557 2261 8601
rect 2209 8549 2218 8557
rect 2218 8549 2252 8557
rect 2252 8549 2261 8557
rect 2409 8753 2418 8761
rect 2418 8753 2452 8761
rect 2452 8753 2461 8761
rect 2409 8709 2461 8753
rect 2609 8927 2661 8971
rect 2609 8919 2618 8927
rect 2618 8919 2652 8927
rect 2652 8919 2661 8927
rect 2809 9033 2818 9041
rect 2818 9033 2852 9041
rect 2852 9033 2861 9041
rect 2809 8989 2861 9033
rect 3009 9207 3061 9251
rect 3009 9199 3018 9207
rect 3018 9199 3052 9207
rect 3052 9199 3061 9207
rect 3209 9313 3218 9321
rect 3218 9313 3252 9321
rect 3252 9313 3261 9321
rect 3209 9269 3261 9313
rect 3409 9487 3461 9531
rect 3409 9479 3418 9487
rect 3418 9479 3452 9487
rect 3452 9479 3461 9487
rect 3609 9593 3618 9601
rect 3618 9593 3652 9601
rect 3652 9593 3661 9601
rect 3609 9549 3661 9593
rect 3809 9767 3861 9811
rect 3809 9759 3818 9767
rect 3818 9759 3852 9767
rect 3852 9759 3861 9767
rect 4009 9874 4061 9883
rect 4009 9840 4018 9874
rect 4018 9840 4052 9874
rect 4052 9840 4061 9874
rect 4009 9831 4061 9840
rect 2409 8664 2461 8673
rect 2409 8630 2418 8664
rect 2418 8630 2452 8664
rect 2452 8630 2461 8664
rect 2409 8621 2461 8630
rect 809 7454 861 7463
rect 809 7420 818 7454
rect 818 7420 852 7454
rect 852 7420 861 7454
rect 809 7411 861 7420
rect 9 6753 18 6761
rect 18 6753 52 6761
rect 52 6753 61 6761
rect 9 6709 61 6753
rect 209 6927 261 6971
rect 209 6919 218 6927
rect 218 6919 252 6927
rect 252 6919 261 6927
rect 409 7033 418 7041
rect 418 7033 452 7041
rect 452 7033 461 7041
rect 409 6989 461 7033
rect 609 7207 661 7251
rect 609 7199 618 7207
rect 618 7199 652 7207
rect 652 7199 661 7207
rect 809 7313 818 7321
rect 818 7313 852 7321
rect 852 7313 861 7321
rect 809 7269 861 7313
rect 1009 7577 1061 7621
rect 1009 7569 1018 7577
rect 1018 7569 1052 7577
rect 1052 7569 1061 7577
rect 1209 7683 1218 7691
rect 1218 7683 1252 7691
rect 1252 7683 1261 7691
rect 1209 7639 1261 7683
rect 1409 7857 1461 7901
rect 1409 7849 1418 7857
rect 1418 7849 1452 7857
rect 1452 7849 1461 7857
rect 1609 7963 1618 7971
rect 1618 7963 1652 7971
rect 1652 7963 1661 7971
rect 1609 7919 1661 7963
rect 1809 8137 1861 8181
rect 1809 8129 1818 8137
rect 1818 8129 1852 8137
rect 1852 8129 1861 8137
rect 2009 8243 2018 8251
rect 2018 8243 2052 8251
rect 2052 8243 2061 8251
rect 2009 8199 2061 8243
rect 2209 8417 2261 8461
rect 2209 8409 2218 8417
rect 2218 8409 2252 8417
rect 2252 8409 2261 8417
rect 2409 8523 2418 8531
rect 2418 8523 2452 8531
rect 2452 8523 2461 8531
rect 2409 8479 2461 8523
rect 2609 8787 2661 8831
rect 2609 8779 2618 8787
rect 2618 8779 2652 8787
rect 2652 8779 2661 8787
rect 2809 8893 2818 8901
rect 2818 8893 2852 8901
rect 2852 8893 2861 8901
rect 2809 8849 2861 8893
rect 3009 9067 3061 9111
rect 3009 9059 3018 9067
rect 3018 9059 3052 9067
rect 3052 9059 3061 9067
rect 3209 9173 3218 9181
rect 3218 9173 3252 9181
rect 3252 9173 3261 9181
rect 3209 9129 3261 9173
rect 3409 9347 3461 9391
rect 3409 9339 3418 9347
rect 3418 9339 3452 9347
rect 3452 9339 3461 9347
rect 3609 9453 3618 9461
rect 3618 9453 3652 9461
rect 3652 9453 3661 9461
rect 3609 9409 3661 9453
rect 3809 9627 3861 9671
rect 3809 9619 3818 9627
rect 3818 9619 3852 9627
rect 3852 9619 3861 9627
rect 4009 9733 4018 9741
rect 4018 9733 4052 9741
rect 4052 9733 4061 9741
rect 4009 9689 4061 9733
rect 4209 9890 4261 9899
rect 4209 9856 4218 9890
rect 4218 9856 4252 9890
rect 4252 9856 4261 9890
rect 4209 9847 4261 9856
rect 2609 8680 2661 8689
rect 2609 8646 2618 8680
rect 2618 8646 2652 8680
rect 2652 8646 2661 8680
rect 2609 8637 2661 8646
rect 1009 7470 1061 7479
rect 1009 7436 1018 7470
rect 1018 7436 1052 7470
rect 1052 7436 1061 7470
rect 1009 7427 1061 7436
rect 9 6613 18 6621
rect 18 6613 52 6621
rect 52 6613 61 6621
rect 9 6569 61 6613
rect 209 6787 261 6831
rect 209 6779 218 6787
rect 218 6779 252 6787
rect 252 6779 261 6787
rect 409 6893 418 6901
rect 418 6893 452 6901
rect 452 6893 461 6901
rect 409 6849 461 6893
rect 609 7067 661 7111
rect 609 7059 618 7067
rect 618 7059 652 7067
rect 652 7059 661 7067
rect 809 7173 818 7181
rect 818 7173 852 7181
rect 852 7173 861 7181
rect 809 7129 861 7173
rect 1009 7347 1061 7391
rect 1009 7339 1018 7347
rect 1018 7339 1052 7347
rect 1052 7339 1061 7347
rect 1209 7543 1218 7551
rect 1218 7543 1252 7551
rect 1252 7543 1261 7551
rect 1209 7499 1261 7543
rect 1409 7717 1461 7761
rect 1409 7709 1418 7717
rect 1418 7709 1452 7717
rect 1452 7709 1461 7717
rect 1609 7823 1618 7831
rect 1618 7823 1652 7831
rect 1652 7823 1661 7831
rect 1609 7779 1661 7823
rect 1809 7997 1861 8041
rect 1809 7989 1818 7997
rect 1818 7989 1852 7997
rect 1852 7989 1861 7997
rect 2009 8103 2018 8111
rect 2018 8103 2052 8111
rect 2052 8103 2061 8111
rect 2009 8059 2061 8103
rect 2209 8277 2261 8321
rect 2209 8269 2218 8277
rect 2218 8269 2252 8277
rect 2252 8269 2261 8277
rect 2409 8383 2418 8391
rect 2418 8383 2452 8391
rect 2452 8383 2461 8391
rect 2409 8339 2461 8383
rect 2609 8557 2661 8601
rect 2609 8549 2618 8557
rect 2618 8549 2652 8557
rect 2652 8549 2661 8557
rect 2809 8753 2818 8761
rect 2818 8753 2852 8761
rect 2852 8753 2861 8761
rect 2809 8709 2861 8753
rect 3009 8927 3061 8971
rect 3009 8919 3018 8927
rect 3018 8919 3052 8927
rect 3052 8919 3061 8927
rect 3209 9033 3218 9041
rect 3218 9033 3252 9041
rect 3252 9033 3261 9041
rect 3209 8989 3261 9033
rect 3409 9207 3461 9251
rect 3409 9199 3418 9207
rect 3418 9199 3452 9207
rect 3452 9199 3461 9207
rect 3609 9313 3618 9321
rect 3618 9313 3652 9321
rect 3652 9313 3661 9321
rect 3609 9269 3661 9313
rect 3809 9487 3861 9531
rect 3809 9479 3818 9487
rect 3818 9479 3852 9487
rect 3852 9479 3861 9487
rect 4009 9593 4018 9601
rect 4018 9593 4052 9601
rect 4052 9593 4061 9601
rect 4009 9549 4061 9593
rect 4209 9767 4261 9811
rect 4209 9759 4218 9767
rect 4218 9759 4252 9767
rect 4252 9759 4261 9767
rect 4409 9874 4461 9883
rect 4409 9840 4418 9874
rect 4418 9840 4452 9874
rect 4452 9840 4461 9874
rect 4409 9831 4461 9840
rect 2809 8664 2861 8673
rect 2809 8630 2818 8664
rect 2818 8630 2852 8664
rect 2852 8630 2861 8664
rect 2809 8621 2861 8630
rect 1209 7454 1261 7463
rect 1209 7420 1218 7454
rect 1218 7420 1252 7454
rect 1252 7420 1261 7454
rect 1209 7411 1261 7420
rect 9 6473 18 6481
rect 18 6473 52 6481
rect 52 6473 61 6481
rect 9 6429 61 6473
rect 209 6647 261 6691
rect 209 6639 218 6647
rect 218 6639 252 6647
rect 252 6639 261 6647
rect 409 6753 418 6761
rect 418 6753 452 6761
rect 452 6753 461 6761
rect 409 6709 461 6753
rect 609 6927 661 6971
rect 609 6919 618 6927
rect 618 6919 652 6927
rect 652 6919 661 6927
rect 809 7033 818 7041
rect 818 7033 852 7041
rect 852 7033 861 7041
rect 809 6989 861 7033
rect 1009 7207 1061 7251
rect 1009 7199 1018 7207
rect 1018 7199 1052 7207
rect 1052 7199 1061 7207
rect 1209 7313 1218 7321
rect 1218 7313 1252 7321
rect 1252 7313 1261 7321
rect 1209 7269 1261 7313
rect 1409 7577 1461 7621
rect 1409 7569 1418 7577
rect 1418 7569 1452 7577
rect 1452 7569 1461 7577
rect 1609 7683 1618 7691
rect 1618 7683 1652 7691
rect 1652 7683 1661 7691
rect 1609 7639 1661 7683
rect 1809 7857 1861 7901
rect 1809 7849 1818 7857
rect 1818 7849 1852 7857
rect 1852 7849 1861 7857
rect 2009 7963 2018 7971
rect 2018 7963 2052 7971
rect 2052 7963 2061 7971
rect 2009 7919 2061 7963
rect 2209 8137 2261 8181
rect 2209 8129 2218 8137
rect 2218 8129 2252 8137
rect 2252 8129 2261 8137
rect 2409 8243 2418 8251
rect 2418 8243 2452 8251
rect 2452 8243 2461 8251
rect 2409 8199 2461 8243
rect 2609 8417 2661 8461
rect 2609 8409 2618 8417
rect 2618 8409 2652 8417
rect 2652 8409 2661 8417
rect 2809 8523 2818 8531
rect 2818 8523 2852 8531
rect 2852 8523 2861 8531
rect 2809 8479 2861 8523
rect 3009 8787 3061 8831
rect 3009 8779 3018 8787
rect 3018 8779 3052 8787
rect 3052 8779 3061 8787
rect 3209 8893 3218 8901
rect 3218 8893 3252 8901
rect 3252 8893 3261 8901
rect 3209 8849 3261 8893
rect 3409 9067 3461 9111
rect 3409 9059 3418 9067
rect 3418 9059 3452 9067
rect 3452 9059 3461 9067
rect 3609 9173 3618 9181
rect 3618 9173 3652 9181
rect 3652 9173 3661 9181
rect 3609 9129 3661 9173
rect 3809 9347 3861 9391
rect 3809 9339 3818 9347
rect 3818 9339 3852 9347
rect 3852 9339 3861 9347
rect 4009 9453 4018 9461
rect 4018 9453 4052 9461
rect 4052 9453 4061 9461
rect 4009 9409 4061 9453
rect 4209 9627 4261 9671
rect 4209 9619 4218 9627
rect 4218 9619 4252 9627
rect 4252 9619 4261 9627
rect 4409 9733 4418 9741
rect 4418 9733 4452 9741
rect 4452 9733 4461 9741
rect 4409 9689 4461 9733
rect 4609 9890 4661 9899
rect 4609 9856 4618 9890
rect 4618 9856 4652 9890
rect 4652 9856 4661 9890
rect 4609 9847 4661 9856
rect 3009 8680 3061 8689
rect 3009 8646 3018 8680
rect 3018 8646 3052 8680
rect 3052 8646 3061 8680
rect 3009 8637 3061 8646
rect 1409 7470 1461 7479
rect 1409 7436 1418 7470
rect 1418 7436 1452 7470
rect 1452 7436 1461 7470
rect 1409 7427 1461 7436
rect 9 6333 18 6341
rect 18 6333 52 6341
rect 52 6333 61 6341
rect 9 6289 61 6333
rect 209 6507 261 6551
rect 209 6499 218 6507
rect 218 6499 252 6507
rect 252 6499 261 6507
rect 409 6613 418 6621
rect 418 6613 452 6621
rect 452 6613 461 6621
rect 409 6569 461 6613
rect 609 6787 661 6831
rect 609 6779 618 6787
rect 618 6779 652 6787
rect 652 6779 661 6787
rect 809 6893 818 6901
rect 818 6893 852 6901
rect 852 6893 861 6901
rect 809 6849 861 6893
rect 1009 7067 1061 7111
rect 1009 7059 1018 7067
rect 1018 7059 1052 7067
rect 1052 7059 1061 7067
rect 1209 7173 1218 7181
rect 1218 7173 1252 7181
rect 1252 7173 1261 7181
rect 1209 7129 1261 7173
rect 1409 7347 1461 7391
rect 1409 7339 1418 7347
rect 1418 7339 1452 7347
rect 1452 7339 1461 7347
rect 1609 7543 1618 7551
rect 1618 7543 1652 7551
rect 1652 7543 1661 7551
rect 1609 7499 1661 7543
rect 1809 7717 1861 7761
rect 1809 7709 1818 7717
rect 1818 7709 1852 7717
rect 1852 7709 1861 7717
rect 2009 7823 2018 7831
rect 2018 7823 2052 7831
rect 2052 7823 2061 7831
rect 2009 7779 2061 7823
rect 2209 7997 2261 8041
rect 2209 7989 2218 7997
rect 2218 7989 2252 7997
rect 2252 7989 2261 7997
rect 2409 8103 2418 8111
rect 2418 8103 2452 8111
rect 2452 8103 2461 8111
rect 2409 8059 2461 8103
rect 2609 8277 2661 8321
rect 2609 8269 2618 8277
rect 2618 8269 2652 8277
rect 2652 8269 2661 8277
rect 2809 8383 2818 8391
rect 2818 8383 2852 8391
rect 2852 8383 2861 8391
rect 2809 8339 2861 8383
rect 3009 8557 3061 8601
rect 3009 8549 3018 8557
rect 3018 8549 3052 8557
rect 3052 8549 3061 8557
rect 3209 8753 3218 8761
rect 3218 8753 3252 8761
rect 3252 8753 3261 8761
rect 3209 8709 3261 8753
rect 3409 8927 3461 8971
rect 3409 8919 3418 8927
rect 3418 8919 3452 8927
rect 3452 8919 3461 8927
rect 3609 9033 3618 9041
rect 3618 9033 3652 9041
rect 3652 9033 3661 9041
rect 3609 8989 3661 9033
rect 3809 9207 3861 9251
rect 3809 9199 3818 9207
rect 3818 9199 3852 9207
rect 3852 9199 3861 9207
rect 4009 9313 4018 9321
rect 4018 9313 4052 9321
rect 4052 9313 4061 9321
rect 4009 9269 4061 9313
rect 4209 9487 4261 9531
rect 4209 9479 4218 9487
rect 4218 9479 4252 9487
rect 4252 9479 4261 9487
rect 4409 9593 4418 9601
rect 4418 9593 4452 9601
rect 4452 9593 4461 9601
rect 4409 9549 4461 9593
rect 4609 9767 4661 9811
rect 4609 9759 4618 9767
rect 4618 9759 4652 9767
rect 4652 9759 4661 9767
rect 4809 9874 4861 9883
rect 4809 9840 4818 9874
rect 4818 9840 4852 9874
rect 4852 9840 4861 9874
rect 4809 9831 4861 9840
rect 3209 8664 3261 8673
rect 3209 8630 3218 8664
rect 3218 8630 3252 8664
rect 3252 8630 3261 8664
rect 3209 8621 3261 8630
rect 1609 7454 1661 7463
rect 1609 7420 1618 7454
rect 1618 7420 1652 7454
rect 1652 7420 1661 7454
rect 1609 7411 1661 7420
rect 9 6244 61 6253
rect 9 6210 18 6244
rect 18 6210 52 6244
rect 52 6210 61 6244
rect 9 6201 61 6210
rect 9 6103 18 6111
rect 18 6103 52 6111
rect 52 6103 61 6111
rect 9 6059 61 6103
rect 209 6367 261 6411
rect 209 6359 218 6367
rect 218 6359 252 6367
rect 252 6359 261 6367
rect 409 6473 418 6481
rect 418 6473 452 6481
rect 452 6473 461 6481
rect 409 6429 461 6473
rect 609 6647 661 6691
rect 609 6639 618 6647
rect 618 6639 652 6647
rect 652 6639 661 6647
rect 809 6753 818 6761
rect 818 6753 852 6761
rect 852 6753 861 6761
rect 809 6709 861 6753
rect 1009 6927 1061 6971
rect 1009 6919 1018 6927
rect 1018 6919 1052 6927
rect 1052 6919 1061 6927
rect 1209 7033 1218 7041
rect 1218 7033 1252 7041
rect 1252 7033 1261 7041
rect 1209 6989 1261 7033
rect 1409 7207 1461 7251
rect 1409 7199 1418 7207
rect 1418 7199 1452 7207
rect 1452 7199 1461 7207
rect 1609 7313 1618 7321
rect 1618 7313 1652 7321
rect 1652 7313 1661 7321
rect 1609 7269 1661 7313
rect 1809 7577 1861 7621
rect 1809 7569 1818 7577
rect 1818 7569 1852 7577
rect 1852 7569 1861 7577
rect 2009 7683 2018 7691
rect 2018 7683 2052 7691
rect 2052 7683 2061 7691
rect 2009 7639 2061 7683
rect 2209 7857 2261 7901
rect 2209 7849 2218 7857
rect 2218 7849 2252 7857
rect 2252 7849 2261 7857
rect 2409 7963 2418 7971
rect 2418 7963 2452 7971
rect 2452 7963 2461 7971
rect 2409 7919 2461 7963
rect 2609 8137 2661 8181
rect 2609 8129 2618 8137
rect 2618 8129 2652 8137
rect 2652 8129 2661 8137
rect 2809 8243 2818 8251
rect 2818 8243 2852 8251
rect 2852 8243 2861 8251
rect 2809 8199 2861 8243
rect 3009 8417 3061 8461
rect 3009 8409 3018 8417
rect 3018 8409 3052 8417
rect 3052 8409 3061 8417
rect 3209 8523 3218 8531
rect 3218 8523 3252 8531
rect 3252 8523 3261 8531
rect 3209 8479 3261 8523
rect 3409 8787 3461 8831
rect 3409 8779 3418 8787
rect 3418 8779 3452 8787
rect 3452 8779 3461 8787
rect 3609 8893 3618 8901
rect 3618 8893 3652 8901
rect 3652 8893 3661 8901
rect 3609 8849 3661 8893
rect 3809 9067 3861 9111
rect 3809 9059 3818 9067
rect 3818 9059 3852 9067
rect 3852 9059 3861 9067
rect 4009 9173 4018 9181
rect 4018 9173 4052 9181
rect 4052 9173 4061 9181
rect 4009 9129 4061 9173
rect 4209 9347 4261 9391
rect 4209 9339 4218 9347
rect 4218 9339 4252 9347
rect 4252 9339 4261 9347
rect 4409 9453 4418 9461
rect 4418 9453 4452 9461
rect 4452 9453 4461 9461
rect 4409 9409 4461 9453
rect 4609 9627 4661 9671
rect 4609 9619 4618 9627
rect 4618 9619 4652 9627
rect 4652 9619 4661 9627
rect 4809 9733 4818 9741
rect 4818 9733 4852 9741
rect 4852 9733 4861 9741
rect 4809 9689 4861 9733
rect 5009 9890 5061 9899
rect 5009 9856 5018 9890
rect 5018 9856 5052 9890
rect 5052 9856 5061 9890
rect 5009 9847 5061 9856
rect 3409 8680 3461 8689
rect 3409 8646 3418 8680
rect 3418 8646 3452 8680
rect 3452 8646 3461 8680
rect 3409 8637 3461 8646
rect 1809 7470 1861 7479
rect 1809 7436 1818 7470
rect 1818 7436 1852 7470
rect 1852 7436 1861 7470
rect 1809 7427 1861 7436
rect 209 6260 261 6269
rect 209 6226 218 6260
rect 218 6226 252 6260
rect 252 6226 261 6260
rect 209 6217 261 6226
rect 9 5963 18 5971
rect 18 5963 52 5971
rect 52 5963 61 5971
rect 9 5919 61 5963
rect 209 6137 261 6181
rect 209 6129 218 6137
rect 218 6129 252 6137
rect 252 6129 261 6137
rect 409 6333 418 6341
rect 418 6333 452 6341
rect 452 6333 461 6341
rect 409 6289 461 6333
rect 609 6507 661 6551
rect 609 6499 618 6507
rect 618 6499 652 6507
rect 652 6499 661 6507
rect 809 6613 818 6621
rect 818 6613 852 6621
rect 852 6613 861 6621
rect 809 6569 861 6613
rect 1009 6787 1061 6831
rect 1009 6779 1018 6787
rect 1018 6779 1052 6787
rect 1052 6779 1061 6787
rect 1209 6893 1218 6901
rect 1218 6893 1252 6901
rect 1252 6893 1261 6901
rect 1209 6849 1261 6893
rect 1409 7067 1461 7111
rect 1409 7059 1418 7067
rect 1418 7059 1452 7067
rect 1452 7059 1461 7067
rect 1609 7173 1618 7181
rect 1618 7173 1652 7181
rect 1652 7173 1661 7181
rect 1609 7129 1661 7173
rect 1809 7347 1861 7391
rect 1809 7339 1818 7347
rect 1818 7339 1852 7347
rect 1852 7339 1861 7347
rect 2009 7543 2018 7551
rect 2018 7543 2052 7551
rect 2052 7543 2061 7551
rect 2009 7499 2061 7543
rect 2209 7717 2261 7761
rect 2209 7709 2218 7717
rect 2218 7709 2252 7717
rect 2252 7709 2261 7717
rect 2409 7823 2418 7831
rect 2418 7823 2452 7831
rect 2452 7823 2461 7831
rect 2409 7779 2461 7823
rect 2609 7997 2661 8041
rect 2609 7989 2618 7997
rect 2618 7989 2652 7997
rect 2652 7989 2661 7997
rect 2809 8103 2818 8111
rect 2818 8103 2852 8111
rect 2852 8103 2861 8111
rect 2809 8059 2861 8103
rect 3009 8277 3061 8321
rect 3009 8269 3018 8277
rect 3018 8269 3052 8277
rect 3052 8269 3061 8277
rect 3209 8383 3218 8391
rect 3218 8383 3252 8391
rect 3252 8383 3261 8391
rect 3209 8339 3261 8383
rect 3409 8557 3461 8601
rect 3409 8549 3418 8557
rect 3418 8549 3452 8557
rect 3452 8549 3461 8557
rect 3609 8753 3618 8761
rect 3618 8753 3652 8761
rect 3652 8753 3661 8761
rect 3609 8709 3661 8753
rect 3809 8927 3861 8971
rect 3809 8919 3818 8927
rect 3818 8919 3852 8927
rect 3852 8919 3861 8927
rect 4009 9033 4018 9041
rect 4018 9033 4052 9041
rect 4052 9033 4061 9041
rect 4009 8989 4061 9033
rect 4209 9207 4261 9251
rect 4209 9199 4218 9207
rect 4218 9199 4252 9207
rect 4252 9199 4261 9207
rect 4409 9313 4418 9321
rect 4418 9313 4452 9321
rect 4452 9313 4461 9321
rect 4409 9269 4461 9313
rect 4609 9487 4661 9531
rect 4609 9479 4618 9487
rect 4618 9479 4652 9487
rect 4652 9479 4661 9487
rect 4809 9593 4818 9601
rect 4818 9593 4852 9601
rect 4852 9593 4861 9601
rect 4809 9549 4861 9593
rect 5009 9767 5061 9811
rect 5009 9759 5018 9767
rect 5018 9759 5052 9767
rect 5052 9759 5061 9767
rect 5209 9874 5261 9883
rect 5209 9840 5218 9874
rect 5218 9840 5252 9874
rect 5252 9840 5261 9874
rect 5209 9831 5261 9840
rect 3609 8664 3661 8673
rect 3609 8630 3618 8664
rect 3618 8630 3652 8664
rect 3652 8630 3661 8664
rect 3609 8621 3661 8630
rect 2009 7454 2061 7463
rect 2009 7420 2018 7454
rect 2018 7420 2052 7454
rect 2052 7420 2061 7454
rect 2009 7411 2061 7420
rect 409 6244 461 6253
rect 409 6210 418 6244
rect 418 6210 452 6244
rect 452 6210 461 6244
rect 409 6201 461 6210
rect 9 5823 18 5831
rect 18 5823 52 5831
rect 52 5823 61 5831
rect 9 5779 61 5823
rect 209 5997 261 6041
rect 209 5989 218 5997
rect 218 5989 252 5997
rect 252 5989 261 5997
rect 409 6103 418 6111
rect 418 6103 452 6111
rect 452 6103 461 6111
rect 409 6059 461 6103
rect 609 6367 661 6411
rect 609 6359 618 6367
rect 618 6359 652 6367
rect 652 6359 661 6367
rect 809 6473 818 6481
rect 818 6473 852 6481
rect 852 6473 861 6481
rect 809 6429 861 6473
rect 1009 6647 1061 6691
rect 1009 6639 1018 6647
rect 1018 6639 1052 6647
rect 1052 6639 1061 6647
rect 1209 6753 1218 6761
rect 1218 6753 1252 6761
rect 1252 6753 1261 6761
rect 1209 6709 1261 6753
rect 1409 6927 1461 6971
rect 1409 6919 1418 6927
rect 1418 6919 1452 6927
rect 1452 6919 1461 6927
rect 1609 7033 1618 7041
rect 1618 7033 1652 7041
rect 1652 7033 1661 7041
rect 1609 6989 1661 7033
rect 1809 7207 1861 7251
rect 1809 7199 1818 7207
rect 1818 7199 1852 7207
rect 1852 7199 1861 7207
rect 2009 7313 2018 7321
rect 2018 7313 2052 7321
rect 2052 7313 2061 7321
rect 2009 7269 2061 7313
rect 2209 7577 2261 7621
rect 2209 7569 2218 7577
rect 2218 7569 2252 7577
rect 2252 7569 2261 7577
rect 2409 7683 2418 7691
rect 2418 7683 2452 7691
rect 2452 7683 2461 7691
rect 2409 7639 2461 7683
rect 2609 7857 2661 7901
rect 2609 7849 2618 7857
rect 2618 7849 2652 7857
rect 2652 7849 2661 7857
rect 2809 7963 2818 7971
rect 2818 7963 2852 7971
rect 2852 7963 2861 7971
rect 2809 7919 2861 7963
rect 3009 8137 3061 8181
rect 3009 8129 3018 8137
rect 3018 8129 3052 8137
rect 3052 8129 3061 8137
rect 3209 8243 3218 8251
rect 3218 8243 3252 8251
rect 3252 8243 3261 8251
rect 3209 8199 3261 8243
rect 3409 8417 3461 8461
rect 3409 8409 3418 8417
rect 3418 8409 3452 8417
rect 3452 8409 3461 8417
rect 3609 8523 3618 8531
rect 3618 8523 3652 8531
rect 3652 8523 3661 8531
rect 3609 8479 3661 8523
rect 3809 8787 3861 8831
rect 3809 8779 3818 8787
rect 3818 8779 3852 8787
rect 3852 8779 3861 8787
rect 4009 8893 4018 8901
rect 4018 8893 4052 8901
rect 4052 8893 4061 8901
rect 4009 8849 4061 8893
rect 4209 9067 4261 9111
rect 4209 9059 4218 9067
rect 4218 9059 4252 9067
rect 4252 9059 4261 9067
rect 4409 9173 4418 9181
rect 4418 9173 4452 9181
rect 4452 9173 4461 9181
rect 4409 9129 4461 9173
rect 4609 9347 4661 9391
rect 4609 9339 4618 9347
rect 4618 9339 4652 9347
rect 4652 9339 4661 9347
rect 4809 9453 4818 9461
rect 4818 9453 4852 9461
rect 4852 9453 4861 9461
rect 4809 9409 4861 9453
rect 5009 9627 5061 9671
rect 5009 9619 5018 9627
rect 5018 9619 5052 9627
rect 5052 9619 5061 9627
rect 5209 9733 5218 9741
rect 5218 9733 5252 9741
rect 5252 9733 5261 9741
rect 5209 9689 5261 9733
rect 5409 9890 5461 9899
rect 5409 9856 5418 9890
rect 5418 9856 5452 9890
rect 5452 9856 5461 9890
rect 5409 9847 5461 9856
rect 3809 8680 3861 8689
rect 3809 8646 3818 8680
rect 3818 8646 3852 8680
rect 3852 8646 3861 8680
rect 3809 8637 3861 8646
rect 2209 7470 2261 7479
rect 2209 7436 2218 7470
rect 2218 7436 2252 7470
rect 2252 7436 2261 7470
rect 2209 7427 2261 7436
rect 609 6260 661 6269
rect 609 6226 618 6260
rect 618 6226 652 6260
rect 652 6226 661 6260
rect 609 6217 661 6226
rect 9 5683 18 5691
rect 18 5683 52 5691
rect 52 5683 61 5691
rect 9 5639 61 5683
rect 209 5857 261 5901
rect 209 5849 218 5857
rect 218 5849 252 5857
rect 252 5849 261 5857
rect 409 5963 418 5971
rect 418 5963 452 5971
rect 452 5963 461 5971
rect 409 5919 461 5963
rect 609 6137 661 6181
rect 609 6129 618 6137
rect 618 6129 652 6137
rect 652 6129 661 6137
rect 809 6333 818 6341
rect 818 6333 852 6341
rect 852 6333 861 6341
rect 809 6289 861 6333
rect 1009 6507 1061 6551
rect 1009 6499 1018 6507
rect 1018 6499 1052 6507
rect 1052 6499 1061 6507
rect 1209 6613 1218 6621
rect 1218 6613 1252 6621
rect 1252 6613 1261 6621
rect 1209 6569 1261 6613
rect 1409 6787 1461 6831
rect 1409 6779 1418 6787
rect 1418 6779 1452 6787
rect 1452 6779 1461 6787
rect 1609 6893 1618 6901
rect 1618 6893 1652 6901
rect 1652 6893 1661 6901
rect 1609 6849 1661 6893
rect 1809 7067 1861 7111
rect 1809 7059 1818 7067
rect 1818 7059 1852 7067
rect 1852 7059 1861 7067
rect 2009 7173 2018 7181
rect 2018 7173 2052 7181
rect 2052 7173 2061 7181
rect 2009 7129 2061 7173
rect 2209 7347 2261 7391
rect 2209 7339 2218 7347
rect 2218 7339 2252 7347
rect 2252 7339 2261 7347
rect 2409 7543 2418 7551
rect 2418 7543 2452 7551
rect 2452 7543 2461 7551
rect 2409 7499 2461 7543
rect 2609 7717 2661 7761
rect 2609 7709 2618 7717
rect 2618 7709 2652 7717
rect 2652 7709 2661 7717
rect 2809 7823 2818 7831
rect 2818 7823 2852 7831
rect 2852 7823 2861 7831
rect 2809 7779 2861 7823
rect 3009 7997 3061 8041
rect 3009 7989 3018 7997
rect 3018 7989 3052 7997
rect 3052 7989 3061 7997
rect 3209 8103 3218 8111
rect 3218 8103 3252 8111
rect 3252 8103 3261 8111
rect 3209 8059 3261 8103
rect 3409 8277 3461 8321
rect 3409 8269 3418 8277
rect 3418 8269 3452 8277
rect 3452 8269 3461 8277
rect 3609 8383 3618 8391
rect 3618 8383 3652 8391
rect 3652 8383 3661 8391
rect 3609 8339 3661 8383
rect 3809 8557 3861 8601
rect 3809 8549 3818 8557
rect 3818 8549 3852 8557
rect 3852 8549 3861 8557
rect 4009 8753 4018 8761
rect 4018 8753 4052 8761
rect 4052 8753 4061 8761
rect 4009 8709 4061 8753
rect 4209 8927 4261 8971
rect 4209 8919 4218 8927
rect 4218 8919 4252 8927
rect 4252 8919 4261 8927
rect 4409 9033 4418 9041
rect 4418 9033 4452 9041
rect 4452 9033 4461 9041
rect 4409 8989 4461 9033
rect 4609 9207 4661 9251
rect 4609 9199 4618 9207
rect 4618 9199 4652 9207
rect 4652 9199 4661 9207
rect 4809 9313 4818 9321
rect 4818 9313 4852 9321
rect 4852 9313 4861 9321
rect 4809 9269 4861 9313
rect 5009 9487 5061 9531
rect 5009 9479 5018 9487
rect 5018 9479 5052 9487
rect 5052 9479 5061 9487
rect 5209 9593 5218 9601
rect 5218 9593 5252 9601
rect 5252 9593 5261 9601
rect 5209 9549 5261 9593
rect 5409 9767 5461 9811
rect 5409 9759 5418 9767
rect 5418 9759 5452 9767
rect 5452 9759 5461 9767
rect 5609 9874 5661 9883
rect 5609 9840 5618 9874
rect 5618 9840 5652 9874
rect 5652 9840 5661 9874
rect 5609 9831 5661 9840
rect 4009 8664 4061 8673
rect 4009 8630 4018 8664
rect 4018 8630 4052 8664
rect 4052 8630 4061 8664
rect 4009 8621 4061 8630
rect 2409 7454 2461 7463
rect 2409 7420 2418 7454
rect 2418 7420 2452 7454
rect 2452 7420 2461 7454
rect 2409 7411 2461 7420
rect 809 6244 861 6253
rect 809 6210 818 6244
rect 818 6210 852 6244
rect 852 6210 861 6244
rect 809 6201 861 6210
rect 9 5543 18 5551
rect 18 5543 52 5551
rect 52 5543 61 5551
rect 9 5499 61 5543
rect 209 5717 261 5761
rect 209 5709 218 5717
rect 218 5709 252 5717
rect 252 5709 261 5717
rect 409 5823 418 5831
rect 418 5823 452 5831
rect 452 5823 461 5831
rect 409 5779 461 5823
rect 609 5997 661 6041
rect 609 5989 618 5997
rect 618 5989 652 5997
rect 652 5989 661 5997
rect 809 6103 818 6111
rect 818 6103 852 6111
rect 852 6103 861 6111
rect 809 6059 861 6103
rect 1009 6367 1061 6411
rect 1009 6359 1018 6367
rect 1018 6359 1052 6367
rect 1052 6359 1061 6367
rect 1209 6473 1218 6481
rect 1218 6473 1252 6481
rect 1252 6473 1261 6481
rect 1209 6429 1261 6473
rect 1409 6647 1461 6691
rect 1409 6639 1418 6647
rect 1418 6639 1452 6647
rect 1452 6639 1461 6647
rect 1609 6753 1618 6761
rect 1618 6753 1652 6761
rect 1652 6753 1661 6761
rect 1609 6709 1661 6753
rect 1809 6927 1861 6971
rect 1809 6919 1818 6927
rect 1818 6919 1852 6927
rect 1852 6919 1861 6927
rect 2009 7033 2018 7041
rect 2018 7033 2052 7041
rect 2052 7033 2061 7041
rect 2009 6989 2061 7033
rect 2209 7207 2261 7251
rect 2209 7199 2218 7207
rect 2218 7199 2252 7207
rect 2252 7199 2261 7207
rect 2409 7313 2418 7321
rect 2418 7313 2452 7321
rect 2452 7313 2461 7321
rect 2409 7269 2461 7313
rect 2609 7577 2661 7621
rect 2609 7569 2618 7577
rect 2618 7569 2652 7577
rect 2652 7569 2661 7577
rect 2809 7683 2818 7691
rect 2818 7683 2852 7691
rect 2852 7683 2861 7691
rect 2809 7639 2861 7683
rect 3009 7857 3061 7901
rect 3009 7849 3018 7857
rect 3018 7849 3052 7857
rect 3052 7849 3061 7857
rect 3209 7963 3218 7971
rect 3218 7963 3252 7971
rect 3252 7963 3261 7971
rect 3209 7919 3261 7963
rect 3409 8137 3461 8181
rect 3409 8129 3418 8137
rect 3418 8129 3452 8137
rect 3452 8129 3461 8137
rect 3609 8243 3618 8251
rect 3618 8243 3652 8251
rect 3652 8243 3661 8251
rect 3609 8199 3661 8243
rect 3809 8417 3861 8461
rect 3809 8409 3818 8417
rect 3818 8409 3852 8417
rect 3852 8409 3861 8417
rect 4009 8523 4018 8531
rect 4018 8523 4052 8531
rect 4052 8523 4061 8531
rect 4009 8479 4061 8523
rect 4209 8787 4261 8831
rect 4209 8779 4218 8787
rect 4218 8779 4252 8787
rect 4252 8779 4261 8787
rect 4409 8893 4418 8901
rect 4418 8893 4452 8901
rect 4452 8893 4461 8901
rect 4409 8849 4461 8893
rect 4609 9067 4661 9111
rect 4609 9059 4618 9067
rect 4618 9059 4652 9067
rect 4652 9059 4661 9067
rect 4809 9173 4818 9181
rect 4818 9173 4852 9181
rect 4852 9173 4861 9181
rect 4809 9129 4861 9173
rect 5009 9347 5061 9391
rect 5009 9339 5018 9347
rect 5018 9339 5052 9347
rect 5052 9339 5061 9347
rect 5209 9453 5218 9461
rect 5218 9453 5252 9461
rect 5252 9453 5261 9461
rect 5209 9409 5261 9453
rect 5409 9627 5461 9671
rect 5409 9619 5418 9627
rect 5418 9619 5452 9627
rect 5452 9619 5461 9627
rect 5609 9733 5618 9741
rect 5618 9733 5652 9741
rect 5652 9733 5661 9741
rect 5609 9689 5661 9733
rect 5809 9890 5861 9899
rect 5809 9856 5818 9890
rect 5818 9856 5852 9890
rect 5852 9856 5861 9890
rect 5809 9847 5861 9856
rect 4209 8680 4261 8689
rect 4209 8646 4218 8680
rect 4218 8646 4252 8680
rect 4252 8646 4261 8680
rect 4209 8637 4261 8646
rect 2609 7470 2661 7479
rect 2609 7436 2618 7470
rect 2618 7436 2652 7470
rect 2652 7436 2661 7470
rect 2609 7427 2661 7436
rect 1009 6260 1061 6269
rect 1009 6226 1018 6260
rect 1018 6226 1052 6260
rect 1052 6226 1061 6260
rect 1009 6217 1061 6226
rect 9 5403 18 5411
rect 18 5403 52 5411
rect 52 5403 61 5411
rect 9 5359 61 5403
rect 209 5577 261 5621
rect 209 5569 218 5577
rect 218 5569 252 5577
rect 252 5569 261 5577
rect 409 5683 418 5691
rect 418 5683 452 5691
rect 452 5683 461 5691
rect 409 5639 461 5683
rect 609 5857 661 5901
rect 609 5849 618 5857
rect 618 5849 652 5857
rect 652 5849 661 5857
rect 809 5963 818 5971
rect 818 5963 852 5971
rect 852 5963 861 5971
rect 809 5919 861 5963
rect 1009 6137 1061 6181
rect 1009 6129 1018 6137
rect 1018 6129 1052 6137
rect 1052 6129 1061 6137
rect 1209 6333 1218 6341
rect 1218 6333 1252 6341
rect 1252 6333 1261 6341
rect 1209 6289 1261 6333
rect 1409 6507 1461 6551
rect 1409 6499 1418 6507
rect 1418 6499 1452 6507
rect 1452 6499 1461 6507
rect 1609 6613 1618 6621
rect 1618 6613 1652 6621
rect 1652 6613 1661 6621
rect 1609 6569 1661 6613
rect 1809 6787 1861 6831
rect 1809 6779 1818 6787
rect 1818 6779 1852 6787
rect 1852 6779 1861 6787
rect 2009 6893 2018 6901
rect 2018 6893 2052 6901
rect 2052 6893 2061 6901
rect 2009 6849 2061 6893
rect 2209 7067 2261 7111
rect 2209 7059 2218 7067
rect 2218 7059 2252 7067
rect 2252 7059 2261 7067
rect 2409 7173 2418 7181
rect 2418 7173 2452 7181
rect 2452 7173 2461 7181
rect 2409 7129 2461 7173
rect 2609 7347 2661 7391
rect 2609 7339 2618 7347
rect 2618 7339 2652 7347
rect 2652 7339 2661 7347
rect 2809 7543 2818 7551
rect 2818 7543 2852 7551
rect 2852 7543 2861 7551
rect 2809 7499 2861 7543
rect 3009 7717 3061 7761
rect 3009 7709 3018 7717
rect 3018 7709 3052 7717
rect 3052 7709 3061 7717
rect 3209 7823 3218 7831
rect 3218 7823 3252 7831
rect 3252 7823 3261 7831
rect 3209 7779 3261 7823
rect 3409 7997 3461 8041
rect 3409 7989 3418 7997
rect 3418 7989 3452 7997
rect 3452 7989 3461 7997
rect 3609 8103 3618 8111
rect 3618 8103 3652 8111
rect 3652 8103 3661 8111
rect 3609 8059 3661 8103
rect 3809 8277 3861 8321
rect 3809 8269 3818 8277
rect 3818 8269 3852 8277
rect 3852 8269 3861 8277
rect 4009 8383 4018 8391
rect 4018 8383 4052 8391
rect 4052 8383 4061 8391
rect 4009 8339 4061 8383
rect 4209 8557 4261 8601
rect 4209 8549 4218 8557
rect 4218 8549 4252 8557
rect 4252 8549 4261 8557
rect 4409 8753 4418 8761
rect 4418 8753 4452 8761
rect 4452 8753 4461 8761
rect 4409 8709 4461 8753
rect 4609 8927 4661 8971
rect 4609 8919 4618 8927
rect 4618 8919 4652 8927
rect 4652 8919 4661 8927
rect 4809 9033 4818 9041
rect 4818 9033 4852 9041
rect 4852 9033 4861 9041
rect 4809 8989 4861 9033
rect 5009 9207 5061 9251
rect 5009 9199 5018 9207
rect 5018 9199 5052 9207
rect 5052 9199 5061 9207
rect 5209 9313 5218 9321
rect 5218 9313 5252 9321
rect 5252 9313 5261 9321
rect 5209 9269 5261 9313
rect 5409 9487 5461 9531
rect 5409 9479 5418 9487
rect 5418 9479 5452 9487
rect 5452 9479 5461 9487
rect 5609 9593 5618 9601
rect 5618 9593 5652 9601
rect 5652 9593 5661 9601
rect 5609 9549 5661 9593
rect 5809 9767 5861 9811
rect 5809 9759 5818 9767
rect 5818 9759 5852 9767
rect 5852 9759 5861 9767
rect 6009 9874 6061 9883
rect 6009 9840 6018 9874
rect 6018 9840 6052 9874
rect 6052 9840 6061 9874
rect 6009 9831 6061 9840
rect 4409 8664 4461 8673
rect 4409 8630 4418 8664
rect 4418 8630 4452 8664
rect 4452 8630 4461 8664
rect 4409 8621 4461 8630
rect 2809 7454 2861 7463
rect 2809 7420 2818 7454
rect 2818 7420 2852 7454
rect 2852 7420 2861 7454
rect 2809 7411 2861 7420
rect 1209 6244 1261 6253
rect 1209 6210 1218 6244
rect 1218 6210 1252 6244
rect 1252 6210 1261 6244
rect 1209 6201 1261 6210
rect 9 5263 18 5271
rect 18 5263 52 5271
rect 52 5263 61 5271
rect 9 5219 61 5263
rect 209 5437 261 5481
rect 209 5429 218 5437
rect 218 5429 252 5437
rect 252 5429 261 5437
rect 409 5543 418 5551
rect 418 5543 452 5551
rect 452 5543 461 5551
rect 409 5499 461 5543
rect 609 5717 661 5761
rect 609 5709 618 5717
rect 618 5709 652 5717
rect 652 5709 661 5717
rect 809 5823 818 5831
rect 818 5823 852 5831
rect 852 5823 861 5831
rect 809 5779 861 5823
rect 1009 5997 1061 6041
rect 1009 5989 1018 5997
rect 1018 5989 1052 5997
rect 1052 5989 1061 5997
rect 1209 6103 1218 6111
rect 1218 6103 1252 6111
rect 1252 6103 1261 6111
rect 1209 6059 1261 6103
rect 1409 6367 1461 6411
rect 1409 6359 1418 6367
rect 1418 6359 1452 6367
rect 1452 6359 1461 6367
rect 1609 6473 1618 6481
rect 1618 6473 1652 6481
rect 1652 6473 1661 6481
rect 1609 6429 1661 6473
rect 1809 6647 1861 6691
rect 1809 6639 1818 6647
rect 1818 6639 1852 6647
rect 1852 6639 1861 6647
rect 2009 6753 2018 6761
rect 2018 6753 2052 6761
rect 2052 6753 2061 6761
rect 2009 6709 2061 6753
rect 2209 6927 2261 6971
rect 2209 6919 2218 6927
rect 2218 6919 2252 6927
rect 2252 6919 2261 6927
rect 2409 7033 2418 7041
rect 2418 7033 2452 7041
rect 2452 7033 2461 7041
rect 2409 6989 2461 7033
rect 2609 7207 2661 7251
rect 2609 7199 2618 7207
rect 2618 7199 2652 7207
rect 2652 7199 2661 7207
rect 2809 7313 2818 7321
rect 2818 7313 2852 7321
rect 2852 7313 2861 7321
rect 2809 7269 2861 7313
rect 3009 7577 3061 7621
rect 3009 7569 3018 7577
rect 3018 7569 3052 7577
rect 3052 7569 3061 7577
rect 3209 7683 3218 7691
rect 3218 7683 3252 7691
rect 3252 7683 3261 7691
rect 3209 7639 3261 7683
rect 3409 7857 3461 7901
rect 3409 7849 3418 7857
rect 3418 7849 3452 7857
rect 3452 7849 3461 7857
rect 3609 7963 3618 7971
rect 3618 7963 3652 7971
rect 3652 7963 3661 7971
rect 3609 7919 3661 7963
rect 3809 8137 3861 8181
rect 3809 8129 3818 8137
rect 3818 8129 3852 8137
rect 3852 8129 3861 8137
rect 4009 8243 4018 8251
rect 4018 8243 4052 8251
rect 4052 8243 4061 8251
rect 4009 8199 4061 8243
rect 4209 8417 4261 8461
rect 4209 8409 4218 8417
rect 4218 8409 4252 8417
rect 4252 8409 4261 8417
rect 4409 8523 4418 8531
rect 4418 8523 4452 8531
rect 4452 8523 4461 8531
rect 4409 8479 4461 8523
rect 4609 8787 4661 8831
rect 4609 8779 4618 8787
rect 4618 8779 4652 8787
rect 4652 8779 4661 8787
rect 4809 8893 4818 8901
rect 4818 8893 4852 8901
rect 4852 8893 4861 8901
rect 4809 8849 4861 8893
rect 5009 9067 5061 9111
rect 5009 9059 5018 9067
rect 5018 9059 5052 9067
rect 5052 9059 5061 9067
rect 5209 9173 5218 9181
rect 5218 9173 5252 9181
rect 5252 9173 5261 9181
rect 5209 9129 5261 9173
rect 5409 9347 5461 9391
rect 5409 9339 5418 9347
rect 5418 9339 5452 9347
rect 5452 9339 5461 9347
rect 5609 9453 5618 9461
rect 5618 9453 5652 9461
rect 5652 9453 5661 9461
rect 5609 9409 5661 9453
rect 5809 9627 5861 9671
rect 5809 9619 5818 9627
rect 5818 9619 5852 9627
rect 5852 9619 5861 9627
rect 6009 9733 6018 9741
rect 6018 9733 6052 9741
rect 6052 9733 6061 9741
rect 6009 9689 6061 9733
rect 6209 9890 6261 9899
rect 6209 9856 6218 9890
rect 6218 9856 6252 9890
rect 6252 9856 6261 9890
rect 6209 9847 6261 9856
rect 4609 8680 4661 8689
rect 4609 8646 4618 8680
rect 4618 8646 4652 8680
rect 4652 8646 4661 8680
rect 4609 8637 4661 8646
rect 3009 7470 3061 7479
rect 3009 7436 3018 7470
rect 3018 7436 3052 7470
rect 3052 7436 3061 7470
rect 3009 7427 3061 7436
rect 1409 6260 1461 6269
rect 1409 6226 1418 6260
rect 1418 6226 1452 6260
rect 1452 6226 1461 6260
rect 1409 6217 1461 6226
rect 9 5123 18 5131
rect 18 5123 52 5131
rect 52 5123 61 5131
rect 9 5079 61 5123
rect 209 5297 261 5341
rect 209 5289 218 5297
rect 218 5289 252 5297
rect 252 5289 261 5297
rect 409 5403 418 5411
rect 418 5403 452 5411
rect 452 5403 461 5411
rect 409 5359 461 5403
rect 609 5577 661 5621
rect 609 5569 618 5577
rect 618 5569 652 5577
rect 652 5569 661 5577
rect 809 5683 818 5691
rect 818 5683 852 5691
rect 852 5683 861 5691
rect 809 5639 861 5683
rect 1009 5857 1061 5901
rect 1009 5849 1018 5857
rect 1018 5849 1052 5857
rect 1052 5849 1061 5857
rect 1209 5963 1218 5971
rect 1218 5963 1252 5971
rect 1252 5963 1261 5971
rect 1209 5919 1261 5963
rect 1409 6137 1461 6181
rect 1409 6129 1418 6137
rect 1418 6129 1452 6137
rect 1452 6129 1461 6137
rect 1609 6333 1618 6341
rect 1618 6333 1652 6341
rect 1652 6333 1661 6341
rect 1609 6289 1661 6333
rect 1809 6507 1861 6551
rect 1809 6499 1818 6507
rect 1818 6499 1852 6507
rect 1852 6499 1861 6507
rect 2009 6613 2018 6621
rect 2018 6613 2052 6621
rect 2052 6613 2061 6621
rect 2009 6569 2061 6613
rect 2209 6787 2261 6831
rect 2209 6779 2218 6787
rect 2218 6779 2252 6787
rect 2252 6779 2261 6787
rect 2409 6893 2418 6901
rect 2418 6893 2452 6901
rect 2452 6893 2461 6901
rect 2409 6849 2461 6893
rect 2609 7067 2661 7111
rect 2609 7059 2618 7067
rect 2618 7059 2652 7067
rect 2652 7059 2661 7067
rect 2809 7173 2818 7181
rect 2818 7173 2852 7181
rect 2852 7173 2861 7181
rect 2809 7129 2861 7173
rect 3009 7347 3061 7391
rect 3009 7339 3018 7347
rect 3018 7339 3052 7347
rect 3052 7339 3061 7347
rect 3209 7543 3218 7551
rect 3218 7543 3252 7551
rect 3252 7543 3261 7551
rect 3209 7499 3261 7543
rect 3409 7717 3461 7761
rect 3409 7709 3418 7717
rect 3418 7709 3452 7717
rect 3452 7709 3461 7717
rect 3609 7823 3618 7831
rect 3618 7823 3652 7831
rect 3652 7823 3661 7831
rect 3609 7779 3661 7823
rect 3809 7997 3861 8041
rect 3809 7989 3818 7997
rect 3818 7989 3852 7997
rect 3852 7989 3861 7997
rect 4009 8103 4018 8111
rect 4018 8103 4052 8111
rect 4052 8103 4061 8111
rect 4009 8059 4061 8103
rect 4209 8277 4261 8321
rect 4209 8269 4218 8277
rect 4218 8269 4252 8277
rect 4252 8269 4261 8277
rect 4409 8383 4418 8391
rect 4418 8383 4452 8391
rect 4452 8383 4461 8391
rect 4409 8339 4461 8383
rect 4609 8557 4661 8601
rect 4609 8549 4618 8557
rect 4618 8549 4652 8557
rect 4652 8549 4661 8557
rect 4809 8753 4818 8761
rect 4818 8753 4852 8761
rect 4852 8753 4861 8761
rect 4809 8709 4861 8753
rect 5009 8927 5061 8971
rect 5009 8919 5018 8927
rect 5018 8919 5052 8927
rect 5052 8919 5061 8927
rect 5209 9033 5218 9041
rect 5218 9033 5252 9041
rect 5252 9033 5261 9041
rect 5209 8989 5261 9033
rect 5409 9207 5461 9251
rect 5409 9199 5418 9207
rect 5418 9199 5452 9207
rect 5452 9199 5461 9207
rect 5609 9313 5618 9321
rect 5618 9313 5652 9321
rect 5652 9313 5661 9321
rect 5609 9269 5661 9313
rect 5809 9487 5861 9531
rect 5809 9479 5818 9487
rect 5818 9479 5852 9487
rect 5852 9479 5861 9487
rect 6009 9593 6018 9601
rect 6018 9593 6052 9601
rect 6052 9593 6061 9601
rect 6009 9549 6061 9593
rect 6209 9767 6261 9811
rect 6209 9759 6218 9767
rect 6218 9759 6252 9767
rect 6252 9759 6261 9767
rect 4809 8664 4861 8673
rect 4809 8630 4818 8664
rect 4818 8630 4852 8664
rect 4852 8630 4861 8664
rect 4809 8621 4861 8630
rect 3209 7454 3261 7463
rect 3209 7420 3218 7454
rect 3218 7420 3252 7454
rect 3252 7420 3261 7454
rect 3209 7411 3261 7420
rect 1609 6244 1661 6253
rect 1609 6210 1618 6244
rect 1618 6210 1652 6244
rect 1652 6210 1661 6244
rect 1609 6201 1661 6210
rect 209 5157 261 5201
rect 209 5149 218 5157
rect 218 5149 252 5157
rect 252 5149 261 5157
rect 409 5263 418 5271
rect 418 5263 452 5271
rect 452 5263 461 5271
rect 409 5219 461 5263
rect 609 5437 661 5481
rect 609 5429 618 5437
rect 618 5429 652 5437
rect 652 5429 661 5437
rect 809 5543 818 5551
rect 818 5543 852 5551
rect 852 5543 861 5551
rect 809 5499 861 5543
rect 1009 5717 1061 5761
rect 1009 5709 1018 5717
rect 1018 5709 1052 5717
rect 1052 5709 1061 5717
rect 1209 5823 1218 5831
rect 1218 5823 1252 5831
rect 1252 5823 1261 5831
rect 1209 5779 1261 5823
rect 1409 5997 1461 6041
rect 1409 5989 1418 5997
rect 1418 5989 1452 5997
rect 1452 5989 1461 5997
rect 1609 6103 1618 6111
rect 1618 6103 1652 6111
rect 1652 6103 1661 6111
rect 1609 6059 1661 6103
rect 1809 6367 1861 6411
rect 1809 6359 1818 6367
rect 1818 6359 1852 6367
rect 1852 6359 1861 6367
rect 2009 6473 2018 6481
rect 2018 6473 2052 6481
rect 2052 6473 2061 6481
rect 2009 6429 2061 6473
rect 2209 6647 2261 6691
rect 2209 6639 2218 6647
rect 2218 6639 2252 6647
rect 2252 6639 2261 6647
rect 2409 6753 2418 6761
rect 2418 6753 2452 6761
rect 2452 6753 2461 6761
rect 2409 6709 2461 6753
rect 2609 6927 2661 6971
rect 2609 6919 2618 6927
rect 2618 6919 2652 6927
rect 2652 6919 2661 6927
rect 2809 7033 2818 7041
rect 2818 7033 2852 7041
rect 2852 7033 2861 7041
rect 2809 6989 2861 7033
rect 3009 7207 3061 7251
rect 3009 7199 3018 7207
rect 3018 7199 3052 7207
rect 3052 7199 3061 7207
rect 3209 7313 3218 7321
rect 3218 7313 3252 7321
rect 3252 7313 3261 7321
rect 3209 7269 3261 7313
rect 3409 7577 3461 7621
rect 3409 7569 3418 7577
rect 3418 7569 3452 7577
rect 3452 7569 3461 7577
rect 3609 7683 3618 7691
rect 3618 7683 3652 7691
rect 3652 7683 3661 7691
rect 3609 7639 3661 7683
rect 3809 7857 3861 7901
rect 3809 7849 3818 7857
rect 3818 7849 3852 7857
rect 3852 7849 3861 7857
rect 4009 7963 4018 7971
rect 4018 7963 4052 7971
rect 4052 7963 4061 7971
rect 4009 7919 4061 7963
rect 4209 8137 4261 8181
rect 4209 8129 4218 8137
rect 4218 8129 4252 8137
rect 4252 8129 4261 8137
rect 4409 8243 4418 8251
rect 4418 8243 4452 8251
rect 4452 8243 4461 8251
rect 4409 8199 4461 8243
rect 4609 8417 4661 8461
rect 4609 8409 4618 8417
rect 4618 8409 4652 8417
rect 4652 8409 4661 8417
rect 4809 8523 4818 8531
rect 4818 8523 4852 8531
rect 4852 8523 4861 8531
rect 4809 8479 4861 8523
rect 5009 8787 5061 8831
rect 5009 8779 5018 8787
rect 5018 8779 5052 8787
rect 5052 8779 5061 8787
rect 5209 8893 5218 8901
rect 5218 8893 5252 8901
rect 5252 8893 5261 8901
rect 5209 8849 5261 8893
rect 5409 9067 5461 9111
rect 5409 9059 5418 9067
rect 5418 9059 5452 9067
rect 5452 9059 5461 9067
rect 5609 9173 5618 9181
rect 5618 9173 5652 9181
rect 5652 9173 5661 9181
rect 5609 9129 5661 9173
rect 5809 9347 5861 9391
rect 5809 9339 5818 9347
rect 5818 9339 5852 9347
rect 5852 9339 5861 9347
rect 6009 9453 6018 9461
rect 6018 9453 6052 9461
rect 6052 9453 6061 9461
rect 6009 9409 6061 9453
rect 6209 9627 6261 9671
rect 6209 9619 6218 9627
rect 6218 9619 6252 9627
rect 6252 9619 6261 9627
rect 6409 9733 6418 9741
rect 6418 9733 6452 9741
rect 6452 9733 6461 9741
rect 6409 9689 6461 9733
rect 6507 9689 6559 9741
rect 5009 8680 5061 8689
rect 5009 8646 5018 8680
rect 5018 8646 5052 8680
rect 5052 8646 5061 8680
rect 5009 8637 5061 8646
rect 3409 7470 3461 7479
rect 3409 7436 3418 7470
rect 3418 7436 3452 7470
rect 3452 7436 3461 7470
rect 3409 7427 3461 7436
rect 1809 6260 1861 6269
rect 1809 6226 1818 6260
rect 1818 6226 1852 6260
rect 1852 6226 1861 6260
rect 1809 6217 1861 6226
rect 409 5123 418 5131
rect 418 5123 452 5131
rect 452 5123 461 5131
rect 409 5079 461 5123
rect 609 5297 661 5341
rect 609 5289 618 5297
rect 618 5289 652 5297
rect 652 5289 661 5297
rect 809 5403 818 5411
rect 818 5403 852 5411
rect 852 5403 861 5411
rect 809 5359 861 5403
rect 1009 5577 1061 5621
rect 1009 5569 1018 5577
rect 1018 5569 1052 5577
rect 1052 5569 1061 5577
rect 1209 5683 1218 5691
rect 1218 5683 1252 5691
rect 1252 5683 1261 5691
rect 1209 5639 1261 5683
rect 1409 5857 1461 5901
rect 1409 5849 1418 5857
rect 1418 5849 1452 5857
rect 1452 5849 1461 5857
rect 1609 5963 1618 5971
rect 1618 5963 1652 5971
rect 1652 5963 1661 5971
rect 1609 5919 1661 5963
rect 1809 6137 1861 6181
rect 1809 6129 1818 6137
rect 1818 6129 1852 6137
rect 1852 6129 1861 6137
rect 2009 6333 2018 6341
rect 2018 6333 2052 6341
rect 2052 6333 2061 6341
rect 2009 6289 2061 6333
rect 2209 6507 2261 6551
rect 2209 6499 2218 6507
rect 2218 6499 2252 6507
rect 2252 6499 2261 6507
rect 2409 6613 2418 6621
rect 2418 6613 2452 6621
rect 2452 6613 2461 6621
rect 2409 6569 2461 6613
rect 2609 6787 2661 6831
rect 2609 6779 2618 6787
rect 2618 6779 2652 6787
rect 2652 6779 2661 6787
rect 2809 6893 2818 6901
rect 2818 6893 2852 6901
rect 2852 6893 2861 6901
rect 2809 6849 2861 6893
rect 3009 7067 3061 7111
rect 3009 7059 3018 7067
rect 3018 7059 3052 7067
rect 3052 7059 3061 7067
rect 3209 7173 3218 7181
rect 3218 7173 3252 7181
rect 3252 7173 3261 7181
rect 3209 7129 3261 7173
rect 3409 7347 3461 7391
rect 3409 7339 3418 7347
rect 3418 7339 3452 7347
rect 3452 7339 3461 7347
rect 3609 7543 3618 7551
rect 3618 7543 3652 7551
rect 3652 7543 3661 7551
rect 3609 7499 3661 7543
rect 3809 7717 3861 7761
rect 3809 7709 3818 7717
rect 3818 7709 3852 7717
rect 3852 7709 3861 7717
rect 4009 7823 4018 7831
rect 4018 7823 4052 7831
rect 4052 7823 4061 7831
rect 4009 7779 4061 7823
rect 4209 7997 4261 8041
rect 4209 7989 4218 7997
rect 4218 7989 4252 7997
rect 4252 7989 4261 7997
rect 4409 8103 4418 8111
rect 4418 8103 4452 8111
rect 4452 8103 4461 8111
rect 4409 8059 4461 8103
rect 4609 8277 4661 8321
rect 4609 8269 4618 8277
rect 4618 8269 4652 8277
rect 4652 8269 4661 8277
rect 4809 8383 4818 8391
rect 4818 8383 4852 8391
rect 4852 8383 4861 8391
rect 4809 8339 4861 8383
rect 5009 8557 5061 8601
rect 5009 8549 5018 8557
rect 5018 8549 5052 8557
rect 5052 8549 5061 8557
rect 5209 8753 5218 8761
rect 5218 8753 5252 8761
rect 5252 8753 5261 8761
rect 5209 8709 5261 8753
rect 5409 8927 5461 8971
rect 5409 8919 5418 8927
rect 5418 8919 5452 8927
rect 5452 8919 5461 8927
rect 5609 9033 5618 9041
rect 5618 9033 5652 9041
rect 5652 9033 5661 9041
rect 5609 8989 5661 9033
rect 5809 9207 5861 9251
rect 5809 9199 5818 9207
rect 5818 9199 5852 9207
rect 5852 9199 5861 9207
rect 6009 9313 6018 9321
rect 6018 9313 6052 9321
rect 6052 9313 6061 9321
rect 6009 9269 6061 9313
rect 6209 9487 6261 9531
rect 6209 9479 6218 9487
rect 6218 9479 6252 9487
rect 6252 9479 6261 9487
rect 6409 9593 6418 9601
rect 6418 9593 6452 9601
rect 6452 9593 6461 9601
rect 6409 9549 6461 9593
rect 6507 9549 6559 9601
rect 5209 8664 5261 8673
rect 5209 8630 5218 8664
rect 5218 8630 5252 8664
rect 5252 8630 5261 8664
rect 5209 8621 5261 8630
rect 3609 7454 3661 7463
rect 3609 7420 3618 7454
rect 3618 7420 3652 7454
rect 3652 7420 3661 7454
rect 3609 7411 3661 7420
rect 2009 6244 2061 6253
rect 2009 6210 2018 6244
rect 2018 6210 2052 6244
rect 2052 6210 2061 6244
rect 2009 6201 2061 6210
rect 609 5157 661 5201
rect 609 5149 618 5157
rect 618 5149 652 5157
rect 652 5149 661 5157
rect 809 5263 818 5271
rect 818 5263 852 5271
rect 852 5263 861 5271
rect 809 5219 861 5263
rect 1009 5437 1061 5481
rect 1009 5429 1018 5437
rect 1018 5429 1052 5437
rect 1052 5429 1061 5437
rect 1209 5543 1218 5551
rect 1218 5543 1252 5551
rect 1252 5543 1261 5551
rect 1209 5499 1261 5543
rect 1409 5717 1461 5761
rect 1409 5709 1418 5717
rect 1418 5709 1452 5717
rect 1452 5709 1461 5717
rect 1609 5823 1618 5831
rect 1618 5823 1652 5831
rect 1652 5823 1661 5831
rect 1609 5779 1661 5823
rect 1809 5997 1861 6041
rect 1809 5989 1818 5997
rect 1818 5989 1852 5997
rect 1852 5989 1861 5997
rect 2009 6103 2018 6111
rect 2018 6103 2052 6111
rect 2052 6103 2061 6111
rect 2009 6059 2061 6103
rect 2209 6367 2261 6411
rect 2209 6359 2218 6367
rect 2218 6359 2252 6367
rect 2252 6359 2261 6367
rect 2409 6473 2418 6481
rect 2418 6473 2452 6481
rect 2452 6473 2461 6481
rect 2409 6429 2461 6473
rect 2609 6647 2661 6691
rect 2609 6639 2618 6647
rect 2618 6639 2652 6647
rect 2652 6639 2661 6647
rect 2809 6753 2818 6761
rect 2818 6753 2852 6761
rect 2852 6753 2861 6761
rect 2809 6709 2861 6753
rect 3009 6927 3061 6971
rect 3009 6919 3018 6927
rect 3018 6919 3052 6927
rect 3052 6919 3061 6927
rect 3209 7033 3218 7041
rect 3218 7033 3252 7041
rect 3252 7033 3261 7041
rect 3209 6989 3261 7033
rect 3409 7207 3461 7251
rect 3409 7199 3418 7207
rect 3418 7199 3452 7207
rect 3452 7199 3461 7207
rect 3609 7313 3618 7321
rect 3618 7313 3652 7321
rect 3652 7313 3661 7321
rect 3609 7269 3661 7313
rect 3809 7577 3861 7621
rect 3809 7569 3818 7577
rect 3818 7569 3852 7577
rect 3852 7569 3861 7577
rect 4009 7683 4018 7691
rect 4018 7683 4052 7691
rect 4052 7683 4061 7691
rect 4009 7639 4061 7683
rect 4209 7857 4261 7901
rect 4209 7849 4218 7857
rect 4218 7849 4252 7857
rect 4252 7849 4261 7857
rect 4409 7963 4418 7971
rect 4418 7963 4452 7971
rect 4452 7963 4461 7971
rect 4409 7919 4461 7963
rect 4609 8137 4661 8181
rect 4609 8129 4618 8137
rect 4618 8129 4652 8137
rect 4652 8129 4661 8137
rect 4809 8243 4818 8251
rect 4818 8243 4852 8251
rect 4852 8243 4861 8251
rect 4809 8199 4861 8243
rect 5009 8417 5061 8461
rect 5009 8409 5018 8417
rect 5018 8409 5052 8417
rect 5052 8409 5061 8417
rect 5209 8523 5218 8531
rect 5218 8523 5252 8531
rect 5252 8523 5261 8531
rect 5209 8479 5261 8523
rect 5409 8787 5461 8831
rect 5409 8779 5418 8787
rect 5418 8779 5452 8787
rect 5452 8779 5461 8787
rect 5609 8893 5618 8901
rect 5618 8893 5652 8901
rect 5652 8893 5661 8901
rect 5609 8849 5661 8893
rect 5809 9067 5861 9111
rect 5809 9059 5818 9067
rect 5818 9059 5852 9067
rect 5852 9059 5861 9067
rect 6009 9173 6018 9181
rect 6018 9173 6052 9181
rect 6052 9173 6061 9181
rect 6009 9129 6061 9173
rect 6209 9347 6261 9391
rect 6209 9339 6218 9347
rect 6218 9339 6252 9347
rect 6252 9339 6261 9347
rect 6409 9453 6418 9461
rect 6418 9453 6452 9461
rect 6452 9453 6461 9461
rect 6409 9409 6461 9453
rect 6507 9409 6559 9461
rect 5409 8680 5461 8689
rect 5409 8646 5418 8680
rect 5418 8646 5452 8680
rect 5452 8646 5461 8680
rect 5409 8637 5461 8646
rect 3809 7470 3861 7479
rect 3809 7436 3818 7470
rect 3818 7436 3852 7470
rect 3852 7436 3861 7470
rect 3809 7427 3861 7436
rect 2209 6260 2261 6269
rect 2209 6226 2218 6260
rect 2218 6226 2252 6260
rect 2252 6226 2261 6260
rect 2209 6217 2261 6226
rect 809 5123 818 5131
rect 818 5123 852 5131
rect 852 5123 861 5131
rect 809 5079 861 5123
rect 1009 5297 1061 5341
rect 1009 5289 1018 5297
rect 1018 5289 1052 5297
rect 1052 5289 1061 5297
rect 1209 5403 1218 5411
rect 1218 5403 1252 5411
rect 1252 5403 1261 5411
rect 1209 5359 1261 5403
rect 1409 5577 1461 5621
rect 1409 5569 1418 5577
rect 1418 5569 1452 5577
rect 1452 5569 1461 5577
rect 1609 5683 1618 5691
rect 1618 5683 1652 5691
rect 1652 5683 1661 5691
rect 1609 5639 1661 5683
rect 1809 5857 1861 5901
rect 1809 5849 1818 5857
rect 1818 5849 1852 5857
rect 1852 5849 1861 5857
rect 2009 5963 2018 5971
rect 2018 5963 2052 5971
rect 2052 5963 2061 5971
rect 2009 5919 2061 5963
rect 2209 6137 2261 6181
rect 2209 6129 2218 6137
rect 2218 6129 2252 6137
rect 2252 6129 2261 6137
rect 2409 6333 2418 6341
rect 2418 6333 2452 6341
rect 2452 6333 2461 6341
rect 2409 6289 2461 6333
rect 2609 6507 2661 6551
rect 2609 6499 2618 6507
rect 2618 6499 2652 6507
rect 2652 6499 2661 6507
rect 2809 6613 2818 6621
rect 2818 6613 2852 6621
rect 2852 6613 2861 6621
rect 2809 6569 2861 6613
rect 3009 6787 3061 6831
rect 3009 6779 3018 6787
rect 3018 6779 3052 6787
rect 3052 6779 3061 6787
rect 3209 6893 3218 6901
rect 3218 6893 3252 6901
rect 3252 6893 3261 6901
rect 3209 6849 3261 6893
rect 3409 7067 3461 7111
rect 3409 7059 3418 7067
rect 3418 7059 3452 7067
rect 3452 7059 3461 7067
rect 3609 7173 3618 7181
rect 3618 7173 3652 7181
rect 3652 7173 3661 7181
rect 3609 7129 3661 7173
rect 3809 7347 3861 7391
rect 3809 7339 3818 7347
rect 3818 7339 3852 7347
rect 3852 7339 3861 7347
rect 4009 7543 4018 7551
rect 4018 7543 4052 7551
rect 4052 7543 4061 7551
rect 4009 7499 4061 7543
rect 4209 7717 4261 7761
rect 4209 7709 4218 7717
rect 4218 7709 4252 7717
rect 4252 7709 4261 7717
rect 4409 7823 4418 7831
rect 4418 7823 4452 7831
rect 4452 7823 4461 7831
rect 4409 7779 4461 7823
rect 4609 7997 4661 8041
rect 4609 7989 4618 7997
rect 4618 7989 4652 7997
rect 4652 7989 4661 7997
rect 4809 8103 4818 8111
rect 4818 8103 4852 8111
rect 4852 8103 4861 8111
rect 4809 8059 4861 8103
rect 5009 8277 5061 8321
rect 5009 8269 5018 8277
rect 5018 8269 5052 8277
rect 5052 8269 5061 8277
rect 5209 8383 5218 8391
rect 5218 8383 5252 8391
rect 5252 8383 5261 8391
rect 5209 8339 5261 8383
rect 5409 8557 5461 8601
rect 5409 8549 5418 8557
rect 5418 8549 5452 8557
rect 5452 8549 5461 8557
rect 5609 8753 5618 8761
rect 5618 8753 5652 8761
rect 5652 8753 5661 8761
rect 5609 8709 5661 8753
rect 5809 8927 5861 8971
rect 5809 8919 5818 8927
rect 5818 8919 5852 8927
rect 5852 8919 5861 8927
rect 6009 9033 6018 9041
rect 6018 9033 6052 9041
rect 6052 9033 6061 9041
rect 6009 8989 6061 9033
rect 6209 9207 6261 9251
rect 6209 9199 6218 9207
rect 6218 9199 6252 9207
rect 6252 9199 6261 9207
rect 6409 9313 6418 9321
rect 6418 9313 6452 9321
rect 6452 9313 6461 9321
rect 6409 9269 6461 9313
rect 6507 9269 6559 9321
rect 5609 8664 5661 8673
rect 5609 8630 5618 8664
rect 5618 8630 5652 8664
rect 5652 8630 5661 8664
rect 5609 8621 5661 8630
rect 4009 7454 4061 7463
rect 4009 7420 4018 7454
rect 4018 7420 4052 7454
rect 4052 7420 4061 7454
rect 4009 7411 4061 7420
rect 2409 6244 2461 6253
rect 2409 6210 2418 6244
rect 2418 6210 2452 6244
rect 2452 6210 2461 6244
rect 2409 6201 2461 6210
rect 1009 5157 1061 5201
rect 1009 5149 1018 5157
rect 1018 5149 1052 5157
rect 1052 5149 1061 5157
rect 1209 5263 1218 5271
rect 1218 5263 1252 5271
rect 1252 5263 1261 5271
rect 1209 5219 1261 5263
rect 1409 5437 1461 5481
rect 1409 5429 1418 5437
rect 1418 5429 1452 5437
rect 1452 5429 1461 5437
rect 1609 5543 1618 5551
rect 1618 5543 1652 5551
rect 1652 5543 1661 5551
rect 1609 5499 1661 5543
rect 1809 5717 1861 5761
rect 1809 5709 1818 5717
rect 1818 5709 1852 5717
rect 1852 5709 1861 5717
rect 2009 5823 2018 5831
rect 2018 5823 2052 5831
rect 2052 5823 2061 5831
rect 2009 5779 2061 5823
rect 2209 5997 2261 6041
rect 2209 5989 2218 5997
rect 2218 5989 2252 5997
rect 2252 5989 2261 5997
rect 2409 6103 2418 6111
rect 2418 6103 2452 6111
rect 2452 6103 2461 6111
rect 2409 6059 2461 6103
rect 2609 6367 2661 6411
rect 2609 6359 2618 6367
rect 2618 6359 2652 6367
rect 2652 6359 2661 6367
rect 2809 6473 2818 6481
rect 2818 6473 2852 6481
rect 2852 6473 2861 6481
rect 2809 6429 2861 6473
rect 3009 6647 3061 6691
rect 3009 6639 3018 6647
rect 3018 6639 3052 6647
rect 3052 6639 3061 6647
rect 3209 6753 3218 6761
rect 3218 6753 3252 6761
rect 3252 6753 3261 6761
rect 3209 6709 3261 6753
rect 3409 6927 3461 6971
rect 3409 6919 3418 6927
rect 3418 6919 3452 6927
rect 3452 6919 3461 6927
rect 3609 7033 3618 7041
rect 3618 7033 3652 7041
rect 3652 7033 3661 7041
rect 3609 6989 3661 7033
rect 3809 7207 3861 7251
rect 3809 7199 3818 7207
rect 3818 7199 3852 7207
rect 3852 7199 3861 7207
rect 4009 7313 4018 7321
rect 4018 7313 4052 7321
rect 4052 7313 4061 7321
rect 4009 7269 4061 7313
rect 4209 7577 4261 7621
rect 4209 7569 4218 7577
rect 4218 7569 4252 7577
rect 4252 7569 4261 7577
rect 4409 7683 4418 7691
rect 4418 7683 4452 7691
rect 4452 7683 4461 7691
rect 4409 7639 4461 7683
rect 4609 7857 4661 7901
rect 4609 7849 4618 7857
rect 4618 7849 4652 7857
rect 4652 7849 4661 7857
rect 4809 7963 4818 7971
rect 4818 7963 4852 7971
rect 4852 7963 4861 7971
rect 4809 7919 4861 7963
rect 5009 8137 5061 8181
rect 5009 8129 5018 8137
rect 5018 8129 5052 8137
rect 5052 8129 5061 8137
rect 5209 8243 5218 8251
rect 5218 8243 5252 8251
rect 5252 8243 5261 8251
rect 5209 8199 5261 8243
rect 5409 8417 5461 8461
rect 5409 8409 5418 8417
rect 5418 8409 5452 8417
rect 5452 8409 5461 8417
rect 5609 8523 5618 8531
rect 5618 8523 5652 8531
rect 5652 8523 5661 8531
rect 5609 8479 5661 8523
rect 5809 8787 5861 8831
rect 5809 8779 5818 8787
rect 5818 8779 5852 8787
rect 5852 8779 5861 8787
rect 6009 8893 6018 8901
rect 6018 8893 6052 8901
rect 6052 8893 6061 8901
rect 6009 8849 6061 8893
rect 6209 9067 6261 9111
rect 6209 9059 6218 9067
rect 6218 9059 6252 9067
rect 6252 9059 6261 9067
rect 6409 9173 6418 9181
rect 6418 9173 6452 9181
rect 6452 9173 6461 9181
rect 6409 9129 6461 9173
rect 6507 9129 6559 9181
rect 5809 8680 5861 8689
rect 5809 8646 5818 8680
rect 5818 8646 5852 8680
rect 5852 8646 5861 8680
rect 5809 8637 5861 8646
rect 4209 7470 4261 7479
rect 4209 7436 4218 7470
rect 4218 7436 4252 7470
rect 4252 7436 4261 7470
rect 4209 7427 4261 7436
rect 2609 6260 2661 6269
rect 2609 6226 2618 6260
rect 2618 6226 2652 6260
rect 2652 6226 2661 6260
rect 2609 6217 2661 6226
rect 1209 5123 1218 5131
rect 1218 5123 1252 5131
rect 1252 5123 1261 5131
rect 1209 5079 1261 5123
rect 1409 5297 1461 5341
rect 1409 5289 1418 5297
rect 1418 5289 1452 5297
rect 1452 5289 1461 5297
rect 1609 5403 1618 5411
rect 1618 5403 1652 5411
rect 1652 5403 1661 5411
rect 1609 5359 1661 5403
rect 1809 5577 1861 5621
rect 1809 5569 1818 5577
rect 1818 5569 1852 5577
rect 1852 5569 1861 5577
rect 2009 5683 2018 5691
rect 2018 5683 2052 5691
rect 2052 5683 2061 5691
rect 2009 5639 2061 5683
rect 2209 5857 2261 5901
rect 2209 5849 2218 5857
rect 2218 5849 2252 5857
rect 2252 5849 2261 5857
rect 2409 5963 2418 5971
rect 2418 5963 2452 5971
rect 2452 5963 2461 5971
rect 2409 5919 2461 5963
rect 2609 6137 2661 6181
rect 2609 6129 2618 6137
rect 2618 6129 2652 6137
rect 2652 6129 2661 6137
rect 2809 6333 2818 6341
rect 2818 6333 2852 6341
rect 2852 6333 2861 6341
rect 2809 6289 2861 6333
rect 3009 6507 3061 6551
rect 3009 6499 3018 6507
rect 3018 6499 3052 6507
rect 3052 6499 3061 6507
rect 3209 6613 3218 6621
rect 3218 6613 3252 6621
rect 3252 6613 3261 6621
rect 3209 6569 3261 6613
rect 3409 6787 3461 6831
rect 3409 6779 3418 6787
rect 3418 6779 3452 6787
rect 3452 6779 3461 6787
rect 3609 6893 3618 6901
rect 3618 6893 3652 6901
rect 3652 6893 3661 6901
rect 3609 6849 3661 6893
rect 3809 7067 3861 7111
rect 3809 7059 3818 7067
rect 3818 7059 3852 7067
rect 3852 7059 3861 7067
rect 4009 7173 4018 7181
rect 4018 7173 4052 7181
rect 4052 7173 4061 7181
rect 4009 7129 4061 7173
rect 4209 7347 4261 7391
rect 4209 7339 4218 7347
rect 4218 7339 4252 7347
rect 4252 7339 4261 7347
rect 4409 7543 4418 7551
rect 4418 7543 4452 7551
rect 4452 7543 4461 7551
rect 4409 7499 4461 7543
rect 4609 7717 4661 7761
rect 4609 7709 4618 7717
rect 4618 7709 4652 7717
rect 4652 7709 4661 7717
rect 4809 7823 4818 7831
rect 4818 7823 4852 7831
rect 4852 7823 4861 7831
rect 4809 7779 4861 7823
rect 5009 7997 5061 8041
rect 5009 7989 5018 7997
rect 5018 7989 5052 7997
rect 5052 7989 5061 7997
rect 5209 8103 5218 8111
rect 5218 8103 5252 8111
rect 5252 8103 5261 8111
rect 5209 8059 5261 8103
rect 5409 8277 5461 8321
rect 5409 8269 5418 8277
rect 5418 8269 5452 8277
rect 5452 8269 5461 8277
rect 5609 8383 5618 8391
rect 5618 8383 5652 8391
rect 5652 8383 5661 8391
rect 5609 8339 5661 8383
rect 5809 8557 5861 8601
rect 5809 8549 5818 8557
rect 5818 8549 5852 8557
rect 5852 8549 5861 8557
rect 6009 8753 6018 8761
rect 6018 8753 6052 8761
rect 6052 8753 6061 8761
rect 6009 8709 6061 8753
rect 6209 8927 6261 8971
rect 6209 8919 6218 8927
rect 6218 8919 6252 8927
rect 6252 8919 6261 8927
rect 6409 9033 6418 9041
rect 6418 9033 6452 9041
rect 6452 9033 6461 9041
rect 6409 8989 6461 9033
rect 6507 8989 6559 9041
rect 6009 8664 6061 8673
rect 6009 8630 6018 8664
rect 6018 8630 6052 8664
rect 6052 8630 6061 8664
rect 6009 8621 6061 8630
rect 4409 7454 4461 7463
rect 4409 7420 4418 7454
rect 4418 7420 4452 7454
rect 4452 7420 4461 7454
rect 4409 7411 4461 7420
rect 2809 6244 2861 6253
rect 2809 6210 2818 6244
rect 2818 6210 2852 6244
rect 2852 6210 2861 6244
rect 2809 6201 2861 6210
rect 1409 5157 1461 5201
rect 1409 5149 1418 5157
rect 1418 5149 1452 5157
rect 1452 5149 1461 5157
rect 1609 5263 1618 5271
rect 1618 5263 1652 5271
rect 1652 5263 1661 5271
rect 1609 5219 1661 5263
rect 1809 5437 1861 5481
rect 1809 5429 1818 5437
rect 1818 5429 1852 5437
rect 1852 5429 1861 5437
rect 2009 5543 2018 5551
rect 2018 5543 2052 5551
rect 2052 5543 2061 5551
rect 2009 5499 2061 5543
rect 2209 5717 2261 5761
rect 2209 5709 2218 5717
rect 2218 5709 2252 5717
rect 2252 5709 2261 5717
rect 2409 5823 2418 5831
rect 2418 5823 2452 5831
rect 2452 5823 2461 5831
rect 2409 5779 2461 5823
rect 2609 5997 2661 6041
rect 2609 5989 2618 5997
rect 2618 5989 2652 5997
rect 2652 5989 2661 5997
rect 2809 6103 2818 6111
rect 2818 6103 2852 6111
rect 2852 6103 2861 6111
rect 2809 6059 2861 6103
rect 3009 6367 3061 6411
rect 3009 6359 3018 6367
rect 3018 6359 3052 6367
rect 3052 6359 3061 6367
rect 3209 6473 3218 6481
rect 3218 6473 3252 6481
rect 3252 6473 3261 6481
rect 3209 6429 3261 6473
rect 3409 6647 3461 6691
rect 3409 6639 3418 6647
rect 3418 6639 3452 6647
rect 3452 6639 3461 6647
rect 3609 6753 3618 6761
rect 3618 6753 3652 6761
rect 3652 6753 3661 6761
rect 3609 6709 3661 6753
rect 3809 6927 3861 6971
rect 3809 6919 3818 6927
rect 3818 6919 3852 6927
rect 3852 6919 3861 6927
rect 4009 7033 4018 7041
rect 4018 7033 4052 7041
rect 4052 7033 4061 7041
rect 4009 6989 4061 7033
rect 4209 7207 4261 7251
rect 4209 7199 4218 7207
rect 4218 7199 4252 7207
rect 4252 7199 4261 7207
rect 4409 7313 4418 7321
rect 4418 7313 4452 7321
rect 4452 7313 4461 7321
rect 4409 7269 4461 7313
rect 4609 7577 4661 7621
rect 4609 7569 4618 7577
rect 4618 7569 4652 7577
rect 4652 7569 4661 7577
rect 4809 7683 4818 7691
rect 4818 7683 4852 7691
rect 4852 7683 4861 7691
rect 4809 7639 4861 7683
rect 5009 7857 5061 7901
rect 5009 7849 5018 7857
rect 5018 7849 5052 7857
rect 5052 7849 5061 7857
rect 5209 7963 5218 7971
rect 5218 7963 5252 7971
rect 5252 7963 5261 7971
rect 5209 7919 5261 7963
rect 5409 8137 5461 8181
rect 5409 8129 5418 8137
rect 5418 8129 5452 8137
rect 5452 8129 5461 8137
rect 5609 8243 5618 8251
rect 5618 8243 5652 8251
rect 5652 8243 5661 8251
rect 5609 8199 5661 8243
rect 5809 8417 5861 8461
rect 5809 8409 5818 8417
rect 5818 8409 5852 8417
rect 5852 8409 5861 8417
rect 6009 8523 6018 8531
rect 6018 8523 6052 8531
rect 6052 8523 6061 8531
rect 6009 8479 6061 8523
rect 6209 8787 6261 8831
rect 6209 8779 6218 8787
rect 6218 8779 6252 8787
rect 6252 8779 6261 8787
rect 6409 8893 6418 8901
rect 6418 8893 6452 8901
rect 6452 8893 6461 8901
rect 6409 8849 6461 8893
rect 6507 8849 6559 8901
rect 6209 8680 6261 8689
rect 6209 8646 6218 8680
rect 6218 8646 6252 8680
rect 6252 8646 6261 8680
rect 6209 8637 6261 8646
rect 4609 7470 4661 7479
rect 4609 7436 4618 7470
rect 4618 7436 4652 7470
rect 4652 7436 4661 7470
rect 4609 7427 4661 7436
rect 3009 6260 3061 6269
rect 3009 6226 3018 6260
rect 3018 6226 3052 6260
rect 3052 6226 3061 6260
rect 3009 6217 3061 6226
rect 1609 5123 1618 5131
rect 1618 5123 1652 5131
rect 1652 5123 1661 5131
rect 1609 5079 1661 5123
rect 1809 5297 1861 5341
rect 1809 5289 1818 5297
rect 1818 5289 1852 5297
rect 1852 5289 1861 5297
rect 2009 5403 2018 5411
rect 2018 5403 2052 5411
rect 2052 5403 2061 5411
rect 2009 5359 2061 5403
rect 2209 5577 2261 5621
rect 2209 5569 2218 5577
rect 2218 5569 2252 5577
rect 2252 5569 2261 5577
rect 2409 5683 2418 5691
rect 2418 5683 2452 5691
rect 2452 5683 2461 5691
rect 2409 5639 2461 5683
rect 2609 5857 2661 5901
rect 2609 5849 2618 5857
rect 2618 5849 2652 5857
rect 2652 5849 2661 5857
rect 2809 5963 2818 5971
rect 2818 5963 2852 5971
rect 2852 5963 2861 5971
rect 2809 5919 2861 5963
rect 3009 6137 3061 6181
rect 3009 6129 3018 6137
rect 3018 6129 3052 6137
rect 3052 6129 3061 6137
rect 3209 6333 3218 6341
rect 3218 6333 3252 6341
rect 3252 6333 3261 6341
rect 3209 6289 3261 6333
rect 3409 6507 3461 6551
rect 3409 6499 3418 6507
rect 3418 6499 3452 6507
rect 3452 6499 3461 6507
rect 3609 6613 3618 6621
rect 3618 6613 3652 6621
rect 3652 6613 3661 6621
rect 3609 6569 3661 6613
rect 3809 6787 3861 6831
rect 3809 6779 3818 6787
rect 3818 6779 3852 6787
rect 3852 6779 3861 6787
rect 4009 6893 4018 6901
rect 4018 6893 4052 6901
rect 4052 6893 4061 6901
rect 4009 6849 4061 6893
rect 4209 7067 4261 7111
rect 4209 7059 4218 7067
rect 4218 7059 4252 7067
rect 4252 7059 4261 7067
rect 4409 7173 4418 7181
rect 4418 7173 4452 7181
rect 4452 7173 4461 7181
rect 4409 7129 4461 7173
rect 4609 7347 4661 7391
rect 4609 7339 4618 7347
rect 4618 7339 4652 7347
rect 4652 7339 4661 7347
rect 4809 7543 4818 7551
rect 4818 7543 4852 7551
rect 4852 7543 4861 7551
rect 4809 7499 4861 7543
rect 5009 7717 5061 7761
rect 5009 7709 5018 7717
rect 5018 7709 5052 7717
rect 5052 7709 5061 7717
rect 5209 7823 5218 7831
rect 5218 7823 5252 7831
rect 5252 7823 5261 7831
rect 5209 7779 5261 7823
rect 5409 7997 5461 8041
rect 5409 7989 5418 7997
rect 5418 7989 5452 7997
rect 5452 7989 5461 7997
rect 5609 8103 5618 8111
rect 5618 8103 5652 8111
rect 5652 8103 5661 8111
rect 5609 8059 5661 8103
rect 5809 8277 5861 8321
rect 5809 8269 5818 8277
rect 5818 8269 5852 8277
rect 5852 8269 5861 8277
rect 6009 8383 6018 8391
rect 6018 8383 6052 8391
rect 6052 8383 6061 8391
rect 6009 8339 6061 8383
rect 6209 8557 6261 8601
rect 6209 8549 6218 8557
rect 6218 8549 6252 8557
rect 6252 8549 6261 8557
rect 6409 8753 6418 8761
rect 6418 8753 6452 8761
rect 6452 8753 6461 8761
rect 6409 8709 6461 8753
rect 6507 8709 6559 8761
rect 4809 7454 4861 7463
rect 4809 7420 4818 7454
rect 4818 7420 4852 7454
rect 4852 7420 4861 7454
rect 4809 7411 4861 7420
rect 3209 6244 3261 6253
rect 3209 6210 3218 6244
rect 3218 6210 3252 6244
rect 3252 6210 3261 6244
rect 3209 6201 3261 6210
rect 1809 5157 1861 5201
rect 1809 5149 1818 5157
rect 1818 5149 1852 5157
rect 1852 5149 1861 5157
rect 2009 5263 2018 5271
rect 2018 5263 2052 5271
rect 2052 5263 2061 5271
rect 2009 5219 2061 5263
rect 2209 5437 2261 5481
rect 2209 5429 2218 5437
rect 2218 5429 2252 5437
rect 2252 5429 2261 5437
rect 2409 5543 2418 5551
rect 2418 5543 2452 5551
rect 2452 5543 2461 5551
rect 2409 5499 2461 5543
rect 2609 5717 2661 5761
rect 2609 5709 2618 5717
rect 2618 5709 2652 5717
rect 2652 5709 2661 5717
rect 2809 5823 2818 5831
rect 2818 5823 2852 5831
rect 2852 5823 2861 5831
rect 2809 5779 2861 5823
rect 3009 5997 3061 6041
rect 3009 5989 3018 5997
rect 3018 5989 3052 5997
rect 3052 5989 3061 5997
rect 3209 6103 3218 6111
rect 3218 6103 3252 6111
rect 3252 6103 3261 6111
rect 3209 6059 3261 6103
rect 3409 6367 3461 6411
rect 3409 6359 3418 6367
rect 3418 6359 3452 6367
rect 3452 6359 3461 6367
rect 3609 6473 3618 6481
rect 3618 6473 3652 6481
rect 3652 6473 3661 6481
rect 3609 6429 3661 6473
rect 3809 6647 3861 6691
rect 3809 6639 3818 6647
rect 3818 6639 3852 6647
rect 3852 6639 3861 6647
rect 4009 6753 4018 6761
rect 4018 6753 4052 6761
rect 4052 6753 4061 6761
rect 4009 6709 4061 6753
rect 4209 6927 4261 6971
rect 4209 6919 4218 6927
rect 4218 6919 4252 6927
rect 4252 6919 4261 6927
rect 4409 7033 4418 7041
rect 4418 7033 4452 7041
rect 4452 7033 4461 7041
rect 4409 6989 4461 7033
rect 4609 7207 4661 7251
rect 4609 7199 4618 7207
rect 4618 7199 4652 7207
rect 4652 7199 4661 7207
rect 4809 7313 4818 7321
rect 4818 7313 4852 7321
rect 4852 7313 4861 7321
rect 4809 7269 4861 7313
rect 5009 7577 5061 7621
rect 5009 7569 5018 7577
rect 5018 7569 5052 7577
rect 5052 7569 5061 7577
rect 5209 7683 5218 7691
rect 5218 7683 5252 7691
rect 5252 7683 5261 7691
rect 5209 7639 5261 7683
rect 5409 7857 5461 7901
rect 5409 7849 5418 7857
rect 5418 7849 5452 7857
rect 5452 7849 5461 7857
rect 5609 7963 5618 7971
rect 5618 7963 5652 7971
rect 5652 7963 5661 7971
rect 5609 7919 5661 7963
rect 5809 8137 5861 8181
rect 5809 8129 5818 8137
rect 5818 8129 5852 8137
rect 5852 8129 5861 8137
rect 6009 8243 6018 8251
rect 6018 8243 6052 8251
rect 6052 8243 6061 8251
rect 6009 8199 6061 8243
rect 6209 8417 6261 8461
rect 6209 8409 6218 8417
rect 6218 8409 6252 8417
rect 6252 8409 6261 8417
rect 6409 8523 6418 8531
rect 6418 8523 6452 8531
rect 6452 8523 6461 8531
rect 6409 8479 6461 8523
rect 6507 8479 6559 8531
rect 5009 7470 5061 7479
rect 5009 7436 5018 7470
rect 5018 7436 5052 7470
rect 5052 7436 5061 7470
rect 5009 7427 5061 7436
rect 3409 6260 3461 6269
rect 3409 6226 3418 6260
rect 3418 6226 3452 6260
rect 3452 6226 3461 6260
rect 3409 6217 3461 6226
rect 2009 5123 2018 5131
rect 2018 5123 2052 5131
rect 2052 5123 2061 5131
rect 2009 5079 2061 5123
rect 2209 5297 2261 5341
rect 2209 5289 2218 5297
rect 2218 5289 2252 5297
rect 2252 5289 2261 5297
rect 2409 5403 2418 5411
rect 2418 5403 2452 5411
rect 2452 5403 2461 5411
rect 2409 5359 2461 5403
rect 2609 5577 2661 5621
rect 2609 5569 2618 5577
rect 2618 5569 2652 5577
rect 2652 5569 2661 5577
rect 2809 5683 2818 5691
rect 2818 5683 2852 5691
rect 2852 5683 2861 5691
rect 2809 5639 2861 5683
rect 3009 5857 3061 5901
rect 3009 5849 3018 5857
rect 3018 5849 3052 5857
rect 3052 5849 3061 5857
rect 3209 5963 3218 5971
rect 3218 5963 3252 5971
rect 3252 5963 3261 5971
rect 3209 5919 3261 5963
rect 3409 6137 3461 6181
rect 3409 6129 3418 6137
rect 3418 6129 3452 6137
rect 3452 6129 3461 6137
rect 3609 6333 3618 6341
rect 3618 6333 3652 6341
rect 3652 6333 3661 6341
rect 3609 6289 3661 6333
rect 3809 6507 3861 6551
rect 3809 6499 3818 6507
rect 3818 6499 3852 6507
rect 3852 6499 3861 6507
rect 4009 6613 4018 6621
rect 4018 6613 4052 6621
rect 4052 6613 4061 6621
rect 4009 6569 4061 6613
rect 4209 6787 4261 6831
rect 4209 6779 4218 6787
rect 4218 6779 4252 6787
rect 4252 6779 4261 6787
rect 4409 6893 4418 6901
rect 4418 6893 4452 6901
rect 4452 6893 4461 6901
rect 4409 6849 4461 6893
rect 4609 7067 4661 7111
rect 4609 7059 4618 7067
rect 4618 7059 4652 7067
rect 4652 7059 4661 7067
rect 4809 7173 4818 7181
rect 4818 7173 4852 7181
rect 4852 7173 4861 7181
rect 4809 7129 4861 7173
rect 5009 7347 5061 7391
rect 5009 7339 5018 7347
rect 5018 7339 5052 7347
rect 5052 7339 5061 7347
rect 5209 7543 5218 7551
rect 5218 7543 5252 7551
rect 5252 7543 5261 7551
rect 5209 7499 5261 7543
rect 5409 7717 5461 7761
rect 5409 7709 5418 7717
rect 5418 7709 5452 7717
rect 5452 7709 5461 7717
rect 5609 7823 5618 7831
rect 5618 7823 5652 7831
rect 5652 7823 5661 7831
rect 5609 7779 5661 7823
rect 5809 7997 5861 8041
rect 5809 7989 5818 7997
rect 5818 7989 5852 7997
rect 5852 7989 5861 7997
rect 6009 8103 6018 8111
rect 6018 8103 6052 8111
rect 6052 8103 6061 8111
rect 6009 8059 6061 8103
rect 6209 8277 6261 8321
rect 6209 8269 6218 8277
rect 6218 8269 6252 8277
rect 6252 8269 6261 8277
rect 6409 8383 6418 8391
rect 6418 8383 6452 8391
rect 6452 8383 6461 8391
rect 6409 8339 6461 8383
rect 6507 8339 6559 8391
rect 5209 7454 5261 7463
rect 5209 7420 5218 7454
rect 5218 7420 5252 7454
rect 5252 7420 5261 7454
rect 5209 7411 5261 7420
rect 3609 6244 3661 6253
rect 3609 6210 3618 6244
rect 3618 6210 3652 6244
rect 3652 6210 3661 6244
rect 3609 6201 3661 6210
rect 2209 5157 2261 5201
rect 2209 5149 2218 5157
rect 2218 5149 2252 5157
rect 2252 5149 2261 5157
rect 2409 5263 2418 5271
rect 2418 5263 2452 5271
rect 2452 5263 2461 5271
rect 2409 5219 2461 5263
rect 2609 5437 2661 5481
rect 2609 5429 2618 5437
rect 2618 5429 2652 5437
rect 2652 5429 2661 5437
rect 2809 5543 2818 5551
rect 2818 5543 2852 5551
rect 2852 5543 2861 5551
rect 2809 5499 2861 5543
rect 3009 5717 3061 5761
rect 3009 5709 3018 5717
rect 3018 5709 3052 5717
rect 3052 5709 3061 5717
rect 3209 5823 3218 5831
rect 3218 5823 3252 5831
rect 3252 5823 3261 5831
rect 3209 5779 3261 5823
rect 3409 5997 3461 6041
rect 3409 5989 3418 5997
rect 3418 5989 3452 5997
rect 3452 5989 3461 5997
rect 3609 6103 3618 6111
rect 3618 6103 3652 6111
rect 3652 6103 3661 6111
rect 3609 6059 3661 6103
rect 3809 6367 3861 6411
rect 3809 6359 3818 6367
rect 3818 6359 3852 6367
rect 3852 6359 3861 6367
rect 4009 6473 4018 6481
rect 4018 6473 4052 6481
rect 4052 6473 4061 6481
rect 4009 6429 4061 6473
rect 4209 6647 4261 6691
rect 4209 6639 4218 6647
rect 4218 6639 4252 6647
rect 4252 6639 4261 6647
rect 4409 6753 4418 6761
rect 4418 6753 4452 6761
rect 4452 6753 4461 6761
rect 4409 6709 4461 6753
rect 4609 6927 4661 6971
rect 4609 6919 4618 6927
rect 4618 6919 4652 6927
rect 4652 6919 4661 6927
rect 4809 7033 4818 7041
rect 4818 7033 4852 7041
rect 4852 7033 4861 7041
rect 4809 6989 4861 7033
rect 5009 7207 5061 7251
rect 5009 7199 5018 7207
rect 5018 7199 5052 7207
rect 5052 7199 5061 7207
rect 5209 7313 5218 7321
rect 5218 7313 5252 7321
rect 5252 7313 5261 7321
rect 5209 7269 5261 7313
rect 5409 7577 5461 7621
rect 5409 7569 5418 7577
rect 5418 7569 5452 7577
rect 5452 7569 5461 7577
rect 5609 7683 5618 7691
rect 5618 7683 5652 7691
rect 5652 7683 5661 7691
rect 5609 7639 5661 7683
rect 5809 7857 5861 7901
rect 5809 7849 5818 7857
rect 5818 7849 5852 7857
rect 5852 7849 5861 7857
rect 6009 7963 6018 7971
rect 6018 7963 6052 7971
rect 6052 7963 6061 7971
rect 6009 7919 6061 7963
rect 6209 8137 6261 8181
rect 6209 8129 6218 8137
rect 6218 8129 6252 8137
rect 6252 8129 6261 8137
rect 6409 8243 6418 8251
rect 6418 8243 6452 8251
rect 6452 8243 6461 8251
rect 6409 8199 6461 8243
rect 6507 8199 6559 8251
rect 5409 7470 5461 7479
rect 5409 7436 5418 7470
rect 5418 7436 5452 7470
rect 5452 7436 5461 7470
rect 5409 7427 5461 7436
rect 3809 6260 3861 6269
rect 3809 6226 3818 6260
rect 3818 6226 3852 6260
rect 3852 6226 3861 6260
rect 3809 6217 3861 6226
rect 2409 5123 2418 5131
rect 2418 5123 2452 5131
rect 2452 5123 2461 5131
rect 2409 5079 2461 5123
rect 2609 5297 2661 5341
rect 2609 5289 2618 5297
rect 2618 5289 2652 5297
rect 2652 5289 2661 5297
rect 2809 5403 2818 5411
rect 2818 5403 2852 5411
rect 2852 5403 2861 5411
rect 2809 5359 2861 5403
rect 3009 5577 3061 5621
rect 3009 5569 3018 5577
rect 3018 5569 3052 5577
rect 3052 5569 3061 5577
rect 3209 5683 3218 5691
rect 3218 5683 3252 5691
rect 3252 5683 3261 5691
rect 3209 5639 3261 5683
rect 3409 5857 3461 5901
rect 3409 5849 3418 5857
rect 3418 5849 3452 5857
rect 3452 5849 3461 5857
rect 3609 5963 3618 5971
rect 3618 5963 3652 5971
rect 3652 5963 3661 5971
rect 3609 5919 3661 5963
rect 3809 6137 3861 6181
rect 3809 6129 3818 6137
rect 3818 6129 3852 6137
rect 3852 6129 3861 6137
rect 4009 6333 4018 6341
rect 4018 6333 4052 6341
rect 4052 6333 4061 6341
rect 4009 6289 4061 6333
rect 4209 6507 4261 6551
rect 4209 6499 4218 6507
rect 4218 6499 4252 6507
rect 4252 6499 4261 6507
rect 4409 6613 4418 6621
rect 4418 6613 4452 6621
rect 4452 6613 4461 6621
rect 4409 6569 4461 6613
rect 4609 6787 4661 6831
rect 4609 6779 4618 6787
rect 4618 6779 4652 6787
rect 4652 6779 4661 6787
rect 4809 6893 4818 6901
rect 4818 6893 4852 6901
rect 4852 6893 4861 6901
rect 4809 6849 4861 6893
rect 5009 7067 5061 7111
rect 5009 7059 5018 7067
rect 5018 7059 5052 7067
rect 5052 7059 5061 7067
rect 5209 7173 5218 7181
rect 5218 7173 5252 7181
rect 5252 7173 5261 7181
rect 5209 7129 5261 7173
rect 5409 7347 5461 7391
rect 5409 7339 5418 7347
rect 5418 7339 5452 7347
rect 5452 7339 5461 7347
rect 5609 7543 5618 7551
rect 5618 7543 5652 7551
rect 5652 7543 5661 7551
rect 5609 7499 5661 7543
rect 5809 7717 5861 7761
rect 5809 7709 5818 7717
rect 5818 7709 5852 7717
rect 5852 7709 5861 7717
rect 6009 7823 6018 7831
rect 6018 7823 6052 7831
rect 6052 7823 6061 7831
rect 6009 7779 6061 7823
rect 6209 7997 6261 8041
rect 6209 7989 6218 7997
rect 6218 7989 6252 7997
rect 6252 7989 6261 7997
rect 6409 8103 6418 8111
rect 6418 8103 6452 8111
rect 6452 8103 6461 8111
rect 6409 8059 6461 8103
rect 6507 8059 6559 8111
rect 5609 7454 5661 7463
rect 5609 7420 5618 7454
rect 5618 7420 5652 7454
rect 5652 7420 5661 7454
rect 5609 7411 5661 7420
rect 4009 6244 4061 6253
rect 4009 6210 4018 6244
rect 4018 6210 4052 6244
rect 4052 6210 4061 6244
rect 4009 6201 4061 6210
rect 2609 5157 2661 5201
rect 2609 5149 2618 5157
rect 2618 5149 2652 5157
rect 2652 5149 2661 5157
rect 2809 5263 2818 5271
rect 2818 5263 2852 5271
rect 2852 5263 2861 5271
rect 2809 5219 2861 5263
rect 3009 5437 3061 5481
rect 3009 5429 3018 5437
rect 3018 5429 3052 5437
rect 3052 5429 3061 5437
rect 3209 5543 3218 5551
rect 3218 5543 3252 5551
rect 3252 5543 3261 5551
rect 3209 5499 3261 5543
rect 3409 5717 3461 5761
rect 3409 5709 3418 5717
rect 3418 5709 3452 5717
rect 3452 5709 3461 5717
rect 3609 5823 3618 5831
rect 3618 5823 3652 5831
rect 3652 5823 3661 5831
rect 3609 5779 3661 5823
rect 3809 5997 3861 6041
rect 3809 5989 3818 5997
rect 3818 5989 3852 5997
rect 3852 5989 3861 5997
rect 4009 6103 4018 6111
rect 4018 6103 4052 6111
rect 4052 6103 4061 6111
rect 4009 6059 4061 6103
rect 4209 6367 4261 6411
rect 4209 6359 4218 6367
rect 4218 6359 4252 6367
rect 4252 6359 4261 6367
rect 4409 6473 4418 6481
rect 4418 6473 4452 6481
rect 4452 6473 4461 6481
rect 4409 6429 4461 6473
rect 4609 6647 4661 6691
rect 4609 6639 4618 6647
rect 4618 6639 4652 6647
rect 4652 6639 4661 6647
rect 4809 6753 4818 6761
rect 4818 6753 4852 6761
rect 4852 6753 4861 6761
rect 4809 6709 4861 6753
rect 5009 6927 5061 6971
rect 5009 6919 5018 6927
rect 5018 6919 5052 6927
rect 5052 6919 5061 6927
rect 5209 7033 5218 7041
rect 5218 7033 5252 7041
rect 5252 7033 5261 7041
rect 5209 6989 5261 7033
rect 5409 7207 5461 7251
rect 5409 7199 5418 7207
rect 5418 7199 5452 7207
rect 5452 7199 5461 7207
rect 5609 7313 5618 7321
rect 5618 7313 5652 7321
rect 5652 7313 5661 7321
rect 5609 7269 5661 7313
rect 5809 7577 5861 7621
rect 5809 7569 5818 7577
rect 5818 7569 5852 7577
rect 5852 7569 5861 7577
rect 6009 7683 6018 7691
rect 6018 7683 6052 7691
rect 6052 7683 6061 7691
rect 6009 7639 6061 7683
rect 6209 7857 6261 7901
rect 6209 7849 6218 7857
rect 6218 7849 6252 7857
rect 6252 7849 6261 7857
rect 6409 7963 6418 7971
rect 6418 7963 6452 7971
rect 6452 7963 6461 7971
rect 6409 7919 6461 7963
rect 6507 7919 6559 7971
rect 5809 7470 5861 7479
rect 5809 7436 5818 7470
rect 5818 7436 5852 7470
rect 5852 7436 5861 7470
rect 5809 7427 5861 7436
rect 4209 6260 4261 6269
rect 4209 6226 4218 6260
rect 4218 6226 4252 6260
rect 4252 6226 4261 6260
rect 4209 6217 4261 6226
rect 2809 5123 2818 5131
rect 2818 5123 2852 5131
rect 2852 5123 2861 5131
rect 2809 5079 2861 5123
rect 3009 5297 3061 5341
rect 3009 5289 3018 5297
rect 3018 5289 3052 5297
rect 3052 5289 3061 5297
rect 3209 5403 3218 5411
rect 3218 5403 3252 5411
rect 3252 5403 3261 5411
rect 3209 5359 3261 5403
rect 3409 5577 3461 5621
rect 3409 5569 3418 5577
rect 3418 5569 3452 5577
rect 3452 5569 3461 5577
rect 3609 5683 3618 5691
rect 3618 5683 3652 5691
rect 3652 5683 3661 5691
rect 3609 5639 3661 5683
rect 3809 5857 3861 5901
rect 3809 5849 3818 5857
rect 3818 5849 3852 5857
rect 3852 5849 3861 5857
rect 4009 5963 4018 5971
rect 4018 5963 4052 5971
rect 4052 5963 4061 5971
rect 4009 5919 4061 5963
rect 4209 6137 4261 6181
rect 4209 6129 4218 6137
rect 4218 6129 4252 6137
rect 4252 6129 4261 6137
rect 4409 6333 4418 6341
rect 4418 6333 4452 6341
rect 4452 6333 4461 6341
rect 4409 6289 4461 6333
rect 4609 6507 4661 6551
rect 4609 6499 4618 6507
rect 4618 6499 4652 6507
rect 4652 6499 4661 6507
rect 4809 6613 4818 6621
rect 4818 6613 4852 6621
rect 4852 6613 4861 6621
rect 4809 6569 4861 6613
rect 5009 6787 5061 6831
rect 5009 6779 5018 6787
rect 5018 6779 5052 6787
rect 5052 6779 5061 6787
rect 5209 6893 5218 6901
rect 5218 6893 5252 6901
rect 5252 6893 5261 6901
rect 5209 6849 5261 6893
rect 5409 7067 5461 7111
rect 5409 7059 5418 7067
rect 5418 7059 5452 7067
rect 5452 7059 5461 7067
rect 5609 7173 5618 7181
rect 5618 7173 5652 7181
rect 5652 7173 5661 7181
rect 5609 7129 5661 7173
rect 5809 7347 5861 7391
rect 5809 7339 5818 7347
rect 5818 7339 5852 7347
rect 5852 7339 5861 7347
rect 6009 7543 6018 7551
rect 6018 7543 6052 7551
rect 6052 7543 6061 7551
rect 6009 7499 6061 7543
rect 6209 7717 6261 7761
rect 6209 7709 6218 7717
rect 6218 7709 6252 7717
rect 6252 7709 6261 7717
rect 6409 7823 6418 7831
rect 6418 7823 6452 7831
rect 6452 7823 6461 7831
rect 6409 7779 6461 7823
rect 6507 7779 6559 7831
rect 6009 7454 6061 7463
rect 6009 7420 6018 7454
rect 6018 7420 6052 7454
rect 6052 7420 6061 7454
rect 6009 7411 6061 7420
rect 4409 6244 4461 6253
rect 4409 6210 4418 6244
rect 4418 6210 4452 6244
rect 4452 6210 4461 6244
rect 4409 6201 4461 6210
rect 3009 5157 3061 5201
rect 3009 5149 3018 5157
rect 3018 5149 3052 5157
rect 3052 5149 3061 5157
rect 3209 5263 3218 5271
rect 3218 5263 3252 5271
rect 3252 5263 3261 5271
rect 3209 5219 3261 5263
rect 3409 5437 3461 5481
rect 3409 5429 3418 5437
rect 3418 5429 3452 5437
rect 3452 5429 3461 5437
rect 3609 5543 3618 5551
rect 3618 5543 3652 5551
rect 3652 5543 3661 5551
rect 3609 5499 3661 5543
rect 3809 5717 3861 5761
rect 3809 5709 3818 5717
rect 3818 5709 3852 5717
rect 3852 5709 3861 5717
rect 4009 5823 4018 5831
rect 4018 5823 4052 5831
rect 4052 5823 4061 5831
rect 4009 5779 4061 5823
rect 4209 5997 4261 6041
rect 4209 5989 4218 5997
rect 4218 5989 4252 5997
rect 4252 5989 4261 5997
rect 4409 6103 4418 6111
rect 4418 6103 4452 6111
rect 4452 6103 4461 6111
rect 4409 6059 4461 6103
rect 4609 6367 4661 6411
rect 4609 6359 4618 6367
rect 4618 6359 4652 6367
rect 4652 6359 4661 6367
rect 4809 6473 4818 6481
rect 4818 6473 4852 6481
rect 4852 6473 4861 6481
rect 4809 6429 4861 6473
rect 5009 6647 5061 6691
rect 5009 6639 5018 6647
rect 5018 6639 5052 6647
rect 5052 6639 5061 6647
rect 5209 6753 5218 6761
rect 5218 6753 5252 6761
rect 5252 6753 5261 6761
rect 5209 6709 5261 6753
rect 5409 6927 5461 6971
rect 5409 6919 5418 6927
rect 5418 6919 5452 6927
rect 5452 6919 5461 6927
rect 5609 7033 5618 7041
rect 5618 7033 5652 7041
rect 5652 7033 5661 7041
rect 5609 6989 5661 7033
rect 5809 7207 5861 7251
rect 5809 7199 5818 7207
rect 5818 7199 5852 7207
rect 5852 7199 5861 7207
rect 6009 7313 6018 7321
rect 6018 7313 6052 7321
rect 6052 7313 6061 7321
rect 6009 7269 6061 7313
rect 6209 7577 6261 7621
rect 6209 7569 6218 7577
rect 6218 7569 6252 7577
rect 6252 7569 6261 7577
rect 6409 7683 6418 7691
rect 6418 7683 6452 7691
rect 6452 7683 6461 7691
rect 6409 7639 6461 7683
rect 6507 7639 6559 7691
rect 6209 7470 6261 7479
rect 6209 7436 6218 7470
rect 6218 7436 6252 7470
rect 6252 7436 6261 7470
rect 6209 7427 6261 7436
rect 4609 6260 4661 6269
rect 4609 6226 4618 6260
rect 4618 6226 4652 6260
rect 4652 6226 4661 6260
rect 4609 6217 4661 6226
rect 3209 5123 3218 5131
rect 3218 5123 3252 5131
rect 3252 5123 3261 5131
rect 3209 5079 3261 5123
rect 3409 5297 3461 5341
rect 3409 5289 3418 5297
rect 3418 5289 3452 5297
rect 3452 5289 3461 5297
rect 3609 5403 3618 5411
rect 3618 5403 3652 5411
rect 3652 5403 3661 5411
rect 3609 5359 3661 5403
rect 3809 5577 3861 5621
rect 3809 5569 3818 5577
rect 3818 5569 3852 5577
rect 3852 5569 3861 5577
rect 4009 5683 4018 5691
rect 4018 5683 4052 5691
rect 4052 5683 4061 5691
rect 4009 5639 4061 5683
rect 4209 5857 4261 5901
rect 4209 5849 4218 5857
rect 4218 5849 4252 5857
rect 4252 5849 4261 5857
rect 4409 5963 4418 5971
rect 4418 5963 4452 5971
rect 4452 5963 4461 5971
rect 4409 5919 4461 5963
rect 4609 6137 4661 6181
rect 4609 6129 4618 6137
rect 4618 6129 4652 6137
rect 4652 6129 4661 6137
rect 4809 6333 4818 6341
rect 4818 6333 4852 6341
rect 4852 6333 4861 6341
rect 4809 6289 4861 6333
rect 5009 6507 5061 6551
rect 5009 6499 5018 6507
rect 5018 6499 5052 6507
rect 5052 6499 5061 6507
rect 5209 6613 5218 6621
rect 5218 6613 5252 6621
rect 5252 6613 5261 6621
rect 5209 6569 5261 6613
rect 5409 6787 5461 6831
rect 5409 6779 5418 6787
rect 5418 6779 5452 6787
rect 5452 6779 5461 6787
rect 5609 6893 5618 6901
rect 5618 6893 5652 6901
rect 5652 6893 5661 6901
rect 5609 6849 5661 6893
rect 5809 7067 5861 7111
rect 5809 7059 5818 7067
rect 5818 7059 5852 7067
rect 5852 7059 5861 7067
rect 6009 7173 6018 7181
rect 6018 7173 6052 7181
rect 6052 7173 6061 7181
rect 6009 7129 6061 7173
rect 6209 7347 6261 7391
rect 6209 7339 6218 7347
rect 6218 7339 6252 7347
rect 6252 7339 6261 7347
rect 6409 7543 6418 7551
rect 6418 7543 6452 7551
rect 6452 7543 6461 7551
rect 6409 7499 6461 7543
rect 6507 7499 6559 7551
rect 4809 6244 4861 6253
rect 4809 6210 4818 6244
rect 4818 6210 4852 6244
rect 4852 6210 4861 6244
rect 4809 6201 4861 6210
rect 3409 5157 3461 5201
rect 3409 5149 3418 5157
rect 3418 5149 3452 5157
rect 3452 5149 3461 5157
rect 3609 5263 3618 5271
rect 3618 5263 3652 5271
rect 3652 5263 3661 5271
rect 3609 5219 3661 5263
rect 3809 5437 3861 5481
rect 3809 5429 3818 5437
rect 3818 5429 3852 5437
rect 3852 5429 3861 5437
rect 4009 5543 4018 5551
rect 4018 5543 4052 5551
rect 4052 5543 4061 5551
rect 4009 5499 4061 5543
rect 4209 5717 4261 5761
rect 4209 5709 4218 5717
rect 4218 5709 4252 5717
rect 4252 5709 4261 5717
rect 4409 5823 4418 5831
rect 4418 5823 4452 5831
rect 4452 5823 4461 5831
rect 4409 5779 4461 5823
rect 4609 5997 4661 6041
rect 4609 5989 4618 5997
rect 4618 5989 4652 5997
rect 4652 5989 4661 5997
rect 4809 6103 4818 6111
rect 4818 6103 4852 6111
rect 4852 6103 4861 6111
rect 4809 6059 4861 6103
rect 5009 6367 5061 6411
rect 5009 6359 5018 6367
rect 5018 6359 5052 6367
rect 5052 6359 5061 6367
rect 5209 6473 5218 6481
rect 5218 6473 5252 6481
rect 5252 6473 5261 6481
rect 5209 6429 5261 6473
rect 5409 6647 5461 6691
rect 5409 6639 5418 6647
rect 5418 6639 5452 6647
rect 5452 6639 5461 6647
rect 5609 6753 5618 6761
rect 5618 6753 5652 6761
rect 5652 6753 5661 6761
rect 5609 6709 5661 6753
rect 5809 6927 5861 6971
rect 5809 6919 5818 6927
rect 5818 6919 5852 6927
rect 5852 6919 5861 6927
rect 6009 7033 6018 7041
rect 6018 7033 6052 7041
rect 6052 7033 6061 7041
rect 6009 6989 6061 7033
rect 6209 7207 6261 7251
rect 6209 7199 6218 7207
rect 6218 7199 6252 7207
rect 6252 7199 6261 7207
rect 6409 7313 6418 7321
rect 6418 7313 6452 7321
rect 6452 7313 6461 7321
rect 6409 7269 6461 7313
rect 6507 7269 6559 7321
rect 5009 6260 5061 6269
rect 5009 6226 5018 6260
rect 5018 6226 5052 6260
rect 5052 6226 5061 6260
rect 5009 6217 5061 6226
rect 3609 5123 3618 5131
rect 3618 5123 3652 5131
rect 3652 5123 3661 5131
rect 3609 5079 3661 5123
rect 3809 5297 3861 5341
rect 3809 5289 3818 5297
rect 3818 5289 3852 5297
rect 3852 5289 3861 5297
rect 4009 5403 4018 5411
rect 4018 5403 4052 5411
rect 4052 5403 4061 5411
rect 4009 5359 4061 5403
rect 4209 5577 4261 5621
rect 4209 5569 4218 5577
rect 4218 5569 4252 5577
rect 4252 5569 4261 5577
rect 4409 5683 4418 5691
rect 4418 5683 4452 5691
rect 4452 5683 4461 5691
rect 4409 5639 4461 5683
rect 4609 5857 4661 5901
rect 4609 5849 4618 5857
rect 4618 5849 4652 5857
rect 4652 5849 4661 5857
rect 4809 5963 4818 5971
rect 4818 5963 4852 5971
rect 4852 5963 4861 5971
rect 4809 5919 4861 5963
rect 5009 6137 5061 6181
rect 5009 6129 5018 6137
rect 5018 6129 5052 6137
rect 5052 6129 5061 6137
rect 5209 6333 5218 6341
rect 5218 6333 5252 6341
rect 5252 6333 5261 6341
rect 5209 6289 5261 6333
rect 5409 6507 5461 6551
rect 5409 6499 5418 6507
rect 5418 6499 5452 6507
rect 5452 6499 5461 6507
rect 5609 6613 5618 6621
rect 5618 6613 5652 6621
rect 5652 6613 5661 6621
rect 5609 6569 5661 6613
rect 5809 6787 5861 6831
rect 5809 6779 5818 6787
rect 5818 6779 5852 6787
rect 5852 6779 5861 6787
rect 6009 6893 6018 6901
rect 6018 6893 6052 6901
rect 6052 6893 6061 6901
rect 6009 6849 6061 6893
rect 6209 7067 6261 7111
rect 6209 7059 6218 7067
rect 6218 7059 6252 7067
rect 6252 7059 6261 7067
rect 6409 7173 6418 7181
rect 6418 7173 6452 7181
rect 6452 7173 6461 7181
rect 6409 7129 6461 7173
rect 6507 7129 6559 7181
rect 5209 6244 5261 6253
rect 5209 6210 5218 6244
rect 5218 6210 5252 6244
rect 5252 6210 5261 6244
rect 5209 6201 5261 6210
rect 3809 5157 3861 5201
rect 3809 5149 3818 5157
rect 3818 5149 3852 5157
rect 3852 5149 3861 5157
rect 4009 5263 4018 5271
rect 4018 5263 4052 5271
rect 4052 5263 4061 5271
rect 4009 5219 4061 5263
rect 4209 5437 4261 5481
rect 4209 5429 4218 5437
rect 4218 5429 4252 5437
rect 4252 5429 4261 5437
rect 4409 5543 4418 5551
rect 4418 5543 4452 5551
rect 4452 5543 4461 5551
rect 4409 5499 4461 5543
rect 4609 5717 4661 5761
rect 4609 5709 4618 5717
rect 4618 5709 4652 5717
rect 4652 5709 4661 5717
rect 4809 5823 4818 5831
rect 4818 5823 4852 5831
rect 4852 5823 4861 5831
rect 4809 5779 4861 5823
rect 5009 5997 5061 6041
rect 5009 5989 5018 5997
rect 5018 5989 5052 5997
rect 5052 5989 5061 5997
rect 5209 6103 5218 6111
rect 5218 6103 5252 6111
rect 5252 6103 5261 6111
rect 5209 6059 5261 6103
rect 5409 6367 5461 6411
rect 5409 6359 5418 6367
rect 5418 6359 5452 6367
rect 5452 6359 5461 6367
rect 5609 6473 5618 6481
rect 5618 6473 5652 6481
rect 5652 6473 5661 6481
rect 5609 6429 5661 6473
rect 5809 6647 5861 6691
rect 5809 6639 5818 6647
rect 5818 6639 5852 6647
rect 5852 6639 5861 6647
rect 6009 6753 6018 6761
rect 6018 6753 6052 6761
rect 6052 6753 6061 6761
rect 6009 6709 6061 6753
rect 6209 6927 6261 6971
rect 6209 6919 6218 6927
rect 6218 6919 6252 6927
rect 6252 6919 6261 6927
rect 6409 7033 6418 7041
rect 6418 7033 6452 7041
rect 6452 7033 6461 7041
rect 6409 6989 6461 7033
rect 6507 6989 6559 7041
rect 5409 6260 5461 6269
rect 5409 6226 5418 6260
rect 5418 6226 5452 6260
rect 5452 6226 5461 6260
rect 5409 6217 5461 6226
rect 4009 5123 4018 5131
rect 4018 5123 4052 5131
rect 4052 5123 4061 5131
rect 4009 5079 4061 5123
rect 4209 5297 4261 5341
rect 4209 5289 4218 5297
rect 4218 5289 4252 5297
rect 4252 5289 4261 5297
rect 4409 5403 4418 5411
rect 4418 5403 4452 5411
rect 4452 5403 4461 5411
rect 4409 5359 4461 5403
rect 4609 5577 4661 5621
rect 4609 5569 4618 5577
rect 4618 5569 4652 5577
rect 4652 5569 4661 5577
rect 4809 5683 4818 5691
rect 4818 5683 4852 5691
rect 4852 5683 4861 5691
rect 4809 5639 4861 5683
rect 5009 5857 5061 5901
rect 5009 5849 5018 5857
rect 5018 5849 5052 5857
rect 5052 5849 5061 5857
rect 5209 5963 5218 5971
rect 5218 5963 5252 5971
rect 5252 5963 5261 5971
rect 5209 5919 5261 5963
rect 5409 6137 5461 6181
rect 5409 6129 5418 6137
rect 5418 6129 5452 6137
rect 5452 6129 5461 6137
rect 5609 6333 5618 6341
rect 5618 6333 5652 6341
rect 5652 6333 5661 6341
rect 5609 6289 5661 6333
rect 5809 6507 5861 6551
rect 5809 6499 5818 6507
rect 5818 6499 5852 6507
rect 5852 6499 5861 6507
rect 6009 6613 6018 6621
rect 6018 6613 6052 6621
rect 6052 6613 6061 6621
rect 6009 6569 6061 6613
rect 6209 6787 6261 6831
rect 6209 6779 6218 6787
rect 6218 6779 6252 6787
rect 6252 6779 6261 6787
rect 6409 6893 6418 6901
rect 6418 6893 6452 6901
rect 6452 6893 6461 6901
rect 6409 6849 6461 6893
rect 6507 6849 6559 6901
rect 5609 6244 5661 6253
rect 5609 6210 5618 6244
rect 5618 6210 5652 6244
rect 5652 6210 5661 6244
rect 5609 6201 5661 6210
rect 4209 5157 4261 5201
rect 4209 5149 4218 5157
rect 4218 5149 4252 5157
rect 4252 5149 4261 5157
rect 4409 5263 4418 5271
rect 4418 5263 4452 5271
rect 4452 5263 4461 5271
rect 4409 5219 4461 5263
rect 4609 5437 4661 5481
rect 4609 5429 4618 5437
rect 4618 5429 4652 5437
rect 4652 5429 4661 5437
rect 4809 5543 4818 5551
rect 4818 5543 4852 5551
rect 4852 5543 4861 5551
rect 4809 5499 4861 5543
rect 5009 5717 5061 5761
rect 5009 5709 5018 5717
rect 5018 5709 5052 5717
rect 5052 5709 5061 5717
rect 5209 5823 5218 5831
rect 5218 5823 5252 5831
rect 5252 5823 5261 5831
rect 5209 5779 5261 5823
rect 5409 5997 5461 6041
rect 5409 5989 5418 5997
rect 5418 5989 5452 5997
rect 5452 5989 5461 5997
rect 5609 6103 5618 6111
rect 5618 6103 5652 6111
rect 5652 6103 5661 6111
rect 5609 6059 5661 6103
rect 5809 6367 5861 6411
rect 5809 6359 5818 6367
rect 5818 6359 5852 6367
rect 5852 6359 5861 6367
rect 6009 6473 6018 6481
rect 6018 6473 6052 6481
rect 6052 6473 6061 6481
rect 6009 6429 6061 6473
rect 6209 6647 6261 6691
rect 6209 6639 6218 6647
rect 6218 6639 6252 6647
rect 6252 6639 6261 6647
rect 6409 6753 6418 6761
rect 6418 6753 6452 6761
rect 6452 6753 6461 6761
rect 6409 6709 6461 6753
rect 6507 6709 6559 6761
rect 5809 6260 5861 6269
rect 5809 6226 5818 6260
rect 5818 6226 5852 6260
rect 5852 6226 5861 6260
rect 5809 6217 5861 6226
rect 4409 5123 4418 5131
rect 4418 5123 4452 5131
rect 4452 5123 4461 5131
rect 4409 5079 4461 5123
rect 4609 5297 4661 5341
rect 4609 5289 4618 5297
rect 4618 5289 4652 5297
rect 4652 5289 4661 5297
rect 4809 5403 4818 5411
rect 4818 5403 4852 5411
rect 4852 5403 4861 5411
rect 4809 5359 4861 5403
rect 5009 5577 5061 5621
rect 5009 5569 5018 5577
rect 5018 5569 5052 5577
rect 5052 5569 5061 5577
rect 5209 5683 5218 5691
rect 5218 5683 5252 5691
rect 5252 5683 5261 5691
rect 5209 5639 5261 5683
rect 5409 5857 5461 5901
rect 5409 5849 5418 5857
rect 5418 5849 5452 5857
rect 5452 5849 5461 5857
rect 5609 5963 5618 5971
rect 5618 5963 5652 5971
rect 5652 5963 5661 5971
rect 5609 5919 5661 5963
rect 5809 6137 5861 6181
rect 5809 6129 5818 6137
rect 5818 6129 5852 6137
rect 5852 6129 5861 6137
rect 6009 6333 6018 6341
rect 6018 6333 6052 6341
rect 6052 6333 6061 6341
rect 6009 6289 6061 6333
rect 6209 6507 6261 6551
rect 6209 6499 6218 6507
rect 6218 6499 6252 6507
rect 6252 6499 6261 6507
rect 6409 6613 6418 6621
rect 6418 6613 6452 6621
rect 6452 6613 6461 6621
rect 6409 6569 6461 6613
rect 6507 6569 6559 6621
rect 6009 6244 6061 6253
rect 6009 6210 6018 6244
rect 6018 6210 6052 6244
rect 6052 6210 6061 6244
rect 6009 6201 6061 6210
rect 4609 5157 4661 5201
rect 4609 5149 4618 5157
rect 4618 5149 4652 5157
rect 4652 5149 4661 5157
rect 4809 5263 4818 5271
rect 4818 5263 4852 5271
rect 4852 5263 4861 5271
rect 4809 5219 4861 5263
rect 5009 5437 5061 5481
rect 5009 5429 5018 5437
rect 5018 5429 5052 5437
rect 5052 5429 5061 5437
rect 5209 5543 5218 5551
rect 5218 5543 5252 5551
rect 5252 5543 5261 5551
rect 5209 5499 5261 5543
rect 5409 5717 5461 5761
rect 5409 5709 5418 5717
rect 5418 5709 5452 5717
rect 5452 5709 5461 5717
rect 5609 5823 5618 5831
rect 5618 5823 5652 5831
rect 5652 5823 5661 5831
rect 5609 5779 5661 5823
rect 5809 5997 5861 6041
rect 5809 5989 5818 5997
rect 5818 5989 5852 5997
rect 5852 5989 5861 5997
rect 6009 6103 6018 6111
rect 6018 6103 6052 6111
rect 6052 6103 6061 6111
rect 6009 6059 6061 6103
rect 6209 6367 6261 6411
rect 6209 6359 6218 6367
rect 6218 6359 6252 6367
rect 6252 6359 6261 6367
rect 6409 6473 6418 6481
rect 6418 6473 6452 6481
rect 6452 6473 6461 6481
rect 6409 6429 6461 6473
rect 6507 6429 6559 6481
rect 6209 6260 6261 6269
rect 6209 6226 6218 6260
rect 6218 6226 6252 6260
rect 6252 6226 6261 6260
rect 6209 6217 6261 6226
rect 4809 5123 4818 5131
rect 4818 5123 4852 5131
rect 4852 5123 4861 5131
rect 4809 5079 4861 5123
rect 5009 5297 5061 5341
rect 5009 5289 5018 5297
rect 5018 5289 5052 5297
rect 5052 5289 5061 5297
rect 5209 5403 5218 5411
rect 5218 5403 5252 5411
rect 5252 5403 5261 5411
rect 5209 5359 5261 5403
rect 5409 5577 5461 5621
rect 5409 5569 5418 5577
rect 5418 5569 5452 5577
rect 5452 5569 5461 5577
rect 5609 5683 5618 5691
rect 5618 5683 5652 5691
rect 5652 5683 5661 5691
rect 5609 5639 5661 5683
rect 5809 5857 5861 5901
rect 5809 5849 5818 5857
rect 5818 5849 5852 5857
rect 5852 5849 5861 5857
rect 6009 5963 6018 5971
rect 6018 5963 6052 5971
rect 6052 5963 6061 5971
rect 6009 5919 6061 5963
rect 6209 6137 6261 6181
rect 6209 6129 6218 6137
rect 6218 6129 6252 6137
rect 6252 6129 6261 6137
rect 6409 6333 6418 6341
rect 6418 6333 6452 6341
rect 6452 6333 6461 6341
rect 6409 6289 6461 6333
rect 6507 6289 6559 6341
rect 5009 5157 5061 5201
rect 5009 5149 5018 5157
rect 5018 5149 5052 5157
rect 5052 5149 5061 5157
rect 5209 5263 5218 5271
rect 5218 5263 5252 5271
rect 5252 5263 5261 5271
rect 5209 5219 5261 5263
rect 5409 5437 5461 5481
rect 5409 5429 5418 5437
rect 5418 5429 5452 5437
rect 5452 5429 5461 5437
rect 5609 5543 5618 5551
rect 5618 5543 5652 5551
rect 5652 5543 5661 5551
rect 5609 5499 5661 5543
rect 5809 5717 5861 5761
rect 5809 5709 5818 5717
rect 5818 5709 5852 5717
rect 5852 5709 5861 5717
rect 6009 5823 6018 5831
rect 6018 5823 6052 5831
rect 6052 5823 6061 5831
rect 6009 5779 6061 5823
rect 6209 5997 6261 6041
rect 6209 5989 6218 5997
rect 6218 5989 6252 5997
rect 6252 5989 6261 5997
rect 6409 6103 6418 6111
rect 6418 6103 6452 6111
rect 6452 6103 6461 6111
rect 6409 6059 6461 6103
rect 6507 6059 6559 6111
rect 5209 5123 5218 5131
rect 5218 5123 5252 5131
rect 5252 5123 5261 5131
rect 5209 5079 5261 5123
rect 5409 5297 5461 5341
rect 5409 5289 5418 5297
rect 5418 5289 5452 5297
rect 5452 5289 5461 5297
rect 5609 5403 5618 5411
rect 5618 5403 5652 5411
rect 5652 5403 5661 5411
rect 5609 5359 5661 5403
rect 5809 5577 5861 5621
rect 5809 5569 5818 5577
rect 5818 5569 5852 5577
rect 5852 5569 5861 5577
rect 6009 5683 6018 5691
rect 6018 5683 6052 5691
rect 6052 5683 6061 5691
rect 6009 5639 6061 5683
rect 6209 5857 6261 5901
rect 6209 5849 6218 5857
rect 6218 5849 6252 5857
rect 6252 5849 6261 5857
rect 6409 5963 6418 5971
rect 6418 5963 6452 5971
rect 6452 5963 6461 5971
rect 6409 5919 6461 5963
rect 6507 5919 6559 5971
rect 5409 5157 5461 5201
rect 5409 5149 5418 5157
rect 5418 5149 5452 5157
rect 5452 5149 5461 5157
rect 5609 5263 5618 5271
rect 5618 5263 5652 5271
rect 5652 5263 5661 5271
rect 5609 5219 5661 5263
rect 5809 5437 5861 5481
rect 5809 5429 5818 5437
rect 5818 5429 5852 5437
rect 5852 5429 5861 5437
rect 6009 5543 6018 5551
rect 6018 5543 6052 5551
rect 6052 5543 6061 5551
rect 6009 5499 6061 5543
rect 6209 5717 6261 5761
rect 6209 5709 6218 5717
rect 6218 5709 6252 5717
rect 6252 5709 6261 5717
rect 6409 5823 6418 5831
rect 6418 5823 6452 5831
rect 6452 5823 6461 5831
rect 6409 5779 6461 5823
rect 6507 5779 6559 5831
rect 5609 5123 5618 5131
rect 5618 5123 5652 5131
rect 5652 5123 5661 5131
rect 5609 5079 5661 5123
rect 5809 5297 5861 5341
rect 5809 5289 5818 5297
rect 5818 5289 5852 5297
rect 5852 5289 5861 5297
rect 6009 5403 6018 5411
rect 6018 5403 6052 5411
rect 6052 5403 6061 5411
rect 6009 5359 6061 5403
rect 6209 5577 6261 5621
rect 6209 5569 6218 5577
rect 6218 5569 6252 5577
rect 6252 5569 6261 5577
rect 6409 5683 6418 5691
rect 6418 5683 6452 5691
rect 6452 5683 6461 5691
rect 6409 5639 6461 5683
rect 6507 5639 6559 5691
rect 5809 5157 5861 5201
rect 5809 5149 5818 5157
rect 5818 5149 5852 5157
rect 5852 5149 5861 5157
rect 6009 5263 6018 5271
rect 6018 5263 6052 5271
rect 6052 5263 6061 5271
rect 6009 5219 6061 5263
rect 6209 5437 6261 5481
rect 6209 5429 6218 5437
rect 6218 5429 6252 5437
rect 6252 5429 6261 5437
rect 6409 5543 6418 5551
rect 6418 5543 6452 5551
rect 6452 5543 6461 5551
rect 6409 5499 6461 5543
rect 6507 5499 6559 5551
rect 6009 5123 6018 5131
rect 6018 5123 6052 5131
rect 6052 5123 6061 5131
rect 6009 5079 6061 5123
rect 6209 5297 6261 5341
rect 6209 5289 6218 5297
rect 6218 5289 6252 5297
rect 6252 5289 6261 5297
rect 6409 5403 6418 5411
rect 6418 5403 6452 5411
rect 6452 5403 6461 5411
rect 6409 5359 6461 5403
rect 6507 5359 6559 5411
rect 6209 5157 6261 5201
rect 6209 5149 6218 5157
rect 6218 5149 6252 5157
rect 6252 5149 6261 5157
rect 6409 5263 6418 5271
rect 6418 5263 6452 5271
rect 6452 5263 6461 5271
rect 6409 5219 6461 5263
rect 6507 5219 6559 5271
rect 6409 5123 6418 5131
rect 6418 5123 6452 5131
rect 6452 5123 6461 5131
rect 6409 5079 6461 5123
rect 6507 5079 6559 5131
rect 9 4894 61 4903
rect 9 4860 18 4894
rect 18 4860 52 4894
rect 52 4860 61 4894
rect 9 4851 61 4860
rect 9 4753 18 4761
rect 18 4753 52 4761
rect 52 4753 61 4761
rect 9 4709 61 4753
rect 209 4910 261 4919
rect 209 4876 218 4910
rect 218 4876 252 4910
rect 252 4876 261 4910
rect 209 4867 261 4876
rect 9 4613 18 4621
rect 18 4613 52 4621
rect 52 4613 61 4621
rect 9 4569 61 4613
rect 209 4787 261 4831
rect 209 4779 218 4787
rect 218 4779 252 4787
rect 252 4779 261 4787
rect 409 4894 461 4903
rect 409 4860 418 4894
rect 418 4860 452 4894
rect 452 4860 461 4894
rect 409 4851 461 4860
rect 9 4473 18 4481
rect 18 4473 52 4481
rect 52 4473 61 4481
rect 9 4429 61 4473
rect 209 4647 261 4691
rect 209 4639 218 4647
rect 218 4639 252 4647
rect 252 4639 261 4647
rect 409 4753 418 4761
rect 418 4753 452 4761
rect 452 4753 461 4761
rect 409 4709 461 4753
rect 609 4910 661 4919
rect 609 4876 618 4910
rect 618 4876 652 4910
rect 652 4876 661 4910
rect 609 4867 661 4876
rect 9 4333 18 4341
rect 18 4333 52 4341
rect 52 4333 61 4341
rect 9 4289 61 4333
rect 209 4507 261 4551
rect 209 4499 218 4507
rect 218 4499 252 4507
rect 252 4499 261 4507
rect 409 4613 418 4621
rect 418 4613 452 4621
rect 452 4613 461 4621
rect 409 4569 461 4613
rect 609 4787 661 4831
rect 609 4779 618 4787
rect 618 4779 652 4787
rect 652 4779 661 4787
rect 809 4894 861 4903
rect 809 4860 818 4894
rect 818 4860 852 4894
rect 852 4860 861 4894
rect 809 4851 861 4860
rect 9 4193 18 4201
rect 18 4193 52 4201
rect 52 4193 61 4201
rect 9 4149 61 4193
rect 209 4367 261 4411
rect 209 4359 218 4367
rect 218 4359 252 4367
rect 252 4359 261 4367
rect 409 4473 418 4481
rect 418 4473 452 4481
rect 452 4473 461 4481
rect 409 4429 461 4473
rect 609 4647 661 4691
rect 609 4639 618 4647
rect 618 4639 652 4647
rect 652 4639 661 4647
rect 809 4753 818 4761
rect 818 4753 852 4761
rect 852 4753 861 4761
rect 809 4709 861 4753
rect 1009 4910 1061 4919
rect 1009 4876 1018 4910
rect 1018 4876 1052 4910
rect 1052 4876 1061 4910
rect 1009 4867 1061 4876
rect 9 4053 18 4061
rect 18 4053 52 4061
rect 52 4053 61 4061
rect 9 4009 61 4053
rect 209 4227 261 4271
rect 209 4219 218 4227
rect 218 4219 252 4227
rect 252 4219 261 4227
rect 409 4333 418 4341
rect 418 4333 452 4341
rect 452 4333 461 4341
rect 409 4289 461 4333
rect 609 4507 661 4551
rect 609 4499 618 4507
rect 618 4499 652 4507
rect 652 4499 661 4507
rect 809 4613 818 4621
rect 818 4613 852 4621
rect 852 4613 861 4621
rect 809 4569 861 4613
rect 1009 4787 1061 4831
rect 1009 4779 1018 4787
rect 1018 4779 1052 4787
rect 1052 4779 1061 4787
rect 1209 4894 1261 4903
rect 1209 4860 1218 4894
rect 1218 4860 1252 4894
rect 1252 4860 1261 4894
rect 1209 4851 1261 4860
rect 9 3913 18 3921
rect 18 3913 52 3921
rect 52 3913 61 3921
rect 9 3869 61 3913
rect 209 4087 261 4131
rect 209 4079 218 4087
rect 218 4079 252 4087
rect 252 4079 261 4087
rect 409 4193 418 4201
rect 418 4193 452 4201
rect 452 4193 461 4201
rect 409 4149 461 4193
rect 609 4367 661 4411
rect 609 4359 618 4367
rect 618 4359 652 4367
rect 652 4359 661 4367
rect 809 4473 818 4481
rect 818 4473 852 4481
rect 852 4473 861 4481
rect 809 4429 861 4473
rect 1009 4647 1061 4691
rect 1009 4639 1018 4647
rect 1018 4639 1052 4647
rect 1052 4639 1061 4647
rect 1209 4753 1218 4761
rect 1218 4753 1252 4761
rect 1252 4753 1261 4761
rect 1209 4709 1261 4753
rect 1409 4910 1461 4919
rect 1409 4876 1418 4910
rect 1418 4876 1452 4910
rect 1452 4876 1461 4910
rect 1409 4867 1461 4876
rect 9 3773 18 3781
rect 18 3773 52 3781
rect 52 3773 61 3781
rect 9 3729 61 3773
rect 209 3947 261 3991
rect 209 3939 218 3947
rect 218 3939 252 3947
rect 252 3939 261 3947
rect 409 4053 418 4061
rect 418 4053 452 4061
rect 452 4053 461 4061
rect 409 4009 461 4053
rect 609 4227 661 4271
rect 609 4219 618 4227
rect 618 4219 652 4227
rect 652 4219 661 4227
rect 809 4333 818 4341
rect 818 4333 852 4341
rect 852 4333 861 4341
rect 809 4289 861 4333
rect 1009 4507 1061 4551
rect 1009 4499 1018 4507
rect 1018 4499 1052 4507
rect 1052 4499 1061 4507
rect 1209 4613 1218 4621
rect 1218 4613 1252 4621
rect 1252 4613 1261 4621
rect 1209 4569 1261 4613
rect 1409 4787 1461 4831
rect 1409 4779 1418 4787
rect 1418 4779 1452 4787
rect 1452 4779 1461 4787
rect 1609 4894 1661 4903
rect 1609 4860 1618 4894
rect 1618 4860 1652 4894
rect 1652 4860 1661 4894
rect 1609 4851 1661 4860
rect 9 3684 61 3693
rect 9 3650 18 3684
rect 18 3650 52 3684
rect 52 3650 61 3684
rect 9 3641 61 3650
rect 9 3543 18 3551
rect 18 3543 52 3551
rect 52 3543 61 3551
rect 9 3499 61 3543
rect 209 3807 261 3851
rect 209 3799 218 3807
rect 218 3799 252 3807
rect 252 3799 261 3807
rect 409 3913 418 3921
rect 418 3913 452 3921
rect 452 3913 461 3921
rect 409 3869 461 3913
rect 609 4087 661 4131
rect 609 4079 618 4087
rect 618 4079 652 4087
rect 652 4079 661 4087
rect 809 4193 818 4201
rect 818 4193 852 4201
rect 852 4193 861 4201
rect 809 4149 861 4193
rect 1009 4367 1061 4411
rect 1009 4359 1018 4367
rect 1018 4359 1052 4367
rect 1052 4359 1061 4367
rect 1209 4473 1218 4481
rect 1218 4473 1252 4481
rect 1252 4473 1261 4481
rect 1209 4429 1261 4473
rect 1409 4647 1461 4691
rect 1409 4639 1418 4647
rect 1418 4639 1452 4647
rect 1452 4639 1461 4647
rect 1609 4753 1618 4761
rect 1618 4753 1652 4761
rect 1652 4753 1661 4761
rect 1609 4709 1661 4753
rect 1809 4910 1861 4919
rect 1809 4876 1818 4910
rect 1818 4876 1852 4910
rect 1852 4876 1861 4910
rect 1809 4867 1861 4876
rect 209 3700 261 3709
rect 209 3666 218 3700
rect 218 3666 252 3700
rect 252 3666 261 3700
rect 209 3657 261 3666
rect 9 3403 18 3411
rect 18 3403 52 3411
rect 52 3403 61 3411
rect 9 3359 61 3403
rect 209 3577 261 3621
rect 209 3569 218 3577
rect 218 3569 252 3577
rect 252 3569 261 3577
rect 409 3773 418 3781
rect 418 3773 452 3781
rect 452 3773 461 3781
rect 409 3729 461 3773
rect 609 3947 661 3991
rect 609 3939 618 3947
rect 618 3939 652 3947
rect 652 3939 661 3947
rect 809 4053 818 4061
rect 818 4053 852 4061
rect 852 4053 861 4061
rect 809 4009 861 4053
rect 1009 4227 1061 4271
rect 1009 4219 1018 4227
rect 1018 4219 1052 4227
rect 1052 4219 1061 4227
rect 1209 4333 1218 4341
rect 1218 4333 1252 4341
rect 1252 4333 1261 4341
rect 1209 4289 1261 4333
rect 1409 4507 1461 4551
rect 1409 4499 1418 4507
rect 1418 4499 1452 4507
rect 1452 4499 1461 4507
rect 1609 4613 1618 4621
rect 1618 4613 1652 4621
rect 1652 4613 1661 4621
rect 1609 4569 1661 4613
rect 1809 4787 1861 4831
rect 1809 4779 1818 4787
rect 1818 4779 1852 4787
rect 1852 4779 1861 4787
rect 2009 4894 2061 4903
rect 2009 4860 2018 4894
rect 2018 4860 2052 4894
rect 2052 4860 2061 4894
rect 2009 4851 2061 4860
rect 409 3684 461 3693
rect 409 3650 418 3684
rect 418 3650 452 3684
rect 452 3650 461 3684
rect 409 3641 461 3650
rect 9 3263 18 3271
rect 18 3263 52 3271
rect 52 3263 61 3271
rect 9 3219 61 3263
rect 209 3437 261 3481
rect 209 3429 218 3437
rect 218 3429 252 3437
rect 252 3429 261 3437
rect 409 3543 418 3551
rect 418 3543 452 3551
rect 452 3543 461 3551
rect 409 3499 461 3543
rect 609 3807 661 3851
rect 609 3799 618 3807
rect 618 3799 652 3807
rect 652 3799 661 3807
rect 809 3913 818 3921
rect 818 3913 852 3921
rect 852 3913 861 3921
rect 809 3869 861 3913
rect 1009 4087 1061 4131
rect 1009 4079 1018 4087
rect 1018 4079 1052 4087
rect 1052 4079 1061 4087
rect 1209 4193 1218 4201
rect 1218 4193 1252 4201
rect 1252 4193 1261 4201
rect 1209 4149 1261 4193
rect 1409 4367 1461 4411
rect 1409 4359 1418 4367
rect 1418 4359 1452 4367
rect 1452 4359 1461 4367
rect 1609 4473 1618 4481
rect 1618 4473 1652 4481
rect 1652 4473 1661 4481
rect 1609 4429 1661 4473
rect 1809 4647 1861 4691
rect 1809 4639 1818 4647
rect 1818 4639 1852 4647
rect 1852 4639 1861 4647
rect 2009 4753 2018 4761
rect 2018 4753 2052 4761
rect 2052 4753 2061 4761
rect 2009 4709 2061 4753
rect 2209 4910 2261 4919
rect 2209 4876 2218 4910
rect 2218 4876 2252 4910
rect 2252 4876 2261 4910
rect 2209 4867 2261 4876
rect 609 3700 661 3709
rect 609 3666 618 3700
rect 618 3666 652 3700
rect 652 3666 661 3700
rect 609 3657 661 3666
rect 9 3123 18 3131
rect 18 3123 52 3131
rect 52 3123 61 3131
rect 9 3079 61 3123
rect 209 3297 261 3341
rect 209 3289 218 3297
rect 218 3289 252 3297
rect 252 3289 261 3297
rect 409 3403 418 3411
rect 418 3403 452 3411
rect 452 3403 461 3411
rect 409 3359 461 3403
rect 609 3577 661 3621
rect 609 3569 618 3577
rect 618 3569 652 3577
rect 652 3569 661 3577
rect 809 3773 818 3781
rect 818 3773 852 3781
rect 852 3773 861 3781
rect 809 3729 861 3773
rect 1009 3947 1061 3991
rect 1009 3939 1018 3947
rect 1018 3939 1052 3947
rect 1052 3939 1061 3947
rect 1209 4053 1218 4061
rect 1218 4053 1252 4061
rect 1252 4053 1261 4061
rect 1209 4009 1261 4053
rect 1409 4227 1461 4271
rect 1409 4219 1418 4227
rect 1418 4219 1452 4227
rect 1452 4219 1461 4227
rect 1609 4333 1618 4341
rect 1618 4333 1652 4341
rect 1652 4333 1661 4341
rect 1609 4289 1661 4333
rect 1809 4507 1861 4551
rect 1809 4499 1818 4507
rect 1818 4499 1852 4507
rect 1852 4499 1861 4507
rect 2009 4613 2018 4621
rect 2018 4613 2052 4621
rect 2052 4613 2061 4621
rect 2009 4569 2061 4613
rect 2209 4787 2261 4831
rect 2209 4779 2218 4787
rect 2218 4779 2252 4787
rect 2252 4779 2261 4787
rect 2409 4894 2461 4903
rect 2409 4860 2418 4894
rect 2418 4860 2452 4894
rect 2452 4860 2461 4894
rect 2409 4851 2461 4860
rect 809 3684 861 3693
rect 809 3650 818 3684
rect 818 3650 852 3684
rect 852 3650 861 3684
rect 809 3641 861 3650
rect 9 2983 18 2991
rect 18 2983 52 2991
rect 52 2983 61 2991
rect 9 2939 61 2983
rect 209 3157 261 3201
rect 209 3149 218 3157
rect 218 3149 252 3157
rect 252 3149 261 3157
rect 409 3263 418 3271
rect 418 3263 452 3271
rect 452 3263 461 3271
rect 409 3219 461 3263
rect 609 3437 661 3481
rect 609 3429 618 3437
rect 618 3429 652 3437
rect 652 3429 661 3437
rect 809 3543 818 3551
rect 818 3543 852 3551
rect 852 3543 861 3551
rect 809 3499 861 3543
rect 1009 3807 1061 3851
rect 1009 3799 1018 3807
rect 1018 3799 1052 3807
rect 1052 3799 1061 3807
rect 1209 3913 1218 3921
rect 1218 3913 1252 3921
rect 1252 3913 1261 3921
rect 1209 3869 1261 3913
rect 1409 4087 1461 4131
rect 1409 4079 1418 4087
rect 1418 4079 1452 4087
rect 1452 4079 1461 4087
rect 1609 4193 1618 4201
rect 1618 4193 1652 4201
rect 1652 4193 1661 4201
rect 1609 4149 1661 4193
rect 1809 4367 1861 4411
rect 1809 4359 1818 4367
rect 1818 4359 1852 4367
rect 1852 4359 1861 4367
rect 2009 4473 2018 4481
rect 2018 4473 2052 4481
rect 2052 4473 2061 4481
rect 2009 4429 2061 4473
rect 2209 4647 2261 4691
rect 2209 4639 2218 4647
rect 2218 4639 2252 4647
rect 2252 4639 2261 4647
rect 2409 4753 2418 4761
rect 2418 4753 2452 4761
rect 2452 4753 2461 4761
rect 2409 4709 2461 4753
rect 2609 4910 2661 4919
rect 2609 4876 2618 4910
rect 2618 4876 2652 4910
rect 2652 4876 2661 4910
rect 2609 4867 2661 4876
rect 1009 3700 1061 3709
rect 1009 3666 1018 3700
rect 1018 3666 1052 3700
rect 1052 3666 1061 3700
rect 1009 3657 1061 3666
rect 9 2843 18 2851
rect 18 2843 52 2851
rect 52 2843 61 2851
rect 9 2799 61 2843
rect 209 3017 261 3061
rect 209 3009 218 3017
rect 218 3009 252 3017
rect 252 3009 261 3017
rect 409 3123 418 3131
rect 418 3123 452 3131
rect 452 3123 461 3131
rect 409 3079 461 3123
rect 609 3297 661 3341
rect 609 3289 618 3297
rect 618 3289 652 3297
rect 652 3289 661 3297
rect 809 3403 818 3411
rect 818 3403 852 3411
rect 852 3403 861 3411
rect 809 3359 861 3403
rect 1009 3577 1061 3621
rect 1009 3569 1018 3577
rect 1018 3569 1052 3577
rect 1052 3569 1061 3577
rect 1209 3773 1218 3781
rect 1218 3773 1252 3781
rect 1252 3773 1261 3781
rect 1209 3729 1261 3773
rect 1409 3947 1461 3991
rect 1409 3939 1418 3947
rect 1418 3939 1452 3947
rect 1452 3939 1461 3947
rect 1609 4053 1618 4061
rect 1618 4053 1652 4061
rect 1652 4053 1661 4061
rect 1609 4009 1661 4053
rect 1809 4227 1861 4271
rect 1809 4219 1818 4227
rect 1818 4219 1852 4227
rect 1852 4219 1861 4227
rect 2009 4333 2018 4341
rect 2018 4333 2052 4341
rect 2052 4333 2061 4341
rect 2009 4289 2061 4333
rect 2209 4507 2261 4551
rect 2209 4499 2218 4507
rect 2218 4499 2252 4507
rect 2252 4499 2261 4507
rect 2409 4613 2418 4621
rect 2418 4613 2452 4621
rect 2452 4613 2461 4621
rect 2409 4569 2461 4613
rect 2609 4787 2661 4831
rect 2609 4779 2618 4787
rect 2618 4779 2652 4787
rect 2652 4779 2661 4787
rect 2809 4894 2861 4903
rect 2809 4860 2818 4894
rect 2818 4860 2852 4894
rect 2852 4860 2861 4894
rect 2809 4851 2861 4860
rect 1209 3684 1261 3693
rect 1209 3650 1218 3684
rect 1218 3650 1252 3684
rect 1252 3650 1261 3684
rect 1209 3641 1261 3650
rect 9 2703 18 2711
rect 18 2703 52 2711
rect 52 2703 61 2711
rect 9 2659 61 2703
rect 209 2877 261 2921
rect 209 2869 218 2877
rect 218 2869 252 2877
rect 252 2869 261 2877
rect 409 2983 418 2991
rect 418 2983 452 2991
rect 452 2983 461 2991
rect 409 2939 461 2983
rect 609 3157 661 3201
rect 609 3149 618 3157
rect 618 3149 652 3157
rect 652 3149 661 3157
rect 809 3263 818 3271
rect 818 3263 852 3271
rect 852 3263 861 3271
rect 809 3219 861 3263
rect 1009 3437 1061 3481
rect 1009 3429 1018 3437
rect 1018 3429 1052 3437
rect 1052 3429 1061 3437
rect 1209 3543 1218 3551
rect 1218 3543 1252 3551
rect 1252 3543 1261 3551
rect 1209 3499 1261 3543
rect 1409 3807 1461 3851
rect 1409 3799 1418 3807
rect 1418 3799 1452 3807
rect 1452 3799 1461 3807
rect 1609 3913 1618 3921
rect 1618 3913 1652 3921
rect 1652 3913 1661 3921
rect 1609 3869 1661 3913
rect 1809 4087 1861 4131
rect 1809 4079 1818 4087
rect 1818 4079 1852 4087
rect 1852 4079 1861 4087
rect 2009 4193 2018 4201
rect 2018 4193 2052 4201
rect 2052 4193 2061 4201
rect 2009 4149 2061 4193
rect 2209 4367 2261 4411
rect 2209 4359 2218 4367
rect 2218 4359 2252 4367
rect 2252 4359 2261 4367
rect 2409 4473 2418 4481
rect 2418 4473 2452 4481
rect 2452 4473 2461 4481
rect 2409 4429 2461 4473
rect 2609 4647 2661 4691
rect 2609 4639 2618 4647
rect 2618 4639 2652 4647
rect 2652 4639 2661 4647
rect 2809 4753 2818 4761
rect 2818 4753 2852 4761
rect 2852 4753 2861 4761
rect 2809 4709 2861 4753
rect 3009 4910 3061 4919
rect 3009 4876 3018 4910
rect 3018 4876 3052 4910
rect 3052 4876 3061 4910
rect 3009 4867 3061 4876
rect 1409 3700 1461 3709
rect 1409 3666 1418 3700
rect 1418 3666 1452 3700
rect 1452 3666 1461 3700
rect 1409 3657 1461 3666
rect 9 2563 18 2571
rect 18 2563 52 2571
rect 52 2563 61 2571
rect 9 2519 61 2563
rect 209 2737 261 2781
rect 209 2729 218 2737
rect 218 2729 252 2737
rect 252 2729 261 2737
rect 409 2843 418 2851
rect 418 2843 452 2851
rect 452 2843 461 2851
rect 409 2799 461 2843
rect 609 3017 661 3061
rect 609 3009 618 3017
rect 618 3009 652 3017
rect 652 3009 661 3017
rect 809 3123 818 3131
rect 818 3123 852 3131
rect 852 3123 861 3131
rect 809 3079 861 3123
rect 1009 3297 1061 3341
rect 1009 3289 1018 3297
rect 1018 3289 1052 3297
rect 1052 3289 1061 3297
rect 1209 3403 1218 3411
rect 1218 3403 1252 3411
rect 1252 3403 1261 3411
rect 1209 3359 1261 3403
rect 1409 3577 1461 3621
rect 1409 3569 1418 3577
rect 1418 3569 1452 3577
rect 1452 3569 1461 3577
rect 1609 3773 1618 3781
rect 1618 3773 1652 3781
rect 1652 3773 1661 3781
rect 1609 3729 1661 3773
rect 1809 3947 1861 3991
rect 1809 3939 1818 3947
rect 1818 3939 1852 3947
rect 1852 3939 1861 3947
rect 2009 4053 2018 4061
rect 2018 4053 2052 4061
rect 2052 4053 2061 4061
rect 2009 4009 2061 4053
rect 2209 4227 2261 4271
rect 2209 4219 2218 4227
rect 2218 4219 2252 4227
rect 2252 4219 2261 4227
rect 2409 4333 2418 4341
rect 2418 4333 2452 4341
rect 2452 4333 2461 4341
rect 2409 4289 2461 4333
rect 2609 4507 2661 4551
rect 2609 4499 2618 4507
rect 2618 4499 2652 4507
rect 2652 4499 2661 4507
rect 2809 4613 2818 4621
rect 2818 4613 2852 4621
rect 2852 4613 2861 4621
rect 2809 4569 2861 4613
rect 3009 4787 3061 4831
rect 3009 4779 3018 4787
rect 3018 4779 3052 4787
rect 3052 4779 3061 4787
rect 3209 4894 3261 4903
rect 3209 4860 3218 4894
rect 3218 4860 3252 4894
rect 3252 4860 3261 4894
rect 3209 4851 3261 4860
rect 1609 3684 1661 3693
rect 1609 3650 1618 3684
rect 1618 3650 1652 3684
rect 1652 3650 1661 3684
rect 1609 3641 1661 3650
rect 9 2474 61 2483
rect 9 2440 18 2474
rect 18 2440 52 2474
rect 52 2440 61 2474
rect 9 2431 61 2440
rect 9 2333 18 2341
rect 18 2333 52 2341
rect 52 2333 61 2341
rect 9 2289 61 2333
rect 209 2597 261 2641
rect 209 2589 218 2597
rect 218 2589 252 2597
rect 252 2589 261 2597
rect 409 2703 418 2711
rect 418 2703 452 2711
rect 452 2703 461 2711
rect 409 2659 461 2703
rect 609 2877 661 2921
rect 609 2869 618 2877
rect 618 2869 652 2877
rect 652 2869 661 2877
rect 809 2983 818 2991
rect 818 2983 852 2991
rect 852 2983 861 2991
rect 809 2939 861 2983
rect 1009 3157 1061 3201
rect 1009 3149 1018 3157
rect 1018 3149 1052 3157
rect 1052 3149 1061 3157
rect 1209 3263 1218 3271
rect 1218 3263 1252 3271
rect 1252 3263 1261 3271
rect 1209 3219 1261 3263
rect 1409 3437 1461 3481
rect 1409 3429 1418 3437
rect 1418 3429 1452 3437
rect 1452 3429 1461 3437
rect 1609 3543 1618 3551
rect 1618 3543 1652 3551
rect 1652 3543 1661 3551
rect 1609 3499 1661 3543
rect 1809 3807 1861 3851
rect 1809 3799 1818 3807
rect 1818 3799 1852 3807
rect 1852 3799 1861 3807
rect 2009 3913 2018 3921
rect 2018 3913 2052 3921
rect 2052 3913 2061 3921
rect 2009 3869 2061 3913
rect 2209 4087 2261 4131
rect 2209 4079 2218 4087
rect 2218 4079 2252 4087
rect 2252 4079 2261 4087
rect 2409 4193 2418 4201
rect 2418 4193 2452 4201
rect 2452 4193 2461 4201
rect 2409 4149 2461 4193
rect 2609 4367 2661 4411
rect 2609 4359 2618 4367
rect 2618 4359 2652 4367
rect 2652 4359 2661 4367
rect 2809 4473 2818 4481
rect 2818 4473 2852 4481
rect 2852 4473 2861 4481
rect 2809 4429 2861 4473
rect 3009 4647 3061 4691
rect 3009 4639 3018 4647
rect 3018 4639 3052 4647
rect 3052 4639 3061 4647
rect 3209 4753 3218 4761
rect 3218 4753 3252 4761
rect 3252 4753 3261 4761
rect 3209 4709 3261 4753
rect 3409 4910 3461 4919
rect 3409 4876 3418 4910
rect 3418 4876 3452 4910
rect 3452 4876 3461 4910
rect 3409 4867 3461 4876
rect 1809 3700 1861 3709
rect 1809 3666 1818 3700
rect 1818 3666 1852 3700
rect 1852 3666 1861 3700
rect 1809 3657 1861 3666
rect 209 2490 261 2499
rect 209 2456 218 2490
rect 218 2456 252 2490
rect 252 2456 261 2490
rect 209 2447 261 2456
rect 9 2193 18 2201
rect 18 2193 52 2201
rect 52 2193 61 2201
rect 9 2149 61 2193
rect 209 2367 261 2411
rect 209 2359 218 2367
rect 218 2359 252 2367
rect 252 2359 261 2367
rect 409 2563 418 2571
rect 418 2563 452 2571
rect 452 2563 461 2571
rect 409 2519 461 2563
rect 609 2737 661 2781
rect 609 2729 618 2737
rect 618 2729 652 2737
rect 652 2729 661 2737
rect 809 2843 818 2851
rect 818 2843 852 2851
rect 852 2843 861 2851
rect 809 2799 861 2843
rect 1009 3017 1061 3061
rect 1009 3009 1018 3017
rect 1018 3009 1052 3017
rect 1052 3009 1061 3017
rect 1209 3123 1218 3131
rect 1218 3123 1252 3131
rect 1252 3123 1261 3131
rect 1209 3079 1261 3123
rect 1409 3297 1461 3341
rect 1409 3289 1418 3297
rect 1418 3289 1452 3297
rect 1452 3289 1461 3297
rect 1609 3403 1618 3411
rect 1618 3403 1652 3411
rect 1652 3403 1661 3411
rect 1609 3359 1661 3403
rect 1809 3577 1861 3621
rect 1809 3569 1818 3577
rect 1818 3569 1852 3577
rect 1852 3569 1861 3577
rect 2009 3773 2018 3781
rect 2018 3773 2052 3781
rect 2052 3773 2061 3781
rect 2009 3729 2061 3773
rect 2209 3947 2261 3991
rect 2209 3939 2218 3947
rect 2218 3939 2252 3947
rect 2252 3939 2261 3947
rect 2409 4053 2418 4061
rect 2418 4053 2452 4061
rect 2452 4053 2461 4061
rect 2409 4009 2461 4053
rect 2609 4227 2661 4271
rect 2609 4219 2618 4227
rect 2618 4219 2652 4227
rect 2652 4219 2661 4227
rect 2809 4333 2818 4341
rect 2818 4333 2852 4341
rect 2852 4333 2861 4341
rect 2809 4289 2861 4333
rect 3009 4507 3061 4551
rect 3009 4499 3018 4507
rect 3018 4499 3052 4507
rect 3052 4499 3061 4507
rect 3209 4613 3218 4621
rect 3218 4613 3252 4621
rect 3252 4613 3261 4621
rect 3209 4569 3261 4613
rect 3409 4787 3461 4831
rect 3409 4779 3418 4787
rect 3418 4779 3452 4787
rect 3452 4779 3461 4787
rect 3609 4894 3661 4903
rect 3609 4860 3618 4894
rect 3618 4860 3652 4894
rect 3652 4860 3661 4894
rect 3609 4851 3661 4860
rect 2009 3684 2061 3693
rect 2009 3650 2018 3684
rect 2018 3650 2052 3684
rect 2052 3650 2061 3684
rect 2009 3641 2061 3650
rect 409 2474 461 2483
rect 409 2440 418 2474
rect 418 2440 452 2474
rect 452 2440 461 2474
rect 409 2431 461 2440
rect 9 2053 18 2061
rect 18 2053 52 2061
rect 52 2053 61 2061
rect 9 2009 61 2053
rect 209 2227 261 2271
rect 209 2219 218 2227
rect 218 2219 252 2227
rect 252 2219 261 2227
rect 409 2333 418 2341
rect 418 2333 452 2341
rect 452 2333 461 2341
rect 409 2289 461 2333
rect 609 2597 661 2641
rect 609 2589 618 2597
rect 618 2589 652 2597
rect 652 2589 661 2597
rect 809 2703 818 2711
rect 818 2703 852 2711
rect 852 2703 861 2711
rect 809 2659 861 2703
rect 1009 2877 1061 2921
rect 1009 2869 1018 2877
rect 1018 2869 1052 2877
rect 1052 2869 1061 2877
rect 1209 2983 1218 2991
rect 1218 2983 1252 2991
rect 1252 2983 1261 2991
rect 1209 2939 1261 2983
rect 1409 3157 1461 3201
rect 1409 3149 1418 3157
rect 1418 3149 1452 3157
rect 1452 3149 1461 3157
rect 1609 3263 1618 3271
rect 1618 3263 1652 3271
rect 1652 3263 1661 3271
rect 1609 3219 1661 3263
rect 1809 3437 1861 3481
rect 1809 3429 1818 3437
rect 1818 3429 1852 3437
rect 1852 3429 1861 3437
rect 2009 3543 2018 3551
rect 2018 3543 2052 3551
rect 2052 3543 2061 3551
rect 2009 3499 2061 3543
rect 2209 3807 2261 3851
rect 2209 3799 2218 3807
rect 2218 3799 2252 3807
rect 2252 3799 2261 3807
rect 2409 3913 2418 3921
rect 2418 3913 2452 3921
rect 2452 3913 2461 3921
rect 2409 3869 2461 3913
rect 2609 4087 2661 4131
rect 2609 4079 2618 4087
rect 2618 4079 2652 4087
rect 2652 4079 2661 4087
rect 2809 4193 2818 4201
rect 2818 4193 2852 4201
rect 2852 4193 2861 4201
rect 2809 4149 2861 4193
rect 3009 4367 3061 4411
rect 3009 4359 3018 4367
rect 3018 4359 3052 4367
rect 3052 4359 3061 4367
rect 3209 4473 3218 4481
rect 3218 4473 3252 4481
rect 3252 4473 3261 4481
rect 3209 4429 3261 4473
rect 3409 4647 3461 4691
rect 3409 4639 3418 4647
rect 3418 4639 3452 4647
rect 3452 4639 3461 4647
rect 3609 4753 3618 4761
rect 3618 4753 3652 4761
rect 3652 4753 3661 4761
rect 3609 4709 3661 4753
rect 3809 4910 3861 4919
rect 3809 4876 3818 4910
rect 3818 4876 3852 4910
rect 3852 4876 3861 4910
rect 3809 4867 3861 4876
rect 2209 3700 2261 3709
rect 2209 3666 2218 3700
rect 2218 3666 2252 3700
rect 2252 3666 2261 3700
rect 2209 3657 2261 3666
rect 609 2490 661 2499
rect 609 2456 618 2490
rect 618 2456 652 2490
rect 652 2456 661 2490
rect 609 2447 661 2456
rect 9 1913 18 1921
rect 18 1913 52 1921
rect 52 1913 61 1921
rect 9 1869 61 1913
rect 209 2087 261 2131
rect 209 2079 218 2087
rect 218 2079 252 2087
rect 252 2079 261 2087
rect 409 2193 418 2201
rect 418 2193 452 2201
rect 452 2193 461 2201
rect 409 2149 461 2193
rect 609 2367 661 2411
rect 609 2359 618 2367
rect 618 2359 652 2367
rect 652 2359 661 2367
rect 809 2563 818 2571
rect 818 2563 852 2571
rect 852 2563 861 2571
rect 809 2519 861 2563
rect 1009 2737 1061 2781
rect 1009 2729 1018 2737
rect 1018 2729 1052 2737
rect 1052 2729 1061 2737
rect 1209 2843 1218 2851
rect 1218 2843 1252 2851
rect 1252 2843 1261 2851
rect 1209 2799 1261 2843
rect 1409 3017 1461 3061
rect 1409 3009 1418 3017
rect 1418 3009 1452 3017
rect 1452 3009 1461 3017
rect 1609 3123 1618 3131
rect 1618 3123 1652 3131
rect 1652 3123 1661 3131
rect 1609 3079 1661 3123
rect 1809 3297 1861 3341
rect 1809 3289 1818 3297
rect 1818 3289 1852 3297
rect 1852 3289 1861 3297
rect 2009 3403 2018 3411
rect 2018 3403 2052 3411
rect 2052 3403 2061 3411
rect 2009 3359 2061 3403
rect 2209 3577 2261 3621
rect 2209 3569 2218 3577
rect 2218 3569 2252 3577
rect 2252 3569 2261 3577
rect 2409 3773 2418 3781
rect 2418 3773 2452 3781
rect 2452 3773 2461 3781
rect 2409 3729 2461 3773
rect 2609 3947 2661 3991
rect 2609 3939 2618 3947
rect 2618 3939 2652 3947
rect 2652 3939 2661 3947
rect 2809 4053 2818 4061
rect 2818 4053 2852 4061
rect 2852 4053 2861 4061
rect 2809 4009 2861 4053
rect 3009 4227 3061 4271
rect 3009 4219 3018 4227
rect 3018 4219 3052 4227
rect 3052 4219 3061 4227
rect 3209 4333 3218 4341
rect 3218 4333 3252 4341
rect 3252 4333 3261 4341
rect 3209 4289 3261 4333
rect 3409 4507 3461 4551
rect 3409 4499 3418 4507
rect 3418 4499 3452 4507
rect 3452 4499 3461 4507
rect 3609 4613 3618 4621
rect 3618 4613 3652 4621
rect 3652 4613 3661 4621
rect 3609 4569 3661 4613
rect 3809 4787 3861 4831
rect 3809 4779 3818 4787
rect 3818 4779 3852 4787
rect 3852 4779 3861 4787
rect 4009 4894 4061 4903
rect 4009 4860 4018 4894
rect 4018 4860 4052 4894
rect 4052 4860 4061 4894
rect 4009 4851 4061 4860
rect 2409 3684 2461 3693
rect 2409 3650 2418 3684
rect 2418 3650 2452 3684
rect 2452 3650 2461 3684
rect 2409 3641 2461 3650
rect 809 2474 861 2483
rect 809 2440 818 2474
rect 818 2440 852 2474
rect 852 2440 861 2474
rect 809 2431 861 2440
rect 9 1773 18 1781
rect 18 1773 52 1781
rect 52 1773 61 1781
rect 9 1729 61 1773
rect 209 1947 261 1991
rect 209 1939 218 1947
rect 218 1939 252 1947
rect 252 1939 261 1947
rect 409 2053 418 2061
rect 418 2053 452 2061
rect 452 2053 461 2061
rect 409 2009 461 2053
rect 609 2227 661 2271
rect 609 2219 618 2227
rect 618 2219 652 2227
rect 652 2219 661 2227
rect 809 2333 818 2341
rect 818 2333 852 2341
rect 852 2333 861 2341
rect 809 2289 861 2333
rect 1009 2597 1061 2641
rect 1009 2589 1018 2597
rect 1018 2589 1052 2597
rect 1052 2589 1061 2597
rect 1209 2703 1218 2711
rect 1218 2703 1252 2711
rect 1252 2703 1261 2711
rect 1209 2659 1261 2703
rect 1409 2877 1461 2921
rect 1409 2869 1418 2877
rect 1418 2869 1452 2877
rect 1452 2869 1461 2877
rect 1609 2983 1618 2991
rect 1618 2983 1652 2991
rect 1652 2983 1661 2991
rect 1609 2939 1661 2983
rect 1809 3157 1861 3201
rect 1809 3149 1818 3157
rect 1818 3149 1852 3157
rect 1852 3149 1861 3157
rect 2009 3263 2018 3271
rect 2018 3263 2052 3271
rect 2052 3263 2061 3271
rect 2009 3219 2061 3263
rect 2209 3437 2261 3481
rect 2209 3429 2218 3437
rect 2218 3429 2252 3437
rect 2252 3429 2261 3437
rect 2409 3543 2418 3551
rect 2418 3543 2452 3551
rect 2452 3543 2461 3551
rect 2409 3499 2461 3543
rect 2609 3807 2661 3851
rect 2609 3799 2618 3807
rect 2618 3799 2652 3807
rect 2652 3799 2661 3807
rect 2809 3913 2818 3921
rect 2818 3913 2852 3921
rect 2852 3913 2861 3921
rect 2809 3869 2861 3913
rect 3009 4087 3061 4131
rect 3009 4079 3018 4087
rect 3018 4079 3052 4087
rect 3052 4079 3061 4087
rect 3209 4193 3218 4201
rect 3218 4193 3252 4201
rect 3252 4193 3261 4201
rect 3209 4149 3261 4193
rect 3409 4367 3461 4411
rect 3409 4359 3418 4367
rect 3418 4359 3452 4367
rect 3452 4359 3461 4367
rect 3609 4473 3618 4481
rect 3618 4473 3652 4481
rect 3652 4473 3661 4481
rect 3609 4429 3661 4473
rect 3809 4647 3861 4691
rect 3809 4639 3818 4647
rect 3818 4639 3852 4647
rect 3852 4639 3861 4647
rect 4009 4753 4018 4761
rect 4018 4753 4052 4761
rect 4052 4753 4061 4761
rect 4009 4709 4061 4753
rect 4209 4910 4261 4919
rect 4209 4876 4218 4910
rect 4218 4876 4252 4910
rect 4252 4876 4261 4910
rect 4209 4867 4261 4876
rect 2609 3700 2661 3709
rect 2609 3666 2618 3700
rect 2618 3666 2652 3700
rect 2652 3666 2661 3700
rect 2609 3657 2661 3666
rect 1009 2490 1061 2499
rect 1009 2456 1018 2490
rect 1018 2456 1052 2490
rect 1052 2456 1061 2490
rect 1009 2447 1061 2456
rect 9 1633 18 1641
rect 18 1633 52 1641
rect 52 1633 61 1641
rect 9 1589 61 1633
rect 209 1807 261 1851
rect 209 1799 218 1807
rect 218 1799 252 1807
rect 252 1799 261 1807
rect 409 1913 418 1921
rect 418 1913 452 1921
rect 452 1913 461 1921
rect 409 1869 461 1913
rect 609 2087 661 2131
rect 609 2079 618 2087
rect 618 2079 652 2087
rect 652 2079 661 2087
rect 809 2193 818 2201
rect 818 2193 852 2201
rect 852 2193 861 2201
rect 809 2149 861 2193
rect 1009 2367 1061 2411
rect 1009 2359 1018 2367
rect 1018 2359 1052 2367
rect 1052 2359 1061 2367
rect 1209 2563 1218 2571
rect 1218 2563 1252 2571
rect 1252 2563 1261 2571
rect 1209 2519 1261 2563
rect 1409 2737 1461 2781
rect 1409 2729 1418 2737
rect 1418 2729 1452 2737
rect 1452 2729 1461 2737
rect 1609 2843 1618 2851
rect 1618 2843 1652 2851
rect 1652 2843 1661 2851
rect 1609 2799 1661 2843
rect 1809 3017 1861 3061
rect 1809 3009 1818 3017
rect 1818 3009 1852 3017
rect 1852 3009 1861 3017
rect 2009 3123 2018 3131
rect 2018 3123 2052 3131
rect 2052 3123 2061 3131
rect 2009 3079 2061 3123
rect 2209 3297 2261 3341
rect 2209 3289 2218 3297
rect 2218 3289 2252 3297
rect 2252 3289 2261 3297
rect 2409 3403 2418 3411
rect 2418 3403 2452 3411
rect 2452 3403 2461 3411
rect 2409 3359 2461 3403
rect 2609 3577 2661 3621
rect 2609 3569 2618 3577
rect 2618 3569 2652 3577
rect 2652 3569 2661 3577
rect 2809 3773 2818 3781
rect 2818 3773 2852 3781
rect 2852 3773 2861 3781
rect 2809 3729 2861 3773
rect 3009 3947 3061 3991
rect 3009 3939 3018 3947
rect 3018 3939 3052 3947
rect 3052 3939 3061 3947
rect 3209 4053 3218 4061
rect 3218 4053 3252 4061
rect 3252 4053 3261 4061
rect 3209 4009 3261 4053
rect 3409 4227 3461 4271
rect 3409 4219 3418 4227
rect 3418 4219 3452 4227
rect 3452 4219 3461 4227
rect 3609 4333 3618 4341
rect 3618 4333 3652 4341
rect 3652 4333 3661 4341
rect 3609 4289 3661 4333
rect 3809 4507 3861 4551
rect 3809 4499 3818 4507
rect 3818 4499 3852 4507
rect 3852 4499 3861 4507
rect 4009 4613 4018 4621
rect 4018 4613 4052 4621
rect 4052 4613 4061 4621
rect 4009 4569 4061 4613
rect 4209 4787 4261 4831
rect 4209 4779 4218 4787
rect 4218 4779 4252 4787
rect 4252 4779 4261 4787
rect 4409 4894 4461 4903
rect 4409 4860 4418 4894
rect 4418 4860 4452 4894
rect 4452 4860 4461 4894
rect 4409 4851 4461 4860
rect 2809 3684 2861 3693
rect 2809 3650 2818 3684
rect 2818 3650 2852 3684
rect 2852 3650 2861 3684
rect 2809 3641 2861 3650
rect 1209 2474 1261 2483
rect 1209 2440 1218 2474
rect 1218 2440 1252 2474
rect 1252 2440 1261 2474
rect 1209 2431 1261 2440
rect 9 1493 18 1501
rect 18 1493 52 1501
rect 52 1493 61 1501
rect 9 1449 61 1493
rect 209 1667 261 1711
rect 209 1659 218 1667
rect 218 1659 252 1667
rect 252 1659 261 1667
rect 409 1773 418 1781
rect 418 1773 452 1781
rect 452 1773 461 1781
rect 409 1729 461 1773
rect 609 1947 661 1991
rect 609 1939 618 1947
rect 618 1939 652 1947
rect 652 1939 661 1947
rect 809 2053 818 2061
rect 818 2053 852 2061
rect 852 2053 861 2061
rect 809 2009 861 2053
rect 1009 2227 1061 2271
rect 1009 2219 1018 2227
rect 1018 2219 1052 2227
rect 1052 2219 1061 2227
rect 1209 2333 1218 2341
rect 1218 2333 1252 2341
rect 1252 2333 1261 2341
rect 1209 2289 1261 2333
rect 1409 2597 1461 2641
rect 1409 2589 1418 2597
rect 1418 2589 1452 2597
rect 1452 2589 1461 2597
rect 1609 2703 1618 2711
rect 1618 2703 1652 2711
rect 1652 2703 1661 2711
rect 1609 2659 1661 2703
rect 1809 2877 1861 2921
rect 1809 2869 1818 2877
rect 1818 2869 1852 2877
rect 1852 2869 1861 2877
rect 2009 2983 2018 2991
rect 2018 2983 2052 2991
rect 2052 2983 2061 2991
rect 2009 2939 2061 2983
rect 2209 3157 2261 3201
rect 2209 3149 2218 3157
rect 2218 3149 2252 3157
rect 2252 3149 2261 3157
rect 2409 3263 2418 3271
rect 2418 3263 2452 3271
rect 2452 3263 2461 3271
rect 2409 3219 2461 3263
rect 2609 3437 2661 3481
rect 2609 3429 2618 3437
rect 2618 3429 2652 3437
rect 2652 3429 2661 3437
rect 2809 3543 2818 3551
rect 2818 3543 2852 3551
rect 2852 3543 2861 3551
rect 2809 3499 2861 3543
rect 3009 3807 3061 3851
rect 3009 3799 3018 3807
rect 3018 3799 3052 3807
rect 3052 3799 3061 3807
rect 3209 3913 3218 3921
rect 3218 3913 3252 3921
rect 3252 3913 3261 3921
rect 3209 3869 3261 3913
rect 3409 4087 3461 4131
rect 3409 4079 3418 4087
rect 3418 4079 3452 4087
rect 3452 4079 3461 4087
rect 3609 4193 3618 4201
rect 3618 4193 3652 4201
rect 3652 4193 3661 4201
rect 3609 4149 3661 4193
rect 3809 4367 3861 4411
rect 3809 4359 3818 4367
rect 3818 4359 3852 4367
rect 3852 4359 3861 4367
rect 4009 4473 4018 4481
rect 4018 4473 4052 4481
rect 4052 4473 4061 4481
rect 4009 4429 4061 4473
rect 4209 4647 4261 4691
rect 4209 4639 4218 4647
rect 4218 4639 4252 4647
rect 4252 4639 4261 4647
rect 4409 4753 4418 4761
rect 4418 4753 4452 4761
rect 4452 4753 4461 4761
rect 4409 4709 4461 4753
rect 4609 4910 4661 4919
rect 4609 4876 4618 4910
rect 4618 4876 4652 4910
rect 4652 4876 4661 4910
rect 4609 4867 4661 4876
rect 3009 3700 3061 3709
rect 3009 3666 3018 3700
rect 3018 3666 3052 3700
rect 3052 3666 3061 3700
rect 3009 3657 3061 3666
rect 1409 2490 1461 2499
rect 1409 2456 1418 2490
rect 1418 2456 1452 2490
rect 1452 2456 1461 2490
rect 1409 2447 1461 2456
rect 9 1353 18 1361
rect 18 1353 52 1361
rect 52 1353 61 1361
rect 9 1309 61 1353
rect 209 1527 261 1571
rect 209 1519 218 1527
rect 218 1519 252 1527
rect 252 1519 261 1527
rect 409 1633 418 1641
rect 418 1633 452 1641
rect 452 1633 461 1641
rect 409 1589 461 1633
rect 609 1807 661 1851
rect 609 1799 618 1807
rect 618 1799 652 1807
rect 652 1799 661 1807
rect 809 1913 818 1921
rect 818 1913 852 1921
rect 852 1913 861 1921
rect 809 1869 861 1913
rect 1009 2087 1061 2131
rect 1009 2079 1018 2087
rect 1018 2079 1052 2087
rect 1052 2079 1061 2087
rect 1209 2193 1218 2201
rect 1218 2193 1252 2201
rect 1252 2193 1261 2201
rect 1209 2149 1261 2193
rect 1409 2367 1461 2411
rect 1409 2359 1418 2367
rect 1418 2359 1452 2367
rect 1452 2359 1461 2367
rect 1609 2563 1618 2571
rect 1618 2563 1652 2571
rect 1652 2563 1661 2571
rect 1609 2519 1661 2563
rect 1809 2737 1861 2781
rect 1809 2729 1818 2737
rect 1818 2729 1852 2737
rect 1852 2729 1861 2737
rect 2009 2843 2018 2851
rect 2018 2843 2052 2851
rect 2052 2843 2061 2851
rect 2009 2799 2061 2843
rect 2209 3017 2261 3061
rect 2209 3009 2218 3017
rect 2218 3009 2252 3017
rect 2252 3009 2261 3017
rect 2409 3123 2418 3131
rect 2418 3123 2452 3131
rect 2452 3123 2461 3131
rect 2409 3079 2461 3123
rect 2609 3297 2661 3341
rect 2609 3289 2618 3297
rect 2618 3289 2652 3297
rect 2652 3289 2661 3297
rect 2809 3403 2818 3411
rect 2818 3403 2852 3411
rect 2852 3403 2861 3411
rect 2809 3359 2861 3403
rect 3009 3577 3061 3621
rect 3009 3569 3018 3577
rect 3018 3569 3052 3577
rect 3052 3569 3061 3577
rect 3209 3773 3218 3781
rect 3218 3773 3252 3781
rect 3252 3773 3261 3781
rect 3209 3729 3261 3773
rect 3409 3947 3461 3991
rect 3409 3939 3418 3947
rect 3418 3939 3452 3947
rect 3452 3939 3461 3947
rect 3609 4053 3618 4061
rect 3618 4053 3652 4061
rect 3652 4053 3661 4061
rect 3609 4009 3661 4053
rect 3809 4227 3861 4271
rect 3809 4219 3818 4227
rect 3818 4219 3852 4227
rect 3852 4219 3861 4227
rect 4009 4333 4018 4341
rect 4018 4333 4052 4341
rect 4052 4333 4061 4341
rect 4009 4289 4061 4333
rect 4209 4507 4261 4551
rect 4209 4499 4218 4507
rect 4218 4499 4252 4507
rect 4252 4499 4261 4507
rect 4409 4613 4418 4621
rect 4418 4613 4452 4621
rect 4452 4613 4461 4621
rect 4409 4569 4461 4613
rect 4609 4787 4661 4831
rect 4609 4779 4618 4787
rect 4618 4779 4652 4787
rect 4652 4779 4661 4787
rect 4809 4894 4861 4903
rect 4809 4860 4818 4894
rect 4818 4860 4852 4894
rect 4852 4860 4861 4894
rect 4809 4851 4861 4860
rect 3209 3684 3261 3693
rect 3209 3650 3218 3684
rect 3218 3650 3252 3684
rect 3252 3650 3261 3684
rect 3209 3641 3261 3650
rect 1609 2474 1661 2483
rect 1609 2440 1618 2474
rect 1618 2440 1652 2474
rect 1652 2440 1661 2474
rect 1609 2431 1661 2440
rect 9 1264 61 1273
rect 9 1230 18 1264
rect 18 1230 52 1264
rect 52 1230 61 1264
rect 9 1221 61 1230
rect 9 1123 18 1131
rect 18 1123 52 1131
rect 52 1123 61 1131
rect 9 1079 61 1123
rect 209 1387 261 1431
rect 209 1379 218 1387
rect 218 1379 252 1387
rect 252 1379 261 1387
rect 409 1493 418 1501
rect 418 1493 452 1501
rect 452 1493 461 1501
rect 409 1449 461 1493
rect 609 1667 661 1711
rect 609 1659 618 1667
rect 618 1659 652 1667
rect 652 1659 661 1667
rect 809 1773 818 1781
rect 818 1773 852 1781
rect 852 1773 861 1781
rect 809 1729 861 1773
rect 1009 1947 1061 1991
rect 1009 1939 1018 1947
rect 1018 1939 1052 1947
rect 1052 1939 1061 1947
rect 1209 2053 1218 2061
rect 1218 2053 1252 2061
rect 1252 2053 1261 2061
rect 1209 2009 1261 2053
rect 1409 2227 1461 2271
rect 1409 2219 1418 2227
rect 1418 2219 1452 2227
rect 1452 2219 1461 2227
rect 1609 2333 1618 2341
rect 1618 2333 1652 2341
rect 1652 2333 1661 2341
rect 1609 2289 1661 2333
rect 1809 2597 1861 2641
rect 1809 2589 1818 2597
rect 1818 2589 1852 2597
rect 1852 2589 1861 2597
rect 2009 2703 2018 2711
rect 2018 2703 2052 2711
rect 2052 2703 2061 2711
rect 2009 2659 2061 2703
rect 2209 2877 2261 2921
rect 2209 2869 2218 2877
rect 2218 2869 2252 2877
rect 2252 2869 2261 2877
rect 2409 2983 2418 2991
rect 2418 2983 2452 2991
rect 2452 2983 2461 2991
rect 2409 2939 2461 2983
rect 2609 3157 2661 3201
rect 2609 3149 2618 3157
rect 2618 3149 2652 3157
rect 2652 3149 2661 3157
rect 2809 3263 2818 3271
rect 2818 3263 2852 3271
rect 2852 3263 2861 3271
rect 2809 3219 2861 3263
rect 3009 3437 3061 3481
rect 3009 3429 3018 3437
rect 3018 3429 3052 3437
rect 3052 3429 3061 3437
rect 3209 3543 3218 3551
rect 3218 3543 3252 3551
rect 3252 3543 3261 3551
rect 3209 3499 3261 3543
rect 3409 3807 3461 3851
rect 3409 3799 3418 3807
rect 3418 3799 3452 3807
rect 3452 3799 3461 3807
rect 3609 3913 3618 3921
rect 3618 3913 3652 3921
rect 3652 3913 3661 3921
rect 3609 3869 3661 3913
rect 3809 4087 3861 4131
rect 3809 4079 3818 4087
rect 3818 4079 3852 4087
rect 3852 4079 3861 4087
rect 4009 4193 4018 4201
rect 4018 4193 4052 4201
rect 4052 4193 4061 4201
rect 4009 4149 4061 4193
rect 4209 4367 4261 4411
rect 4209 4359 4218 4367
rect 4218 4359 4252 4367
rect 4252 4359 4261 4367
rect 4409 4473 4418 4481
rect 4418 4473 4452 4481
rect 4452 4473 4461 4481
rect 4409 4429 4461 4473
rect 4609 4647 4661 4691
rect 4609 4639 4618 4647
rect 4618 4639 4652 4647
rect 4652 4639 4661 4647
rect 4809 4753 4818 4761
rect 4818 4753 4852 4761
rect 4852 4753 4861 4761
rect 4809 4709 4861 4753
rect 5009 4910 5061 4919
rect 5009 4876 5018 4910
rect 5018 4876 5052 4910
rect 5052 4876 5061 4910
rect 5009 4867 5061 4876
rect 3409 3700 3461 3709
rect 3409 3666 3418 3700
rect 3418 3666 3452 3700
rect 3452 3666 3461 3700
rect 3409 3657 3461 3666
rect 1809 2490 1861 2499
rect 1809 2456 1818 2490
rect 1818 2456 1852 2490
rect 1852 2456 1861 2490
rect 1809 2447 1861 2456
rect 209 1280 261 1289
rect 209 1246 218 1280
rect 218 1246 252 1280
rect 252 1246 261 1280
rect 209 1237 261 1246
rect 9 983 18 991
rect 18 983 52 991
rect 52 983 61 991
rect 9 939 61 983
rect 209 1157 261 1201
rect 209 1149 218 1157
rect 218 1149 252 1157
rect 252 1149 261 1157
rect 409 1353 418 1361
rect 418 1353 452 1361
rect 452 1353 461 1361
rect 409 1309 461 1353
rect 609 1527 661 1571
rect 609 1519 618 1527
rect 618 1519 652 1527
rect 652 1519 661 1527
rect 809 1633 818 1641
rect 818 1633 852 1641
rect 852 1633 861 1641
rect 809 1589 861 1633
rect 1009 1807 1061 1851
rect 1009 1799 1018 1807
rect 1018 1799 1052 1807
rect 1052 1799 1061 1807
rect 1209 1913 1218 1921
rect 1218 1913 1252 1921
rect 1252 1913 1261 1921
rect 1209 1869 1261 1913
rect 1409 2087 1461 2131
rect 1409 2079 1418 2087
rect 1418 2079 1452 2087
rect 1452 2079 1461 2087
rect 1609 2193 1618 2201
rect 1618 2193 1652 2201
rect 1652 2193 1661 2201
rect 1609 2149 1661 2193
rect 1809 2367 1861 2411
rect 1809 2359 1818 2367
rect 1818 2359 1852 2367
rect 1852 2359 1861 2367
rect 2009 2563 2018 2571
rect 2018 2563 2052 2571
rect 2052 2563 2061 2571
rect 2009 2519 2061 2563
rect 2209 2737 2261 2781
rect 2209 2729 2218 2737
rect 2218 2729 2252 2737
rect 2252 2729 2261 2737
rect 2409 2843 2418 2851
rect 2418 2843 2452 2851
rect 2452 2843 2461 2851
rect 2409 2799 2461 2843
rect 2609 3017 2661 3061
rect 2609 3009 2618 3017
rect 2618 3009 2652 3017
rect 2652 3009 2661 3017
rect 2809 3123 2818 3131
rect 2818 3123 2852 3131
rect 2852 3123 2861 3131
rect 2809 3079 2861 3123
rect 3009 3297 3061 3341
rect 3009 3289 3018 3297
rect 3018 3289 3052 3297
rect 3052 3289 3061 3297
rect 3209 3403 3218 3411
rect 3218 3403 3252 3411
rect 3252 3403 3261 3411
rect 3209 3359 3261 3403
rect 3409 3577 3461 3621
rect 3409 3569 3418 3577
rect 3418 3569 3452 3577
rect 3452 3569 3461 3577
rect 3609 3773 3618 3781
rect 3618 3773 3652 3781
rect 3652 3773 3661 3781
rect 3609 3729 3661 3773
rect 3809 3947 3861 3991
rect 3809 3939 3818 3947
rect 3818 3939 3852 3947
rect 3852 3939 3861 3947
rect 4009 4053 4018 4061
rect 4018 4053 4052 4061
rect 4052 4053 4061 4061
rect 4009 4009 4061 4053
rect 4209 4227 4261 4271
rect 4209 4219 4218 4227
rect 4218 4219 4252 4227
rect 4252 4219 4261 4227
rect 4409 4333 4418 4341
rect 4418 4333 4452 4341
rect 4452 4333 4461 4341
rect 4409 4289 4461 4333
rect 4609 4507 4661 4551
rect 4609 4499 4618 4507
rect 4618 4499 4652 4507
rect 4652 4499 4661 4507
rect 4809 4613 4818 4621
rect 4818 4613 4852 4621
rect 4852 4613 4861 4621
rect 4809 4569 4861 4613
rect 5009 4787 5061 4831
rect 5009 4779 5018 4787
rect 5018 4779 5052 4787
rect 5052 4779 5061 4787
rect 5209 4894 5261 4903
rect 5209 4860 5218 4894
rect 5218 4860 5252 4894
rect 5252 4860 5261 4894
rect 5209 4851 5261 4860
rect 3609 3684 3661 3693
rect 3609 3650 3618 3684
rect 3618 3650 3652 3684
rect 3652 3650 3661 3684
rect 3609 3641 3661 3650
rect 2009 2474 2061 2483
rect 2009 2440 2018 2474
rect 2018 2440 2052 2474
rect 2052 2440 2061 2474
rect 2009 2431 2061 2440
rect 409 1264 461 1273
rect 409 1230 418 1264
rect 418 1230 452 1264
rect 452 1230 461 1264
rect 409 1221 461 1230
rect 9 843 18 851
rect 18 843 52 851
rect 52 843 61 851
rect 9 799 61 843
rect 209 1017 261 1061
rect 209 1009 218 1017
rect 218 1009 252 1017
rect 252 1009 261 1017
rect 409 1123 418 1131
rect 418 1123 452 1131
rect 452 1123 461 1131
rect 409 1079 461 1123
rect 609 1387 661 1431
rect 609 1379 618 1387
rect 618 1379 652 1387
rect 652 1379 661 1387
rect 809 1493 818 1501
rect 818 1493 852 1501
rect 852 1493 861 1501
rect 809 1449 861 1493
rect 1009 1667 1061 1711
rect 1009 1659 1018 1667
rect 1018 1659 1052 1667
rect 1052 1659 1061 1667
rect 1209 1773 1218 1781
rect 1218 1773 1252 1781
rect 1252 1773 1261 1781
rect 1209 1729 1261 1773
rect 1409 1947 1461 1991
rect 1409 1939 1418 1947
rect 1418 1939 1452 1947
rect 1452 1939 1461 1947
rect 1609 2053 1618 2061
rect 1618 2053 1652 2061
rect 1652 2053 1661 2061
rect 1609 2009 1661 2053
rect 1809 2227 1861 2271
rect 1809 2219 1818 2227
rect 1818 2219 1852 2227
rect 1852 2219 1861 2227
rect 2009 2333 2018 2341
rect 2018 2333 2052 2341
rect 2052 2333 2061 2341
rect 2009 2289 2061 2333
rect 2209 2597 2261 2641
rect 2209 2589 2218 2597
rect 2218 2589 2252 2597
rect 2252 2589 2261 2597
rect 2409 2703 2418 2711
rect 2418 2703 2452 2711
rect 2452 2703 2461 2711
rect 2409 2659 2461 2703
rect 2609 2877 2661 2921
rect 2609 2869 2618 2877
rect 2618 2869 2652 2877
rect 2652 2869 2661 2877
rect 2809 2983 2818 2991
rect 2818 2983 2852 2991
rect 2852 2983 2861 2991
rect 2809 2939 2861 2983
rect 3009 3157 3061 3201
rect 3009 3149 3018 3157
rect 3018 3149 3052 3157
rect 3052 3149 3061 3157
rect 3209 3263 3218 3271
rect 3218 3263 3252 3271
rect 3252 3263 3261 3271
rect 3209 3219 3261 3263
rect 3409 3437 3461 3481
rect 3409 3429 3418 3437
rect 3418 3429 3452 3437
rect 3452 3429 3461 3437
rect 3609 3543 3618 3551
rect 3618 3543 3652 3551
rect 3652 3543 3661 3551
rect 3609 3499 3661 3543
rect 3809 3807 3861 3851
rect 3809 3799 3818 3807
rect 3818 3799 3852 3807
rect 3852 3799 3861 3807
rect 4009 3913 4018 3921
rect 4018 3913 4052 3921
rect 4052 3913 4061 3921
rect 4009 3869 4061 3913
rect 4209 4087 4261 4131
rect 4209 4079 4218 4087
rect 4218 4079 4252 4087
rect 4252 4079 4261 4087
rect 4409 4193 4418 4201
rect 4418 4193 4452 4201
rect 4452 4193 4461 4201
rect 4409 4149 4461 4193
rect 4609 4367 4661 4411
rect 4609 4359 4618 4367
rect 4618 4359 4652 4367
rect 4652 4359 4661 4367
rect 4809 4473 4818 4481
rect 4818 4473 4852 4481
rect 4852 4473 4861 4481
rect 4809 4429 4861 4473
rect 5009 4647 5061 4691
rect 5009 4639 5018 4647
rect 5018 4639 5052 4647
rect 5052 4639 5061 4647
rect 5209 4753 5218 4761
rect 5218 4753 5252 4761
rect 5252 4753 5261 4761
rect 5209 4709 5261 4753
rect 5409 4910 5461 4919
rect 5409 4876 5418 4910
rect 5418 4876 5452 4910
rect 5452 4876 5461 4910
rect 5409 4867 5461 4876
rect 3809 3700 3861 3709
rect 3809 3666 3818 3700
rect 3818 3666 3852 3700
rect 3852 3666 3861 3700
rect 3809 3657 3861 3666
rect 2209 2490 2261 2499
rect 2209 2456 2218 2490
rect 2218 2456 2252 2490
rect 2252 2456 2261 2490
rect 2209 2447 2261 2456
rect 609 1280 661 1289
rect 609 1246 618 1280
rect 618 1246 652 1280
rect 652 1246 661 1280
rect 609 1237 661 1246
rect 9 703 18 711
rect 18 703 52 711
rect 52 703 61 711
rect 9 659 61 703
rect 209 877 261 921
rect 209 869 218 877
rect 218 869 252 877
rect 252 869 261 877
rect 409 983 418 991
rect 418 983 452 991
rect 452 983 461 991
rect 409 939 461 983
rect 609 1157 661 1201
rect 609 1149 618 1157
rect 618 1149 652 1157
rect 652 1149 661 1157
rect 809 1353 818 1361
rect 818 1353 852 1361
rect 852 1353 861 1361
rect 809 1309 861 1353
rect 1009 1527 1061 1571
rect 1009 1519 1018 1527
rect 1018 1519 1052 1527
rect 1052 1519 1061 1527
rect 1209 1633 1218 1641
rect 1218 1633 1252 1641
rect 1252 1633 1261 1641
rect 1209 1589 1261 1633
rect 1409 1807 1461 1851
rect 1409 1799 1418 1807
rect 1418 1799 1452 1807
rect 1452 1799 1461 1807
rect 1609 1913 1618 1921
rect 1618 1913 1652 1921
rect 1652 1913 1661 1921
rect 1609 1869 1661 1913
rect 1809 2087 1861 2131
rect 1809 2079 1818 2087
rect 1818 2079 1852 2087
rect 1852 2079 1861 2087
rect 2009 2193 2018 2201
rect 2018 2193 2052 2201
rect 2052 2193 2061 2201
rect 2009 2149 2061 2193
rect 2209 2367 2261 2411
rect 2209 2359 2218 2367
rect 2218 2359 2252 2367
rect 2252 2359 2261 2367
rect 2409 2563 2418 2571
rect 2418 2563 2452 2571
rect 2452 2563 2461 2571
rect 2409 2519 2461 2563
rect 2609 2737 2661 2781
rect 2609 2729 2618 2737
rect 2618 2729 2652 2737
rect 2652 2729 2661 2737
rect 2809 2843 2818 2851
rect 2818 2843 2852 2851
rect 2852 2843 2861 2851
rect 2809 2799 2861 2843
rect 3009 3017 3061 3061
rect 3009 3009 3018 3017
rect 3018 3009 3052 3017
rect 3052 3009 3061 3017
rect 3209 3123 3218 3131
rect 3218 3123 3252 3131
rect 3252 3123 3261 3131
rect 3209 3079 3261 3123
rect 3409 3297 3461 3341
rect 3409 3289 3418 3297
rect 3418 3289 3452 3297
rect 3452 3289 3461 3297
rect 3609 3403 3618 3411
rect 3618 3403 3652 3411
rect 3652 3403 3661 3411
rect 3609 3359 3661 3403
rect 3809 3577 3861 3621
rect 3809 3569 3818 3577
rect 3818 3569 3852 3577
rect 3852 3569 3861 3577
rect 4009 3773 4018 3781
rect 4018 3773 4052 3781
rect 4052 3773 4061 3781
rect 4009 3729 4061 3773
rect 4209 3947 4261 3991
rect 4209 3939 4218 3947
rect 4218 3939 4252 3947
rect 4252 3939 4261 3947
rect 4409 4053 4418 4061
rect 4418 4053 4452 4061
rect 4452 4053 4461 4061
rect 4409 4009 4461 4053
rect 4609 4227 4661 4271
rect 4609 4219 4618 4227
rect 4618 4219 4652 4227
rect 4652 4219 4661 4227
rect 4809 4333 4818 4341
rect 4818 4333 4852 4341
rect 4852 4333 4861 4341
rect 4809 4289 4861 4333
rect 5009 4507 5061 4551
rect 5009 4499 5018 4507
rect 5018 4499 5052 4507
rect 5052 4499 5061 4507
rect 5209 4613 5218 4621
rect 5218 4613 5252 4621
rect 5252 4613 5261 4621
rect 5209 4569 5261 4613
rect 5409 4787 5461 4831
rect 5409 4779 5418 4787
rect 5418 4779 5452 4787
rect 5452 4779 5461 4787
rect 5609 4894 5661 4903
rect 5609 4860 5618 4894
rect 5618 4860 5652 4894
rect 5652 4860 5661 4894
rect 5609 4851 5661 4860
rect 4009 3684 4061 3693
rect 4009 3650 4018 3684
rect 4018 3650 4052 3684
rect 4052 3650 4061 3684
rect 4009 3641 4061 3650
rect 2409 2474 2461 2483
rect 2409 2440 2418 2474
rect 2418 2440 2452 2474
rect 2452 2440 2461 2474
rect 2409 2431 2461 2440
rect 809 1264 861 1273
rect 809 1230 818 1264
rect 818 1230 852 1264
rect 852 1230 861 1264
rect 809 1221 861 1230
rect 9 563 18 571
rect 18 563 52 571
rect 52 563 61 571
rect 9 519 61 563
rect 209 737 261 781
rect 209 729 218 737
rect 218 729 252 737
rect 252 729 261 737
rect 409 843 418 851
rect 418 843 452 851
rect 452 843 461 851
rect 409 799 461 843
rect 609 1017 661 1061
rect 609 1009 618 1017
rect 618 1009 652 1017
rect 652 1009 661 1017
rect 809 1123 818 1131
rect 818 1123 852 1131
rect 852 1123 861 1131
rect 809 1079 861 1123
rect 1009 1387 1061 1431
rect 1009 1379 1018 1387
rect 1018 1379 1052 1387
rect 1052 1379 1061 1387
rect 1209 1493 1218 1501
rect 1218 1493 1252 1501
rect 1252 1493 1261 1501
rect 1209 1449 1261 1493
rect 1409 1667 1461 1711
rect 1409 1659 1418 1667
rect 1418 1659 1452 1667
rect 1452 1659 1461 1667
rect 1609 1773 1618 1781
rect 1618 1773 1652 1781
rect 1652 1773 1661 1781
rect 1609 1729 1661 1773
rect 1809 1947 1861 1991
rect 1809 1939 1818 1947
rect 1818 1939 1852 1947
rect 1852 1939 1861 1947
rect 2009 2053 2018 2061
rect 2018 2053 2052 2061
rect 2052 2053 2061 2061
rect 2009 2009 2061 2053
rect 2209 2227 2261 2271
rect 2209 2219 2218 2227
rect 2218 2219 2252 2227
rect 2252 2219 2261 2227
rect 2409 2333 2418 2341
rect 2418 2333 2452 2341
rect 2452 2333 2461 2341
rect 2409 2289 2461 2333
rect 2609 2597 2661 2641
rect 2609 2589 2618 2597
rect 2618 2589 2652 2597
rect 2652 2589 2661 2597
rect 2809 2703 2818 2711
rect 2818 2703 2852 2711
rect 2852 2703 2861 2711
rect 2809 2659 2861 2703
rect 3009 2877 3061 2921
rect 3009 2869 3018 2877
rect 3018 2869 3052 2877
rect 3052 2869 3061 2877
rect 3209 2983 3218 2991
rect 3218 2983 3252 2991
rect 3252 2983 3261 2991
rect 3209 2939 3261 2983
rect 3409 3157 3461 3201
rect 3409 3149 3418 3157
rect 3418 3149 3452 3157
rect 3452 3149 3461 3157
rect 3609 3263 3618 3271
rect 3618 3263 3652 3271
rect 3652 3263 3661 3271
rect 3609 3219 3661 3263
rect 3809 3437 3861 3481
rect 3809 3429 3818 3437
rect 3818 3429 3852 3437
rect 3852 3429 3861 3437
rect 4009 3543 4018 3551
rect 4018 3543 4052 3551
rect 4052 3543 4061 3551
rect 4009 3499 4061 3543
rect 4209 3807 4261 3851
rect 4209 3799 4218 3807
rect 4218 3799 4252 3807
rect 4252 3799 4261 3807
rect 4409 3913 4418 3921
rect 4418 3913 4452 3921
rect 4452 3913 4461 3921
rect 4409 3869 4461 3913
rect 4609 4087 4661 4131
rect 4609 4079 4618 4087
rect 4618 4079 4652 4087
rect 4652 4079 4661 4087
rect 4809 4193 4818 4201
rect 4818 4193 4852 4201
rect 4852 4193 4861 4201
rect 4809 4149 4861 4193
rect 5009 4367 5061 4411
rect 5009 4359 5018 4367
rect 5018 4359 5052 4367
rect 5052 4359 5061 4367
rect 5209 4473 5218 4481
rect 5218 4473 5252 4481
rect 5252 4473 5261 4481
rect 5209 4429 5261 4473
rect 5409 4647 5461 4691
rect 5409 4639 5418 4647
rect 5418 4639 5452 4647
rect 5452 4639 5461 4647
rect 5609 4753 5618 4761
rect 5618 4753 5652 4761
rect 5652 4753 5661 4761
rect 5609 4709 5661 4753
rect 5809 4910 5861 4919
rect 5809 4876 5818 4910
rect 5818 4876 5852 4910
rect 5852 4876 5861 4910
rect 5809 4867 5861 4876
rect 4209 3700 4261 3709
rect 4209 3666 4218 3700
rect 4218 3666 4252 3700
rect 4252 3666 4261 3700
rect 4209 3657 4261 3666
rect 2609 2490 2661 2499
rect 2609 2456 2618 2490
rect 2618 2456 2652 2490
rect 2652 2456 2661 2490
rect 2609 2447 2661 2456
rect 1009 1280 1061 1289
rect 1009 1246 1018 1280
rect 1018 1246 1052 1280
rect 1052 1246 1061 1280
rect 1009 1237 1061 1246
rect 9 423 18 431
rect 18 423 52 431
rect 52 423 61 431
rect 9 379 61 423
rect 209 597 261 641
rect 209 589 218 597
rect 218 589 252 597
rect 252 589 261 597
rect 409 703 418 711
rect 418 703 452 711
rect 452 703 461 711
rect 409 659 461 703
rect 609 877 661 921
rect 609 869 618 877
rect 618 869 652 877
rect 652 869 661 877
rect 809 983 818 991
rect 818 983 852 991
rect 852 983 861 991
rect 809 939 861 983
rect 1009 1157 1061 1201
rect 1009 1149 1018 1157
rect 1018 1149 1052 1157
rect 1052 1149 1061 1157
rect 1209 1353 1218 1361
rect 1218 1353 1252 1361
rect 1252 1353 1261 1361
rect 1209 1309 1261 1353
rect 1409 1527 1461 1571
rect 1409 1519 1418 1527
rect 1418 1519 1452 1527
rect 1452 1519 1461 1527
rect 1609 1633 1618 1641
rect 1618 1633 1652 1641
rect 1652 1633 1661 1641
rect 1609 1589 1661 1633
rect 1809 1807 1861 1851
rect 1809 1799 1818 1807
rect 1818 1799 1852 1807
rect 1852 1799 1861 1807
rect 2009 1913 2018 1921
rect 2018 1913 2052 1921
rect 2052 1913 2061 1921
rect 2009 1869 2061 1913
rect 2209 2087 2261 2131
rect 2209 2079 2218 2087
rect 2218 2079 2252 2087
rect 2252 2079 2261 2087
rect 2409 2193 2418 2201
rect 2418 2193 2452 2201
rect 2452 2193 2461 2201
rect 2409 2149 2461 2193
rect 2609 2367 2661 2411
rect 2609 2359 2618 2367
rect 2618 2359 2652 2367
rect 2652 2359 2661 2367
rect 2809 2563 2818 2571
rect 2818 2563 2852 2571
rect 2852 2563 2861 2571
rect 2809 2519 2861 2563
rect 3009 2737 3061 2781
rect 3009 2729 3018 2737
rect 3018 2729 3052 2737
rect 3052 2729 3061 2737
rect 3209 2843 3218 2851
rect 3218 2843 3252 2851
rect 3252 2843 3261 2851
rect 3209 2799 3261 2843
rect 3409 3017 3461 3061
rect 3409 3009 3418 3017
rect 3418 3009 3452 3017
rect 3452 3009 3461 3017
rect 3609 3123 3618 3131
rect 3618 3123 3652 3131
rect 3652 3123 3661 3131
rect 3609 3079 3661 3123
rect 3809 3297 3861 3341
rect 3809 3289 3818 3297
rect 3818 3289 3852 3297
rect 3852 3289 3861 3297
rect 4009 3403 4018 3411
rect 4018 3403 4052 3411
rect 4052 3403 4061 3411
rect 4009 3359 4061 3403
rect 4209 3577 4261 3621
rect 4209 3569 4218 3577
rect 4218 3569 4252 3577
rect 4252 3569 4261 3577
rect 4409 3773 4418 3781
rect 4418 3773 4452 3781
rect 4452 3773 4461 3781
rect 4409 3729 4461 3773
rect 4609 3947 4661 3991
rect 4609 3939 4618 3947
rect 4618 3939 4652 3947
rect 4652 3939 4661 3947
rect 4809 4053 4818 4061
rect 4818 4053 4852 4061
rect 4852 4053 4861 4061
rect 4809 4009 4861 4053
rect 5009 4227 5061 4271
rect 5009 4219 5018 4227
rect 5018 4219 5052 4227
rect 5052 4219 5061 4227
rect 5209 4333 5218 4341
rect 5218 4333 5252 4341
rect 5252 4333 5261 4341
rect 5209 4289 5261 4333
rect 5409 4507 5461 4551
rect 5409 4499 5418 4507
rect 5418 4499 5452 4507
rect 5452 4499 5461 4507
rect 5609 4613 5618 4621
rect 5618 4613 5652 4621
rect 5652 4613 5661 4621
rect 5609 4569 5661 4613
rect 5809 4787 5861 4831
rect 5809 4779 5818 4787
rect 5818 4779 5852 4787
rect 5852 4779 5861 4787
rect 6009 4894 6061 4903
rect 6009 4860 6018 4894
rect 6018 4860 6052 4894
rect 6052 4860 6061 4894
rect 6009 4851 6061 4860
rect 4409 3684 4461 3693
rect 4409 3650 4418 3684
rect 4418 3650 4452 3684
rect 4452 3650 4461 3684
rect 4409 3641 4461 3650
rect 2809 2474 2861 2483
rect 2809 2440 2818 2474
rect 2818 2440 2852 2474
rect 2852 2440 2861 2474
rect 2809 2431 2861 2440
rect 1209 1264 1261 1273
rect 1209 1230 1218 1264
rect 1218 1230 1252 1264
rect 1252 1230 1261 1264
rect 1209 1221 1261 1230
rect 9 283 18 291
rect 18 283 52 291
rect 52 283 61 291
rect 9 239 61 283
rect 209 457 261 501
rect 209 449 218 457
rect 218 449 252 457
rect 252 449 261 457
rect 409 563 418 571
rect 418 563 452 571
rect 452 563 461 571
rect 409 519 461 563
rect 609 737 661 781
rect 609 729 618 737
rect 618 729 652 737
rect 652 729 661 737
rect 809 843 818 851
rect 818 843 852 851
rect 852 843 861 851
rect 809 799 861 843
rect 1009 1017 1061 1061
rect 1009 1009 1018 1017
rect 1018 1009 1052 1017
rect 1052 1009 1061 1017
rect 1209 1123 1218 1131
rect 1218 1123 1252 1131
rect 1252 1123 1261 1131
rect 1209 1079 1261 1123
rect 1409 1387 1461 1431
rect 1409 1379 1418 1387
rect 1418 1379 1452 1387
rect 1452 1379 1461 1387
rect 1609 1493 1618 1501
rect 1618 1493 1652 1501
rect 1652 1493 1661 1501
rect 1609 1449 1661 1493
rect 1809 1667 1861 1711
rect 1809 1659 1818 1667
rect 1818 1659 1852 1667
rect 1852 1659 1861 1667
rect 2009 1773 2018 1781
rect 2018 1773 2052 1781
rect 2052 1773 2061 1781
rect 2009 1729 2061 1773
rect 2209 1947 2261 1991
rect 2209 1939 2218 1947
rect 2218 1939 2252 1947
rect 2252 1939 2261 1947
rect 2409 2053 2418 2061
rect 2418 2053 2452 2061
rect 2452 2053 2461 2061
rect 2409 2009 2461 2053
rect 2609 2227 2661 2271
rect 2609 2219 2618 2227
rect 2618 2219 2652 2227
rect 2652 2219 2661 2227
rect 2809 2333 2818 2341
rect 2818 2333 2852 2341
rect 2852 2333 2861 2341
rect 2809 2289 2861 2333
rect 3009 2597 3061 2641
rect 3009 2589 3018 2597
rect 3018 2589 3052 2597
rect 3052 2589 3061 2597
rect 3209 2703 3218 2711
rect 3218 2703 3252 2711
rect 3252 2703 3261 2711
rect 3209 2659 3261 2703
rect 3409 2877 3461 2921
rect 3409 2869 3418 2877
rect 3418 2869 3452 2877
rect 3452 2869 3461 2877
rect 3609 2983 3618 2991
rect 3618 2983 3652 2991
rect 3652 2983 3661 2991
rect 3609 2939 3661 2983
rect 3809 3157 3861 3201
rect 3809 3149 3818 3157
rect 3818 3149 3852 3157
rect 3852 3149 3861 3157
rect 4009 3263 4018 3271
rect 4018 3263 4052 3271
rect 4052 3263 4061 3271
rect 4009 3219 4061 3263
rect 4209 3437 4261 3481
rect 4209 3429 4218 3437
rect 4218 3429 4252 3437
rect 4252 3429 4261 3437
rect 4409 3543 4418 3551
rect 4418 3543 4452 3551
rect 4452 3543 4461 3551
rect 4409 3499 4461 3543
rect 4609 3807 4661 3851
rect 4609 3799 4618 3807
rect 4618 3799 4652 3807
rect 4652 3799 4661 3807
rect 4809 3913 4818 3921
rect 4818 3913 4852 3921
rect 4852 3913 4861 3921
rect 4809 3869 4861 3913
rect 5009 4087 5061 4131
rect 5009 4079 5018 4087
rect 5018 4079 5052 4087
rect 5052 4079 5061 4087
rect 5209 4193 5218 4201
rect 5218 4193 5252 4201
rect 5252 4193 5261 4201
rect 5209 4149 5261 4193
rect 5409 4367 5461 4411
rect 5409 4359 5418 4367
rect 5418 4359 5452 4367
rect 5452 4359 5461 4367
rect 5609 4473 5618 4481
rect 5618 4473 5652 4481
rect 5652 4473 5661 4481
rect 5609 4429 5661 4473
rect 5809 4647 5861 4691
rect 5809 4639 5818 4647
rect 5818 4639 5852 4647
rect 5852 4639 5861 4647
rect 6009 4753 6018 4761
rect 6018 4753 6052 4761
rect 6052 4753 6061 4761
rect 6009 4709 6061 4753
rect 6209 4910 6261 4919
rect 6209 4876 6218 4910
rect 6218 4876 6252 4910
rect 6252 4876 6261 4910
rect 6209 4867 6261 4876
rect 4609 3700 4661 3709
rect 4609 3666 4618 3700
rect 4618 3666 4652 3700
rect 4652 3666 4661 3700
rect 4609 3657 4661 3666
rect 3009 2490 3061 2499
rect 3009 2456 3018 2490
rect 3018 2456 3052 2490
rect 3052 2456 3061 2490
rect 3009 2447 3061 2456
rect 1409 1280 1461 1289
rect 1409 1246 1418 1280
rect 1418 1246 1452 1280
rect 1452 1246 1461 1280
rect 1409 1237 1461 1246
rect 9 143 18 151
rect 18 143 52 151
rect 52 143 61 151
rect 9 99 61 143
rect 209 317 261 361
rect 209 309 218 317
rect 218 309 252 317
rect 252 309 261 317
rect 409 423 418 431
rect 418 423 452 431
rect 452 423 461 431
rect 409 379 461 423
rect 609 597 661 641
rect 609 589 618 597
rect 618 589 652 597
rect 652 589 661 597
rect 809 703 818 711
rect 818 703 852 711
rect 852 703 861 711
rect 809 659 861 703
rect 1009 877 1061 921
rect 1009 869 1018 877
rect 1018 869 1052 877
rect 1052 869 1061 877
rect 1209 983 1218 991
rect 1218 983 1252 991
rect 1252 983 1261 991
rect 1209 939 1261 983
rect 1409 1157 1461 1201
rect 1409 1149 1418 1157
rect 1418 1149 1452 1157
rect 1452 1149 1461 1157
rect 1609 1353 1618 1361
rect 1618 1353 1652 1361
rect 1652 1353 1661 1361
rect 1609 1309 1661 1353
rect 1809 1527 1861 1571
rect 1809 1519 1818 1527
rect 1818 1519 1852 1527
rect 1852 1519 1861 1527
rect 2009 1633 2018 1641
rect 2018 1633 2052 1641
rect 2052 1633 2061 1641
rect 2009 1589 2061 1633
rect 2209 1807 2261 1851
rect 2209 1799 2218 1807
rect 2218 1799 2252 1807
rect 2252 1799 2261 1807
rect 2409 1913 2418 1921
rect 2418 1913 2452 1921
rect 2452 1913 2461 1921
rect 2409 1869 2461 1913
rect 2609 2087 2661 2131
rect 2609 2079 2618 2087
rect 2618 2079 2652 2087
rect 2652 2079 2661 2087
rect 2809 2193 2818 2201
rect 2818 2193 2852 2201
rect 2852 2193 2861 2201
rect 2809 2149 2861 2193
rect 3009 2367 3061 2411
rect 3009 2359 3018 2367
rect 3018 2359 3052 2367
rect 3052 2359 3061 2367
rect 3209 2563 3218 2571
rect 3218 2563 3252 2571
rect 3252 2563 3261 2571
rect 3209 2519 3261 2563
rect 3409 2737 3461 2781
rect 3409 2729 3418 2737
rect 3418 2729 3452 2737
rect 3452 2729 3461 2737
rect 3609 2843 3618 2851
rect 3618 2843 3652 2851
rect 3652 2843 3661 2851
rect 3609 2799 3661 2843
rect 3809 3017 3861 3061
rect 3809 3009 3818 3017
rect 3818 3009 3852 3017
rect 3852 3009 3861 3017
rect 4009 3123 4018 3131
rect 4018 3123 4052 3131
rect 4052 3123 4061 3131
rect 4009 3079 4061 3123
rect 4209 3297 4261 3341
rect 4209 3289 4218 3297
rect 4218 3289 4252 3297
rect 4252 3289 4261 3297
rect 4409 3403 4418 3411
rect 4418 3403 4452 3411
rect 4452 3403 4461 3411
rect 4409 3359 4461 3403
rect 4609 3577 4661 3621
rect 4609 3569 4618 3577
rect 4618 3569 4652 3577
rect 4652 3569 4661 3577
rect 4809 3773 4818 3781
rect 4818 3773 4852 3781
rect 4852 3773 4861 3781
rect 4809 3729 4861 3773
rect 5009 3947 5061 3991
rect 5009 3939 5018 3947
rect 5018 3939 5052 3947
rect 5052 3939 5061 3947
rect 5209 4053 5218 4061
rect 5218 4053 5252 4061
rect 5252 4053 5261 4061
rect 5209 4009 5261 4053
rect 5409 4227 5461 4271
rect 5409 4219 5418 4227
rect 5418 4219 5452 4227
rect 5452 4219 5461 4227
rect 5609 4333 5618 4341
rect 5618 4333 5652 4341
rect 5652 4333 5661 4341
rect 5609 4289 5661 4333
rect 5809 4507 5861 4551
rect 5809 4499 5818 4507
rect 5818 4499 5852 4507
rect 5852 4499 5861 4507
rect 6009 4613 6018 4621
rect 6018 4613 6052 4621
rect 6052 4613 6061 4621
rect 6009 4569 6061 4613
rect 6209 4787 6261 4831
rect 6209 4779 6218 4787
rect 6218 4779 6252 4787
rect 6252 4779 6261 4787
rect 4809 3684 4861 3693
rect 4809 3650 4818 3684
rect 4818 3650 4852 3684
rect 4852 3650 4861 3684
rect 4809 3641 4861 3650
rect 3209 2474 3261 2483
rect 3209 2440 3218 2474
rect 3218 2440 3252 2474
rect 3252 2440 3261 2474
rect 3209 2431 3261 2440
rect 1609 1264 1661 1273
rect 1609 1230 1618 1264
rect 1618 1230 1652 1264
rect 1652 1230 1661 1264
rect 1609 1221 1661 1230
rect 9 54 61 63
rect 9 20 18 54
rect 18 20 52 54
rect 52 20 61 54
rect 9 11 61 20
rect -91 -60 -39 -15
rect -91 -67 -82 -60
rect -82 -67 -48 -60
rect -48 -67 -39 -60
rect -91 -94 -82 -79
rect -82 -94 -48 -79
rect -48 -94 -39 -79
rect -91 -131 -39 -94
rect 9 -74 61 -22
rect 209 177 261 221
rect 209 169 218 177
rect 218 169 252 177
rect 252 169 261 177
rect 409 283 418 291
rect 418 283 452 291
rect 452 283 461 291
rect 409 239 461 283
rect 609 457 661 501
rect 609 449 618 457
rect 618 449 652 457
rect 652 449 661 457
rect 809 563 818 571
rect 818 563 852 571
rect 852 563 861 571
rect 809 519 861 563
rect 1009 737 1061 781
rect 1009 729 1018 737
rect 1018 729 1052 737
rect 1052 729 1061 737
rect 1209 843 1218 851
rect 1218 843 1252 851
rect 1252 843 1261 851
rect 1209 799 1261 843
rect 1409 1017 1461 1061
rect 1409 1009 1418 1017
rect 1418 1009 1452 1017
rect 1452 1009 1461 1017
rect 1609 1123 1618 1131
rect 1618 1123 1652 1131
rect 1652 1123 1661 1131
rect 1609 1079 1661 1123
rect 1809 1387 1861 1431
rect 1809 1379 1818 1387
rect 1818 1379 1852 1387
rect 1852 1379 1861 1387
rect 2009 1493 2018 1501
rect 2018 1493 2052 1501
rect 2052 1493 2061 1501
rect 2009 1449 2061 1493
rect 2209 1667 2261 1711
rect 2209 1659 2218 1667
rect 2218 1659 2252 1667
rect 2252 1659 2261 1667
rect 2409 1773 2418 1781
rect 2418 1773 2452 1781
rect 2452 1773 2461 1781
rect 2409 1729 2461 1773
rect 2609 1947 2661 1991
rect 2609 1939 2618 1947
rect 2618 1939 2652 1947
rect 2652 1939 2661 1947
rect 2809 2053 2818 2061
rect 2818 2053 2852 2061
rect 2852 2053 2861 2061
rect 2809 2009 2861 2053
rect 3009 2227 3061 2271
rect 3009 2219 3018 2227
rect 3018 2219 3052 2227
rect 3052 2219 3061 2227
rect 3209 2333 3218 2341
rect 3218 2333 3252 2341
rect 3252 2333 3261 2341
rect 3209 2289 3261 2333
rect 3409 2597 3461 2641
rect 3409 2589 3418 2597
rect 3418 2589 3452 2597
rect 3452 2589 3461 2597
rect 3609 2703 3618 2711
rect 3618 2703 3652 2711
rect 3652 2703 3661 2711
rect 3609 2659 3661 2703
rect 3809 2877 3861 2921
rect 3809 2869 3818 2877
rect 3818 2869 3852 2877
rect 3852 2869 3861 2877
rect 4009 2983 4018 2991
rect 4018 2983 4052 2991
rect 4052 2983 4061 2991
rect 4009 2939 4061 2983
rect 4209 3157 4261 3201
rect 4209 3149 4218 3157
rect 4218 3149 4252 3157
rect 4252 3149 4261 3157
rect 4409 3263 4418 3271
rect 4418 3263 4452 3271
rect 4452 3263 4461 3271
rect 4409 3219 4461 3263
rect 4609 3437 4661 3481
rect 4609 3429 4618 3437
rect 4618 3429 4652 3437
rect 4652 3429 4661 3437
rect 4809 3543 4818 3551
rect 4818 3543 4852 3551
rect 4852 3543 4861 3551
rect 4809 3499 4861 3543
rect 5009 3807 5061 3851
rect 5009 3799 5018 3807
rect 5018 3799 5052 3807
rect 5052 3799 5061 3807
rect 5209 3913 5218 3921
rect 5218 3913 5252 3921
rect 5252 3913 5261 3921
rect 5209 3869 5261 3913
rect 5409 4087 5461 4131
rect 5409 4079 5418 4087
rect 5418 4079 5452 4087
rect 5452 4079 5461 4087
rect 5609 4193 5618 4201
rect 5618 4193 5652 4201
rect 5652 4193 5661 4201
rect 5609 4149 5661 4193
rect 5809 4367 5861 4411
rect 5809 4359 5818 4367
rect 5818 4359 5852 4367
rect 5852 4359 5861 4367
rect 6009 4473 6018 4481
rect 6018 4473 6052 4481
rect 6052 4473 6061 4481
rect 6009 4429 6061 4473
rect 6209 4647 6261 4691
rect 6209 4639 6218 4647
rect 6218 4639 6252 4647
rect 6252 4639 6261 4647
rect 6409 4753 6418 4761
rect 6418 4753 6452 4761
rect 6452 4753 6461 4761
rect 6409 4709 6461 4753
rect 6507 4709 6559 4761
rect 5009 3700 5061 3709
rect 5009 3666 5018 3700
rect 5018 3666 5052 3700
rect 5052 3666 5061 3700
rect 5009 3657 5061 3666
rect 3409 2490 3461 2499
rect 3409 2456 3418 2490
rect 3418 2456 3452 2490
rect 3452 2456 3461 2490
rect 3409 2447 3461 2456
rect 1809 1280 1861 1289
rect 1809 1246 1818 1280
rect 1818 1246 1852 1280
rect 1852 1246 1861 1280
rect 1809 1237 1861 1246
rect 209 70 261 79
rect 209 36 218 70
rect 218 36 252 70
rect 252 36 261 70
rect 209 27 261 36
rect 109 -60 161 -15
rect 109 -67 118 -60
rect 118 -67 152 -60
rect 152 -67 161 -60
rect -91 -166 -82 -143
rect -82 -166 -48 -143
rect -48 -166 -39 -143
rect -91 -195 -39 -166
rect -75 -248 -23 -239
rect -75 -282 -66 -248
rect -66 -282 -32 -248
rect -32 -282 -23 -248
rect -75 -291 -23 -282
rect -91 -363 -39 -326
rect -91 -378 -82 -363
rect -82 -378 -48 -363
rect -48 -378 -39 -363
rect -91 -397 -82 -390
rect -82 -397 -48 -390
rect -48 -397 -39 -390
rect -91 -435 -39 -397
rect -91 -442 -82 -435
rect -82 -442 -48 -435
rect -48 -442 -39 -435
rect -91 -469 -82 -454
rect -82 -469 -48 -454
rect -48 -469 -39 -454
rect -91 -506 -39 -469
rect 109 -94 118 -79
rect 118 -94 152 -79
rect 152 -94 161 -79
rect 109 -131 161 -94
rect 209 -74 261 -22
rect 409 143 418 151
rect 418 143 452 151
rect 452 143 461 151
rect 409 99 461 143
rect 609 317 661 361
rect 609 309 618 317
rect 618 309 652 317
rect 652 309 661 317
rect 809 423 818 431
rect 818 423 852 431
rect 852 423 861 431
rect 809 379 861 423
rect 1009 597 1061 641
rect 1009 589 1018 597
rect 1018 589 1052 597
rect 1052 589 1061 597
rect 1209 703 1218 711
rect 1218 703 1252 711
rect 1252 703 1261 711
rect 1209 659 1261 703
rect 1409 877 1461 921
rect 1409 869 1418 877
rect 1418 869 1452 877
rect 1452 869 1461 877
rect 1609 983 1618 991
rect 1618 983 1652 991
rect 1652 983 1661 991
rect 1609 939 1661 983
rect 1809 1157 1861 1201
rect 1809 1149 1818 1157
rect 1818 1149 1852 1157
rect 1852 1149 1861 1157
rect 2009 1353 2018 1361
rect 2018 1353 2052 1361
rect 2052 1353 2061 1361
rect 2009 1309 2061 1353
rect 2209 1527 2261 1571
rect 2209 1519 2218 1527
rect 2218 1519 2252 1527
rect 2252 1519 2261 1527
rect 2409 1633 2418 1641
rect 2418 1633 2452 1641
rect 2452 1633 2461 1641
rect 2409 1589 2461 1633
rect 2609 1807 2661 1851
rect 2609 1799 2618 1807
rect 2618 1799 2652 1807
rect 2652 1799 2661 1807
rect 2809 1913 2818 1921
rect 2818 1913 2852 1921
rect 2852 1913 2861 1921
rect 2809 1869 2861 1913
rect 3009 2087 3061 2131
rect 3009 2079 3018 2087
rect 3018 2079 3052 2087
rect 3052 2079 3061 2087
rect 3209 2193 3218 2201
rect 3218 2193 3252 2201
rect 3252 2193 3261 2201
rect 3209 2149 3261 2193
rect 3409 2367 3461 2411
rect 3409 2359 3418 2367
rect 3418 2359 3452 2367
rect 3452 2359 3461 2367
rect 3609 2563 3618 2571
rect 3618 2563 3652 2571
rect 3652 2563 3661 2571
rect 3609 2519 3661 2563
rect 3809 2737 3861 2781
rect 3809 2729 3818 2737
rect 3818 2729 3852 2737
rect 3852 2729 3861 2737
rect 4009 2843 4018 2851
rect 4018 2843 4052 2851
rect 4052 2843 4061 2851
rect 4009 2799 4061 2843
rect 4209 3017 4261 3061
rect 4209 3009 4218 3017
rect 4218 3009 4252 3017
rect 4252 3009 4261 3017
rect 4409 3123 4418 3131
rect 4418 3123 4452 3131
rect 4452 3123 4461 3131
rect 4409 3079 4461 3123
rect 4609 3297 4661 3341
rect 4609 3289 4618 3297
rect 4618 3289 4652 3297
rect 4652 3289 4661 3297
rect 4809 3403 4818 3411
rect 4818 3403 4852 3411
rect 4852 3403 4861 3411
rect 4809 3359 4861 3403
rect 5009 3577 5061 3621
rect 5009 3569 5018 3577
rect 5018 3569 5052 3577
rect 5052 3569 5061 3577
rect 5209 3773 5218 3781
rect 5218 3773 5252 3781
rect 5252 3773 5261 3781
rect 5209 3729 5261 3773
rect 5409 3947 5461 3991
rect 5409 3939 5418 3947
rect 5418 3939 5452 3947
rect 5452 3939 5461 3947
rect 5609 4053 5618 4061
rect 5618 4053 5652 4061
rect 5652 4053 5661 4061
rect 5609 4009 5661 4053
rect 5809 4227 5861 4271
rect 5809 4219 5818 4227
rect 5818 4219 5852 4227
rect 5852 4219 5861 4227
rect 6009 4333 6018 4341
rect 6018 4333 6052 4341
rect 6052 4333 6061 4341
rect 6009 4289 6061 4333
rect 6209 4507 6261 4551
rect 6209 4499 6218 4507
rect 6218 4499 6252 4507
rect 6252 4499 6261 4507
rect 6409 4613 6418 4621
rect 6418 4613 6452 4621
rect 6452 4613 6461 4621
rect 6409 4569 6461 4613
rect 6507 4569 6559 4621
rect 5209 3684 5261 3693
rect 5209 3650 5218 3684
rect 5218 3650 5252 3684
rect 5252 3650 5261 3684
rect 5209 3641 5261 3650
rect 3609 2474 3661 2483
rect 3609 2440 3618 2474
rect 3618 2440 3652 2474
rect 3652 2440 3661 2474
rect 3609 2431 3661 2440
rect 2009 1264 2061 1273
rect 2009 1230 2018 1264
rect 2018 1230 2052 1264
rect 2052 1230 2061 1264
rect 2009 1221 2061 1230
rect 409 54 461 63
rect 409 20 418 54
rect 418 20 452 54
rect 452 20 461 54
rect 409 11 461 20
rect 309 -60 361 -15
rect 309 -67 318 -60
rect 318 -67 352 -60
rect 352 -67 361 -60
rect 109 -166 118 -143
rect 118 -166 152 -143
rect 152 -166 161 -143
rect 109 -195 161 -166
rect 125 -248 177 -239
rect 125 -282 134 -248
rect 134 -282 168 -248
rect 168 -282 177 -248
rect 125 -291 177 -282
rect 109 -363 161 -326
rect 109 -378 118 -363
rect 118 -378 152 -363
rect 152 -378 161 -363
rect 109 -397 118 -390
rect 118 -397 152 -390
rect 152 -397 161 -390
rect 109 -435 161 -397
rect 109 -442 118 -435
rect 118 -442 152 -435
rect 152 -442 161 -435
rect 109 -469 118 -454
rect 118 -469 152 -454
rect 152 -469 161 -454
rect 109 -506 161 -469
rect 309 -94 318 -79
rect 318 -94 352 -79
rect 352 -94 361 -79
rect 309 -131 361 -94
rect 409 -74 461 -22
rect 609 177 661 221
rect 609 169 618 177
rect 618 169 652 177
rect 652 169 661 177
rect 809 283 818 291
rect 818 283 852 291
rect 852 283 861 291
rect 809 239 861 283
rect 1009 457 1061 501
rect 1009 449 1018 457
rect 1018 449 1052 457
rect 1052 449 1061 457
rect 1209 563 1218 571
rect 1218 563 1252 571
rect 1252 563 1261 571
rect 1209 519 1261 563
rect 1409 737 1461 781
rect 1409 729 1418 737
rect 1418 729 1452 737
rect 1452 729 1461 737
rect 1609 843 1618 851
rect 1618 843 1652 851
rect 1652 843 1661 851
rect 1609 799 1661 843
rect 1809 1017 1861 1061
rect 1809 1009 1818 1017
rect 1818 1009 1852 1017
rect 1852 1009 1861 1017
rect 2009 1123 2018 1131
rect 2018 1123 2052 1131
rect 2052 1123 2061 1131
rect 2009 1079 2061 1123
rect 2209 1387 2261 1431
rect 2209 1379 2218 1387
rect 2218 1379 2252 1387
rect 2252 1379 2261 1387
rect 2409 1493 2418 1501
rect 2418 1493 2452 1501
rect 2452 1493 2461 1501
rect 2409 1449 2461 1493
rect 2609 1667 2661 1711
rect 2609 1659 2618 1667
rect 2618 1659 2652 1667
rect 2652 1659 2661 1667
rect 2809 1773 2818 1781
rect 2818 1773 2852 1781
rect 2852 1773 2861 1781
rect 2809 1729 2861 1773
rect 3009 1947 3061 1991
rect 3009 1939 3018 1947
rect 3018 1939 3052 1947
rect 3052 1939 3061 1947
rect 3209 2053 3218 2061
rect 3218 2053 3252 2061
rect 3252 2053 3261 2061
rect 3209 2009 3261 2053
rect 3409 2227 3461 2271
rect 3409 2219 3418 2227
rect 3418 2219 3452 2227
rect 3452 2219 3461 2227
rect 3609 2333 3618 2341
rect 3618 2333 3652 2341
rect 3652 2333 3661 2341
rect 3609 2289 3661 2333
rect 3809 2597 3861 2641
rect 3809 2589 3818 2597
rect 3818 2589 3852 2597
rect 3852 2589 3861 2597
rect 4009 2703 4018 2711
rect 4018 2703 4052 2711
rect 4052 2703 4061 2711
rect 4009 2659 4061 2703
rect 4209 2877 4261 2921
rect 4209 2869 4218 2877
rect 4218 2869 4252 2877
rect 4252 2869 4261 2877
rect 4409 2983 4418 2991
rect 4418 2983 4452 2991
rect 4452 2983 4461 2991
rect 4409 2939 4461 2983
rect 4609 3157 4661 3201
rect 4609 3149 4618 3157
rect 4618 3149 4652 3157
rect 4652 3149 4661 3157
rect 4809 3263 4818 3271
rect 4818 3263 4852 3271
rect 4852 3263 4861 3271
rect 4809 3219 4861 3263
rect 5009 3437 5061 3481
rect 5009 3429 5018 3437
rect 5018 3429 5052 3437
rect 5052 3429 5061 3437
rect 5209 3543 5218 3551
rect 5218 3543 5252 3551
rect 5252 3543 5261 3551
rect 5209 3499 5261 3543
rect 5409 3807 5461 3851
rect 5409 3799 5418 3807
rect 5418 3799 5452 3807
rect 5452 3799 5461 3807
rect 5609 3913 5618 3921
rect 5618 3913 5652 3921
rect 5652 3913 5661 3921
rect 5609 3869 5661 3913
rect 5809 4087 5861 4131
rect 5809 4079 5818 4087
rect 5818 4079 5852 4087
rect 5852 4079 5861 4087
rect 6009 4193 6018 4201
rect 6018 4193 6052 4201
rect 6052 4193 6061 4201
rect 6009 4149 6061 4193
rect 6209 4367 6261 4411
rect 6209 4359 6218 4367
rect 6218 4359 6252 4367
rect 6252 4359 6261 4367
rect 6409 4473 6418 4481
rect 6418 4473 6452 4481
rect 6452 4473 6461 4481
rect 6409 4429 6461 4473
rect 6507 4429 6559 4481
rect 5409 3700 5461 3709
rect 5409 3666 5418 3700
rect 5418 3666 5452 3700
rect 5452 3666 5461 3700
rect 5409 3657 5461 3666
rect 3809 2490 3861 2499
rect 3809 2456 3818 2490
rect 3818 2456 3852 2490
rect 3852 2456 3861 2490
rect 3809 2447 3861 2456
rect 2209 1280 2261 1289
rect 2209 1246 2218 1280
rect 2218 1246 2252 1280
rect 2252 1246 2261 1280
rect 2209 1237 2261 1246
rect 609 70 661 79
rect 609 36 618 70
rect 618 36 652 70
rect 652 36 661 70
rect 609 27 661 36
rect 509 -60 561 -15
rect 509 -67 518 -60
rect 518 -67 552 -60
rect 552 -67 561 -60
rect 309 -166 318 -143
rect 318 -166 352 -143
rect 352 -166 361 -143
rect 309 -195 361 -166
rect 325 -248 377 -239
rect 325 -282 334 -248
rect 334 -282 368 -248
rect 368 -282 377 -248
rect 325 -291 377 -282
rect 309 -363 361 -326
rect 309 -378 318 -363
rect 318 -378 352 -363
rect 352 -378 361 -363
rect 309 -397 318 -390
rect 318 -397 352 -390
rect 352 -397 361 -390
rect 309 -435 361 -397
rect 309 -442 318 -435
rect 318 -442 352 -435
rect 352 -442 361 -435
rect 309 -469 318 -454
rect 318 -469 352 -454
rect 352 -469 361 -454
rect 309 -506 361 -469
rect 509 -94 518 -79
rect 518 -94 552 -79
rect 552 -94 561 -79
rect 509 -131 561 -94
rect 609 -74 661 -22
rect 809 143 818 151
rect 818 143 852 151
rect 852 143 861 151
rect 809 99 861 143
rect 1009 317 1061 361
rect 1009 309 1018 317
rect 1018 309 1052 317
rect 1052 309 1061 317
rect 1209 423 1218 431
rect 1218 423 1252 431
rect 1252 423 1261 431
rect 1209 379 1261 423
rect 1409 597 1461 641
rect 1409 589 1418 597
rect 1418 589 1452 597
rect 1452 589 1461 597
rect 1609 703 1618 711
rect 1618 703 1652 711
rect 1652 703 1661 711
rect 1609 659 1661 703
rect 1809 877 1861 921
rect 1809 869 1818 877
rect 1818 869 1852 877
rect 1852 869 1861 877
rect 2009 983 2018 991
rect 2018 983 2052 991
rect 2052 983 2061 991
rect 2009 939 2061 983
rect 2209 1157 2261 1201
rect 2209 1149 2218 1157
rect 2218 1149 2252 1157
rect 2252 1149 2261 1157
rect 2409 1353 2418 1361
rect 2418 1353 2452 1361
rect 2452 1353 2461 1361
rect 2409 1309 2461 1353
rect 2609 1527 2661 1571
rect 2609 1519 2618 1527
rect 2618 1519 2652 1527
rect 2652 1519 2661 1527
rect 2809 1633 2818 1641
rect 2818 1633 2852 1641
rect 2852 1633 2861 1641
rect 2809 1589 2861 1633
rect 3009 1807 3061 1851
rect 3009 1799 3018 1807
rect 3018 1799 3052 1807
rect 3052 1799 3061 1807
rect 3209 1913 3218 1921
rect 3218 1913 3252 1921
rect 3252 1913 3261 1921
rect 3209 1869 3261 1913
rect 3409 2087 3461 2131
rect 3409 2079 3418 2087
rect 3418 2079 3452 2087
rect 3452 2079 3461 2087
rect 3609 2193 3618 2201
rect 3618 2193 3652 2201
rect 3652 2193 3661 2201
rect 3609 2149 3661 2193
rect 3809 2367 3861 2411
rect 3809 2359 3818 2367
rect 3818 2359 3852 2367
rect 3852 2359 3861 2367
rect 4009 2563 4018 2571
rect 4018 2563 4052 2571
rect 4052 2563 4061 2571
rect 4009 2519 4061 2563
rect 4209 2737 4261 2781
rect 4209 2729 4218 2737
rect 4218 2729 4252 2737
rect 4252 2729 4261 2737
rect 4409 2843 4418 2851
rect 4418 2843 4452 2851
rect 4452 2843 4461 2851
rect 4409 2799 4461 2843
rect 4609 3017 4661 3061
rect 4609 3009 4618 3017
rect 4618 3009 4652 3017
rect 4652 3009 4661 3017
rect 4809 3123 4818 3131
rect 4818 3123 4852 3131
rect 4852 3123 4861 3131
rect 4809 3079 4861 3123
rect 5009 3297 5061 3341
rect 5009 3289 5018 3297
rect 5018 3289 5052 3297
rect 5052 3289 5061 3297
rect 5209 3403 5218 3411
rect 5218 3403 5252 3411
rect 5252 3403 5261 3411
rect 5209 3359 5261 3403
rect 5409 3577 5461 3621
rect 5409 3569 5418 3577
rect 5418 3569 5452 3577
rect 5452 3569 5461 3577
rect 5609 3773 5618 3781
rect 5618 3773 5652 3781
rect 5652 3773 5661 3781
rect 5609 3729 5661 3773
rect 5809 3947 5861 3991
rect 5809 3939 5818 3947
rect 5818 3939 5852 3947
rect 5852 3939 5861 3947
rect 6009 4053 6018 4061
rect 6018 4053 6052 4061
rect 6052 4053 6061 4061
rect 6009 4009 6061 4053
rect 6209 4227 6261 4271
rect 6209 4219 6218 4227
rect 6218 4219 6252 4227
rect 6252 4219 6261 4227
rect 6409 4333 6418 4341
rect 6418 4333 6452 4341
rect 6452 4333 6461 4341
rect 6409 4289 6461 4333
rect 6507 4289 6559 4341
rect 5609 3684 5661 3693
rect 5609 3650 5618 3684
rect 5618 3650 5652 3684
rect 5652 3650 5661 3684
rect 5609 3641 5661 3650
rect 4009 2474 4061 2483
rect 4009 2440 4018 2474
rect 4018 2440 4052 2474
rect 4052 2440 4061 2474
rect 4009 2431 4061 2440
rect 2409 1264 2461 1273
rect 2409 1230 2418 1264
rect 2418 1230 2452 1264
rect 2452 1230 2461 1264
rect 2409 1221 2461 1230
rect 809 54 861 63
rect 809 20 818 54
rect 818 20 852 54
rect 852 20 861 54
rect 809 11 861 20
rect 709 -60 761 -15
rect 709 -67 718 -60
rect 718 -67 752 -60
rect 752 -67 761 -60
rect 509 -166 518 -143
rect 518 -166 552 -143
rect 552 -166 561 -143
rect 509 -195 561 -166
rect 525 -248 577 -239
rect 525 -282 534 -248
rect 534 -282 568 -248
rect 568 -282 577 -248
rect 525 -291 577 -282
rect 509 -363 561 -326
rect 509 -378 518 -363
rect 518 -378 552 -363
rect 552 -378 561 -363
rect 509 -397 518 -390
rect 518 -397 552 -390
rect 552 -397 561 -390
rect 509 -435 561 -397
rect 509 -442 518 -435
rect 518 -442 552 -435
rect 552 -442 561 -435
rect 509 -469 518 -454
rect 518 -469 552 -454
rect 552 -469 561 -454
rect 509 -506 561 -469
rect 709 -94 718 -79
rect 718 -94 752 -79
rect 752 -94 761 -79
rect 709 -131 761 -94
rect 809 -74 861 -22
rect 1009 177 1061 221
rect 1009 169 1018 177
rect 1018 169 1052 177
rect 1052 169 1061 177
rect 1209 283 1218 291
rect 1218 283 1252 291
rect 1252 283 1261 291
rect 1209 239 1261 283
rect 1409 457 1461 501
rect 1409 449 1418 457
rect 1418 449 1452 457
rect 1452 449 1461 457
rect 1609 563 1618 571
rect 1618 563 1652 571
rect 1652 563 1661 571
rect 1609 519 1661 563
rect 1809 737 1861 781
rect 1809 729 1818 737
rect 1818 729 1852 737
rect 1852 729 1861 737
rect 2009 843 2018 851
rect 2018 843 2052 851
rect 2052 843 2061 851
rect 2009 799 2061 843
rect 2209 1017 2261 1061
rect 2209 1009 2218 1017
rect 2218 1009 2252 1017
rect 2252 1009 2261 1017
rect 2409 1123 2418 1131
rect 2418 1123 2452 1131
rect 2452 1123 2461 1131
rect 2409 1079 2461 1123
rect 2609 1387 2661 1431
rect 2609 1379 2618 1387
rect 2618 1379 2652 1387
rect 2652 1379 2661 1387
rect 2809 1493 2818 1501
rect 2818 1493 2852 1501
rect 2852 1493 2861 1501
rect 2809 1449 2861 1493
rect 3009 1667 3061 1711
rect 3009 1659 3018 1667
rect 3018 1659 3052 1667
rect 3052 1659 3061 1667
rect 3209 1773 3218 1781
rect 3218 1773 3252 1781
rect 3252 1773 3261 1781
rect 3209 1729 3261 1773
rect 3409 1947 3461 1991
rect 3409 1939 3418 1947
rect 3418 1939 3452 1947
rect 3452 1939 3461 1947
rect 3609 2053 3618 2061
rect 3618 2053 3652 2061
rect 3652 2053 3661 2061
rect 3609 2009 3661 2053
rect 3809 2227 3861 2271
rect 3809 2219 3818 2227
rect 3818 2219 3852 2227
rect 3852 2219 3861 2227
rect 4009 2333 4018 2341
rect 4018 2333 4052 2341
rect 4052 2333 4061 2341
rect 4009 2289 4061 2333
rect 4209 2597 4261 2641
rect 4209 2589 4218 2597
rect 4218 2589 4252 2597
rect 4252 2589 4261 2597
rect 4409 2703 4418 2711
rect 4418 2703 4452 2711
rect 4452 2703 4461 2711
rect 4409 2659 4461 2703
rect 4609 2877 4661 2921
rect 4609 2869 4618 2877
rect 4618 2869 4652 2877
rect 4652 2869 4661 2877
rect 4809 2983 4818 2991
rect 4818 2983 4852 2991
rect 4852 2983 4861 2991
rect 4809 2939 4861 2983
rect 5009 3157 5061 3201
rect 5009 3149 5018 3157
rect 5018 3149 5052 3157
rect 5052 3149 5061 3157
rect 5209 3263 5218 3271
rect 5218 3263 5252 3271
rect 5252 3263 5261 3271
rect 5209 3219 5261 3263
rect 5409 3437 5461 3481
rect 5409 3429 5418 3437
rect 5418 3429 5452 3437
rect 5452 3429 5461 3437
rect 5609 3543 5618 3551
rect 5618 3543 5652 3551
rect 5652 3543 5661 3551
rect 5609 3499 5661 3543
rect 5809 3807 5861 3851
rect 5809 3799 5818 3807
rect 5818 3799 5852 3807
rect 5852 3799 5861 3807
rect 6009 3913 6018 3921
rect 6018 3913 6052 3921
rect 6052 3913 6061 3921
rect 6009 3869 6061 3913
rect 6209 4087 6261 4131
rect 6209 4079 6218 4087
rect 6218 4079 6252 4087
rect 6252 4079 6261 4087
rect 6409 4193 6418 4201
rect 6418 4193 6452 4201
rect 6452 4193 6461 4201
rect 6409 4149 6461 4193
rect 6507 4149 6559 4201
rect 5809 3700 5861 3709
rect 5809 3666 5818 3700
rect 5818 3666 5852 3700
rect 5852 3666 5861 3700
rect 5809 3657 5861 3666
rect 4209 2490 4261 2499
rect 4209 2456 4218 2490
rect 4218 2456 4252 2490
rect 4252 2456 4261 2490
rect 4209 2447 4261 2456
rect 2609 1280 2661 1289
rect 2609 1246 2618 1280
rect 2618 1246 2652 1280
rect 2652 1246 2661 1280
rect 2609 1237 2661 1246
rect 1009 70 1061 79
rect 1009 36 1018 70
rect 1018 36 1052 70
rect 1052 36 1061 70
rect 1009 27 1061 36
rect 909 -60 961 -15
rect 909 -67 918 -60
rect 918 -67 952 -60
rect 952 -67 961 -60
rect 709 -166 718 -143
rect 718 -166 752 -143
rect 752 -166 761 -143
rect 709 -195 761 -166
rect 725 -248 777 -239
rect 725 -282 734 -248
rect 734 -282 768 -248
rect 768 -282 777 -248
rect 725 -291 777 -282
rect 709 -363 761 -326
rect 709 -378 718 -363
rect 718 -378 752 -363
rect 752 -378 761 -363
rect 709 -397 718 -390
rect 718 -397 752 -390
rect 752 -397 761 -390
rect 709 -435 761 -397
rect 709 -442 718 -435
rect 718 -442 752 -435
rect 752 -442 761 -435
rect 709 -469 718 -454
rect 718 -469 752 -454
rect 752 -469 761 -454
rect 709 -506 761 -469
rect 909 -94 918 -79
rect 918 -94 952 -79
rect 952 -94 961 -79
rect 909 -131 961 -94
rect 1009 -74 1061 -22
rect 1209 143 1218 151
rect 1218 143 1252 151
rect 1252 143 1261 151
rect 1209 99 1261 143
rect 1409 317 1461 361
rect 1409 309 1418 317
rect 1418 309 1452 317
rect 1452 309 1461 317
rect 1609 423 1618 431
rect 1618 423 1652 431
rect 1652 423 1661 431
rect 1609 379 1661 423
rect 1809 597 1861 641
rect 1809 589 1818 597
rect 1818 589 1852 597
rect 1852 589 1861 597
rect 2009 703 2018 711
rect 2018 703 2052 711
rect 2052 703 2061 711
rect 2009 659 2061 703
rect 2209 877 2261 921
rect 2209 869 2218 877
rect 2218 869 2252 877
rect 2252 869 2261 877
rect 2409 983 2418 991
rect 2418 983 2452 991
rect 2452 983 2461 991
rect 2409 939 2461 983
rect 2609 1157 2661 1201
rect 2609 1149 2618 1157
rect 2618 1149 2652 1157
rect 2652 1149 2661 1157
rect 2809 1353 2818 1361
rect 2818 1353 2852 1361
rect 2852 1353 2861 1361
rect 2809 1309 2861 1353
rect 3009 1527 3061 1571
rect 3009 1519 3018 1527
rect 3018 1519 3052 1527
rect 3052 1519 3061 1527
rect 3209 1633 3218 1641
rect 3218 1633 3252 1641
rect 3252 1633 3261 1641
rect 3209 1589 3261 1633
rect 3409 1807 3461 1851
rect 3409 1799 3418 1807
rect 3418 1799 3452 1807
rect 3452 1799 3461 1807
rect 3609 1913 3618 1921
rect 3618 1913 3652 1921
rect 3652 1913 3661 1921
rect 3609 1869 3661 1913
rect 3809 2087 3861 2131
rect 3809 2079 3818 2087
rect 3818 2079 3852 2087
rect 3852 2079 3861 2087
rect 4009 2193 4018 2201
rect 4018 2193 4052 2201
rect 4052 2193 4061 2201
rect 4009 2149 4061 2193
rect 4209 2367 4261 2411
rect 4209 2359 4218 2367
rect 4218 2359 4252 2367
rect 4252 2359 4261 2367
rect 4409 2563 4418 2571
rect 4418 2563 4452 2571
rect 4452 2563 4461 2571
rect 4409 2519 4461 2563
rect 4609 2737 4661 2781
rect 4609 2729 4618 2737
rect 4618 2729 4652 2737
rect 4652 2729 4661 2737
rect 4809 2843 4818 2851
rect 4818 2843 4852 2851
rect 4852 2843 4861 2851
rect 4809 2799 4861 2843
rect 5009 3017 5061 3061
rect 5009 3009 5018 3017
rect 5018 3009 5052 3017
rect 5052 3009 5061 3017
rect 5209 3123 5218 3131
rect 5218 3123 5252 3131
rect 5252 3123 5261 3131
rect 5209 3079 5261 3123
rect 5409 3297 5461 3341
rect 5409 3289 5418 3297
rect 5418 3289 5452 3297
rect 5452 3289 5461 3297
rect 5609 3403 5618 3411
rect 5618 3403 5652 3411
rect 5652 3403 5661 3411
rect 5609 3359 5661 3403
rect 5809 3577 5861 3621
rect 5809 3569 5818 3577
rect 5818 3569 5852 3577
rect 5852 3569 5861 3577
rect 6009 3773 6018 3781
rect 6018 3773 6052 3781
rect 6052 3773 6061 3781
rect 6009 3729 6061 3773
rect 6209 3947 6261 3991
rect 6209 3939 6218 3947
rect 6218 3939 6252 3947
rect 6252 3939 6261 3947
rect 6409 4053 6418 4061
rect 6418 4053 6452 4061
rect 6452 4053 6461 4061
rect 6409 4009 6461 4053
rect 6507 4009 6559 4061
rect 6009 3684 6061 3693
rect 6009 3650 6018 3684
rect 6018 3650 6052 3684
rect 6052 3650 6061 3684
rect 6009 3641 6061 3650
rect 4409 2474 4461 2483
rect 4409 2440 4418 2474
rect 4418 2440 4452 2474
rect 4452 2440 4461 2474
rect 4409 2431 4461 2440
rect 2809 1264 2861 1273
rect 2809 1230 2818 1264
rect 2818 1230 2852 1264
rect 2852 1230 2861 1264
rect 2809 1221 2861 1230
rect 1209 54 1261 63
rect 1209 20 1218 54
rect 1218 20 1252 54
rect 1252 20 1261 54
rect 1209 11 1261 20
rect 1109 -60 1161 -15
rect 1109 -67 1118 -60
rect 1118 -67 1152 -60
rect 1152 -67 1161 -60
rect 909 -166 918 -143
rect 918 -166 952 -143
rect 952 -166 961 -143
rect 909 -195 961 -166
rect 925 -248 977 -239
rect 925 -282 934 -248
rect 934 -282 968 -248
rect 968 -282 977 -248
rect 925 -291 977 -282
rect 909 -363 961 -326
rect 909 -378 918 -363
rect 918 -378 952 -363
rect 952 -378 961 -363
rect 909 -397 918 -390
rect 918 -397 952 -390
rect 952 -397 961 -390
rect 909 -435 961 -397
rect 909 -442 918 -435
rect 918 -442 952 -435
rect 952 -442 961 -435
rect 909 -469 918 -454
rect 918 -469 952 -454
rect 952 -469 961 -454
rect 909 -506 961 -469
rect 1109 -94 1118 -79
rect 1118 -94 1152 -79
rect 1152 -94 1161 -79
rect 1109 -131 1161 -94
rect 1209 -74 1261 -22
rect 1409 177 1461 221
rect 1409 169 1418 177
rect 1418 169 1452 177
rect 1452 169 1461 177
rect 1609 283 1618 291
rect 1618 283 1652 291
rect 1652 283 1661 291
rect 1609 239 1661 283
rect 1809 457 1861 501
rect 1809 449 1818 457
rect 1818 449 1852 457
rect 1852 449 1861 457
rect 2009 563 2018 571
rect 2018 563 2052 571
rect 2052 563 2061 571
rect 2009 519 2061 563
rect 2209 737 2261 781
rect 2209 729 2218 737
rect 2218 729 2252 737
rect 2252 729 2261 737
rect 2409 843 2418 851
rect 2418 843 2452 851
rect 2452 843 2461 851
rect 2409 799 2461 843
rect 2609 1017 2661 1061
rect 2609 1009 2618 1017
rect 2618 1009 2652 1017
rect 2652 1009 2661 1017
rect 2809 1123 2818 1131
rect 2818 1123 2852 1131
rect 2852 1123 2861 1131
rect 2809 1079 2861 1123
rect 3009 1387 3061 1431
rect 3009 1379 3018 1387
rect 3018 1379 3052 1387
rect 3052 1379 3061 1387
rect 3209 1493 3218 1501
rect 3218 1493 3252 1501
rect 3252 1493 3261 1501
rect 3209 1449 3261 1493
rect 3409 1667 3461 1711
rect 3409 1659 3418 1667
rect 3418 1659 3452 1667
rect 3452 1659 3461 1667
rect 3609 1773 3618 1781
rect 3618 1773 3652 1781
rect 3652 1773 3661 1781
rect 3609 1729 3661 1773
rect 3809 1947 3861 1991
rect 3809 1939 3818 1947
rect 3818 1939 3852 1947
rect 3852 1939 3861 1947
rect 4009 2053 4018 2061
rect 4018 2053 4052 2061
rect 4052 2053 4061 2061
rect 4009 2009 4061 2053
rect 4209 2227 4261 2271
rect 4209 2219 4218 2227
rect 4218 2219 4252 2227
rect 4252 2219 4261 2227
rect 4409 2333 4418 2341
rect 4418 2333 4452 2341
rect 4452 2333 4461 2341
rect 4409 2289 4461 2333
rect 4609 2597 4661 2641
rect 4609 2589 4618 2597
rect 4618 2589 4652 2597
rect 4652 2589 4661 2597
rect 4809 2703 4818 2711
rect 4818 2703 4852 2711
rect 4852 2703 4861 2711
rect 4809 2659 4861 2703
rect 5009 2877 5061 2921
rect 5009 2869 5018 2877
rect 5018 2869 5052 2877
rect 5052 2869 5061 2877
rect 5209 2983 5218 2991
rect 5218 2983 5252 2991
rect 5252 2983 5261 2991
rect 5209 2939 5261 2983
rect 5409 3157 5461 3201
rect 5409 3149 5418 3157
rect 5418 3149 5452 3157
rect 5452 3149 5461 3157
rect 5609 3263 5618 3271
rect 5618 3263 5652 3271
rect 5652 3263 5661 3271
rect 5609 3219 5661 3263
rect 5809 3437 5861 3481
rect 5809 3429 5818 3437
rect 5818 3429 5852 3437
rect 5852 3429 5861 3437
rect 6009 3543 6018 3551
rect 6018 3543 6052 3551
rect 6052 3543 6061 3551
rect 6009 3499 6061 3543
rect 6209 3807 6261 3851
rect 6209 3799 6218 3807
rect 6218 3799 6252 3807
rect 6252 3799 6261 3807
rect 6409 3913 6418 3921
rect 6418 3913 6452 3921
rect 6452 3913 6461 3921
rect 6409 3869 6461 3913
rect 6507 3869 6559 3921
rect 6209 3700 6261 3709
rect 6209 3666 6218 3700
rect 6218 3666 6252 3700
rect 6252 3666 6261 3700
rect 6209 3657 6261 3666
rect 4609 2490 4661 2499
rect 4609 2456 4618 2490
rect 4618 2456 4652 2490
rect 4652 2456 4661 2490
rect 4609 2447 4661 2456
rect 3009 1280 3061 1289
rect 3009 1246 3018 1280
rect 3018 1246 3052 1280
rect 3052 1246 3061 1280
rect 3009 1237 3061 1246
rect 1409 70 1461 79
rect 1409 36 1418 70
rect 1418 36 1452 70
rect 1452 36 1461 70
rect 1409 27 1461 36
rect 1309 -60 1361 -15
rect 1309 -67 1318 -60
rect 1318 -67 1352 -60
rect 1352 -67 1361 -60
rect 1109 -166 1118 -143
rect 1118 -166 1152 -143
rect 1152 -166 1161 -143
rect 1109 -195 1161 -166
rect 1125 -248 1177 -239
rect 1125 -282 1134 -248
rect 1134 -282 1168 -248
rect 1168 -282 1177 -248
rect 1125 -291 1177 -282
rect 1109 -363 1161 -326
rect 1109 -378 1118 -363
rect 1118 -378 1152 -363
rect 1152 -378 1161 -363
rect 1109 -397 1118 -390
rect 1118 -397 1152 -390
rect 1152 -397 1161 -390
rect 1109 -435 1161 -397
rect 1109 -442 1118 -435
rect 1118 -442 1152 -435
rect 1152 -442 1161 -435
rect 1109 -469 1118 -454
rect 1118 -469 1152 -454
rect 1152 -469 1161 -454
rect 1109 -506 1161 -469
rect 1309 -94 1318 -79
rect 1318 -94 1352 -79
rect 1352 -94 1361 -79
rect 1309 -131 1361 -94
rect 1409 -74 1461 -22
rect 1609 143 1618 151
rect 1618 143 1652 151
rect 1652 143 1661 151
rect 1609 99 1661 143
rect 1809 317 1861 361
rect 1809 309 1818 317
rect 1818 309 1852 317
rect 1852 309 1861 317
rect 2009 423 2018 431
rect 2018 423 2052 431
rect 2052 423 2061 431
rect 2009 379 2061 423
rect 2209 597 2261 641
rect 2209 589 2218 597
rect 2218 589 2252 597
rect 2252 589 2261 597
rect 2409 703 2418 711
rect 2418 703 2452 711
rect 2452 703 2461 711
rect 2409 659 2461 703
rect 2609 877 2661 921
rect 2609 869 2618 877
rect 2618 869 2652 877
rect 2652 869 2661 877
rect 2809 983 2818 991
rect 2818 983 2852 991
rect 2852 983 2861 991
rect 2809 939 2861 983
rect 3009 1157 3061 1201
rect 3009 1149 3018 1157
rect 3018 1149 3052 1157
rect 3052 1149 3061 1157
rect 3209 1353 3218 1361
rect 3218 1353 3252 1361
rect 3252 1353 3261 1361
rect 3209 1309 3261 1353
rect 3409 1527 3461 1571
rect 3409 1519 3418 1527
rect 3418 1519 3452 1527
rect 3452 1519 3461 1527
rect 3609 1633 3618 1641
rect 3618 1633 3652 1641
rect 3652 1633 3661 1641
rect 3609 1589 3661 1633
rect 3809 1807 3861 1851
rect 3809 1799 3818 1807
rect 3818 1799 3852 1807
rect 3852 1799 3861 1807
rect 4009 1913 4018 1921
rect 4018 1913 4052 1921
rect 4052 1913 4061 1921
rect 4009 1869 4061 1913
rect 4209 2087 4261 2131
rect 4209 2079 4218 2087
rect 4218 2079 4252 2087
rect 4252 2079 4261 2087
rect 4409 2193 4418 2201
rect 4418 2193 4452 2201
rect 4452 2193 4461 2201
rect 4409 2149 4461 2193
rect 4609 2367 4661 2411
rect 4609 2359 4618 2367
rect 4618 2359 4652 2367
rect 4652 2359 4661 2367
rect 4809 2563 4818 2571
rect 4818 2563 4852 2571
rect 4852 2563 4861 2571
rect 4809 2519 4861 2563
rect 5009 2737 5061 2781
rect 5009 2729 5018 2737
rect 5018 2729 5052 2737
rect 5052 2729 5061 2737
rect 5209 2843 5218 2851
rect 5218 2843 5252 2851
rect 5252 2843 5261 2851
rect 5209 2799 5261 2843
rect 5409 3017 5461 3061
rect 5409 3009 5418 3017
rect 5418 3009 5452 3017
rect 5452 3009 5461 3017
rect 5609 3123 5618 3131
rect 5618 3123 5652 3131
rect 5652 3123 5661 3131
rect 5609 3079 5661 3123
rect 5809 3297 5861 3341
rect 5809 3289 5818 3297
rect 5818 3289 5852 3297
rect 5852 3289 5861 3297
rect 6009 3403 6018 3411
rect 6018 3403 6052 3411
rect 6052 3403 6061 3411
rect 6009 3359 6061 3403
rect 6209 3577 6261 3621
rect 6209 3569 6218 3577
rect 6218 3569 6252 3577
rect 6252 3569 6261 3577
rect 6409 3773 6418 3781
rect 6418 3773 6452 3781
rect 6452 3773 6461 3781
rect 6409 3729 6461 3773
rect 6507 3729 6559 3781
rect 4809 2474 4861 2483
rect 4809 2440 4818 2474
rect 4818 2440 4852 2474
rect 4852 2440 4861 2474
rect 4809 2431 4861 2440
rect 3209 1264 3261 1273
rect 3209 1230 3218 1264
rect 3218 1230 3252 1264
rect 3252 1230 3261 1264
rect 3209 1221 3261 1230
rect 1609 54 1661 63
rect 1609 20 1618 54
rect 1618 20 1652 54
rect 1652 20 1661 54
rect 1609 11 1661 20
rect 1509 -60 1561 -15
rect 1509 -67 1518 -60
rect 1518 -67 1552 -60
rect 1552 -67 1561 -60
rect 1309 -166 1318 -143
rect 1318 -166 1352 -143
rect 1352 -166 1361 -143
rect 1309 -195 1361 -166
rect 1325 -248 1377 -239
rect 1325 -282 1334 -248
rect 1334 -282 1368 -248
rect 1368 -282 1377 -248
rect 1325 -291 1377 -282
rect 1309 -363 1361 -326
rect 1309 -378 1318 -363
rect 1318 -378 1352 -363
rect 1352 -378 1361 -363
rect 1309 -397 1318 -390
rect 1318 -397 1352 -390
rect 1352 -397 1361 -390
rect 1309 -435 1361 -397
rect 1309 -442 1318 -435
rect 1318 -442 1352 -435
rect 1352 -442 1361 -435
rect 1309 -469 1318 -454
rect 1318 -469 1352 -454
rect 1352 -469 1361 -454
rect 1309 -506 1361 -469
rect 1509 -94 1518 -79
rect 1518 -94 1552 -79
rect 1552 -94 1561 -79
rect 1509 -131 1561 -94
rect 1609 -74 1661 -22
rect 1809 177 1861 221
rect 1809 169 1818 177
rect 1818 169 1852 177
rect 1852 169 1861 177
rect 2009 283 2018 291
rect 2018 283 2052 291
rect 2052 283 2061 291
rect 2009 239 2061 283
rect 2209 457 2261 501
rect 2209 449 2218 457
rect 2218 449 2252 457
rect 2252 449 2261 457
rect 2409 563 2418 571
rect 2418 563 2452 571
rect 2452 563 2461 571
rect 2409 519 2461 563
rect 2609 737 2661 781
rect 2609 729 2618 737
rect 2618 729 2652 737
rect 2652 729 2661 737
rect 2809 843 2818 851
rect 2818 843 2852 851
rect 2852 843 2861 851
rect 2809 799 2861 843
rect 3009 1017 3061 1061
rect 3009 1009 3018 1017
rect 3018 1009 3052 1017
rect 3052 1009 3061 1017
rect 3209 1123 3218 1131
rect 3218 1123 3252 1131
rect 3252 1123 3261 1131
rect 3209 1079 3261 1123
rect 3409 1387 3461 1431
rect 3409 1379 3418 1387
rect 3418 1379 3452 1387
rect 3452 1379 3461 1387
rect 3609 1493 3618 1501
rect 3618 1493 3652 1501
rect 3652 1493 3661 1501
rect 3609 1449 3661 1493
rect 3809 1667 3861 1711
rect 3809 1659 3818 1667
rect 3818 1659 3852 1667
rect 3852 1659 3861 1667
rect 4009 1773 4018 1781
rect 4018 1773 4052 1781
rect 4052 1773 4061 1781
rect 4009 1729 4061 1773
rect 4209 1947 4261 1991
rect 4209 1939 4218 1947
rect 4218 1939 4252 1947
rect 4252 1939 4261 1947
rect 4409 2053 4418 2061
rect 4418 2053 4452 2061
rect 4452 2053 4461 2061
rect 4409 2009 4461 2053
rect 4609 2227 4661 2271
rect 4609 2219 4618 2227
rect 4618 2219 4652 2227
rect 4652 2219 4661 2227
rect 4809 2333 4818 2341
rect 4818 2333 4852 2341
rect 4852 2333 4861 2341
rect 4809 2289 4861 2333
rect 5009 2597 5061 2641
rect 5009 2589 5018 2597
rect 5018 2589 5052 2597
rect 5052 2589 5061 2597
rect 5209 2703 5218 2711
rect 5218 2703 5252 2711
rect 5252 2703 5261 2711
rect 5209 2659 5261 2703
rect 5409 2877 5461 2921
rect 5409 2869 5418 2877
rect 5418 2869 5452 2877
rect 5452 2869 5461 2877
rect 5609 2983 5618 2991
rect 5618 2983 5652 2991
rect 5652 2983 5661 2991
rect 5609 2939 5661 2983
rect 5809 3157 5861 3201
rect 5809 3149 5818 3157
rect 5818 3149 5852 3157
rect 5852 3149 5861 3157
rect 6009 3263 6018 3271
rect 6018 3263 6052 3271
rect 6052 3263 6061 3271
rect 6009 3219 6061 3263
rect 6209 3437 6261 3481
rect 6209 3429 6218 3437
rect 6218 3429 6252 3437
rect 6252 3429 6261 3437
rect 6409 3543 6418 3551
rect 6418 3543 6452 3551
rect 6452 3543 6461 3551
rect 6409 3499 6461 3543
rect 6507 3499 6559 3551
rect 5009 2490 5061 2499
rect 5009 2456 5018 2490
rect 5018 2456 5052 2490
rect 5052 2456 5061 2490
rect 5009 2447 5061 2456
rect 3409 1280 3461 1289
rect 3409 1246 3418 1280
rect 3418 1246 3452 1280
rect 3452 1246 3461 1280
rect 3409 1237 3461 1246
rect 1809 70 1861 79
rect 1809 36 1818 70
rect 1818 36 1852 70
rect 1852 36 1861 70
rect 1809 27 1861 36
rect 1709 -60 1761 -15
rect 1709 -67 1718 -60
rect 1718 -67 1752 -60
rect 1752 -67 1761 -60
rect 1509 -166 1518 -143
rect 1518 -166 1552 -143
rect 1552 -166 1561 -143
rect 1509 -195 1561 -166
rect 1525 -248 1577 -239
rect 1525 -282 1534 -248
rect 1534 -282 1568 -248
rect 1568 -282 1577 -248
rect 1525 -291 1577 -282
rect 1509 -363 1561 -326
rect 1509 -378 1518 -363
rect 1518 -378 1552 -363
rect 1552 -378 1561 -363
rect 1509 -397 1518 -390
rect 1518 -397 1552 -390
rect 1552 -397 1561 -390
rect 1509 -435 1561 -397
rect 1509 -442 1518 -435
rect 1518 -442 1552 -435
rect 1552 -442 1561 -435
rect 1509 -469 1518 -454
rect 1518 -469 1552 -454
rect 1552 -469 1561 -454
rect 1509 -506 1561 -469
rect 1709 -94 1718 -79
rect 1718 -94 1752 -79
rect 1752 -94 1761 -79
rect 1709 -131 1761 -94
rect 1809 -74 1861 -22
rect 2009 143 2018 151
rect 2018 143 2052 151
rect 2052 143 2061 151
rect 2009 99 2061 143
rect 2209 317 2261 361
rect 2209 309 2218 317
rect 2218 309 2252 317
rect 2252 309 2261 317
rect 2409 423 2418 431
rect 2418 423 2452 431
rect 2452 423 2461 431
rect 2409 379 2461 423
rect 2609 597 2661 641
rect 2609 589 2618 597
rect 2618 589 2652 597
rect 2652 589 2661 597
rect 2809 703 2818 711
rect 2818 703 2852 711
rect 2852 703 2861 711
rect 2809 659 2861 703
rect 3009 877 3061 921
rect 3009 869 3018 877
rect 3018 869 3052 877
rect 3052 869 3061 877
rect 3209 983 3218 991
rect 3218 983 3252 991
rect 3252 983 3261 991
rect 3209 939 3261 983
rect 3409 1157 3461 1201
rect 3409 1149 3418 1157
rect 3418 1149 3452 1157
rect 3452 1149 3461 1157
rect 3609 1353 3618 1361
rect 3618 1353 3652 1361
rect 3652 1353 3661 1361
rect 3609 1309 3661 1353
rect 3809 1527 3861 1571
rect 3809 1519 3818 1527
rect 3818 1519 3852 1527
rect 3852 1519 3861 1527
rect 4009 1633 4018 1641
rect 4018 1633 4052 1641
rect 4052 1633 4061 1641
rect 4009 1589 4061 1633
rect 4209 1807 4261 1851
rect 4209 1799 4218 1807
rect 4218 1799 4252 1807
rect 4252 1799 4261 1807
rect 4409 1913 4418 1921
rect 4418 1913 4452 1921
rect 4452 1913 4461 1921
rect 4409 1869 4461 1913
rect 4609 2087 4661 2131
rect 4609 2079 4618 2087
rect 4618 2079 4652 2087
rect 4652 2079 4661 2087
rect 4809 2193 4818 2201
rect 4818 2193 4852 2201
rect 4852 2193 4861 2201
rect 4809 2149 4861 2193
rect 5009 2367 5061 2411
rect 5009 2359 5018 2367
rect 5018 2359 5052 2367
rect 5052 2359 5061 2367
rect 5209 2563 5218 2571
rect 5218 2563 5252 2571
rect 5252 2563 5261 2571
rect 5209 2519 5261 2563
rect 5409 2737 5461 2781
rect 5409 2729 5418 2737
rect 5418 2729 5452 2737
rect 5452 2729 5461 2737
rect 5609 2843 5618 2851
rect 5618 2843 5652 2851
rect 5652 2843 5661 2851
rect 5609 2799 5661 2843
rect 5809 3017 5861 3061
rect 5809 3009 5818 3017
rect 5818 3009 5852 3017
rect 5852 3009 5861 3017
rect 6009 3123 6018 3131
rect 6018 3123 6052 3131
rect 6052 3123 6061 3131
rect 6009 3079 6061 3123
rect 6209 3297 6261 3341
rect 6209 3289 6218 3297
rect 6218 3289 6252 3297
rect 6252 3289 6261 3297
rect 6409 3403 6418 3411
rect 6418 3403 6452 3411
rect 6452 3403 6461 3411
rect 6409 3359 6461 3403
rect 6507 3359 6559 3411
rect 5209 2474 5261 2483
rect 5209 2440 5218 2474
rect 5218 2440 5252 2474
rect 5252 2440 5261 2474
rect 5209 2431 5261 2440
rect 3609 1264 3661 1273
rect 3609 1230 3618 1264
rect 3618 1230 3652 1264
rect 3652 1230 3661 1264
rect 3609 1221 3661 1230
rect 2009 54 2061 63
rect 2009 20 2018 54
rect 2018 20 2052 54
rect 2052 20 2061 54
rect 2009 11 2061 20
rect 1909 -60 1961 -15
rect 1909 -67 1918 -60
rect 1918 -67 1952 -60
rect 1952 -67 1961 -60
rect 1709 -166 1718 -143
rect 1718 -166 1752 -143
rect 1752 -166 1761 -143
rect 1709 -195 1761 -166
rect 1725 -248 1777 -239
rect 1725 -282 1734 -248
rect 1734 -282 1768 -248
rect 1768 -282 1777 -248
rect 1725 -291 1777 -282
rect 1709 -363 1761 -326
rect 1709 -378 1718 -363
rect 1718 -378 1752 -363
rect 1752 -378 1761 -363
rect 1709 -397 1718 -390
rect 1718 -397 1752 -390
rect 1752 -397 1761 -390
rect 1709 -435 1761 -397
rect 1709 -442 1718 -435
rect 1718 -442 1752 -435
rect 1752 -442 1761 -435
rect 1709 -469 1718 -454
rect 1718 -469 1752 -454
rect 1752 -469 1761 -454
rect 1709 -506 1761 -469
rect 1909 -94 1918 -79
rect 1918 -94 1952 -79
rect 1952 -94 1961 -79
rect 1909 -131 1961 -94
rect 2009 -74 2061 -22
rect 2209 177 2261 221
rect 2209 169 2218 177
rect 2218 169 2252 177
rect 2252 169 2261 177
rect 2409 283 2418 291
rect 2418 283 2452 291
rect 2452 283 2461 291
rect 2409 239 2461 283
rect 2609 457 2661 501
rect 2609 449 2618 457
rect 2618 449 2652 457
rect 2652 449 2661 457
rect 2809 563 2818 571
rect 2818 563 2852 571
rect 2852 563 2861 571
rect 2809 519 2861 563
rect 3009 737 3061 781
rect 3009 729 3018 737
rect 3018 729 3052 737
rect 3052 729 3061 737
rect 3209 843 3218 851
rect 3218 843 3252 851
rect 3252 843 3261 851
rect 3209 799 3261 843
rect 3409 1017 3461 1061
rect 3409 1009 3418 1017
rect 3418 1009 3452 1017
rect 3452 1009 3461 1017
rect 3609 1123 3618 1131
rect 3618 1123 3652 1131
rect 3652 1123 3661 1131
rect 3609 1079 3661 1123
rect 3809 1387 3861 1431
rect 3809 1379 3818 1387
rect 3818 1379 3852 1387
rect 3852 1379 3861 1387
rect 4009 1493 4018 1501
rect 4018 1493 4052 1501
rect 4052 1493 4061 1501
rect 4009 1449 4061 1493
rect 4209 1667 4261 1711
rect 4209 1659 4218 1667
rect 4218 1659 4252 1667
rect 4252 1659 4261 1667
rect 4409 1773 4418 1781
rect 4418 1773 4452 1781
rect 4452 1773 4461 1781
rect 4409 1729 4461 1773
rect 4609 1947 4661 1991
rect 4609 1939 4618 1947
rect 4618 1939 4652 1947
rect 4652 1939 4661 1947
rect 4809 2053 4818 2061
rect 4818 2053 4852 2061
rect 4852 2053 4861 2061
rect 4809 2009 4861 2053
rect 5009 2227 5061 2271
rect 5009 2219 5018 2227
rect 5018 2219 5052 2227
rect 5052 2219 5061 2227
rect 5209 2333 5218 2341
rect 5218 2333 5252 2341
rect 5252 2333 5261 2341
rect 5209 2289 5261 2333
rect 5409 2597 5461 2641
rect 5409 2589 5418 2597
rect 5418 2589 5452 2597
rect 5452 2589 5461 2597
rect 5609 2703 5618 2711
rect 5618 2703 5652 2711
rect 5652 2703 5661 2711
rect 5609 2659 5661 2703
rect 5809 2877 5861 2921
rect 5809 2869 5818 2877
rect 5818 2869 5852 2877
rect 5852 2869 5861 2877
rect 6009 2983 6018 2991
rect 6018 2983 6052 2991
rect 6052 2983 6061 2991
rect 6009 2939 6061 2983
rect 6209 3157 6261 3201
rect 6209 3149 6218 3157
rect 6218 3149 6252 3157
rect 6252 3149 6261 3157
rect 6409 3263 6418 3271
rect 6418 3263 6452 3271
rect 6452 3263 6461 3271
rect 6409 3219 6461 3263
rect 6507 3219 6559 3271
rect 5409 2490 5461 2499
rect 5409 2456 5418 2490
rect 5418 2456 5452 2490
rect 5452 2456 5461 2490
rect 5409 2447 5461 2456
rect 3809 1280 3861 1289
rect 3809 1246 3818 1280
rect 3818 1246 3852 1280
rect 3852 1246 3861 1280
rect 3809 1237 3861 1246
rect 2209 70 2261 79
rect 2209 36 2218 70
rect 2218 36 2252 70
rect 2252 36 2261 70
rect 2209 27 2261 36
rect 2109 -60 2161 -15
rect 2109 -67 2118 -60
rect 2118 -67 2152 -60
rect 2152 -67 2161 -60
rect 1909 -166 1918 -143
rect 1918 -166 1952 -143
rect 1952 -166 1961 -143
rect 1909 -195 1961 -166
rect 1925 -248 1977 -239
rect 1925 -282 1934 -248
rect 1934 -282 1968 -248
rect 1968 -282 1977 -248
rect 1925 -291 1977 -282
rect 1909 -363 1961 -326
rect 1909 -378 1918 -363
rect 1918 -378 1952 -363
rect 1952 -378 1961 -363
rect 1909 -397 1918 -390
rect 1918 -397 1952 -390
rect 1952 -397 1961 -390
rect 1909 -435 1961 -397
rect 1909 -442 1918 -435
rect 1918 -442 1952 -435
rect 1952 -442 1961 -435
rect 1909 -469 1918 -454
rect 1918 -469 1952 -454
rect 1952 -469 1961 -454
rect 1909 -506 1961 -469
rect 2109 -94 2118 -79
rect 2118 -94 2152 -79
rect 2152 -94 2161 -79
rect 2109 -131 2161 -94
rect 2209 -74 2261 -22
rect 2409 143 2418 151
rect 2418 143 2452 151
rect 2452 143 2461 151
rect 2409 99 2461 143
rect 2609 317 2661 361
rect 2609 309 2618 317
rect 2618 309 2652 317
rect 2652 309 2661 317
rect 2809 423 2818 431
rect 2818 423 2852 431
rect 2852 423 2861 431
rect 2809 379 2861 423
rect 3009 597 3061 641
rect 3009 589 3018 597
rect 3018 589 3052 597
rect 3052 589 3061 597
rect 3209 703 3218 711
rect 3218 703 3252 711
rect 3252 703 3261 711
rect 3209 659 3261 703
rect 3409 877 3461 921
rect 3409 869 3418 877
rect 3418 869 3452 877
rect 3452 869 3461 877
rect 3609 983 3618 991
rect 3618 983 3652 991
rect 3652 983 3661 991
rect 3609 939 3661 983
rect 3809 1157 3861 1201
rect 3809 1149 3818 1157
rect 3818 1149 3852 1157
rect 3852 1149 3861 1157
rect 4009 1353 4018 1361
rect 4018 1353 4052 1361
rect 4052 1353 4061 1361
rect 4009 1309 4061 1353
rect 4209 1527 4261 1571
rect 4209 1519 4218 1527
rect 4218 1519 4252 1527
rect 4252 1519 4261 1527
rect 4409 1633 4418 1641
rect 4418 1633 4452 1641
rect 4452 1633 4461 1641
rect 4409 1589 4461 1633
rect 4609 1807 4661 1851
rect 4609 1799 4618 1807
rect 4618 1799 4652 1807
rect 4652 1799 4661 1807
rect 4809 1913 4818 1921
rect 4818 1913 4852 1921
rect 4852 1913 4861 1921
rect 4809 1869 4861 1913
rect 5009 2087 5061 2131
rect 5009 2079 5018 2087
rect 5018 2079 5052 2087
rect 5052 2079 5061 2087
rect 5209 2193 5218 2201
rect 5218 2193 5252 2201
rect 5252 2193 5261 2201
rect 5209 2149 5261 2193
rect 5409 2367 5461 2411
rect 5409 2359 5418 2367
rect 5418 2359 5452 2367
rect 5452 2359 5461 2367
rect 5609 2563 5618 2571
rect 5618 2563 5652 2571
rect 5652 2563 5661 2571
rect 5609 2519 5661 2563
rect 5809 2737 5861 2781
rect 5809 2729 5818 2737
rect 5818 2729 5852 2737
rect 5852 2729 5861 2737
rect 6009 2843 6018 2851
rect 6018 2843 6052 2851
rect 6052 2843 6061 2851
rect 6009 2799 6061 2843
rect 6209 3017 6261 3061
rect 6209 3009 6218 3017
rect 6218 3009 6252 3017
rect 6252 3009 6261 3017
rect 6409 3123 6418 3131
rect 6418 3123 6452 3131
rect 6452 3123 6461 3131
rect 6409 3079 6461 3123
rect 6507 3079 6559 3131
rect 5609 2474 5661 2483
rect 5609 2440 5618 2474
rect 5618 2440 5652 2474
rect 5652 2440 5661 2474
rect 5609 2431 5661 2440
rect 4009 1264 4061 1273
rect 4009 1230 4018 1264
rect 4018 1230 4052 1264
rect 4052 1230 4061 1264
rect 4009 1221 4061 1230
rect 2409 54 2461 63
rect 2409 20 2418 54
rect 2418 20 2452 54
rect 2452 20 2461 54
rect 2409 11 2461 20
rect 2309 -60 2361 -15
rect 2309 -67 2318 -60
rect 2318 -67 2352 -60
rect 2352 -67 2361 -60
rect 2109 -166 2118 -143
rect 2118 -166 2152 -143
rect 2152 -166 2161 -143
rect 2109 -195 2161 -166
rect 2125 -248 2177 -239
rect 2125 -282 2134 -248
rect 2134 -282 2168 -248
rect 2168 -282 2177 -248
rect 2125 -291 2177 -282
rect 2109 -363 2161 -326
rect 2109 -378 2118 -363
rect 2118 -378 2152 -363
rect 2152 -378 2161 -363
rect 2109 -397 2118 -390
rect 2118 -397 2152 -390
rect 2152 -397 2161 -390
rect 2109 -435 2161 -397
rect 2109 -442 2118 -435
rect 2118 -442 2152 -435
rect 2152 -442 2161 -435
rect 2109 -469 2118 -454
rect 2118 -469 2152 -454
rect 2152 -469 2161 -454
rect 2109 -506 2161 -469
rect 2309 -94 2318 -79
rect 2318 -94 2352 -79
rect 2352 -94 2361 -79
rect 2309 -131 2361 -94
rect 2409 -74 2461 -22
rect 2609 177 2661 221
rect 2609 169 2618 177
rect 2618 169 2652 177
rect 2652 169 2661 177
rect 2809 283 2818 291
rect 2818 283 2852 291
rect 2852 283 2861 291
rect 2809 239 2861 283
rect 3009 457 3061 501
rect 3009 449 3018 457
rect 3018 449 3052 457
rect 3052 449 3061 457
rect 3209 563 3218 571
rect 3218 563 3252 571
rect 3252 563 3261 571
rect 3209 519 3261 563
rect 3409 737 3461 781
rect 3409 729 3418 737
rect 3418 729 3452 737
rect 3452 729 3461 737
rect 3609 843 3618 851
rect 3618 843 3652 851
rect 3652 843 3661 851
rect 3609 799 3661 843
rect 3809 1017 3861 1061
rect 3809 1009 3818 1017
rect 3818 1009 3852 1017
rect 3852 1009 3861 1017
rect 4009 1123 4018 1131
rect 4018 1123 4052 1131
rect 4052 1123 4061 1131
rect 4009 1079 4061 1123
rect 4209 1387 4261 1431
rect 4209 1379 4218 1387
rect 4218 1379 4252 1387
rect 4252 1379 4261 1387
rect 4409 1493 4418 1501
rect 4418 1493 4452 1501
rect 4452 1493 4461 1501
rect 4409 1449 4461 1493
rect 4609 1667 4661 1711
rect 4609 1659 4618 1667
rect 4618 1659 4652 1667
rect 4652 1659 4661 1667
rect 4809 1773 4818 1781
rect 4818 1773 4852 1781
rect 4852 1773 4861 1781
rect 4809 1729 4861 1773
rect 5009 1947 5061 1991
rect 5009 1939 5018 1947
rect 5018 1939 5052 1947
rect 5052 1939 5061 1947
rect 5209 2053 5218 2061
rect 5218 2053 5252 2061
rect 5252 2053 5261 2061
rect 5209 2009 5261 2053
rect 5409 2227 5461 2271
rect 5409 2219 5418 2227
rect 5418 2219 5452 2227
rect 5452 2219 5461 2227
rect 5609 2333 5618 2341
rect 5618 2333 5652 2341
rect 5652 2333 5661 2341
rect 5609 2289 5661 2333
rect 5809 2597 5861 2641
rect 5809 2589 5818 2597
rect 5818 2589 5852 2597
rect 5852 2589 5861 2597
rect 6009 2703 6018 2711
rect 6018 2703 6052 2711
rect 6052 2703 6061 2711
rect 6009 2659 6061 2703
rect 6209 2877 6261 2921
rect 6209 2869 6218 2877
rect 6218 2869 6252 2877
rect 6252 2869 6261 2877
rect 6409 2983 6418 2991
rect 6418 2983 6452 2991
rect 6452 2983 6461 2991
rect 6409 2939 6461 2983
rect 6507 2939 6559 2991
rect 5809 2490 5861 2499
rect 5809 2456 5818 2490
rect 5818 2456 5852 2490
rect 5852 2456 5861 2490
rect 5809 2447 5861 2456
rect 4209 1280 4261 1289
rect 4209 1246 4218 1280
rect 4218 1246 4252 1280
rect 4252 1246 4261 1280
rect 4209 1237 4261 1246
rect 2609 70 2661 79
rect 2609 36 2618 70
rect 2618 36 2652 70
rect 2652 36 2661 70
rect 2609 27 2661 36
rect 2509 -60 2561 -15
rect 2509 -67 2518 -60
rect 2518 -67 2552 -60
rect 2552 -67 2561 -60
rect 2309 -166 2318 -143
rect 2318 -166 2352 -143
rect 2352 -166 2361 -143
rect 2309 -195 2361 -166
rect 2325 -248 2377 -239
rect 2325 -282 2334 -248
rect 2334 -282 2368 -248
rect 2368 -282 2377 -248
rect 2325 -291 2377 -282
rect 2309 -363 2361 -326
rect 2309 -378 2318 -363
rect 2318 -378 2352 -363
rect 2352 -378 2361 -363
rect 2309 -397 2318 -390
rect 2318 -397 2352 -390
rect 2352 -397 2361 -390
rect 2309 -435 2361 -397
rect 2309 -442 2318 -435
rect 2318 -442 2352 -435
rect 2352 -442 2361 -435
rect 2309 -469 2318 -454
rect 2318 -469 2352 -454
rect 2352 -469 2361 -454
rect 2309 -506 2361 -469
rect 2509 -94 2518 -79
rect 2518 -94 2552 -79
rect 2552 -94 2561 -79
rect 2509 -131 2561 -94
rect 2609 -74 2661 -22
rect 2809 143 2818 151
rect 2818 143 2852 151
rect 2852 143 2861 151
rect 2809 99 2861 143
rect 3009 317 3061 361
rect 3009 309 3018 317
rect 3018 309 3052 317
rect 3052 309 3061 317
rect 3209 423 3218 431
rect 3218 423 3252 431
rect 3252 423 3261 431
rect 3209 379 3261 423
rect 3409 597 3461 641
rect 3409 589 3418 597
rect 3418 589 3452 597
rect 3452 589 3461 597
rect 3609 703 3618 711
rect 3618 703 3652 711
rect 3652 703 3661 711
rect 3609 659 3661 703
rect 3809 877 3861 921
rect 3809 869 3818 877
rect 3818 869 3852 877
rect 3852 869 3861 877
rect 4009 983 4018 991
rect 4018 983 4052 991
rect 4052 983 4061 991
rect 4009 939 4061 983
rect 4209 1157 4261 1201
rect 4209 1149 4218 1157
rect 4218 1149 4252 1157
rect 4252 1149 4261 1157
rect 4409 1353 4418 1361
rect 4418 1353 4452 1361
rect 4452 1353 4461 1361
rect 4409 1309 4461 1353
rect 4609 1527 4661 1571
rect 4609 1519 4618 1527
rect 4618 1519 4652 1527
rect 4652 1519 4661 1527
rect 4809 1633 4818 1641
rect 4818 1633 4852 1641
rect 4852 1633 4861 1641
rect 4809 1589 4861 1633
rect 5009 1807 5061 1851
rect 5009 1799 5018 1807
rect 5018 1799 5052 1807
rect 5052 1799 5061 1807
rect 5209 1913 5218 1921
rect 5218 1913 5252 1921
rect 5252 1913 5261 1921
rect 5209 1869 5261 1913
rect 5409 2087 5461 2131
rect 5409 2079 5418 2087
rect 5418 2079 5452 2087
rect 5452 2079 5461 2087
rect 5609 2193 5618 2201
rect 5618 2193 5652 2201
rect 5652 2193 5661 2201
rect 5609 2149 5661 2193
rect 5809 2367 5861 2411
rect 5809 2359 5818 2367
rect 5818 2359 5852 2367
rect 5852 2359 5861 2367
rect 6009 2563 6018 2571
rect 6018 2563 6052 2571
rect 6052 2563 6061 2571
rect 6009 2519 6061 2563
rect 6209 2737 6261 2781
rect 6209 2729 6218 2737
rect 6218 2729 6252 2737
rect 6252 2729 6261 2737
rect 6409 2843 6418 2851
rect 6418 2843 6452 2851
rect 6452 2843 6461 2851
rect 6409 2799 6461 2843
rect 6507 2799 6559 2851
rect 6009 2474 6061 2483
rect 6009 2440 6018 2474
rect 6018 2440 6052 2474
rect 6052 2440 6061 2474
rect 6009 2431 6061 2440
rect 4409 1264 4461 1273
rect 4409 1230 4418 1264
rect 4418 1230 4452 1264
rect 4452 1230 4461 1264
rect 4409 1221 4461 1230
rect 2809 54 2861 63
rect 2809 20 2818 54
rect 2818 20 2852 54
rect 2852 20 2861 54
rect 2809 11 2861 20
rect 2709 -60 2761 -15
rect 2709 -67 2718 -60
rect 2718 -67 2752 -60
rect 2752 -67 2761 -60
rect 2509 -166 2518 -143
rect 2518 -166 2552 -143
rect 2552 -166 2561 -143
rect 2509 -195 2561 -166
rect 2525 -248 2577 -239
rect 2525 -282 2534 -248
rect 2534 -282 2568 -248
rect 2568 -282 2577 -248
rect 2525 -291 2577 -282
rect 2509 -363 2561 -326
rect 2509 -378 2518 -363
rect 2518 -378 2552 -363
rect 2552 -378 2561 -363
rect 2509 -397 2518 -390
rect 2518 -397 2552 -390
rect 2552 -397 2561 -390
rect 2509 -435 2561 -397
rect 2509 -442 2518 -435
rect 2518 -442 2552 -435
rect 2552 -442 2561 -435
rect 2509 -469 2518 -454
rect 2518 -469 2552 -454
rect 2552 -469 2561 -454
rect 2509 -506 2561 -469
rect 2709 -94 2718 -79
rect 2718 -94 2752 -79
rect 2752 -94 2761 -79
rect 2709 -131 2761 -94
rect 2809 -74 2861 -22
rect 3009 177 3061 221
rect 3009 169 3018 177
rect 3018 169 3052 177
rect 3052 169 3061 177
rect 3209 283 3218 291
rect 3218 283 3252 291
rect 3252 283 3261 291
rect 3209 239 3261 283
rect 3409 457 3461 501
rect 3409 449 3418 457
rect 3418 449 3452 457
rect 3452 449 3461 457
rect 3609 563 3618 571
rect 3618 563 3652 571
rect 3652 563 3661 571
rect 3609 519 3661 563
rect 3809 737 3861 781
rect 3809 729 3818 737
rect 3818 729 3852 737
rect 3852 729 3861 737
rect 4009 843 4018 851
rect 4018 843 4052 851
rect 4052 843 4061 851
rect 4009 799 4061 843
rect 4209 1017 4261 1061
rect 4209 1009 4218 1017
rect 4218 1009 4252 1017
rect 4252 1009 4261 1017
rect 4409 1123 4418 1131
rect 4418 1123 4452 1131
rect 4452 1123 4461 1131
rect 4409 1079 4461 1123
rect 4609 1387 4661 1431
rect 4609 1379 4618 1387
rect 4618 1379 4652 1387
rect 4652 1379 4661 1387
rect 4809 1493 4818 1501
rect 4818 1493 4852 1501
rect 4852 1493 4861 1501
rect 4809 1449 4861 1493
rect 5009 1667 5061 1711
rect 5009 1659 5018 1667
rect 5018 1659 5052 1667
rect 5052 1659 5061 1667
rect 5209 1773 5218 1781
rect 5218 1773 5252 1781
rect 5252 1773 5261 1781
rect 5209 1729 5261 1773
rect 5409 1947 5461 1991
rect 5409 1939 5418 1947
rect 5418 1939 5452 1947
rect 5452 1939 5461 1947
rect 5609 2053 5618 2061
rect 5618 2053 5652 2061
rect 5652 2053 5661 2061
rect 5609 2009 5661 2053
rect 5809 2227 5861 2271
rect 5809 2219 5818 2227
rect 5818 2219 5852 2227
rect 5852 2219 5861 2227
rect 6009 2333 6018 2341
rect 6018 2333 6052 2341
rect 6052 2333 6061 2341
rect 6009 2289 6061 2333
rect 6209 2597 6261 2641
rect 6209 2589 6218 2597
rect 6218 2589 6252 2597
rect 6252 2589 6261 2597
rect 6409 2703 6418 2711
rect 6418 2703 6452 2711
rect 6452 2703 6461 2711
rect 6409 2659 6461 2703
rect 6507 2659 6559 2711
rect 6209 2490 6261 2499
rect 6209 2456 6218 2490
rect 6218 2456 6252 2490
rect 6252 2456 6261 2490
rect 6209 2447 6261 2456
rect 4609 1280 4661 1289
rect 4609 1246 4618 1280
rect 4618 1246 4652 1280
rect 4652 1246 4661 1280
rect 4609 1237 4661 1246
rect 3009 70 3061 79
rect 3009 36 3018 70
rect 3018 36 3052 70
rect 3052 36 3061 70
rect 3009 27 3061 36
rect 2909 -60 2961 -15
rect 2909 -67 2918 -60
rect 2918 -67 2952 -60
rect 2952 -67 2961 -60
rect 2709 -166 2718 -143
rect 2718 -166 2752 -143
rect 2752 -166 2761 -143
rect 2709 -195 2761 -166
rect 2725 -248 2777 -239
rect 2725 -282 2734 -248
rect 2734 -282 2768 -248
rect 2768 -282 2777 -248
rect 2725 -291 2777 -282
rect 2709 -363 2761 -326
rect 2709 -378 2718 -363
rect 2718 -378 2752 -363
rect 2752 -378 2761 -363
rect 2709 -397 2718 -390
rect 2718 -397 2752 -390
rect 2752 -397 2761 -390
rect 2709 -435 2761 -397
rect 2709 -442 2718 -435
rect 2718 -442 2752 -435
rect 2752 -442 2761 -435
rect 2709 -469 2718 -454
rect 2718 -469 2752 -454
rect 2752 -469 2761 -454
rect 2709 -506 2761 -469
rect 2909 -94 2918 -79
rect 2918 -94 2952 -79
rect 2952 -94 2961 -79
rect 2909 -131 2961 -94
rect 3009 -74 3061 -22
rect 3209 143 3218 151
rect 3218 143 3252 151
rect 3252 143 3261 151
rect 3209 99 3261 143
rect 3409 317 3461 361
rect 3409 309 3418 317
rect 3418 309 3452 317
rect 3452 309 3461 317
rect 3609 423 3618 431
rect 3618 423 3652 431
rect 3652 423 3661 431
rect 3609 379 3661 423
rect 3809 597 3861 641
rect 3809 589 3818 597
rect 3818 589 3852 597
rect 3852 589 3861 597
rect 4009 703 4018 711
rect 4018 703 4052 711
rect 4052 703 4061 711
rect 4009 659 4061 703
rect 4209 877 4261 921
rect 4209 869 4218 877
rect 4218 869 4252 877
rect 4252 869 4261 877
rect 4409 983 4418 991
rect 4418 983 4452 991
rect 4452 983 4461 991
rect 4409 939 4461 983
rect 4609 1157 4661 1201
rect 4609 1149 4618 1157
rect 4618 1149 4652 1157
rect 4652 1149 4661 1157
rect 4809 1353 4818 1361
rect 4818 1353 4852 1361
rect 4852 1353 4861 1361
rect 4809 1309 4861 1353
rect 5009 1527 5061 1571
rect 5009 1519 5018 1527
rect 5018 1519 5052 1527
rect 5052 1519 5061 1527
rect 5209 1633 5218 1641
rect 5218 1633 5252 1641
rect 5252 1633 5261 1641
rect 5209 1589 5261 1633
rect 5409 1807 5461 1851
rect 5409 1799 5418 1807
rect 5418 1799 5452 1807
rect 5452 1799 5461 1807
rect 5609 1913 5618 1921
rect 5618 1913 5652 1921
rect 5652 1913 5661 1921
rect 5609 1869 5661 1913
rect 5809 2087 5861 2131
rect 5809 2079 5818 2087
rect 5818 2079 5852 2087
rect 5852 2079 5861 2087
rect 6009 2193 6018 2201
rect 6018 2193 6052 2201
rect 6052 2193 6061 2201
rect 6009 2149 6061 2193
rect 6209 2367 6261 2411
rect 6209 2359 6218 2367
rect 6218 2359 6252 2367
rect 6252 2359 6261 2367
rect 6409 2563 6418 2571
rect 6418 2563 6452 2571
rect 6452 2563 6461 2571
rect 6409 2519 6461 2563
rect 6507 2519 6559 2571
rect 4809 1264 4861 1273
rect 4809 1230 4818 1264
rect 4818 1230 4852 1264
rect 4852 1230 4861 1264
rect 4809 1221 4861 1230
rect 3209 54 3261 63
rect 3209 20 3218 54
rect 3218 20 3252 54
rect 3252 20 3261 54
rect 3209 11 3261 20
rect 3109 -60 3161 -15
rect 3109 -67 3118 -60
rect 3118 -67 3152 -60
rect 3152 -67 3161 -60
rect 2909 -166 2918 -143
rect 2918 -166 2952 -143
rect 2952 -166 2961 -143
rect 2909 -195 2961 -166
rect 2925 -248 2977 -239
rect 2925 -282 2934 -248
rect 2934 -282 2968 -248
rect 2968 -282 2977 -248
rect 2925 -291 2977 -282
rect 2909 -363 2961 -326
rect 2909 -378 2918 -363
rect 2918 -378 2952 -363
rect 2952 -378 2961 -363
rect 2909 -397 2918 -390
rect 2918 -397 2952 -390
rect 2952 -397 2961 -390
rect 2909 -435 2961 -397
rect 2909 -442 2918 -435
rect 2918 -442 2952 -435
rect 2952 -442 2961 -435
rect 2909 -469 2918 -454
rect 2918 -469 2952 -454
rect 2952 -469 2961 -454
rect 2909 -506 2961 -469
rect 3109 -94 3118 -79
rect 3118 -94 3152 -79
rect 3152 -94 3161 -79
rect 3109 -131 3161 -94
rect 3209 -74 3261 -22
rect 3409 177 3461 221
rect 3409 169 3418 177
rect 3418 169 3452 177
rect 3452 169 3461 177
rect 3609 283 3618 291
rect 3618 283 3652 291
rect 3652 283 3661 291
rect 3609 239 3661 283
rect 3809 457 3861 501
rect 3809 449 3818 457
rect 3818 449 3852 457
rect 3852 449 3861 457
rect 4009 563 4018 571
rect 4018 563 4052 571
rect 4052 563 4061 571
rect 4009 519 4061 563
rect 4209 737 4261 781
rect 4209 729 4218 737
rect 4218 729 4252 737
rect 4252 729 4261 737
rect 4409 843 4418 851
rect 4418 843 4452 851
rect 4452 843 4461 851
rect 4409 799 4461 843
rect 4609 1017 4661 1061
rect 4609 1009 4618 1017
rect 4618 1009 4652 1017
rect 4652 1009 4661 1017
rect 4809 1123 4818 1131
rect 4818 1123 4852 1131
rect 4852 1123 4861 1131
rect 4809 1079 4861 1123
rect 5009 1387 5061 1431
rect 5009 1379 5018 1387
rect 5018 1379 5052 1387
rect 5052 1379 5061 1387
rect 5209 1493 5218 1501
rect 5218 1493 5252 1501
rect 5252 1493 5261 1501
rect 5209 1449 5261 1493
rect 5409 1667 5461 1711
rect 5409 1659 5418 1667
rect 5418 1659 5452 1667
rect 5452 1659 5461 1667
rect 5609 1773 5618 1781
rect 5618 1773 5652 1781
rect 5652 1773 5661 1781
rect 5609 1729 5661 1773
rect 5809 1947 5861 1991
rect 5809 1939 5818 1947
rect 5818 1939 5852 1947
rect 5852 1939 5861 1947
rect 6009 2053 6018 2061
rect 6018 2053 6052 2061
rect 6052 2053 6061 2061
rect 6009 2009 6061 2053
rect 6209 2227 6261 2271
rect 6209 2219 6218 2227
rect 6218 2219 6252 2227
rect 6252 2219 6261 2227
rect 6409 2333 6418 2341
rect 6418 2333 6452 2341
rect 6452 2333 6461 2341
rect 6409 2289 6461 2333
rect 6507 2289 6559 2341
rect 5009 1280 5061 1289
rect 5009 1246 5018 1280
rect 5018 1246 5052 1280
rect 5052 1246 5061 1280
rect 5009 1237 5061 1246
rect 3409 70 3461 79
rect 3409 36 3418 70
rect 3418 36 3452 70
rect 3452 36 3461 70
rect 3409 27 3461 36
rect 3309 -60 3361 -15
rect 3309 -67 3318 -60
rect 3318 -67 3352 -60
rect 3352 -67 3361 -60
rect 3109 -166 3118 -143
rect 3118 -166 3152 -143
rect 3152 -166 3161 -143
rect 3109 -195 3161 -166
rect 3125 -248 3177 -239
rect 3125 -282 3134 -248
rect 3134 -282 3168 -248
rect 3168 -282 3177 -248
rect 3125 -291 3177 -282
rect 3109 -363 3161 -326
rect 3109 -378 3118 -363
rect 3118 -378 3152 -363
rect 3152 -378 3161 -363
rect 3109 -397 3118 -390
rect 3118 -397 3152 -390
rect 3152 -397 3161 -390
rect 3109 -435 3161 -397
rect 3109 -442 3118 -435
rect 3118 -442 3152 -435
rect 3152 -442 3161 -435
rect 3109 -469 3118 -454
rect 3118 -469 3152 -454
rect 3152 -469 3161 -454
rect 3109 -506 3161 -469
rect 3309 -94 3318 -79
rect 3318 -94 3352 -79
rect 3352 -94 3361 -79
rect 3309 -131 3361 -94
rect 3409 -74 3461 -22
rect 3609 143 3618 151
rect 3618 143 3652 151
rect 3652 143 3661 151
rect 3609 99 3661 143
rect 3809 317 3861 361
rect 3809 309 3818 317
rect 3818 309 3852 317
rect 3852 309 3861 317
rect 4009 423 4018 431
rect 4018 423 4052 431
rect 4052 423 4061 431
rect 4009 379 4061 423
rect 4209 597 4261 641
rect 4209 589 4218 597
rect 4218 589 4252 597
rect 4252 589 4261 597
rect 4409 703 4418 711
rect 4418 703 4452 711
rect 4452 703 4461 711
rect 4409 659 4461 703
rect 4609 877 4661 921
rect 4609 869 4618 877
rect 4618 869 4652 877
rect 4652 869 4661 877
rect 4809 983 4818 991
rect 4818 983 4852 991
rect 4852 983 4861 991
rect 4809 939 4861 983
rect 5009 1157 5061 1201
rect 5009 1149 5018 1157
rect 5018 1149 5052 1157
rect 5052 1149 5061 1157
rect 5209 1353 5218 1361
rect 5218 1353 5252 1361
rect 5252 1353 5261 1361
rect 5209 1309 5261 1353
rect 5409 1527 5461 1571
rect 5409 1519 5418 1527
rect 5418 1519 5452 1527
rect 5452 1519 5461 1527
rect 5609 1633 5618 1641
rect 5618 1633 5652 1641
rect 5652 1633 5661 1641
rect 5609 1589 5661 1633
rect 5809 1807 5861 1851
rect 5809 1799 5818 1807
rect 5818 1799 5852 1807
rect 5852 1799 5861 1807
rect 6009 1913 6018 1921
rect 6018 1913 6052 1921
rect 6052 1913 6061 1921
rect 6009 1869 6061 1913
rect 6209 2087 6261 2131
rect 6209 2079 6218 2087
rect 6218 2079 6252 2087
rect 6252 2079 6261 2087
rect 6409 2193 6418 2201
rect 6418 2193 6452 2201
rect 6452 2193 6461 2201
rect 6409 2149 6461 2193
rect 6507 2149 6559 2201
rect 5209 1264 5261 1273
rect 5209 1230 5218 1264
rect 5218 1230 5252 1264
rect 5252 1230 5261 1264
rect 5209 1221 5261 1230
rect 3609 54 3661 63
rect 3609 20 3618 54
rect 3618 20 3652 54
rect 3652 20 3661 54
rect 3609 11 3661 20
rect 3509 -60 3561 -15
rect 3509 -67 3518 -60
rect 3518 -67 3552 -60
rect 3552 -67 3561 -60
rect 3309 -166 3318 -143
rect 3318 -166 3352 -143
rect 3352 -166 3361 -143
rect 3309 -195 3361 -166
rect 3325 -248 3377 -239
rect 3325 -282 3334 -248
rect 3334 -282 3368 -248
rect 3368 -282 3377 -248
rect 3325 -291 3377 -282
rect 3309 -363 3361 -326
rect 3309 -378 3318 -363
rect 3318 -378 3352 -363
rect 3352 -378 3361 -363
rect 3309 -397 3318 -390
rect 3318 -397 3352 -390
rect 3352 -397 3361 -390
rect 3309 -435 3361 -397
rect 3309 -442 3318 -435
rect 3318 -442 3352 -435
rect 3352 -442 3361 -435
rect 3309 -469 3318 -454
rect 3318 -469 3352 -454
rect 3352 -469 3361 -454
rect 3309 -506 3361 -469
rect 3509 -94 3518 -79
rect 3518 -94 3552 -79
rect 3552 -94 3561 -79
rect 3509 -131 3561 -94
rect 3609 -74 3661 -22
rect 3809 177 3861 221
rect 3809 169 3818 177
rect 3818 169 3852 177
rect 3852 169 3861 177
rect 4009 283 4018 291
rect 4018 283 4052 291
rect 4052 283 4061 291
rect 4009 239 4061 283
rect 4209 457 4261 501
rect 4209 449 4218 457
rect 4218 449 4252 457
rect 4252 449 4261 457
rect 4409 563 4418 571
rect 4418 563 4452 571
rect 4452 563 4461 571
rect 4409 519 4461 563
rect 4609 737 4661 781
rect 4609 729 4618 737
rect 4618 729 4652 737
rect 4652 729 4661 737
rect 4809 843 4818 851
rect 4818 843 4852 851
rect 4852 843 4861 851
rect 4809 799 4861 843
rect 5009 1017 5061 1061
rect 5009 1009 5018 1017
rect 5018 1009 5052 1017
rect 5052 1009 5061 1017
rect 5209 1123 5218 1131
rect 5218 1123 5252 1131
rect 5252 1123 5261 1131
rect 5209 1079 5261 1123
rect 5409 1387 5461 1431
rect 5409 1379 5418 1387
rect 5418 1379 5452 1387
rect 5452 1379 5461 1387
rect 5609 1493 5618 1501
rect 5618 1493 5652 1501
rect 5652 1493 5661 1501
rect 5609 1449 5661 1493
rect 5809 1667 5861 1711
rect 5809 1659 5818 1667
rect 5818 1659 5852 1667
rect 5852 1659 5861 1667
rect 6009 1773 6018 1781
rect 6018 1773 6052 1781
rect 6052 1773 6061 1781
rect 6009 1729 6061 1773
rect 6209 1947 6261 1991
rect 6209 1939 6218 1947
rect 6218 1939 6252 1947
rect 6252 1939 6261 1947
rect 6409 2053 6418 2061
rect 6418 2053 6452 2061
rect 6452 2053 6461 2061
rect 6409 2009 6461 2053
rect 6507 2009 6559 2061
rect 5409 1280 5461 1289
rect 5409 1246 5418 1280
rect 5418 1246 5452 1280
rect 5452 1246 5461 1280
rect 5409 1237 5461 1246
rect 3809 70 3861 79
rect 3809 36 3818 70
rect 3818 36 3852 70
rect 3852 36 3861 70
rect 3809 27 3861 36
rect 3709 -60 3761 -15
rect 3709 -67 3718 -60
rect 3718 -67 3752 -60
rect 3752 -67 3761 -60
rect 3509 -166 3518 -143
rect 3518 -166 3552 -143
rect 3552 -166 3561 -143
rect 3509 -195 3561 -166
rect 3525 -248 3577 -239
rect 3525 -282 3534 -248
rect 3534 -282 3568 -248
rect 3568 -282 3577 -248
rect 3525 -291 3577 -282
rect 3509 -363 3561 -326
rect 3509 -378 3518 -363
rect 3518 -378 3552 -363
rect 3552 -378 3561 -363
rect 3509 -397 3518 -390
rect 3518 -397 3552 -390
rect 3552 -397 3561 -390
rect 3509 -435 3561 -397
rect 3509 -442 3518 -435
rect 3518 -442 3552 -435
rect 3552 -442 3561 -435
rect 3509 -469 3518 -454
rect 3518 -469 3552 -454
rect 3552 -469 3561 -454
rect 3509 -506 3561 -469
rect 3709 -94 3718 -79
rect 3718 -94 3752 -79
rect 3752 -94 3761 -79
rect 3709 -131 3761 -94
rect 3809 -74 3861 -22
rect 4009 143 4018 151
rect 4018 143 4052 151
rect 4052 143 4061 151
rect 4009 99 4061 143
rect 4209 317 4261 361
rect 4209 309 4218 317
rect 4218 309 4252 317
rect 4252 309 4261 317
rect 4409 423 4418 431
rect 4418 423 4452 431
rect 4452 423 4461 431
rect 4409 379 4461 423
rect 4609 597 4661 641
rect 4609 589 4618 597
rect 4618 589 4652 597
rect 4652 589 4661 597
rect 4809 703 4818 711
rect 4818 703 4852 711
rect 4852 703 4861 711
rect 4809 659 4861 703
rect 5009 877 5061 921
rect 5009 869 5018 877
rect 5018 869 5052 877
rect 5052 869 5061 877
rect 5209 983 5218 991
rect 5218 983 5252 991
rect 5252 983 5261 991
rect 5209 939 5261 983
rect 5409 1157 5461 1201
rect 5409 1149 5418 1157
rect 5418 1149 5452 1157
rect 5452 1149 5461 1157
rect 5609 1353 5618 1361
rect 5618 1353 5652 1361
rect 5652 1353 5661 1361
rect 5609 1309 5661 1353
rect 5809 1527 5861 1571
rect 5809 1519 5818 1527
rect 5818 1519 5852 1527
rect 5852 1519 5861 1527
rect 6009 1633 6018 1641
rect 6018 1633 6052 1641
rect 6052 1633 6061 1641
rect 6009 1589 6061 1633
rect 6209 1807 6261 1851
rect 6209 1799 6218 1807
rect 6218 1799 6252 1807
rect 6252 1799 6261 1807
rect 6409 1913 6418 1921
rect 6418 1913 6452 1921
rect 6452 1913 6461 1921
rect 6409 1869 6461 1913
rect 6507 1869 6559 1921
rect 5609 1264 5661 1273
rect 5609 1230 5618 1264
rect 5618 1230 5652 1264
rect 5652 1230 5661 1264
rect 5609 1221 5661 1230
rect 4009 54 4061 63
rect 4009 20 4018 54
rect 4018 20 4052 54
rect 4052 20 4061 54
rect 4009 11 4061 20
rect 3909 -60 3961 -15
rect 3909 -67 3918 -60
rect 3918 -67 3952 -60
rect 3952 -67 3961 -60
rect 3709 -166 3718 -143
rect 3718 -166 3752 -143
rect 3752 -166 3761 -143
rect 3709 -195 3761 -166
rect 3725 -248 3777 -239
rect 3725 -282 3734 -248
rect 3734 -282 3768 -248
rect 3768 -282 3777 -248
rect 3725 -291 3777 -282
rect 3709 -363 3761 -326
rect 3709 -378 3718 -363
rect 3718 -378 3752 -363
rect 3752 -378 3761 -363
rect 3709 -397 3718 -390
rect 3718 -397 3752 -390
rect 3752 -397 3761 -390
rect 3709 -435 3761 -397
rect 3709 -442 3718 -435
rect 3718 -442 3752 -435
rect 3752 -442 3761 -435
rect 3709 -469 3718 -454
rect 3718 -469 3752 -454
rect 3752 -469 3761 -454
rect 3709 -506 3761 -469
rect 3909 -94 3918 -79
rect 3918 -94 3952 -79
rect 3952 -94 3961 -79
rect 3909 -131 3961 -94
rect 4009 -74 4061 -22
rect 4209 177 4261 221
rect 4209 169 4218 177
rect 4218 169 4252 177
rect 4252 169 4261 177
rect 4409 283 4418 291
rect 4418 283 4452 291
rect 4452 283 4461 291
rect 4409 239 4461 283
rect 4609 457 4661 501
rect 4609 449 4618 457
rect 4618 449 4652 457
rect 4652 449 4661 457
rect 4809 563 4818 571
rect 4818 563 4852 571
rect 4852 563 4861 571
rect 4809 519 4861 563
rect 5009 737 5061 781
rect 5009 729 5018 737
rect 5018 729 5052 737
rect 5052 729 5061 737
rect 5209 843 5218 851
rect 5218 843 5252 851
rect 5252 843 5261 851
rect 5209 799 5261 843
rect 5409 1017 5461 1061
rect 5409 1009 5418 1017
rect 5418 1009 5452 1017
rect 5452 1009 5461 1017
rect 5609 1123 5618 1131
rect 5618 1123 5652 1131
rect 5652 1123 5661 1131
rect 5609 1079 5661 1123
rect 5809 1387 5861 1431
rect 5809 1379 5818 1387
rect 5818 1379 5852 1387
rect 5852 1379 5861 1387
rect 6009 1493 6018 1501
rect 6018 1493 6052 1501
rect 6052 1493 6061 1501
rect 6009 1449 6061 1493
rect 6209 1667 6261 1711
rect 6209 1659 6218 1667
rect 6218 1659 6252 1667
rect 6252 1659 6261 1667
rect 6409 1773 6418 1781
rect 6418 1773 6452 1781
rect 6452 1773 6461 1781
rect 6409 1729 6461 1773
rect 6507 1729 6559 1781
rect 5809 1280 5861 1289
rect 5809 1246 5818 1280
rect 5818 1246 5852 1280
rect 5852 1246 5861 1280
rect 5809 1237 5861 1246
rect 4209 70 4261 79
rect 4209 36 4218 70
rect 4218 36 4252 70
rect 4252 36 4261 70
rect 4209 27 4261 36
rect 4109 -60 4161 -15
rect 4109 -67 4118 -60
rect 4118 -67 4152 -60
rect 4152 -67 4161 -60
rect 3909 -166 3918 -143
rect 3918 -166 3952 -143
rect 3952 -166 3961 -143
rect 3909 -195 3961 -166
rect 3925 -248 3977 -239
rect 3925 -282 3934 -248
rect 3934 -282 3968 -248
rect 3968 -282 3977 -248
rect 3925 -291 3977 -282
rect 3909 -363 3961 -326
rect 3909 -378 3918 -363
rect 3918 -378 3952 -363
rect 3952 -378 3961 -363
rect 3909 -397 3918 -390
rect 3918 -397 3952 -390
rect 3952 -397 3961 -390
rect 3909 -435 3961 -397
rect 3909 -442 3918 -435
rect 3918 -442 3952 -435
rect 3952 -442 3961 -435
rect 3909 -469 3918 -454
rect 3918 -469 3952 -454
rect 3952 -469 3961 -454
rect 3909 -506 3961 -469
rect 4109 -94 4118 -79
rect 4118 -94 4152 -79
rect 4152 -94 4161 -79
rect 4109 -131 4161 -94
rect 4209 -74 4261 -22
rect 4409 143 4418 151
rect 4418 143 4452 151
rect 4452 143 4461 151
rect 4409 99 4461 143
rect 4609 317 4661 361
rect 4609 309 4618 317
rect 4618 309 4652 317
rect 4652 309 4661 317
rect 4809 423 4818 431
rect 4818 423 4852 431
rect 4852 423 4861 431
rect 4809 379 4861 423
rect 5009 597 5061 641
rect 5009 589 5018 597
rect 5018 589 5052 597
rect 5052 589 5061 597
rect 5209 703 5218 711
rect 5218 703 5252 711
rect 5252 703 5261 711
rect 5209 659 5261 703
rect 5409 877 5461 921
rect 5409 869 5418 877
rect 5418 869 5452 877
rect 5452 869 5461 877
rect 5609 983 5618 991
rect 5618 983 5652 991
rect 5652 983 5661 991
rect 5609 939 5661 983
rect 5809 1157 5861 1201
rect 5809 1149 5818 1157
rect 5818 1149 5852 1157
rect 5852 1149 5861 1157
rect 6009 1353 6018 1361
rect 6018 1353 6052 1361
rect 6052 1353 6061 1361
rect 6009 1309 6061 1353
rect 6209 1527 6261 1571
rect 6209 1519 6218 1527
rect 6218 1519 6252 1527
rect 6252 1519 6261 1527
rect 6409 1633 6418 1641
rect 6418 1633 6452 1641
rect 6452 1633 6461 1641
rect 6409 1589 6461 1633
rect 6507 1589 6559 1641
rect 6009 1264 6061 1273
rect 6009 1230 6018 1264
rect 6018 1230 6052 1264
rect 6052 1230 6061 1264
rect 6009 1221 6061 1230
rect 4409 54 4461 63
rect 4409 20 4418 54
rect 4418 20 4452 54
rect 4452 20 4461 54
rect 4409 11 4461 20
rect 4309 -60 4361 -15
rect 4309 -67 4318 -60
rect 4318 -67 4352 -60
rect 4352 -67 4361 -60
rect 4109 -166 4118 -143
rect 4118 -166 4152 -143
rect 4152 -166 4161 -143
rect 4109 -195 4161 -166
rect 4125 -248 4177 -239
rect 4125 -282 4134 -248
rect 4134 -282 4168 -248
rect 4168 -282 4177 -248
rect 4125 -291 4177 -282
rect 4109 -363 4161 -326
rect 4109 -378 4118 -363
rect 4118 -378 4152 -363
rect 4152 -378 4161 -363
rect 4109 -397 4118 -390
rect 4118 -397 4152 -390
rect 4152 -397 4161 -390
rect 4109 -435 4161 -397
rect 4109 -442 4118 -435
rect 4118 -442 4152 -435
rect 4152 -442 4161 -435
rect 4109 -469 4118 -454
rect 4118 -469 4152 -454
rect 4152 -469 4161 -454
rect 4109 -506 4161 -469
rect 4309 -94 4318 -79
rect 4318 -94 4352 -79
rect 4352 -94 4361 -79
rect 4309 -131 4361 -94
rect 4409 -74 4461 -22
rect 4609 177 4661 221
rect 4609 169 4618 177
rect 4618 169 4652 177
rect 4652 169 4661 177
rect 4809 283 4818 291
rect 4818 283 4852 291
rect 4852 283 4861 291
rect 4809 239 4861 283
rect 5009 457 5061 501
rect 5009 449 5018 457
rect 5018 449 5052 457
rect 5052 449 5061 457
rect 5209 563 5218 571
rect 5218 563 5252 571
rect 5252 563 5261 571
rect 5209 519 5261 563
rect 5409 737 5461 781
rect 5409 729 5418 737
rect 5418 729 5452 737
rect 5452 729 5461 737
rect 5609 843 5618 851
rect 5618 843 5652 851
rect 5652 843 5661 851
rect 5609 799 5661 843
rect 5809 1017 5861 1061
rect 5809 1009 5818 1017
rect 5818 1009 5852 1017
rect 5852 1009 5861 1017
rect 6009 1123 6018 1131
rect 6018 1123 6052 1131
rect 6052 1123 6061 1131
rect 6009 1079 6061 1123
rect 6209 1387 6261 1431
rect 6209 1379 6218 1387
rect 6218 1379 6252 1387
rect 6252 1379 6261 1387
rect 6409 1493 6418 1501
rect 6418 1493 6452 1501
rect 6452 1493 6461 1501
rect 6409 1449 6461 1493
rect 6507 1449 6559 1501
rect 6209 1280 6261 1289
rect 6209 1246 6218 1280
rect 6218 1246 6252 1280
rect 6252 1246 6261 1280
rect 6209 1237 6261 1246
rect 4609 70 4661 79
rect 4609 36 4618 70
rect 4618 36 4652 70
rect 4652 36 4661 70
rect 4609 27 4661 36
rect 4509 -60 4561 -15
rect 4509 -67 4518 -60
rect 4518 -67 4552 -60
rect 4552 -67 4561 -60
rect 4309 -166 4318 -143
rect 4318 -166 4352 -143
rect 4352 -166 4361 -143
rect 4309 -195 4361 -166
rect 4325 -248 4377 -239
rect 4325 -282 4334 -248
rect 4334 -282 4368 -248
rect 4368 -282 4377 -248
rect 4325 -291 4377 -282
rect 4309 -363 4361 -326
rect 4309 -378 4318 -363
rect 4318 -378 4352 -363
rect 4352 -378 4361 -363
rect 4309 -397 4318 -390
rect 4318 -397 4352 -390
rect 4352 -397 4361 -390
rect 4309 -435 4361 -397
rect 4309 -442 4318 -435
rect 4318 -442 4352 -435
rect 4352 -442 4361 -435
rect 4309 -469 4318 -454
rect 4318 -469 4352 -454
rect 4352 -469 4361 -454
rect 4309 -506 4361 -469
rect 4509 -94 4518 -79
rect 4518 -94 4552 -79
rect 4552 -94 4561 -79
rect 4509 -131 4561 -94
rect 4609 -74 4661 -22
rect 4809 143 4818 151
rect 4818 143 4852 151
rect 4852 143 4861 151
rect 4809 99 4861 143
rect 5009 317 5061 361
rect 5009 309 5018 317
rect 5018 309 5052 317
rect 5052 309 5061 317
rect 5209 423 5218 431
rect 5218 423 5252 431
rect 5252 423 5261 431
rect 5209 379 5261 423
rect 5409 597 5461 641
rect 5409 589 5418 597
rect 5418 589 5452 597
rect 5452 589 5461 597
rect 5609 703 5618 711
rect 5618 703 5652 711
rect 5652 703 5661 711
rect 5609 659 5661 703
rect 5809 877 5861 921
rect 5809 869 5818 877
rect 5818 869 5852 877
rect 5852 869 5861 877
rect 6009 983 6018 991
rect 6018 983 6052 991
rect 6052 983 6061 991
rect 6009 939 6061 983
rect 6209 1157 6261 1201
rect 6209 1149 6218 1157
rect 6218 1149 6252 1157
rect 6252 1149 6261 1157
rect 6409 1353 6418 1361
rect 6418 1353 6452 1361
rect 6452 1353 6461 1361
rect 6409 1309 6461 1353
rect 6507 1309 6559 1361
rect 4809 54 4861 63
rect 4809 20 4818 54
rect 4818 20 4852 54
rect 4852 20 4861 54
rect 4809 11 4861 20
rect 4709 -60 4761 -15
rect 4709 -67 4718 -60
rect 4718 -67 4752 -60
rect 4752 -67 4761 -60
rect 4509 -166 4518 -143
rect 4518 -166 4552 -143
rect 4552 -166 4561 -143
rect 4509 -195 4561 -166
rect 4525 -248 4577 -239
rect 4525 -282 4534 -248
rect 4534 -282 4568 -248
rect 4568 -282 4577 -248
rect 4525 -291 4577 -282
rect 4509 -363 4561 -326
rect 4509 -378 4518 -363
rect 4518 -378 4552 -363
rect 4552 -378 4561 -363
rect 4509 -397 4518 -390
rect 4518 -397 4552 -390
rect 4552 -397 4561 -390
rect 4509 -435 4561 -397
rect 4509 -442 4518 -435
rect 4518 -442 4552 -435
rect 4552 -442 4561 -435
rect 4509 -469 4518 -454
rect 4518 -469 4552 -454
rect 4552 -469 4561 -454
rect 4509 -506 4561 -469
rect 4709 -94 4718 -79
rect 4718 -94 4752 -79
rect 4752 -94 4761 -79
rect 4709 -131 4761 -94
rect 4809 -74 4861 -22
rect 5009 177 5061 221
rect 5009 169 5018 177
rect 5018 169 5052 177
rect 5052 169 5061 177
rect 5209 283 5218 291
rect 5218 283 5252 291
rect 5252 283 5261 291
rect 5209 239 5261 283
rect 5409 457 5461 501
rect 5409 449 5418 457
rect 5418 449 5452 457
rect 5452 449 5461 457
rect 5609 563 5618 571
rect 5618 563 5652 571
rect 5652 563 5661 571
rect 5609 519 5661 563
rect 5809 737 5861 781
rect 5809 729 5818 737
rect 5818 729 5852 737
rect 5852 729 5861 737
rect 6009 843 6018 851
rect 6018 843 6052 851
rect 6052 843 6061 851
rect 6009 799 6061 843
rect 6209 1017 6261 1061
rect 6209 1009 6218 1017
rect 6218 1009 6252 1017
rect 6252 1009 6261 1017
rect 6409 1123 6418 1131
rect 6418 1123 6452 1131
rect 6452 1123 6461 1131
rect 6409 1079 6461 1123
rect 6507 1079 6559 1131
rect 5009 70 5061 79
rect 5009 36 5018 70
rect 5018 36 5052 70
rect 5052 36 5061 70
rect 5009 27 5061 36
rect 4909 -60 4961 -15
rect 4909 -67 4918 -60
rect 4918 -67 4952 -60
rect 4952 -67 4961 -60
rect 4709 -166 4718 -143
rect 4718 -166 4752 -143
rect 4752 -166 4761 -143
rect 4709 -195 4761 -166
rect 4725 -248 4777 -239
rect 4725 -282 4734 -248
rect 4734 -282 4768 -248
rect 4768 -282 4777 -248
rect 4725 -291 4777 -282
rect 4709 -363 4761 -326
rect 4709 -378 4718 -363
rect 4718 -378 4752 -363
rect 4752 -378 4761 -363
rect 4709 -397 4718 -390
rect 4718 -397 4752 -390
rect 4752 -397 4761 -390
rect 4709 -435 4761 -397
rect 4709 -442 4718 -435
rect 4718 -442 4752 -435
rect 4752 -442 4761 -435
rect 4709 -469 4718 -454
rect 4718 -469 4752 -454
rect 4752 -469 4761 -454
rect 4709 -506 4761 -469
rect 4909 -94 4918 -79
rect 4918 -94 4952 -79
rect 4952 -94 4961 -79
rect 4909 -131 4961 -94
rect 5009 -74 5061 -22
rect 5209 143 5218 151
rect 5218 143 5252 151
rect 5252 143 5261 151
rect 5209 99 5261 143
rect 5409 317 5461 361
rect 5409 309 5418 317
rect 5418 309 5452 317
rect 5452 309 5461 317
rect 5609 423 5618 431
rect 5618 423 5652 431
rect 5652 423 5661 431
rect 5609 379 5661 423
rect 5809 597 5861 641
rect 5809 589 5818 597
rect 5818 589 5852 597
rect 5852 589 5861 597
rect 6009 703 6018 711
rect 6018 703 6052 711
rect 6052 703 6061 711
rect 6009 659 6061 703
rect 6209 877 6261 921
rect 6209 869 6218 877
rect 6218 869 6252 877
rect 6252 869 6261 877
rect 6409 983 6418 991
rect 6418 983 6452 991
rect 6452 983 6461 991
rect 6409 939 6461 983
rect 6507 939 6559 991
rect 5209 54 5261 63
rect 5209 20 5218 54
rect 5218 20 5252 54
rect 5252 20 5261 54
rect 5209 11 5261 20
rect 5109 -60 5161 -15
rect 5109 -67 5118 -60
rect 5118 -67 5152 -60
rect 5152 -67 5161 -60
rect 4909 -166 4918 -143
rect 4918 -166 4952 -143
rect 4952 -166 4961 -143
rect 4909 -195 4961 -166
rect 4925 -248 4977 -239
rect 4925 -282 4934 -248
rect 4934 -282 4968 -248
rect 4968 -282 4977 -248
rect 4925 -291 4977 -282
rect 4909 -363 4961 -326
rect 4909 -378 4918 -363
rect 4918 -378 4952 -363
rect 4952 -378 4961 -363
rect 4909 -397 4918 -390
rect 4918 -397 4952 -390
rect 4952 -397 4961 -390
rect 4909 -435 4961 -397
rect 4909 -442 4918 -435
rect 4918 -442 4952 -435
rect 4952 -442 4961 -435
rect 4909 -469 4918 -454
rect 4918 -469 4952 -454
rect 4952 -469 4961 -454
rect 4909 -506 4961 -469
rect 5109 -94 5118 -79
rect 5118 -94 5152 -79
rect 5152 -94 5161 -79
rect 5109 -131 5161 -94
rect 5209 -74 5261 -22
rect 5409 177 5461 221
rect 5409 169 5418 177
rect 5418 169 5452 177
rect 5452 169 5461 177
rect 5609 283 5618 291
rect 5618 283 5652 291
rect 5652 283 5661 291
rect 5609 239 5661 283
rect 5809 457 5861 501
rect 5809 449 5818 457
rect 5818 449 5852 457
rect 5852 449 5861 457
rect 6009 563 6018 571
rect 6018 563 6052 571
rect 6052 563 6061 571
rect 6009 519 6061 563
rect 6209 737 6261 781
rect 6209 729 6218 737
rect 6218 729 6252 737
rect 6252 729 6261 737
rect 6409 843 6418 851
rect 6418 843 6452 851
rect 6452 843 6461 851
rect 6409 799 6461 843
rect 6507 799 6559 851
rect 5409 70 5461 79
rect 5409 36 5418 70
rect 5418 36 5452 70
rect 5452 36 5461 70
rect 5409 27 5461 36
rect 5309 -60 5361 -15
rect 5309 -67 5318 -60
rect 5318 -67 5352 -60
rect 5352 -67 5361 -60
rect 5109 -166 5118 -143
rect 5118 -166 5152 -143
rect 5152 -166 5161 -143
rect 5109 -195 5161 -166
rect 5125 -248 5177 -239
rect 5125 -282 5134 -248
rect 5134 -282 5168 -248
rect 5168 -282 5177 -248
rect 5125 -291 5177 -282
rect 5109 -363 5161 -326
rect 5109 -378 5118 -363
rect 5118 -378 5152 -363
rect 5152 -378 5161 -363
rect 5109 -397 5118 -390
rect 5118 -397 5152 -390
rect 5152 -397 5161 -390
rect 5109 -435 5161 -397
rect 5109 -442 5118 -435
rect 5118 -442 5152 -435
rect 5152 -442 5161 -435
rect 5109 -469 5118 -454
rect 5118 -469 5152 -454
rect 5152 -469 5161 -454
rect 5109 -506 5161 -469
rect 5309 -94 5318 -79
rect 5318 -94 5352 -79
rect 5352 -94 5361 -79
rect 5309 -131 5361 -94
rect 5409 -74 5461 -22
rect 5609 143 5618 151
rect 5618 143 5652 151
rect 5652 143 5661 151
rect 5609 99 5661 143
rect 5809 317 5861 361
rect 5809 309 5818 317
rect 5818 309 5852 317
rect 5852 309 5861 317
rect 6009 423 6018 431
rect 6018 423 6052 431
rect 6052 423 6061 431
rect 6009 379 6061 423
rect 6209 597 6261 641
rect 6209 589 6218 597
rect 6218 589 6252 597
rect 6252 589 6261 597
rect 6409 703 6418 711
rect 6418 703 6452 711
rect 6452 703 6461 711
rect 6409 659 6461 703
rect 6507 659 6559 711
rect 5609 54 5661 63
rect 5609 20 5618 54
rect 5618 20 5652 54
rect 5652 20 5661 54
rect 5609 11 5661 20
rect 5509 -60 5561 -15
rect 5509 -67 5518 -60
rect 5518 -67 5552 -60
rect 5552 -67 5561 -60
rect 5309 -166 5318 -143
rect 5318 -166 5352 -143
rect 5352 -166 5361 -143
rect 5309 -195 5361 -166
rect 5325 -248 5377 -239
rect 5325 -282 5334 -248
rect 5334 -282 5368 -248
rect 5368 -282 5377 -248
rect 5325 -291 5377 -282
rect 5309 -363 5361 -326
rect 5309 -378 5318 -363
rect 5318 -378 5352 -363
rect 5352 -378 5361 -363
rect 5309 -397 5318 -390
rect 5318 -397 5352 -390
rect 5352 -397 5361 -390
rect 5309 -435 5361 -397
rect 5309 -442 5318 -435
rect 5318 -442 5352 -435
rect 5352 -442 5361 -435
rect 5309 -469 5318 -454
rect 5318 -469 5352 -454
rect 5352 -469 5361 -454
rect 5309 -506 5361 -469
rect 5509 -94 5518 -79
rect 5518 -94 5552 -79
rect 5552 -94 5561 -79
rect 5509 -131 5561 -94
rect 5609 -74 5661 -22
rect 5809 177 5861 221
rect 5809 169 5818 177
rect 5818 169 5852 177
rect 5852 169 5861 177
rect 6009 283 6018 291
rect 6018 283 6052 291
rect 6052 283 6061 291
rect 6009 239 6061 283
rect 6209 457 6261 501
rect 6209 449 6218 457
rect 6218 449 6252 457
rect 6252 449 6261 457
rect 6409 563 6418 571
rect 6418 563 6452 571
rect 6452 563 6461 571
rect 6409 519 6461 563
rect 6507 519 6559 571
rect 5809 70 5861 79
rect 5809 36 5818 70
rect 5818 36 5852 70
rect 5852 36 5861 70
rect 5809 27 5861 36
rect 5709 -60 5761 -15
rect 5709 -67 5718 -60
rect 5718 -67 5752 -60
rect 5752 -67 5761 -60
rect 5509 -166 5518 -143
rect 5518 -166 5552 -143
rect 5552 -166 5561 -143
rect 5509 -195 5561 -166
rect 5525 -248 5577 -239
rect 5525 -282 5534 -248
rect 5534 -282 5568 -248
rect 5568 -282 5577 -248
rect 5525 -291 5577 -282
rect 5509 -363 5561 -326
rect 5509 -378 5518 -363
rect 5518 -378 5552 -363
rect 5552 -378 5561 -363
rect 5509 -397 5518 -390
rect 5518 -397 5552 -390
rect 5552 -397 5561 -390
rect 5509 -435 5561 -397
rect 5509 -442 5518 -435
rect 5518 -442 5552 -435
rect 5552 -442 5561 -435
rect 5509 -469 5518 -454
rect 5518 -469 5552 -454
rect 5552 -469 5561 -454
rect 5509 -506 5561 -469
rect 5709 -94 5718 -79
rect 5718 -94 5752 -79
rect 5752 -94 5761 -79
rect 5709 -131 5761 -94
rect 5809 -74 5861 -22
rect 6009 143 6018 151
rect 6018 143 6052 151
rect 6052 143 6061 151
rect 6009 99 6061 143
rect 6209 317 6261 361
rect 6209 309 6218 317
rect 6218 309 6252 317
rect 6252 309 6261 317
rect 6409 423 6418 431
rect 6418 423 6452 431
rect 6452 423 6461 431
rect 6409 379 6461 423
rect 6507 379 6559 431
rect 6009 54 6061 63
rect 6009 20 6018 54
rect 6018 20 6052 54
rect 6052 20 6061 54
rect 6009 11 6061 20
rect 5909 -60 5961 -15
rect 5909 -67 5918 -60
rect 5918 -67 5952 -60
rect 5952 -67 5961 -60
rect 5709 -166 5718 -143
rect 5718 -166 5752 -143
rect 5752 -166 5761 -143
rect 5709 -195 5761 -166
rect 5725 -248 5777 -239
rect 5725 -282 5734 -248
rect 5734 -282 5768 -248
rect 5768 -282 5777 -248
rect 5725 -291 5777 -282
rect 5709 -363 5761 -326
rect 5709 -378 5718 -363
rect 5718 -378 5752 -363
rect 5752 -378 5761 -363
rect 5709 -397 5718 -390
rect 5718 -397 5752 -390
rect 5752 -397 5761 -390
rect 5709 -435 5761 -397
rect 5709 -442 5718 -435
rect 5718 -442 5752 -435
rect 5752 -442 5761 -435
rect 5709 -469 5718 -454
rect 5718 -469 5752 -454
rect 5752 -469 5761 -454
rect 5709 -506 5761 -469
rect 5909 -94 5918 -79
rect 5918 -94 5952 -79
rect 5952 -94 5961 -79
rect 5909 -131 5961 -94
rect 6009 -74 6061 -22
rect 6209 177 6261 221
rect 6209 169 6218 177
rect 6218 169 6252 177
rect 6252 169 6261 177
rect 6409 283 6418 291
rect 6418 283 6452 291
rect 6452 283 6461 291
rect 6409 239 6461 283
rect 6507 239 6559 291
rect 6209 70 6261 79
rect 6209 36 6218 70
rect 6218 36 6252 70
rect 6252 36 6261 70
rect 6209 27 6261 36
rect 6109 -60 6161 -15
rect 6109 -67 6118 -60
rect 6118 -67 6152 -60
rect 6152 -67 6161 -60
rect 5909 -166 5918 -143
rect 5918 -166 5952 -143
rect 5952 -166 5961 -143
rect 5909 -195 5961 -166
rect 5925 -248 5977 -239
rect 5925 -282 5934 -248
rect 5934 -282 5968 -248
rect 5968 -282 5977 -248
rect 5925 -291 5977 -282
rect 5909 -363 5961 -326
rect 5909 -378 5918 -363
rect 5918 -378 5952 -363
rect 5952 -378 5961 -363
rect 5909 -397 5918 -390
rect 5918 -397 5952 -390
rect 5952 -397 5961 -390
rect 5909 -435 5961 -397
rect 5909 -442 5918 -435
rect 5918 -442 5952 -435
rect 5952 -442 5961 -435
rect 5909 -469 5918 -454
rect 5918 -469 5952 -454
rect 5952 -469 5961 -454
rect 5909 -506 5961 -469
rect 6109 -94 6118 -79
rect 6118 -94 6152 -79
rect 6152 -94 6161 -79
rect 6109 -131 6161 -94
rect 6209 -74 6261 -22
rect 6409 143 6418 151
rect 6418 143 6452 151
rect 6452 143 6461 151
rect 6409 99 6461 143
rect 6507 99 6559 151
rect 6711 9759 6763 9811
rect 6711 9619 6763 9671
rect 6711 9479 6763 9531
rect 6711 9339 6763 9391
rect 6711 9199 6763 9251
rect 6711 9059 6763 9111
rect 6711 8919 6763 8971
rect 6711 8779 6763 8831
rect 6711 8549 6763 8601
rect 6711 8409 6763 8461
rect 6711 8269 6763 8321
rect 6711 8129 6763 8181
rect 6711 7989 6763 8041
rect 6711 7849 6763 7901
rect 6711 7709 6763 7761
rect 6711 7569 6763 7621
rect 6711 7339 6763 7391
rect 6711 7199 6763 7251
rect 6711 7059 6763 7111
rect 6711 6919 6763 6971
rect 6711 6779 6763 6831
rect 6711 6639 6763 6691
rect 6711 6499 6763 6551
rect 6711 6359 6763 6411
rect 6711 6129 6763 6181
rect 6711 5989 6763 6041
rect 6711 5849 6763 5901
rect 6711 5709 6763 5761
rect 6711 5569 6763 5621
rect 6711 5429 6763 5481
rect 6711 5289 6763 5341
rect 6711 5149 6763 5201
rect 6711 4779 6763 4831
rect 6711 4639 6763 4691
rect 6711 4499 6763 4551
rect 6711 4359 6763 4411
rect 6711 4219 6763 4271
rect 6711 4079 6763 4131
rect 6711 3939 6763 3991
rect 6711 3799 6763 3851
rect 6711 3569 6763 3621
rect 6711 3429 6763 3481
rect 6711 3289 6763 3341
rect 6711 3149 6763 3201
rect 6711 3009 6763 3061
rect 6711 2869 6763 2921
rect 6711 2729 6763 2781
rect 6711 2589 6763 2641
rect 6711 2359 6763 2411
rect 6711 2219 6763 2271
rect 6711 2079 6763 2131
rect 6711 1939 6763 1991
rect 6711 1799 6763 1851
rect 6711 1659 6763 1711
rect 6711 1519 6763 1571
rect 6711 1379 6763 1431
rect 6711 1149 6763 1201
rect 6711 1009 6763 1061
rect 6711 869 6763 921
rect 6711 729 6763 781
rect 6711 589 6763 641
rect 6711 449 6763 501
rect 6711 309 6763 361
rect 6711 169 6763 221
rect 6309 -60 6361 -15
rect 6309 -67 6318 -60
rect 6318 -67 6352 -60
rect 6352 -67 6361 -60
rect 8153 -8 8205 1
rect 8153 -42 8158 -8
rect 8158 -42 8192 -8
rect 8192 -42 8205 -8
rect 8153 -51 8205 -42
rect 8217 -8 8269 1
rect 8217 -42 8230 -8
rect 8230 -42 8264 -8
rect 8264 -42 8269 -8
rect 8217 -51 8269 -42
rect 8416 -8 8468 1
rect 8480 -8 8532 1
rect 8544 -8 8596 1
rect 8608 -8 8660 1
rect 8672 -8 8724 1
rect 8416 -42 8442 -8
rect 8442 -42 8468 -8
rect 8480 -42 8514 -8
rect 8514 -42 8532 -8
rect 8544 -42 8548 -8
rect 8548 -42 8586 -8
rect 8586 -42 8596 -8
rect 8608 -42 8620 -8
rect 8620 -42 8658 -8
rect 8658 -42 8660 -8
rect 8672 -42 8692 -8
rect 8692 -42 8724 -8
rect 8416 -51 8468 -42
rect 8480 -51 8532 -42
rect 8544 -51 8596 -42
rect 8608 -51 8660 -42
rect 8672 -51 8724 -42
rect 8817 -8 8869 1
rect 8881 -8 8933 1
rect 8945 -8 8997 1
rect 9009 -8 9061 1
rect 9073 -8 9125 1
rect 8817 -42 8849 -8
rect 8849 -42 8869 -8
rect 8881 -42 8883 -8
rect 8883 -42 8921 -8
rect 8921 -42 8933 -8
rect 8945 -42 8955 -8
rect 8955 -42 8993 -8
rect 8993 -42 8997 -8
rect 9009 -42 9027 -8
rect 9027 -42 9061 -8
rect 9073 -42 9099 -8
rect 9099 -42 9125 -8
rect 8817 -51 8869 -42
rect 8881 -51 8933 -42
rect 8945 -51 8997 -42
rect 9009 -51 9061 -42
rect 9073 -51 9125 -42
rect 9272 -8 9324 1
rect 9272 -42 9277 -8
rect 9277 -42 9311 -8
rect 9311 -42 9324 -8
rect 9272 -51 9324 -42
rect 9336 -8 9388 1
rect 9336 -42 9349 -8
rect 9349 -42 9383 -8
rect 9383 -42 9388 -8
rect 9336 -51 9388 -42
rect 6109 -166 6118 -143
rect 6118 -166 6152 -143
rect 6152 -166 6161 -143
rect 6109 -195 6161 -166
rect 6125 -248 6177 -239
rect 6125 -282 6134 -248
rect 6134 -282 6168 -248
rect 6168 -282 6177 -248
rect 6125 -291 6177 -282
rect 6109 -363 6161 -326
rect 6109 -378 6118 -363
rect 6118 -378 6152 -363
rect 6152 -378 6161 -363
rect 6109 -397 6118 -390
rect 6118 -397 6152 -390
rect 6152 -397 6161 -390
rect 6109 -435 6161 -397
rect 6109 -442 6118 -435
rect 6118 -442 6152 -435
rect 6152 -442 6161 -435
rect 6109 -469 6118 -454
rect 6118 -469 6152 -454
rect 6152 -469 6161 -454
rect 6109 -506 6161 -469
rect 6309 -94 6318 -79
rect 6318 -94 6352 -79
rect 6352 -94 6361 -79
rect 6309 -131 6361 -94
rect 6309 -166 6318 -143
rect 6318 -166 6352 -143
rect 6352 -166 6361 -143
rect 6309 -195 6361 -166
rect 8812 -108 8864 -99
rect 8812 -142 8851 -108
rect 8851 -142 8864 -108
rect 8812 -151 8864 -142
rect 8040 -251 8092 -199
rect 8153 -208 8205 -199
rect 8153 -242 8158 -208
rect 8158 -242 8192 -208
rect 8192 -242 8205 -208
rect 8153 -251 8205 -242
rect 8217 -208 8269 -199
rect 8217 -242 8230 -208
rect 8230 -242 8264 -208
rect 8264 -242 8269 -208
rect 8217 -251 8269 -242
rect 8325 -208 8377 -199
rect 8325 -242 8334 -208
rect 8334 -242 8368 -208
rect 8368 -242 8377 -208
rect 8325 -251 8377 -242
rect 8416 -208 8468 -199
rect 8480 -208 8532 -199
rect 8544 -208 8596 -199
rect 8608 -208 8660 -199
rect 8672 -208 8724 -199
rect 8416 -242 8442 -208
rect 8442 -242 8468 -208
rect 8480 -242 8514 -208
rect 8514 -242 8532 -208
rect 8544 -242 8548 -208
rect 8548 -242 8586 -208
rect 8586 -242 8596 -208
rect 8608 -242 8620 -208
rect 8620 -242 8658 -208
rect 8658 -242 8660 -208
rect 8672 -242 8692 -208
rect 8692 -242 8724 -208
rect 8416 -251 8468 -242
rect 8480 -251 8532 -242
rect 8544 -251 8596 -242
rect 8608 -251 8660 -242
rect 8672 -251 8724 -242
rect 8817 -208 8869 -199
rect 8881 -208 8933 -199
rect 8945 -208 8997 -199
rect 9009 -208 9061 -199
rect 9073 -208 9125 -199
rect 8817 -242 8849 -208
rect 8849 -242 8869 -208
rect 8881 -242 8883 -208
rect 8883 -242 8921 -208
rect 8921 -242 8933 -208
rect 8945 -242 8955 -208
rect 8955 -242 8993 -208
rect 8993 -242 8997 -208
rect 9009 -242 9027 -208
rect 9027 -242 9061 -208
rect 9073 -242 9099 -208
rect 9099 -242 9125 -208
rect 8817 -251 8869 -242
rect 8881 -251 8933 -242
rect 8945 -251 8997 -242
rect 9009 -251 9061 -242
rect 9073 -251 9125 -242
rect 9165 -208 9217 -199
rect 9165 -242 9174 -208
rect 9174 -242 9208 -208
rect 9208 -242 9217 -208
rect 9165 -251 9217 -242
rect 9272 -208 9324 -199
rect 9272 -242 9277 -208
rect 9277 -242 9311 -208
rect 9311 -242 9324 -208
rect 9272 -251 9324 -242
rect 9336 -208 9388 -199
rect 9336 -242 9349 -208
rect 9349 -242 9383 -208
rect 9383 -242 9388 -208
rect 9336 -251 9388 -242
rect 6309 -363 6361 -326
rect 8812 -308 8864 -299
rect 8812 -342 8851 -308
rect 8851 -342 8864 -308
rect 8812 -351 8864 -342
rect 6309 -378 6318 -363
rect 6318 -378 6352 -363
rect 6352 -378 6361 -363
rect 6309 -397 6318 -390
rect 6318 -397 6352 -390
rect 6352 -397 6361 -390
rect 6309 -435 6361 -397
rect 6309 -442 6318 -435
rect 6318 -442 6352 -435
rect 6352 -442 6361 -435
rect 8040 -451 8092 -399
rect 8153 -408 8205 -399
rect 8153 -442 8158 -408
rect 8158 -442 8192 -408
rect 8192 -442 8205 -408
rect 8153 -451 8205 -442
rect 8217 -408 8269 -399
rect 8217 -442 8230 -408
rect 8230 -442 8264 -408
rect 8264 -442 8269 -408
rect 8217 -451 8269 -442
rect 6309 -469 6318 -454
rect 6318 -469 6352 -454
rect 6352 -469 6361 -454
rect 8325 -408 8377 -399
rect 8325 -442 8334 -408
rect 8334 -442 8368 -408
rect 8368 -442 8377 -408
rect 8325 -451 8377 -442
rect 8416 -408 8468 -399
rect 8480 -408 8532 -399
rect 8544 -408 8596 -399
rect 8608 -408 8660 -399
rect 8672 -408 8724 -399
rect 8416 -442 8442 -408
rect 8442 -442 8468 -408
rect 8480 -442 8514 -408
rect 8514 -442 8532 -408
rect 8544 -442 8548 -408
rect 8548 -442 8586 -408
rect 8586 -442 8596 -408
rect 8608 -442 8620 -408
rect 8620 -442 8658 -408
rect 8658 -442 8660 -408
rect 8672 -442 8692 -408
rect 8692 -442 8724 -408
rect 8416 -451 8468 -442
rect 8480 -451 8532 -442
rect 8544 -451 8596 -442
rect 8608 -451 8660 -442
rect 8672 -451 8724 -442
rect 8817 -408 8869 -399
rect 8881 -408 8933 -399
rect 8945 -408 8997 -399
rect 9009 -408 9061 -399
rect 9073 -408 9125 -399
rect 8817 -442 8849 -408
rect 8849 -442 8869 -408
rect 8881 -442 8883 -408
rect 8883 -442 8921 -408
rect 8921 -442 8933 -408
rect 8945 -442 8955 -408
rect 8955 -442 8993 -408
rect 8993 -442 8997 -408
rect 9009 -442 9027 -408
rect 9027 -442 9061 -408
rect 9073 -442 9099 -408
rect 9099 -442 9125 -408
rect 8817 -451 8869 -442
rect 8881 -451 8933 -442
rect 8945 -451 8997 -442
rect 9009 -451 9061 -442
rect 9073 -451 9125 -442
rect 9165 -408 9217 -399
rect 9165 -442 9174 -408
rect 9174 -442 9208 -408
rect 9208 -442 9217 -408
rect 9165 -451 9217 -442
rect 9272 -408 9324 -399
rect 9272 -442 9277 -408
rect 9277 -442 9311 -408
rect 9311 -442 9324 -408
rect 9272 -451 9324 -442
rect 9336 -408 9388 -399
rect 9336 -442 9349 -408
rect 9349 -442 9383 -408
rect 9383 -442 9388 -408
rect 9336 -451 9388 -442
rect 6309 -506 6361 -469
rect 8812 -508 8864 -499
rect 8812 -542 8851 -508
rect 8851 -542 8864 -508
rect 8812 -551 8864 -542
rect 8040 -651 8092 -599
rect 8153 -608 8205 -599
rect 8153 -642 8158 -608
rect 8158 -642 8192 -608
rect 8192 -642 8205 -608
rect 8153 -651 8205 -642
rect 8217 -608 8269 -599
rect 8217 -642 8230 -608
rect 8230 -642 8264 -608
rect 8264 -642 8269 -608
rect 8217 -651 8269 -642
rect 8325 -608 8377 -599
rect 8325 -642 8334 -608
rect 8334 -642 8368 -608
rect 8368 -642 8377 -608
rect 8325 -651 8377 -642
rect 8416 -608 8468 -599
rect 8480 -608 8532 -599
rect 8544 -608 8596 -599
rect 8608 -608 8660 -599
rect 8672 -608 8724 -599
rect 8416 -642 8442 -608
rect 8442 -642 8468 -608
rect 8480 -642 8514 -608
rect 8514 -642 8532 -608
rect 8544 -642 8548 -608
rect 8548 -642 8586 -608
rect 8586 -642 8596 -608
rect 8608 -642 8620 -608
rect 8620 -642 8658 -608
rect 8658 -642 8660 -608
rect 8672 -642 8692 -608
rect 8692 -642 8724 -608
rect 8416 -651 8468 -642
rect 8480 -651 8532 -642
rect 8544 -651 8596 -642
rect 8608 -651 8660 -642
rect 8672 -651 8724 -642
rect 8817 -608 8869 -599
rect 8881 -608 8933 -599
rect 8945 -608 8997 -599
rect 9009 -608 9061 -599
rect 9073 -608 9125 -599
rect 8817 -642 8849 -608
rect 8849 -642 8869 -608
rect 8881 -642 8883 -608
rect 8883 -642 8921 -608
rect 8921 -642 8933 -608
rect 8945 -642 8955 -608
rect 8955 -642 8993 -608
rect 8993 -642 8997 -608
rect 9009 -642 9027 -608
rect 9027 -642 9061 -608
rect 9073 -642 9099 -608
rect 9099 -642 9125 -608
rect 8817 -651 8869 -642
rect 8881 -651 8933 -642
rect 8945 -651 8997 -642
rect 9009 -651 9061 -642
rect 9073 -651 9125 -642
rect 9165 -608 9217 -599
rect 9165 -642 9174 -608
rect 9174 -642 9208 -608
rect 9208 -642 9217 -608
rect 9165 -651 9217 -642
rect 9272 -608 9324 -599
rect 9272 -642 9277 -608
rect 9277 -642 9311 -608
rect 9311 -642 9324 -608
rect 9272 -651 9324 -642
rect 9336 -608 9388 -599
rect 9336 -642 9349 -608
rect 9349 -642 9383 -608
rect 9383 -642 9388 -608
rect 9336 -651 9388 -642
rect 8812 -708 8864 -699
rect 8812 -742 8851 -708
rect 8851 -742 8864 -708
rect 8812 -751 8864 -742
rect -9 -837 43 -828
rect -9 -871 -4 -837
rect -4 -871 30 -837
rect 30 -871 43 -837
rect -9 -880 43 -871
rect 55 -837 107 -828
rect 55 -871 68 -837
rect 68 -871 102 -837
rect 102 -871 107 -837
rect 55 -880 107 -871
rect 163 -837 215 -828
rect 163 -871 168 -837
rect 168 -871 202 -837
rect 202 -871 215 -837
rect 163 -880 215 -871
rect 227 -837 279 -828
rect 227 -871 240 -837
rect 240 -871 274 -837
rect 274 -871 279 -837
rect 227 -880 279 -871
rect 391 -837 443 -828
rect 391 -871 396 -837
rect 396 -871 430 -837
rect 430 -871 443 -837
rect 391 -880 443 -871
rect 455 -837 507 -828
rect 455 -871 468 -837
rect 468 -871 502 -837
rect 502 -871 507 -837
rect 455 -880 507 -871
rect 563 -837 615 -828
rect 563 -871 568 -837
rect 568 -871 602 -837
rect 602 -871 615 -837
rect 563 -880 615 -871
rect 627 -837 679 -828
rect 627 -871 640 -837
rect 640 -871 674 -837
rect 674 -871 679 -837
rect 627 -880 679 -871
rect 791 -837 843 -828
rect 791 -871 796 -837
rect 796 -871 830 -837
rect 830 -871 843 -837
rect 791 -880 843 -871
rect 855 -837 907 -828
rect 855 -871 868 -837
rect 868 -871 902 -837
rect 902 -871 907 -837
rect 855 -880 907 -871
rect 963 -837 1015 -828
rect 963 -871 968 -837
rect 968 -871 1002 -837
rect 1002 -871 1015 -837
rect 963 -880 1015 -871
rect 1027 -837 1079 -828
rect 1027 -871 1040 -837
rect 1040 -871 1074 -837
rect 1074 -871 1079 -837
rect 1027 -880 1079 -871
rect 1191 -837 1243 -828
rect 1191 -871 1196 -837
rect 1196 -871 1230 -837
rect 1230 -871 1243 -837
rect 1191 -880 1243 -871
rect 1255 -837 1307 -828
rect 1255 -871 1268 -837
rect 1268 -871 1302 -837
rect 1302 -871 1307 -837
rect 1255 -880 1307 -871
rect 1363 -837 1415 -828
rect 1363 -871 1368 -837
rect 1368 -871 1402 -837
rect 1402 -871 1415 -837
rect 1363 -880 1415 -871
rect 1427 -837 1479 -828
rect 1427 -871 1440 -837
rect 1440 -871 1474 -837
rect 1474 -871 1479 -837
rect 1427 -880 1479 -871
rect 1591 -837 1643 -828
rect 1591 -871 1596 -837
rect 1596 -871 1630 -837
rect 1630 -871 1643 -837
rect 1591 -880 1643 -871
rect 1655 -837 1707 -828
rect 1655 -871 1668 -837
rect 1668 -871 1702 -837
rect 1702 -871 1707 -837
rect 1655 -880 1707 -871
rect 1763 -837 1815 -828
rect 1763 -871 1768 -837
rect 1768 -871 1802 -837
rect 1802 -871 1815 -837
rect 1763 -880 1815 -871
rect 1827 -837 1879 -828
rect 1827 -871 1840 -837
rect 1840 -871 1874 -837
rect 1874 -871 1879 -837
rect 1827 -880 1879 -871
rect 1991 -837 2043 -828
rect 1991 -871 1996 -837
rect 1996 -871 2030 -837
rect 2030 -871 2043 -837
rect 1991 -880 2043 -871
rect 2055 -837 2107 -828
rect 2055 -871 2068 -837
rect 2068 -871 2102 -837
rect 2102 -871 2107 -837
rect 2055 -880 2107 -871
rect 2163 -837 2215 -828
rect 2163 -871 2168 -837
rect 2168 -871 2202 -837
rect 2202 -871 2215 -837
rect 2163 -880 2215 -871
rect 2227 -837 2279 -828
rect 2227 -871 2240 -837
rect 2240 -871 2274 -837
rect 2274 -871 2279 -837
rect 2227 -880 2279 -871
rect 2391 -837 2443 -828
rect 2391 -871 2396 -837
rect 2396 -871 2430 -837
rect 2430 -871 2443 -837
rect 2391 -880 2443 -871
rect 2455 -837 2507 -828
rect 2455 -871 2468 -837
rect 2468 -871 2502 -837
rect 2502 -871 2507 -837
rect 2455 -880 2507 -871
rect 2563 -837 2615 -828
rect 2563 -871 2568 -837
rect 2568 -871 2602 -837
rect 2602 -871 2615 -837
rect 2563 -880 2615 -871
rect 2627 -837 2679 -828
rect 2627 -871 2640 -837
rect 2640 -871 2674 -837
rect 2674 -871 2679 -837
rect 2627 -880 2679 -871
rect 2791 -837 2843 -828
rect 2791 -871 2796 -837
rect 2796 -871 2830 -837
rect 2830 -871 2843 -837
rect 2791 -880 2843 -871
rect 2855 -837 2907 -828
rect 2855 -871 2868 -837
rect 2868 -871 2902 -837
rect 2902 -871 2907 -837
rect 2855 -880 2907 -871
rect 2963 -837 3015 -828
rect 2963 -871 2968 -837
rect 2968 -871 3002 -837
rect 3002 -871 3015 -837
rect 2963 -880 3015 -871
rect 3027 -837 3079 -828
rect 3027 -871 3040 -837
rect 3040 -871 3074 -837
rect 3074 -871 3079 -837
rect 3027 -880 3079 -871
rect 3191 -837 3243 -828
rect 3191 -871 3196 -837
rect 3196 -871 3230 -837
rect 3230 -871 3243 -837
rect 3191 -880 3243 -871
rect 3255 -837 3307 -828
rect 3255 -871 3268 -837
rect 3268 -871 3302 -837
rect 3302 -871 3307 -837
rect 3255 -880 3307 -871
rect 3363 -837 3415 -828
rect 3363 -871 3368 -837
rect 3368 -871 3402 -837
rect 3402 -871 3415 -837
rect 3363 -880 3415 -871
rect 3427 -837 3479 -828
rect 3427 -871 3440 -837
rect 3440 -871 3474 -837
rect 3474 -871 3479 -837
rect 3427 -880 3479 -871
rect 3591 -837 3643 -828
rect 3591 -871 3596 -837
rect 3596 -871 3630 -837
rect 3630 -871 3643 -837
rect 3591 -880 3643 -871
rect 3655 -837 3707 -828
rect 3655 -871 3668 -837
rect 3668 -871 3702 -837
rect 3702 -871 3707 -837
rect 3655 -880 3707 -871
rect 3763 -837 3815 -828
rect 3763 -871 3768 -837
rect 3768 -871 3802 -837
rect 3802 -871 3815 -837
rect 3763 -880 3815 -871
rect 3827 -837 3879 -828
rect 3827 -871 3840 -837
rect 3840 -871 3874 -837
rect 3874 -871 3879 -837
rect 3827 -880 3879 -871
rect 3991 -837 4043 -828
rect 3991 -871 3996 -837
rect 3996 -871 4030 -837
rect 4030 -871 4043 -837
rect 3991 -880 4043 -871
rect 4055 -837 4107 -828
rect 4055 -871 4068 -837
rect 4068 -871 4102 -837
rect 4102 -871 4107 -837
rect 4055 -880 4107 -871
rect 4163 -837 4215 -828
rect 4163 -871 4168 -837
rect 4168 -871 4202 -837
rect 4202 -871 4215 -837
rect 4163 -880 4215 -871
rect 4227 -837 4279 -828
rect 4227 -871 4240 -837
rect 4240 -871 4274 -837
rect 4274 -871 4279 -837
rect 4227 -880 4279 -871
rect 4391 -837 4443 -828
rect 4391 -871 4396 -837
rect 4396 -871 4430 -837
rect 4430 -871 4443 -837
rect 4391 -880 4443 -871
rect 4455 -837 4507 -828
rect 4455 -871 4468 -837
rect 4468 -871 4502 -837
rect 4502 -871 4507 -837
rect 4455 -880 4507 -871
rect 4563 -837 4615 -828
rect 4563 -871 4568 -837
rect 4568 -871 4602 -837
rect 4602 -871 4615 -837
rect 4563 -880 4615 -871
rect 4627 -837 4679 -828
rect 4627 -871 4640 -837
rect 4640 -871 4674 -837
rect 4674 -871 4679 -837
rect 4627 -880 4679 -871
rect 4791 -837 4843 -828
rect 4791 -871 4796 -837
rect 4796 -871 4830 -837
rect 4830 -871 4843 -837
rect 4791 -880 4843 -871
rect 4855 -837 4907 -828
rect 4855 -871 4868 -837
rect 4868 -871 4902 -837
rect 4902 -871 4907 -837
rect 4855 -880 4907 -871
rect 4963 -837 5015 -828
rect 4963 -871 4968 -837
rect 4968 -871 5002 -837
rect 5002 -871 5015 -837
rect 4963 -880 5015 -871
rect 5027 -837 5079 -828
rect 5027 -871 5040 -837
rect 5040 -871 5074 -837
rect 5074 -871 5079 -837
rect 5027 -880 5079 -871
rect 5191 -837 5243 -828
rect 5191 -871 5196 -837
rect 5196 -871 5230 -837
rect 5230 -871 5243 -837
rect 5191 -880 5243 -871
rect 5255 -837 5307 -828
rect 5255 -871 5268 -837
rect 5268 -871 5302 -837
rect 5302 -871 5307 -837
rect 5255 -880 5307 -871
rect 5363 -837 5415 -828
rect 5363 -871 5368 -837
rect 5368 -871 5402 -837
rect 5402 -871 5415 -837
rect 5363 -880 5415 -871
rect 5427 -837 5479 -828
rect 5427 -871 5440 -837
rect 5440 -871 5474 -837
rect 5474 -871 5479 -837
rect 5427 -880 5479 -871
rect 5591 -837 5643 -828
rect 5591 -871 5596 -837
rect 5596 -871 5630 -837
rect 5630 -871 5643 -837
rect 5591 -880 5643 -871
rect 5655 -837 5707 -828
rect 5655 -871 5668 -837
rect 5668 -871 5702 -837
rect 5702 -871 5707 -837
rect 5655 -880 5707 -871
rect 5763 -837 5815 -828
rect 5763 -871 5768 -837
rect 5768 -871 5802 -837
rect 5802 -871 5815 -837
rect 5763 -880 5815 -871
rect 5827 -837 5879 -828
rect 5827 -871 5840 -837
rect 5840 -871 5874 -837
rect 5874 -871 5879 -837
rect 5827 -880 5879 -871
rect 5991 -837 6043 -828
rect 5991 -871 5996 -837
rect 5996 -871 6030 -837
rect 6030 -871 6043 -837
rect 5991 -880 6043 -871
rect 6055 -837 6107 -828
rect 6055 -871 6068 -837
rect 6068 -871 6102 -837
rect 6102 -871 6107 -837
rect 6055 -880 6107 -871
rect 6163 -837 6215 -828
rect 6163 -871 6168 -837
rect 6168 -871 6202 -837
rect 6202 -871 6215 -837
rect 6163 -880 6215 -871
rect 6227 -837 6279 -828
rect 6227 -871 6240 -837
rect 6240 -871 6274 -837
rect 6274 -871 6279 -837
rect 6227 -880 6279 -871
rect 8040 -851 8092 -799
rect 8153 -808 8205 -799
rect 8153 -842 8158 -808
rect 8158 -842 8192 -808
rect 8192 -842 8205 -808
rect 8153 -851 8205 -842
rect 8217 -808 8269 -799
rect 8217 -842 8230 -808
rect 8230 -842 8264 -808
rect 8264 -842 8269 -808
rect 8217 -851 8269 -842
rect 8325 -808 8377 -799
rect 8325 -842 8334 -808
rect 8334 -842 8368 -808
rect 8368 -842 8377 -808
rect 8325 -851 8377 -842
rect 8416 -808 8468 -799
rect 8480 -808 8532 -799
rect 8544 -808 8596 -799
rect 8608 -808 8660 -799
rect 8672 -808 8724 -799
rect 8416 -842 8442 -808
rect 8442 -842 8468 -808
rect 8480 -842 8514 -808
rect 8514 -842 8532 -808
rect 8544 -842 8548 -808
rect 8548 -842 8586 -808
rect 8586 -842 8596 -808
rect 8608 -842 8620 -808
rect 8620 -842 8658 -808
rect 8658 -842 8660 -808
rect 8672 -842 8692 -808
rect 8692 -842 8724 -808
rect 8416 -851 8468 -842
rect 8480 -851 8532 -842
rect 8544 -851 8596 -842
rect 8608 -851 8660 -842
rect 8672 -851 8724 -842
rect 8817 -808 8869 -799
rect 8881 -808 8933 -799
rect 8945 -808 8997 -799
rect 9009 -808 9061 -799
rect 9073 -808 9125 -799
rect 8817 -842 8849 -808
rect 8849 -842 8869 -808
rect 8881 -842 8883 -808
rect 8883 -842 8921 -808
rect 8921 -842 8933 -808
rect 8945 -842 8955 -808
rect 8955 -842 8993 -808
rect 8993 -842 8997 -808
rect 9009 -842 9027 -808
rect 9027 -842 9061 -808
rect 9073 -842 9099 -808
rect 9099 -842 9125 -808
rect 8817 -851 8869 -842
rect 8881 -851 8933 -842
rect 8945 -851 8997 -842
rect 9009 -851 9061 -842
rect 9073 -851 9125 -842
rect 9165 -808 9217 -799
rect 9165 -842 9174 -808
rect 9174 -842 9208 -808
rect 9208 -842 9217 -808
rect 9165 -851 9217 -842
rect 9272 -808 9324 -799
rect 9272 -842 9277 -808
rect 9277 -842 9311 -808
rect 9311 -842 9324 -808
rect 9272 -851 9324 -842
rect 9336 -808 9388 -799
rect 9336 -842 9349 -808
rect 9349 -842 9383 -808
rect 9383 -842 9388 -808
rect 9336 -851 9388 -842
rect 8812 -908 8864 -899
rect 8812 -942 8851 -908
rect 8851 -942 8864 -908
rect 8812 -951 8864 -942
rect 8040 -1051 8092 -999
rect 8153 -1008 8205 -999
rect 8153 -1042 8158 -1008
rect 8158 -1042 8192 -1008
rect 8192 -1042 8205 -1008
rect 8153 -1051 8205 -1042
rect 8217 -1008 8269 -999
rect 8217 -1042 8230 -1008
rect 8230 -1042 8264 -1008
rect 8264 -1042 8269 -1008
rect 8217 -1051 8269 -1042
rect 8325 -1008 8377 -999
rect 8325 -1042 8334 -1008
rect 8334 -1042 8368 -1008
rect 8368 -1042 8377 -1008
rect 8325 -1051 8377 -1042
rect 8416 -1008 8468 -999
rect 8480 -1008 8532 -999
rect 8544 -1008 8596 -999
rect 8608 -1008 8660 -999
rect 8672 -1008 8724 -999
rect 8416 -1042 8442 -1008
rect 8442 -1042 8468 -1008
rect 8480 -1042 8514 -1008
rect 8514 -1042 8532 -1008
rect 8544 -1042 8548 -1008
rect 8548 -1042 8586 -1008
rect 8586 -1042 8596 -1008
rect 8608 -1042 8620 -1008
rect 8620 -1042 8658 -1008
rect 8658 -1042 8660 -1008
rect 8672 -1042 8692 -1008
rect 8692 -1042 8724 -1008
rect 8416 -1051 8468 -1042
rect 8480 -1051 8532 -1042
rect 8544 -1051 8596 -1042
rect 8608 -1051 8660 -1042
rect 8672 -1051 8724 -1042
rect 8817 -1008 8869 -999
rect 8881 -1008 8933 -999
rect 8945 -1008 8997 -999
rect 9009 -1008 9061 -999
rect 9073 -1008 9125 -999
rect 8817 -1042 8849 -1008
rect 8849 -1042 8869 -1008
rect 8881 -1042 8883 -1008
rect 8883 -1042 8921 -1008
rect 8921 -1042 8933 -1008
rect 8945 -1042 8955 -1008
rect 8955 -1042 8993 -1008
rect 8993 -1042 8997 -1008
rect 9009 -1042 9027 -1008
rect 9027 -1042 9061 -1008
rect 9073 -1042 9099 -1008
rect 9099 -1042 9125 -1008
rect 8817 -1051 8869 -1042
rect 8881 -1051 8933 -1042
rect 8945 -1051 8997 -1042
rect 9009 -1051 9061 -1042
rect 9073 -1051 9125 -1042
rect 9165 -1008 9217 -999
rect 9165 -1042 9174 -1008
rect 9174 -1042 9208 -1008
rect 9208 -1042 9217 -1008
rect 9165 -1051 9217 -1042
rect 9272 -1008 9324 -999
rect 9272 -1042 9277 -1008
rect 9277 -1042 9311 -1008
rect 9311 -1042 9324 -1008
rect 9272 -1051 9324 -1042
rect 9336 -1008 9388 -999
rect 9336 -1042 9349 -1008
rect 9349 -1042 9383 -1008
rect 9383 -1042 9388 -1008
rect 9336 -1051 9388 -1042
rect 8812 -1108 8864 -1099
rect 8812 -1142 8851 -1108
rect 8851 -1142 8864 -1108
rect 8812 -1151 8864 -1142
rect 8040 -1251 8092 -1199
rect 8153 -1208 8205 -1199
rect 8153 -1242 8158 -1208
rect 8158 -1242 8192 -1208
rect 8192 -1242 8205 -1208
rect 8153 -1251 8205 -1242
rect 8217 -1208 8269 -1199
rect 8217 -1242 8230 -1208
rect 8230 -1242 8264 -1208
rect 8264 -1242 8269 -1208
rect 8217 -1251 8269 -1242
rect 8325 -1208 8377 -1199
rect 8325 -1242 8334 -1208
rect 8334 -1242 8368 -1208
rect 8368 -1242 8377 -1208
rect 8325 -1251 8377 -1242
rect 8416 -1208 8468 -1199
rect 8480 -1208 8532 -1199
rect 8544 -1208 8596 -1199
rect 8608 -1208 8660 -1199
rect 8672 -1208 8724 -1199
rect 8416 -1242 8442 -1208
rect 8442 -1242 8468 -1208
rect 8480 -1242 8514 -1208
rect 8514 -1242 8532 -1208
rect 8544 -1242 8548 -1208
rect 8548 -1242 8586 -1208
rect 8586 -1242 8596 -1208
rect 8608 -1242 8620 -1208
rect 8620 -1242 8658 -1208
rect 8658 -1242 8660 -1208
rect 8672 -1242 8692 -1208
rect 8692 -1242 8724 -1208
rect 8416 -1251 8468 -1242
rect 8480 -1251 8532 -1242
rect 8544 -1251 8596 -1242
rect 8608 -1251 8660 -1242
rect 8672 -1251 8724 -1242
rect 8817 -1208 8869 -1199
rect 8881 -1208 8933 -1199
rect 8945 -1208 8997 -1199
rect 9009 -1208 9061 -1199
rect 9073 -1208 9125 -1199
rect 8817 -1242 8849 -1208
rect 8849 -1242 8869 -1208
rect 8881 -1242 8883 -1208
rect 8883 -1242 8921 -1208
rect 8921 -1242 8933 -1208
rect 8945 -1242 8955 -1208
rect 8955 -1242 8993 -1208
rect 8993 -1242 8997 -1208
rect 9009 -1242 9027 -1208
rect 9027 -1242 9061 -1208
rect 9073 -1242 9099 -1208
rect 9099 -1242 9125 -1208
rect 8817 -1251 8869 -1242
rect 8881 -1251 8933 -1242
rect 8945 -1251 8997 -1242
rect 9009 -1251 9061 -1242
rect 9073 -1251 9125 -1242
rect 9165 -1208 9217 -1199
rect 9165 -1242 9174 -1208
rect 9174 -1242 9208 -1208
rect 9208 -1242 9217 -1208
rect 9165 -1251 9217 -1242
rect 9272 -1208 9324 -1199
rect 9272 -1242 9277 -1208
rect 9277 -1242 9311 -1208
rect 9311 -1242 9324 -1208
rect 9272 -1251 9324 -1242
rect 9336 -1208 9388 -1199
rect 9336 -1242 9349 -1208
rect 9349 -1242 9383 -1208
rect 9383 -1242 9388 -1208
rect 9336 -1251 9388 -1242
rect 8812 -1308 8864 -1299
rect 8812 -1342 8851 -1308
rect 8851 -1342 8864 -1308
rect 8812 -1351 8864 -1342
rect 8040 -1451 8092 -1399
rect 8153 -1408 8205 -1399
rect 8153 -1442 8158 -1408
rect 8158 -1442 8192 -1408
rect 8192 -1442 8205 -1408
rect 8153 -1451 8205 -1442
rect 8217 -1408 8269 -1399
rect 8217 -1442 8230 -1408
rect 8230 -1442 8264 -1408
rect 8264 -1442 8269 -1408
rect 8217 -1451 8269 -1442
rect 8325 -1408 8377 -1399
rect 8325 -1442 8334 -1408
rect 8334 -1442 8368 -1408
rect 8368 -1442 8377 -1408
rect 8325 -1451 8377 -1442
rect 8416 -1408 8468 -1399
rect 8480 -1408 8532 -1399
rect 8544 -1408 8596 -1399
rect 8608 -1408 8660 -1399
rect 8672 -1408 8724 -1399
rect 8416 -1442 8442 -1408
rect 8442 -1442 8468 -1408
rect 8480 -1442 8514 -1408
rect 8514 -1442 8532 -1408
rect 8544 -1442 8548 -1408
rect 8548 -1442 8586 -1408
rect 8586 -1442 8596 -1408
rect 8608 -1442 8620 -1408
rect 8620 -1442 8658 -1408
rect 8658 -1442 8660 -1408
rect 8672 -1442 8692 -1408
rect 8692 -1442 8724 -1408
rect 8416 -1451 8468 -1442
rect 8480 -1451 8532 -1442
rect 8544 -1451 8596 -1442
rect 8608 -1451 8660 -1442
rect 8672 -1451 8724 -1442
rect 8817 -1408 8869 -1399
rect 8881 -1408 8933 -1399
rect 8945 -1408 8997 -1399
rect 9009 -1408 9061 -1399
rect 9073 -1408 9125 -1399
rect 8817 -1442 8849 -1408
rect 8849 -1442 8869 -1408
rect 8881 -1442 8883 -1408
rect 8883 -1442 8921 -1408
rect 8921 -1442 8933 -1408
rect 8945 -1442 8955 -1408
rect 8955 -1442 8993 -1408
rect 8993 -1442 8997 -1408
rect 9009 -1442 9027 -1408
rect 9027 -1442 9061 -1408
rect 9073 -1442 9099 -1408
rect 9099 -1442 9125 -1408
rect 8817 -1451 8869 -1442
rect 8881 -1451 8933 -1442
rect 8945 -1451 8997 -1442
rect 9009 -1451 9061 -1442
rect 9073 -1451 9125 -1442
rect 9165 -1408 9217 -1399
rect 9165 -1442 9174 -1408
rect 9174 -1442 9208 -1408
rect 9208 -1442 9217 -1408
rect 9165 -1451 9217 -1442
rect 9272 -1408 9324 -1399
rect 9272 -1442 9277 -1408
rect 9277 -1442 9311 -1408
rect 9311 -1442 9324 -1408
rect 9272 -1451 9324 -1442
rect 9336 -1408 9388 -1399
rect 9336 -1442 9349 -1408
rect 9349 -1442 9383 -1408
rect 9383 -1442 9388 -1408
rect 9336 -1451 9388 -1442
rect 8812 -1508 8864 -1499
rect 8812 -1542 8851 -1508
rect 8851 -1542 8864 -1508
rect 8812 -1551 8864 -1542
rect 8040 -1651 8092 -1599
rect 8153 -1608 8205 -1599
rect 8153 -1642 8158 -1608
rect 8158 -1642 8192 -1608
rect 8192 -1642 8205 -1608
rect 8153 -1651 8205 -1642
rect 8217 -1608 8269 -1599
rect 8217 -1642 8230 -1608
rect 8230 -1642 8264 -1608
rect 8264 -1642 8269 -1608
rect 8217 -1651 8269 -1642
rect 8325 -1608 8377 -1599
rect 8325 -1642 8334 -1608
rect 8334 -1642 8368 -1608
rect 8368 -1642 8377 -1608
rect 8325 -1651 8377 -1642
rect 8416 -1608 8468 -1599
rect 8480 -1608 8532 -1599
rect 8544 -1608 8596 -1599
rect 8608 -1608 8660 -1599
rect 8672 -1608 8724 -1599
rect 8416 -1642 8442 -1608
rect 8442 -1642 8468 -1608
rect 8480 -1642 8514 -1608
rect 8514 -1642 8532 -1608
rect 8544 -1642 8548 -1608
rect 8548 -1642 8586 -1608
rect 8586 -1642 8596 -1608
rect 8608 -1642 8620 -1608
rect 8620 -1642 8658 -1608
rect 8658 -1642 8660 -1608
rect 8672 -1642 8692 -1608
rect 8692 -1642 8724 -1608
rect 8416 -1651 8468 -1642
rect 8480 -1651 8532 -1642
rect 8544 -1651 8596 -1642
rect 8608 -1651 8660 -1642
rect 8672 -1651 8724 -1642
rect 8817 -1608 8869 -1599
rect 8881 -1608 8933 -1599
rect 8945 -1608 8997 -1599
rect 9009 -1608 9061 -1599
rect 9073 -1608 9125 -1599
rect 8817 -1642 8849 -1608
rect 8849 -1642 8869 -1608
rect 8881 -1642 8883 -1608
rect 8883 -1642 8921 -1608
rect 8921 -1642 8933 -1608
rect 8945 -1642 8955 -1608
rect 8955 -1642 8993 -1608
rect 8993 -1642 8997 -1608
rect 9009 -1642 9027 -1608
rect 9027 -1642 9061 -1608
rect 9073 -1642 9099 -1608
rect 9099 -1642 9125 -1608
rect 8817 -1651 8869 -1642
rect 8881 -1651 8933 -1642
rect 8945 -1651 8997 -1642
rect 9009 -1651 9061 -1642
rect 9073 -1651 9125 -1642
rect 9165 -1608 9217 -1599
rect 9165 -1642 9174 -1608
rect 9174 -1642 9208 -1608
rect 9208 -1642 9217 -1608
rect 9165 -1651 9217 -1642
rect 9272 -1608 9324 -1599
rect 9272 -1642 9277 -1608
rect 9277 -1642 9311 -1608
rect 9311 -1642 9324 -1608
rect 9272 -1651 9324 -1642
rect 9336 -1608 9388 -1599
rect 9336 -1642 9349 -1608
rect 9349 -1642 9383 -1608
rect 9383 -1642 9388 -1608
rect 9336 -1651 9388 -1642
rect 8812 -1708 8864 -1699
rect 8812 -1742 8851 -1708
rect 8851 -1742 8864 -1708
rect 8812 -1751 8864 -1742
rect 8040 -1851 8092 -1799
rect 8153 -1808 8205 -1799
rect 8153 -1842 8158 -1808
rect 8158 -1842 8192 -1808
rect 8192 -1842 8205 -1808
rect 8153 -1851 8205 -1842
rect 8217 -1808 8269 -1799
rect 8217 -1842 8230 -1808
rect 8230 -1842 8264 -1808
rect 8264 -1842 8269 -1808
rect 8217 -1851 8269 -1842
rect 8325 -1808 8377 -1799
rect 8325 -1842 8334 -1808
rect 8334 -1842 8368 -1808
rect 8368 -1842 8377 -1808
rect 8325 -1851 8377 -1842
rect 8416 -1808 8468 -1799
rect 8480 -1808 8532 -1799
rect 8544 -1808 8596 -1799
rect 8608 -1808 8660 -1799
rect 8672 -1808 8724 -1799
rect 8416 -1842 8442 -1808
rect 8442 -1842 8468 -1808
rect 8480 -1842 8514 -1808
rect 8514 -1842 8532 -1808
rect 8544 -1842 8548 -1808
rect 8548 -1842 8586 -1808
rect 8586 -1842 8596 -1808
rect 8608 -1842 8620 -1808
rect 8620 -1842 8658 -1808
rect 8658 -1842 8660 -1808
rect 8672 -1842 8692 -1808
rect 8692 -1842 8724 -1808
rect 8416 -1851 8468 -1842
rect 8480 -1851 8532 -1842
rect 8544 -1851 8596 -1842
rect 8608 -1851 8660 -1842
rect 8672 -1851 8724 -1842
rect 8817 -1808 8869 -1799
rect 8881 -1808 8933 -1799
rect 8945 -1808 8997 -1799
rect 9009 -1808 9061 -1799
rect 9073 -1808 9125 -1799
rect 8817 -1842 8849 -1808
rect 8849 -1842 8869 -1808
rect 8881 -1842 8883 -1808
rect 8883 -1842 8921 -1808
rect 8921 -1842 8933 -1808
rect 8945 -1842 8955 -1808
rect 8955 -1842 8993 -1808
rect 8993 -1842 8997 -1808
rect 9009 -1842 9027 -1808
rect 9027 -1842 9061 -1808
rect 9073 -1842 9099 -1808
rect 9099 -1842 9125 -1808
rect 8817 -1851 8869 -1842
rect 8881 -1851 8933 -1842
rect 8945 -1851 8997 -1842
rect 9009 -1851 9061 -1842
rect 9073 -1851 9125 -1842
rect 9165 -1808 9217 -1799
rect 9165 -1842 9174 -1808
rect 9174 -1842 9208 -1808
rect 9208 -1842 9217 -1808
rect 9165 -1851 9217 -1842
rect 9272 -1808 9324 -1799
rect 9272 -1842 9277 -1808
rect 9277 -1842 9311 -1808
rect 9311 -1842 9324 -1808
rect 9272 -1851 9324 -1842
rect 9336 -1808 9388 -1799
rect 9336 -1842 9349 -1808
rect 9349 -1842 9383 -1808
rect 9383 -1842 9388 -1808
rect 9336 -1851 9388 -1842
<< metal2 >>
rect 196 9901 274 9902
rect -4 9885 74 9886
rect -4 9829 7 9885
rect 63 9829 74 9885
rect 196 9845 207 9901
rect 263 9845 274 9901
rect 596 9901 674 9902
rect 196 9844 274 9845
rect 396 9885 474 9886
rect -4 9828 74 9829
rect 396 9829 407 9885
rect 463 9829 474 9885
rect 596 9845 607 9901
rect 663 9845 674 9901
rect 996 9901 1074 9902
rect 596 9844 674 9845
rect 796 9885 874 9886
rect 396 9828 474 9829
rect 796 9829 807 9885
rect 863 9829 874 9885
rect 996 9845 1007 9901
rect 1063 9845 1074 9901
rect 1396 9901 1474 9902
rect 996 9844 1074 9845
rect 1196 9885 1274 9886
rect 796 9828 874 9829
rect 1196 9829 1207 9885
rect 1263 9829 1274 9885
rect 1396 9845 1407 9901
rect 1463 9845 1474 9901
rect 1796 9901 1874 9902
rect 1396 9844 1474 9845
rect 1596 9885 1674 9886
rect 1196 9828 1274 9829
rect 1596 9829 1607 9885
rect 1663 9829 1674 9885
rect 1796 9845 1807 9901
rect 1863 9845 1874 9901
rect 2196 9901 2274 9902
rect 1796 9844 1874 9845
rect 1996 9885 2074 9886
rect 1596 9828 1674 9829
rect 1996 9829 2007 9885
rect 2063 9829 2074 9885
rect 2196 9845 2207 9901
rect 2263 9845 2274 9901
rect 2596 9901 2674 9902
rect 2196 9844 2274 9845
rect 2396 9885 2474 9886
rect 1996 9828 2074 9829
rect 2396 9829 2407 9885
rect 2463 9829 2474 9885
rect 2596 9845 2607 9901
rect 2663 9845 2674 9901
rect 2996 9901 3074 9902
rect 2596 9844 2674 9845
rect 2796 9885 2874 9886
rect 2396 9828 2474 9829
rect 2796 9829 2807 9885
rect 2863 9829 2874 9885
rect 2996 9845 3007 9901
rect 3063 9845 3074 9901
rect 3396 9901 3474 9902
rect 2996 9844 3074 9845
rect 3196 9885 3274 9886
rect 2796 9828 2874 9829
rect 3196 9829 3207 9885
rect 3263 9829 3274 9885
rect 3396 9845 3407 9901
rect 3463 9845 3474 9901
rect 3796 9901 3874 9902
rect 3396 9844 3474 9845
rect 3596 9885 3674 9886
rect 3196 9828 3274 9829
rect 3596 9829 3607 9885
rect 3663 9829 3674 9885
rect 3796 9845 3807 9901
rect 3863 9845 3874 9901
rect 4196 9901 4274 9902
rect 3796 9844 3874 9845
rect 3996 9885 4074 9886
rect 3596 9828 3674 9829
rect 3996 9829 4007 9885
rect 4063 9829 4074 9885
rect 4196 9845 4207 9901
rect 4263 9845 4274 9901
rect 4596 9901 4674 9902
rect 4196 9844 4274 9845
rect 4396 9885 4474 9886
rect 3996 9828 4074 9829
rect 4396 9829 4407 9885
rect 4463 9829 4474 9885
rect 4596 9845 4607 9901
rect 4663 9845 4674 9901
rect 4996 9901 5074 9902
rect 4596 9844 4674 9845
rect 4796 9885 4874 9886
rect 4396 9828 4474 9829
rect 4796 9829 4807 9885
rect 4863 9829 4874 9885
rect 4996 9845 5007 9901
rect 5063 9845 5074 9901
rect 5396 9901 5474 9902
rect 4996 9844 5074 9845
rect 5196 9885 5274 9886
rect 4796 9828 4874 9829
rect 5196 9829 5207 9885
rect 5263 9829 5274 9885
rect 5396 9845 5407 9901
rect 5463 9845 5474 9901
rect 5796 9901 5874 9902
rect 5396 9844 5474 9845
rect 5596 9885 5674 9886
rect 5196 9828 5274 9829
rect 5596 9829 5607 9885
rect 5663 9829 5674 9885
rect 5796 9845 5807 9901
rect 5863 9845 5874 9901
rect 6196 9901 6274 9902
rect 5796 9844 5874 9845
rect 5996 9885 6074 9886
rect 5596 9828 5674 9829
rect 5996 9829 6007 9885
rect 6063 9829 6074 9885
rect 6196 9845 6207 9901
rect 6263 9845 6274 9901
rect 6196 9844 6274 9845
rect 5996 9828 6074 9829
rect 202 9811 268 9812
rect 202 9800 209 9811
rect 0 9770 209 9800
rect 202 9759 209 9770
rect 261 9800 268 9811
rect 602 9811 668 9812
rect 602 9800 609 9811
rect 261 9770 609 9800
rect 261 9759 268 9770
rect 202 9758 268 9759
rect 602 9759 609 9770
rect 661 9800 668 9811
rect 1002 9811 1068 9812
rect 1002 9800 1009 9811
rect 661 9770 1009 9800
rect 661 9759 668 9770
rect 602 9758 668 9759
rect 1002 9759 1009 9770
rect 1061 9800 1068 9811
rect 1402 9811 1468 9812
rect 1402 9800 1409 9811
rect 1061 9770 1409 9800
rect 1061 9759 1068 9770
rect 1002 9758 1068 9759
rect 1402 9759 1409 9770
rect 1461 9800 1468 9811
rect 1802 9811 1868 9812
rect 1802 9800 1809 9811
rect 1461 9770 1809 9800
rect 1461 9759 1468 9770
rect 1402 9758 1468 9759
rect 1802 9759 1809 9770
rect 1861 9800 1868 9811
rect 2202 9811 2268 9812
rect 2202 9800 2209 9811
rect 1861 9770 2209 9800
rect 1861 9759 1868 9770
rect 1802 9758 1868 9759
rect 2202 9759 2209 9770
rect 2261 9800 2268 9811
rect 2602 9811 2668 9812
rect 2602 9800 2609 9811
rect 2261 9770 2609 9800
rect 2261 9759 2268 9770
rect 2202 9758 2268 9759
rect 2602 9759 2609 9770
rect 2661 9800 2668 9811
rect 3002 9811 3068 9812
rect 3002 9800 3009 9811
rect 2661 9770 3009 9800
rect 2661 9759 2668 9770
rect 2602 9758 2668 9759
rect 3002 9759 3009 9770
rect 3061 9800 3068 9811
rect 3402 9811 3468 9812
rect 3402 9800 3409 9811
rect 3061 9770 3409 9800
rect 3061 9759 3068 9770
rect 3002 9758 3068 9759
rect 3402 9759 3409 9770
rect 3461 9800 3468 9811
rect 3802 9811 3868 9812
rect 3802 9800 3809 9811
rect 3461 9770 3809 9800
rect 3461 9759 3468 9770
rect 3402 9758 3468 9759
rect 3802 9759 3809 9770
rect 3861 9800 3868 9811
rect 4202 9811 4268 9812
rect 4202 9800 4209 9811
rect 3861 9770 4209 9800
rect 3861 9759 3868 9770
rect 3802 9758 3868 9759
rect 4202 9759 4209 9770
rect 4261 9800 4268 9811
rect 4602 9811 4668 9812
rect 4602 9800 4609 9811
rect 4261 9770 4609 9800
rect 4261 9759 4268 9770
rect 4202 9758 4268 9759
rect 4602 9759 4609 9770
rect 4661 9800 4668 9811
rect 5002 9811 5068 9812
rect 5002 9800 5009 9811
rect 4661 9770 5009 9800
rect 4661 9759 4668 9770
rect 4602 9758 4668 9759
rect 5002 9759 5009 9770
rect 5061 9800 5068 9811
rect 5402 9811 5468 9812
rect 5402 9800 5409 9811
rect 5061 9770 5409 9800
rect 5061 9759 5068 9770
rect 5002 9758 5068 9759
rect 5402 9759 5409 9770
rect 5461 9800 5468 9811
rect 5802 9811 5868 9812
rect 5802 9800 5809 9811
rect 5461 9770 5809 9800
rect 5461 9759 5468 9770
rect 5402 9758 5468 9759
rect 5802 9759 5809 9770
rect 5861 9800 5868 9811
rect 6202 9811 6268 9812
rect 6202 9800 6209 9811
rect 5861 9770 6209 9800
rect 5861 9759 5868 9770
rect 5802 9758 5868 9759
rect 6202 9759 6209 9770
rect 6261 9800 6268 9811
rect 6704 9811 6770 9812
rect 6704 9800 6711 9811
rect 6261 9770 6711 9800
rect 6261 9759 6268 9770
rect 6202 9758 6268 9759
rect 6704 9759 6711 9770
rect 6763 9759 6770 9811
rect 6704 9758 6770 9759
rect 2 9741 68 9742
rect 2 9730 9 9741
rect 0 9700 9 9730
rect 2 9689 9 9700
rect 61 9730 68 9741
rect 402 9741 468 9742
rect 402 9730 409 9741
rect 61 9700 409 9730
rect 61 9689 68 9700
rect 2 9688 68 9689
rect 402 9689 409 9700
rect 461 9730 468 9741
rect 802 9741 868 9742
rect 802 9730 809 9741
rect 461 9700 809 9730
rect 461 9689 468 9700
rect 402 9688 468 9689
rect 802 9689 809 9700
rect 861 9730 868 9741
rect 1202 9741 1268 9742
rect 1202 9730 1209 9741
rect 861 9700 1209 9730
rect 861 9689 868 9700
rect 802 9688 868 9689
rect 1202 9689 1209 9700
rect 1261 9730 1268 9741
rect 1602 9741 1668 9742
rect 1602 9730 1609 9741
rect 1261 9700 1609 9730
rect 1261 9689 1268 9700
rect 1202 9688 1268 9689
rect 1602 9689 1609 9700
rect 1661 9730 1668 9741
rect 2002 9741 2068 9742
rect 2002 9730 2009 9741
rect 1661 9700 2009 9730
rect 1661 9689 1668 9700
rect 1602 9688 1668 9689
rect 2002 9689 2009 9700
rect 2061 9730 2068 9741
rect 2402 9741 2468 9742
rect 2402 9730 2409 9741
rect 2061 9700 2409 9730
rect 2061 9689 2068 9700
rect 2002 9688 2068 9689
rect 2402 9689 2409 9700
rect 2461 9730 2468 9741
rect 2802 9741 2868 9742
rect 2802 9730 2809 9741
rect 2461 9700 2809 9730
rect 2461 9689 2468 9700
rect 2402 9688 2468 9689
rect 2802 9689 2809 9700
rect 2861 9730 2868 9741
rect 3202 9741 3268 9742
rect 3202 9730 3209 9741
rect 2861 9700 3209 9730
rect 2861 9689 2868 9700
rect 2802 9688 2868 9689
rect 3202 9689 3209 9700
rect 3261 9730 3268 9741
rect 3602 9741 3668 9742
rect 3602 9730 3609 9741
rect 3261 9700 3609 9730
rect 3261 9689 3268 9700
rect 3202 9688 3268 9689
rect 3602 9689 3609 9700
rect 3661 9730 3668 9741
rect 4002 9741 4068 9742
rect 4002 9730 4009 9741
rect 3661 9700 4009 9730
rect 3661 9689 3668 9700
rect 3602 9688 3668 9689
rect 4002 9689 4009 9700
rect 4061 9730 4068 9741
rect 4402 9741 4468 9742
rect 4402 9730 4409 9741
rect 4061 9700 4409 9730
rect 4061 9689 4068 9700
rect 4002 9688 4068 9689
rect 4402 9689 4409 9700
rect 4461 9730 4468 9741
rect 4802 9741 4868 9742
rect 4802 9730 4809 9741
rect 4461 9700 4809 9730
rect 4461 9689 4468 9700
rect 4402 9688 4468 9689
rect 4802 9689 4809 9700
rect 4861 9730 4868 9741
rect 5202 9741 5268 9742
rect 5202 9730 5209 9741
rect 4861 9700 5209 9730
rect 4861 9689 4868 9700
rect 4802 9688 4868 9689
rect 5202 9689 5209 9700
rect 5261 9730 5268 9741
rect 5602 9741 5668 9742
rect 5602 9730 5609 9741
rect 5261 9700 5609 9730
rect 5261 9689 5268 9700
rect 5202 9688 5268 9689
rect 5602 9689 5609 9700
rect 5661 9730 5668 9741
rect 6002 9741 6068 9742
rect 6002 9730 6009 9741
rect 5661 9700 6009 9730
rect 5661 9689 5668 9700
rect 5602 9688 5668 9689
rect 6002 9689 6009 9700
rect 6061 9730 6068 9741
rect 6402 9741 6468 9742
rect 6402 9730 6409 9741
rect 6061 9700 6409 9730
rect 6061 9689 6068 9700
rect 6002 9688 6068 9689
rect 6402 9689 6409 9700
rect 6461 9730 6468 9741
rect 6500 9741 6566 9742
rect 6500 9730 6507 9741
rect 6461 9700 6507 9730
rect 6461 9689 6468 9700
rect 6402 9688 6468 9689
rect 6500 9689 6507 9700
rect 6559 9689 6566 9741
rect 6500 9688 6566 9689
rect 202 9671 268 9672
rect 202 9660 209 9671
rect 0 9630 209 9660
rect 202 9619 209 9630
rect 261 9660 268 9671
rect 602 9671 668 9672
rect 602 9660 609 9671
rect 261 9630 609 9660
rect 261 9619 268 9630
rect 202 9618 268 9619
rect 602 9619 609 9630
rect 661 9660 668 9671
rect 1002 9671 1068 9672
rect 1002 9660 1009 9671
rect 661 9630 1009 9660
rect 661 9619 668 9630
rect 602 9618 668 9619
rect 1002 9619 1009 9630
rect 1061 9660 1068 9671
rect 1402 9671 1468 9672
rect 1402 9660 1409 9671
rect 1061 9630 1409 9660
rect 1061 9619 1068 9630
rect 1002 9618 1068 9619
rect 1402 9619 1409 9630
rect 1461 9660 1468 9671
rect 1802 9671 1868 9672
rect 1802 9660 1809 9671
rect 1461 9630 1809 9660
rect 1461 9619 1468 9630
rect 1402 9618 1468 9619
rect 1802 9619 1809 9630
rect 1861 9660 1868 9671
rect 2202 9671 2268 9672
rect 2202 9660 2209 9671
rect 1861 9630 2209 9660
rect 1861 9619 1868 9630
rect 1802 9618 1868 9619
rect 2202 9619 2209 9630
rect 2261 9660 2268 9671
rect 2602 9671 2668 9672
rect 2602 9660 2609 9671
rect 2261 9630 2609 9660
rect 2261 9619 2268 9630
rect 2202 9618 2268 9619
rect 2602 9619 2609 9630
rect 2661 9660 2668 9671
rect 3002 9671 3068 9672
rect 3002 9660 3009 9671
rect 2661 9630 3009 9660
rect 2661 9619 2668 9630
rect 2602 9618 2668 9619
rect 3002 9619 3009 9630
rect 3061 9660 3068 9671
rect 3402 9671 3468 9672
rect 3402 9660 3409 9671
rect 3061 9630 3409 9660
rect 3061 9619 3068 9630
rect 3002 9618 3068 9619
rect 3402 9619 3409 9630
rect 3461 9660 3468 9671
rect 3802 9671 3868 9672
rect 3802 9660 3809 9671
rect 3461 9630 3809 9660
rect 3461 9619 3468 9630
rect 3402 9618 3468 9619
rect 3802 9619 3809 9630
rect 3861 9660 3868 9671
rect 4202 9671 4268 9672
rect 4202 9660 4209 9671
rect 3861 9630 4209 9660
rect 3861 9619 3868 9630
rect 3802 9618 3868 9619
rect 4202 9619 4209 9630
rect 4261 9660 4268 9671
rect 4602 9671 4668 9672
rect 4602 9660 4609 9671
rect 4261 9630 4609 9660
rect 4261 9619 4268 9630
rect 4202 9618 4268 9619
rect 4602 9619 4609 9630
rect 4661 9660 4668 9671
rect 5002 9671 5068 9672
rect 5002 9660 5009 9671
rect 4661 9630 5009 9660
rect 4661 9619 4668 9630
rect 4602 9618 4668 9619
rect 5002 9619 5009 9630
rect 5061 9660 5068 9671
rect 5402 9671 5468 9672
rect 5402 9660 5409 9671
rect 5061 9630 5409 9660
rect 5061 9619 5068 9630
rect 5002 9618 5068 9619
rect 5402 9619 5409 9630
rect 5461 9660 5468 9671
rect 5802 9671 5868 9672
rect 5802 9660 5809 9671
rect 5461 9630 5809 9660
rect 5461 9619 5468 9630
rect 5402 9618 5468 9619
rect 5802 9619 5809 9630
rect 5861 9660 5868 9671
rect 6202 9671 6268 9672
rect 6202 9660 6209 9671
rect 5861 9630 6209 9660
rect 5861 9619 5868 9630
rect 5802 9618 5868 9619
rect 6202 9619 6209 9630
rect 6261 9660 6268 9671
rect 6704 9671 6770 9672
rect 6704 9660 6711 9671
rect 6261 9630 6711 9660
rect 6261 9619 6268 9630
rect 6202 9618 6268 9619
rect 6704 9619 6711 9630
rect 6763 9619 6770 9671
rect 6704 9618 6770 9619
rect 2 9601 68 9602
rect 2 9590 9 9601
rect 0 9560 9 9590
rect 2 9549 9 9560
rect 61 9590 68 9601
rect 402 9601 468 9602
rect 402 9590 409 9601
rect 61 9560 409 9590
rect 61 9549 68 9560
rect 2 9548 68 9549
rect 402 9549 409 9560
rect 461 9590 468 9601
rect 802 9601 868 9602
rect 802 9590 809 9601
rect 461 9560 809 9590
rect 461 9549 468 9560
rect 402 9548 468 9549
rect 802 9549 809 9560
rect 861 9590 868 9601
rect 1202 9601 1268 9602
rect 1202 9590 1209 9601
rect 861 9560 1209 9590
rect 861 9549 868 9560
rect 802 9548 868 9549
rect 1202 9549 1209 9560
rect 1261 9590 1268 9601
rect 1602 9601 1668 9602
rect 1602 9590 1609 9601
rect 1261 9560 1609 9590
rect 1261 9549 1268 9560
rect 1202 9548 1268 9549
rect 1602 9549 1609 9560
rect 1661 9590 1668 9601
rect 2002 9601 2068 9602
rect 2002 9590 2009 9601
rect 1661 9560 2009 9590
rect 1661 9549 1668 9560
rect 1602 9548 1668 9549
rect 2002 9549 2009 9560
rect 2061 9590 2068 9601
rect 2402 9601 2468 9602
rect 2402 9590 2409 9601
rect 2061 9560 2409 9590
rect 2061 9549 2068 9560
rect 2002 9548 2068 9549
rect 2402 9549 2409 9560
rect 2461 9590 2468 9601
rect 2802 9601 2868 9602
rect 2802 9590 2809 9601
rect 2461 9560 2809 9590
rect 2461 9549 2468 9560
rect 2402 9548 2468 9549
rect 2802 9549 2809 9560
rect 2861 9590 2868 9601
rect 3202 9601 3268 9602
rect 3202 9590 3209 9601
rect 2861 9560 3209 9590
rect 2861 9549 2868 9560
rect 2802 9548 2868 9549
rect 3202 9549 3209 9560
rect 3261 9590 3268 9601
rect 3602 9601 3668 9602
rect 3602 9590 3609 9601
rect 3261 9560 3609 9590
rect 3261 9549 3268 9560
rect 3202 9548 3268 9549
rect 3602 9549 3609 9560
rect 3661 9590 3668 9601
rect 4002 9601 4068 9602
rect 4002 9590 4009 9601
rect 3661 9560 4009 9590
rect 3661 9549 3668 9560
rect 3602 9548 3668 9549
rect 4002 9549 4009 9560
rect 4061 9590 4068 9601
rect 4402 9601 4468 9602
rect 4402 9590 4409 9601
rect 4061 9560 4409 9590
rect 4061 9549 4068 9560
rect 4002 9548 4068 9549
rect 4402 9549 4409 9560
rect 4461 9590 4468 9601
rect 4802 9601 4868 9602
rect 4802 9590 4809 9601
rect 4461 9560 4809 9590
rect 4461 9549 4468 9560
rect 4402 9548 4468 9549
rect 4802 9549 4809 9560
rect 4861 9590 4868 9601
rect 5202 9601 5268 9602
rect 5202 9590 5209 9601
rect 4861 9560 5209 9590
rect 4861 9549 4868 9560
rect 4802 9548 4868 9549
rect 5202 9549 5209 9560
rect 5261 9590 5268 9601
rect 5602 9601 5668 9602
rect 5602 9590 5609 9601
rect 5261 9560 5609 9590
rect 5261 9549 5268 9560
rect 5202 9548 5268 9549
rect 5602 9549 5609 9560
rect 5661 9590 5668 9601
rect 6002 9601 6068 9602
rect 6002 9590 6009 9601
rect 5661 9560 6009 9590
rect 5661 9549 5668 9560
rect 5602 9548 5668 9549
rect 6002 9549 6009 9560
rect 6061 9590 6068 9601
rect 6402 9601 6468 9602
rect 6402 9590 6409 9601
rect 6061 9560 6409 9590
rect 6061 9549 6068 9560
rect 6002 9548 6068 9549
rect 6402 9549 6409 9560
rect 6461 9590 6468 9601
rect 6500 9601 6566 9602
rect 6500 9590 6507 9601
rect 6461 9560 6507 9590
rect 6461 9549 6468 9560
rect 6402 9548 6468 9549
rect 6500 9549 6507 9560
rect 6559 9549 6566 9601
rect 6500 9548 6566 9549
rect 202 9531 268 9532
rect 202 9520 209 9531
rect 0 9490 209 9520
rect 202 9479 209 9490
rect 261 9520 268 9531
rect 602 9531 668 9532
rect 602 9520 609 9531
rect 261 9490 609 9520
rect 261 9479 268 9490
rect 202 9478 268 9479
rect 602 9479 609 9490
rect 661 9520 668 9531
rect 1002 9531 1068 9532
rect 1002 9520 1009 9531
rect 661 9490 1009 9520
rect 661 9479 668 9490
rect 602 9478 668 9479
rect 1002 9479 1009 9490
rect 1061 9520 1068 9531
rect 1402 9531 1468 9532
rect 1402 9520 1409 9531
rect 1061 9490 1409 9520
rect 1061 9479 1068 9490
rect 1002 9478 1068 9479
rect 1402 9479 1409 9490
rect 1461 9520 1468 9531
rect 1802 9531 1868 9532
rect 1802 9520 1809 9531
rect 1461 9490 1809 9520
rect 1461 9479 1468 9490
rect 1402 9478 1468 9479
rect 1802 9479 1809 9490
rect 1861 9520 1868 9531
rect 2202 9531 2268 9532
rect 2202 9520 2209 9531
rect 1861 9490 2209 9520
rect 1861 9479 1868 9490
rect 1802 9478 1868 9479
rect 2202 9479 2209 9490
rect 2261 9520 2268 9531
rect 2602 9531 2668 9532
rect 2602 9520 2609 9531
rect 2261 9490 2609 9520
rect 2261 9479 2268 9490
rect 2202 9478 2268 9479
rect 2602 9479 2609 9490
rect 2661 9520 2668 9531
rect 3002 9531 3068 9532
rect 3002 9520 3009 9531
rect 2661 9490 3009 9520
rect 2661 9479 2668 9490
rect 2602 9478 2668 9479
rect 3002 9479 3009 9490
rect 3061 9520 3068 9531
rect 3402 9531 3468 9532
rect 3402 9520 3409 9531
rect 3061 9490 3409 9520
rect 3061 9479 3068 9490
rect 3002 9478 3068 9479
rect 3402 9479 3409 9490
rect 3461 9520 3468 9531
rect 3802 9531 3868 9532
rect 3802 9520 3809 9531
rect 3461 9490 3809 9520
rect 3461 9479 3468 9490
rect 3402 9478 3468 9479
rect 3802 9479 3809 9490
rect 3861 9520 3868 9531
rect 4202 9531 4268 9532
rect 4202 9520 4209 9531
rect 3861 9490 4209 9520
rect 3861 9479 3868 9490
rect 3802 9478 3868 9479
rect 4202 9479 4209 9490
rect 4261 9520 4268 9531
rect 4602 9531 4668 9532
rect 4602 9520 4609 9531
rect 4261 9490 4609 9520
rect 4261 9479 4268 9490
rect 4202 9478 4268 9479
rect 4602 9479 4609 9490
rect 4661 9520 4668 9531
rect 5002 9531 5068 9532
rect 5002 9520 5009 9531
rect 4661 9490 5009 9520
rect 4661 9479 4668 9490
rect 4602 9478 4668 9479
rect 5002 9479 5009 9490
rect 5061 9520 5068 9531
rect 5402 9531 5468 9532
rect 5402 9520 5409 9531
rect 5061 9490 5409 9520
rect 5061 9479 5068 9490
rect 5002 9478 5068 9479
rect 5402 9479 5409 9490
rect 5461 9520 5468 9531
rect 5802 9531 5868 9532
rect 5802 9520 5809 9531
rect 5461 9490 5809 9520
rect 5461 9479 5468 9490
rect 5402 9478 5468 9479
rect 5802 9479 5809 9490
rect 5861 9520 5868 9531
rect 6202 9531 6268 9532
rect 6202 9520 6209 9531
rect 5861 9490 6209 9520
rect 5861 9479 5868 9490
rect 5802 9478 5868 9479
rect 6202 9479 6209 9490
rect 6261 9520 6268 9531
rect 6704 9531 6770 9532
rect 6704 9520 6711 9531
rect 6261 9490 6711 9520
rect 6261 9479 6268 9490
rect 6202 9478 6268 9479
rect 6704 9479 6711 9490
rect 6763 9479 6770 9531
rect 6704 9478 6770 9479
rect 2 9461 68 9462
rect 2 9450 9 9461
rect 0 9420 9 9450
rect 2 9409 9 9420
rect 61 9450 68 9461
rect 402 9461 468 9462
rect 402 9450 409 9461
rect 61 9420 409 9450
rect 61 9409 68 9420
rect 2 9408 68 9409
rect 402 9409 409 9420
rect 461 9450 468 9461
rect 802 9461 868 9462
rect 802 9450 809 9461
rect 461 9420 809 9450
rect 461 9409 468 9420
rect 402 9408 468 9409
rect 802 9409 809 9420
rect 861 9450 868 9461
rect 1202 9461 1268 9462
rect 1202 9450 1209 9461
rect 861 9420 1209 9450
rect 861 9409 868 9420
rect 802 9408 868 9409
rect 1202 9409 1209 9420
rect 1261 9450 1268 9461
rect 1602 9461 1668 9462
rect 1602 9450 1609 9461
rect 1261 9420 1609 9450
rect 1261 9409 1268 9420
rect 1202 9408 1268 9409
rect 1602 9409 1609 9420
rect 1661 9450 1668 9461
rect 2002 9461 2068 9462
rect 2002 9450 2009 9461
rect 1661 9420 2009 9450
rect 1661 9409 1668 9420
rect 1602 9408 1668 9409
rect 2002 9409 2009 9420
rect 2061 9450 2068 9461
rect 2402 9461 2468 9462
rect 2402 9450 2409 9461
rect 2061 9420 2409 9450
rect 2061 9409 2068 9420
rect 2002 9408 2068 9409
rect 2402 9409 2409 9420
rect 2461 9450 2468 9461
rect 2802 9461 2868 9462
rect 2802 9450 2809 9461
rect 2461 9420 2809 9450
rect 2461 9409 2468 9420
rect 2402 9408 2468 9409
rect 2802 9409 2809 9420
rect 2861 9450 2868 9461
rect 3202 9461 3268 9462
rect 3202 9450 3209 9461
rect 2861 9420 3209 9450
rect 2861 9409 2868 9420
rect 2802 9408 2868 9409
rect 3202 9409 3209 9420
rect 3261 9450 3268 9461
rect 3602 9461 3668 9462
rect 3602 9450 3609 9461
rect 3261 9420 3609 9450
rect 3261 9409 3268 9420
rect 3202 9408 3268 9409
rect 3602 9409 3609 9420
rect 3661 9450 3668 9461
rect 4002 9461 4068 9462
rect 4002 9450 4009 9461
rect 3661 9420 4009 9450
rect 3661 9409 3668 9420
rect 3602 9408 3668 9409
rect 4002 9409 4009 9420
rect 4061 9450 4068 9461
rect 4402 9461 4468 9462
rect 4402 9450 4409 9461
rect 4061 9420 4409 9450
rect 4061 9409 4068 9420
rect 4002 9408 4068 9409
rect 4402 9409 4409 9420
rect 4461 9450 4468 9461
rect 4802 9461 4868 9462
rect 4802 9450 4809 9461
rect 4461 9420 4809 9450
rect 4461 9409 4468 9420
rect 4402 9408 4468 9409
rect 4802 9409 4809 9420
rect 4861 9450 4868 9461
rect 5202 9461 5268 9462
rect 5202 9450 5209 9461
rect 4861 9420 5209 9450
rect 4861 9409 4868 9420
rect 4802 9408 4868 9409
rect 5202 9409 5209 9420
rect 5261 9450 5268 9461
rect 5602 9461 5668 9462
rect 5602 9450 5609 9461
rect 5261 9420 5609 9450
rect 5261 9409 5268 9420
rect 5202 9408 5268 9409
rect 5602 9409 5609 9420
rect 5661 9450 5668 9461
rect 6002 9461 6068 9462
rect 6002 9450 6009 9461
rect 5661 9420 6009 9450
rect 5661 9409 5668 9420
rect 5602 9408 5668 9409
rect 6002 9409 6009 9420
rect 6061 9450 6068 9461
rect 6402 9461 6468 9462
rect 6402 9450 6409 9461
rect 6061 9420 6409 9450
rect 6061 9409 6068 9420
rect 6002 9408 6068 9409
rect 6402 9409 6409 9420
rect 6461 9450 6468 9461
rect 6500 9461 6566 9462
rect 6500 9450 6507 9461
rect 6461 9420 6507 9450
rect 6461 9409 6468 9420
rect 6402 9408 6468 9409
rect 6500 9409 6507 9420
rect 6559 9409 6566 9461
rect 6500 9408 6566 9409
rect 202 9391 268 9392
rect 202 9380 209 9391
rect 0 9350 209 9380
rect 202 9339 209 9350
rect 261 9380 268 9391
rect 602 9391 668 9392
rect 602 9380 609 9391
rect 261 9350 609 9380
rect 261 9339 268 9350
rect 202 9338 268 9339
rect 602 9339 609 9350
rect 661 9380 668 9391
rect 1002 9391 1068 9392
rect 1002 9380 1009 9391
rect 661 9350 1009 9380
rect 661 9339 668 9350
rect 602 9338 668 9339
rect 1002 9339 1009 9350
rect 1061 9380 1068 9391
rect 1402 9391 1468 9392
rect 1402 9380 1409 9391
rect 1061 9350 1409 9380
rect 1061 9339 1068 9350
rect 1002 9338 1068 9339
rect 1402 9339 1409 9350
rect 1461 9380 1468 9391
rect 1802 9391 1868 9392
rect 1802 9380 1809 9391
rect 1461 9350 1809 9380
rect 1461 9339 1468 9350
rect 1402 9338 1468 9339
rect 1802 9339 1809 9350
rect 1861 9380 1868 9391
rect 2202 9391 2268 9392
rect 2202 9380 2209 9391
rect 1861 9350 2209 9380
rect 1861 9339 1868 9350
rect 1802 9338 1868 9339
rect 2202 9339 2209 9350
rect 2261 9380 2268 9391
rect 2602 9391 2668 9392
rect 2602 9380 2609 9391
rect 2261 9350 2609 9380
rect 2261 9339 2268 9350
rect 2202 9338 2268 9339
rect 2602 9339 2609 9350
rect 2661 9380 2668 9391
rect 3002 9391 3068 9392
rect 3002 9380 3009 9391
rect 2661 9350 3009 9380
rect 2661 9339 2668 9350
rect 2602 9338 2668 9339
rect 3002 9339 3009 9350
rect 3061 9380 3068 9391
rect 3402 9391 3468 9392
rect 3402 9380 3409 9391
rect 3061 9350 3409 9380
rect 3061 9339 3068 9350
rect 3002 9338 3068 9339
rect 3402 9339 3409 9350
rect 3461 9380 3468 9391
rect 3802 9391 3868 9392
rect 3802 9380 3809 9391
rect 3461 9350 3809 9380
rect 3461 9339 3468 9350
rect 3402 9338 3468 9339
rect 3802 9339 3809 9350
rect 3861 9380 3868 9391
rect 4202 9391 4268 9392
rect 4202 9380 4209 9391
rect 3861 9350 4209 9380
rect 3861 9339 3868 9350
rect 3802 9338 3868 9339
rect 4202 9339 4209 9350
rect 4261 9380 4268 9391
rect 4602 9391 4668 9392
rect 4602 9380 4609 9391
rect 4261 9350 4609 9380
rect 4261 9339 4268 9350
rect 4202 9338 4268 9339
rect 4602 9339 4609 9350
rect 4661 9380 4668 9391
rect 5002 9391 5068 9392
rect 5002 9380 5009 9391
rect 4661 9350 5009 9380
rect 4661 9339 4668 9350
rect 4602 9338 4668 9339
rect 5002 9339 5009 9350
rect 5061 9380 5068 9391
rect 5402 9391 5468 9392
rect 5402 9380 5409 9391
rect 5061 9350 5409 9380
rect 5061 9339 5068 9350
rect 5002 9338 5068 9339
rect 5402 9339 5409 9350
rect 5461 9380 5468 9391
rect 5802 9391 5868 9392
rect 5802 9380 5809 9391
rect 5461 9350 5809 9380
rect 5461 9339 5468 9350
rect 5402 9338 5468 9339
rect 5802 9339 5809 9350
rect 5861 9380 5868 9391
rect 6202 9391 6268 9392
rect 6202 9380 6209 9391
rect 5861 9350 6209 9380
rect 5861 9339 5868 9350
rect 5802 9338 5868 9339
rect 6202 9339 6209 9350
rect 6261 9380 6268 9391
rect 6704 9391 6770 9392
rect 6704 9380 6711 9391
rect 6261 9350 6711 9380
rect 6261 9339 6268 9350
rect 6202 9338 6268 9339
rect 6704 9339 6711 9350
rect 6763 9339 6770 9391
rect 6704 9338 6770 9339
rect 2 9321 68 9322
rect 2 9310 9 9321
rect 0 9280 9 9310
rect 2 9269 9 9280
rect 61 9310 68 9321
rect 402 9321 468 9322
rect 402 9310 409 9321
rect 61 9280 409 9310
rect 61 9269 68 9280
rect 2 9268 68 9269
rect 402 9269 409 9280
rect 461 9310 468 9321
rect 802 9321 868 9322
rect 802 9310 809 9321
rect 461 9280 809 9310
rect 461 9269 468 9280
rect 402 9268 468 9269
rect 802 9269 809 9280
rect 861 9310 868 9321
rect 1202 9321 1268 9322
rect 1202 9310 1209 9321
rect 861 9280 1209 9310
rect 861 9269 868 9280
rect 802 9268 868 9269
rect 1202 9269 1209 9280
rect 1261 9310 1268 9321
rect 1602 9321 1668 9322
rect 1602 9310 1609 9321
rect 1261 9280 1609 9310
rect 1261 9269 1268 9280
rect 1202 9268 1268 9269
rect 1602 9269 1609 9280
rect 1661 9310 1668 9321
rect 2002 9321 2068 9322
rect 2002 9310 2009 9321
rect 1661 9280 2009 9310
rect 1661 9269 1668 9280
rect 1602 9268 1668 9269
rect 2002 9269 2009 9280
rect 2061 9310 2068 9321
rect 2402 9321 2468 9322
rect 2402 9310 2409 9321
rect 2061 9280 2409 9310
rect 2061 9269 2068 9280
rect 2002 9268 2068 9269
rect 2402 9269 2409 9280
rect 2461 9310 2468 9321
rect 2802 9321 2868 9322
rect 2802 9310 2809 9321
rect 2461 9280 2809 9310
rect 2461 9269 2468 9280
rect 2402 9268 2468 9269
rect 2802 9269 2809 9280
rect 2861 9310 2868 9321
rect 3202 9321 3268 9322
rect 3202 9310 3209 9321
rect 2861 9280 3209 9310
rect 2861 9269 2868 9280
rect 2802 9268 2868 9269
rect 3202 9269 3209 9280
rect 3261 9310 3268 9321
rect 3602 9321 3668 9322
rect 3602 9310 3609 9321
rect 3261 9280 3609 9310
rect 3261 9269 3268 9280
rect 3202 9268 3268 9269
rect 3602 9269 3609 9280
rect 3661 9310 3668 9321
rect 4002 9321 4068 9322
rect 4002 9310 4009 9321
rect 3661 9280 4009 9310
rect 3661 9269 3668 9280
rect 3602 9268 3668 9269
rect 4002 9269 4009 9280
rect 4061 9310 4068 9321
rect 4402 9321 4468 9322
rect 4402 9310 4409 9321
rect 4061 9280 4409 9310
rect 4061 9269 4068 9280
rect 4002 9268 4068 9269
rect 4402 9269 4409 9280
rect 4461 9310 4468 9321
rect 4802 9321 4868 9322
rect 4802 9310 4809 9321
rect 4461 9280 4809 9310
rect 4461 9269 4468 9280
rect 4402 9268 4468 9269
rect 4802 9269 4809 9280
rect 4861 9310 4868 9321
rect 5202 9321 5268 9322
rect 5202 9310 5209 9321
rect 4861 9280 5209 9310
rect 4861 9269 4868 9280
rect 4802 9268 4868 9269
rect 5202 9269 5209 9280
rect 5261 9310 5268 9321
rect 5602 9321 5668 9322
rect 5602 9310 5609 9321
rect 5261 9280 5609 9310
rect 5261 9269 5268 9280
rect 5202 9268 5268 9269
rect 5602 9269 5609 9280
rect 5661 9310 5668 9321
rect 6002 9321 6068 9322
rect 6002 9310 6009 9321
rect 5661 9280 6009 9310
rect 5661 9269 5668 9280
rect 5602 9268 5668 9269
rect 6002 9269 6009 9280
rect 6061 9310 6068 9321
rect 6402 9321 6468 9322
rect 6402 9310 6409 9321
rect 6061 9280 6409 9310
rect 6061 9269 6068 9280
rect 6002 9268 6068 9269
rect 6402 9269 6409 9280
rect 6461 9310 6468 9321
rect 6500 9321 6566 9322
rect 6500 9310 6507 9321
rect 6461 9280 6507 9310
rect 6461 9269 6468 9280
rect 6402 9268 6468 9269
rect 6500 9269 6507 9280
rect 6559 9269 6566 9321
rect 6500 9268 6566 9269
rect 202 9251 268 9252
rect 202 9240 209 9251
rect 0 9210 209 9240
rect 202 9199 209 9210
rect 261 9240 268 9251
rect 602 9251 668 9252
rect 602 9240 609 9251
rect 261 9210 609 9240
rect 261 9199 268 9210
rect 202 9198 268 9199
rect 602 9199 609 9210
rect 661 9240 668 9251
rect 1002 9251 1068 9252
rect 1002 9240 1009 9251
rect 661 9210 1009 9240
rect 661 9199 668 9210
rect 602 9198 668 9199
rect 1002 9199 1009 9210
rect 1061 9240 1068 9251
rect 1402 9251 1468 9252
rect 1402 9240 1409 9251
rect 1061 9210 1409 9240
rect 1061 9199 1068 9210
rect 1002 9198 1068 9199
rect 1402 9199 1409 9210
rect 1461 9240 1468 9251
rect 1802 9251 1868 9252
rect 1802 9240 1809 9251
rect 1461 9210 1809 9240
rect 1461 9199 1468 9210
rect 1402 9198 1468 9199
rect 1802 9199 1809 9210
rect 1861 9240 1868 9251
rect 2202 9251 2268 9252
rect 2202 9240 2209 9251
rect 1861 9210 2209 9240
rect 1861 9199 1868 9210
rect 1802 9198 1868 9199
rect 2202 9199 2209 9210
rect 2261 9240 2268 9251
rect 2602 9251 2668 9252
rect 2602 9240 2609 9251
rect 2261 9210 2609 9240
rect 2261 9199 2268 9210
rect 2202 9198 2268 9199
rect 2602 9199 2609 9210
rect 2661 9240 2668 9251
rect 3002 9251 3068 9252
rect 3002 9240 3009 9251
rect 2661 9210 3009 9240
rect 2661 9199 2668 9210
rect 2602 9198 2668 9199
rect 3002 9199 3009 9210
rect 3061 9240 3068 9251
rect 3402 9251 3468 9252
rect 3402 9240 3409 9251
rect 3061 9210 3409 9240
rect 3061 9199 3068 9210
rect 3002 9198 3068 9199
rect 3402 9199 3409 9210
rect 3461 9240 3468 9251
rect 3802 9251 3868 9252
rect 3802 9240 3809 9251
rect 3461 9210 3809 9240
rect 3461 9199 3468 9210
rect 3402 9198 3468 9199
rect 3802 9199 3809 9210
rect 3861 9240 3868 9251
rect 4202 9251 4268 9252
rect 4202 9240 4209 9251
rect 3861 9210 4209 9240
rect 3861 9199 3868 9210
rect 3802 9198 3868 9199
rect 4202 9199 4209 9210
rect 4261 9240 4268 9251
rect 4602 9251 4668 9252
rect 4602 9240 4609 9251
rect 4261 9210 4609 9240
rect 4261 9199 4268 9210
rect 4202 9198 4268 9199
rect 4602 9199 4609 9210
rect 4661 9240 4668 9251
rect 5002 9251 5068 9252
rect 5002 9240 5009 9251
rect 4661 9210 5009 9240
rect 4661 9199 4668 9210
rect 4602 9198 4668 9199
rect 5002 9199 5009 9210
rect 5061 9240 5068 9251
rect 5402 9251 5468 9252
rect 5402 9240 5409 9251
rect 5061 9210 5409 9240
rect 5061 9199 5068 9210
rect 5002 9198 5068 9199
rect 5402 9199 5409 9210
rect 5461 9240 5468 9251
rect 5802 9251 5868 9252
rect 5802 9240 5809 9251
rect 5461 9210 5809 9240
rect 5461 9199 5468 9210
rect 5402 9198 5468 9199
rect 5802 9199 5809 9210
rect 5861 9240 5868 9251
rect 6202 9251 6268 9252
rect 6202 9240 6209 9251
rect 5861 9210 6209 9240
rect 5861 9199 5868 9210
rect 5802 9198 5868 9199
rect 6202 9199 6209 9210
rect 6261 9240 6268 9251
rect 6704 9251 6770 9252
rect 6704 9240 6711 9251
rect 6261 9210 6711 9240
rect 6261 9199 6268 9210
rect 6202 9198 6268 9199
rect 6704 9199 6711 9210
rect 6763 9199 6770 9251
rect 6704 9198 6770 9199
rect 2 9181 68 9182
rect 2 9170 9 9181
rect 0 9140 9 9170
rect 2 9129 9 9140
rect 61 9170 68 9181
rect 402 9181 468 9182
rect 402 9170 409 9181
rect 61 9140 409 9170
rect 61 9129 68 9140
rect 2 9128 68 9129
rect 402 9129 409 9140
rect 461 9170 468 9181
rect 802 9181 868 9182
rect 802 9170 809 9181
rect 461 9140 809 9170
rect 461 9129 468 9140
rect 402 9128 468 9129
rect 802 9129 809 9140
rect 861 9170 868 9181
rect 1202 9181 1268 9182
rect 1202 9170 1209 9181
rect 861 9140 1209 9170
rect 861 9129 868 9140
rect 802 9128 868 9129
rect 1202 9129 1209 9140
rect 1261 9170 1268 9181
rect 1602 9181 1668 9182
rect 1602 9170 1609 9181
rect 1261 9140 1609 9170
rect 1261 9129 1268 9140
rect 1202 9128 1268 9129
rect 1602 9129 1609 9140
rect 1661 9170 1668 9181
rect 2002 9181 2068 9182
rect 2002 9170 2009 9181
rect 1661 9140 2009 9170
rect 1661 9129 1668 9140
rect 1602 9128 1668 9129
rect 2002 9129 2009 9140
rect 2061 9170 2068 9181
rect 2402 9181 2468 9182
rect 2402 9170 2409 9181
rect 2061 9140 2409 9170
rect 2061 9129 2068 9140
rect 2002 9128 2068 9129
rect 2402 9129 2409 9140
rect 2461 9170 2468 9181
rect 2802 9181 2868 9182
rect 2802 9170 2809 9181
rect 2461 9140 2809 9170
rect 2461 9129 2468 9140
rect 2402 9128 2468 9129
rect 2802 9129 2809 9140
rect 2861 9170 2868 9181
rect 3202 9181 3268 9182
rect 3202 9170 3209 9181
rect 2861 9140 3209 9170
rect 2861 9129 2868 9140
rect 2802 9128 2868 9129
rect 3202 9129 3209 9140
rect 3261 9170 3268 9181
rect 3602 9181 3668 9182
rect 3602 9170 3609 9181
rect 3261 9140 3609 9170
rect 3261 9129 3268 9140
rect 3202 9128 3268 9129
rect 3602 9129 3609 9140
rect 3661 9170 3668 9181
rect 4002 9181 4068 9182
rect 4002 9170 4009 9181
rect 3661 9140 4009 9170
rect 3661 9129 3668 9140
rect 3602 9128 3668 9129
rect 4002 9129 4009 9140
rect 4061 9170 4068 9181
rect 4402 9181 4468 9182
rect 4402 9170 4409 9181
rect 4061 9140 4409 9170
rect 4061 9129 4068 9140
rect 4002 9128 4068 9129
rect 4402 9129 4409 9140
rect 4461 9170 4468 9181
rect 4802 9181 4868 9182
rect 4802 9170 4809 9181
rect 4461 9140 4809 9170
rect 4461 9129 4468 9140
rect 4402 9128 4468 9129
rect 4802 9129 4809 9140
rect 4861 9170 4868 9181
rect 5202 9181 5268 9182
rect 5202 9170 5209 9181
rect 4861 9140 5209 9170
rect 4861 9129 4868 9140
rect 4802 9128 4868 9129
rect 5202 9129 5209 9140
rect 5261 9170 5268 9181
rect 5602 9181 5668 9182
rect 5602 9170 5609 9181
rect 5261 9140 5609 9170
rect 5261 9129 5268 9140
rect 5202 9128 5268 9129
rect 5602 9129 5609 9140
rect 5661 9170 5668 9181
rect 6002 9181 6068 9182
rect 6002 9170 6009 9181
rect 5661 9140 6009 9170
rect 5661 9129 5668 9140
rect 5602 9128 5668 9129
rect 6002 9129 6009 9140
rect 6061 9170 6068 9181
rect 6402 9181 6468 9182
rect 6402 9170 6409 9181
rect 6061 9140 6409 9170
rect 6061 9129 6068 9140
rect 6002 9128 6068 9129
rect 6402 9129 6409 9140
rect 6461 9170 6468 9181
rect 6500 9181 6566 9182
rect 6500 9170 6507 9181
rect 6461 9140 6507 9170
rect 6461 9129 6468 9140
rect 6402 9128 6468 9129
rect 6500 9129 6507 9140
rect 6559 9129 6566 9181
rect 6500 9128 6566 9129
rect 202 9111 268 9112
rect 202 9100 209 9111
rect 0 9070 209 9100
rect 202 9059 209 9070
rect 261 9100 268 9111
rect 602 9111 668 9112
rect 602 9100 609 9111
rect 261 9070 609 9100
rect 261 9059 268 9070
rect 202 9058 268 9059
rect 602 9059 609 9070
rect 661 9100 668 9111
rect 1002 9111 1068 9112
rect 1002 9100 1009 9111
rect 661 9070 1009 9100
rect 661 9059 668 9070
rect 602 9058 668 9059
rect 1002 9059 1009 9070
rect 1061 9100 1068 9111
rect 1402 9111 1468 9112
rect 1402 9100 1409 9111
rect 1061 9070 1409 9100
rect 1061 9059 1068 9070
rect 1002 9058 1068 9059
rect 1402 9059 1409 9070
rect 1461 9100 1468 9111
rect 1802 9111 1868 9112
rect 1802 9100 1809 9111
rect 1461 9070 1809 9100
rect 1461 9059 1468 9070
rect 1402 9058 1468 9059
rect 1802 9059 1809 9070
rect 1861 9100 1868 9111
rect 2202 9111 2268 9112
rect 2202 9100 2209 9111
rect 1861 9070 2209 9100
rect 1861 9059 1868 9070
rect 1802 9058 1868 9059
rect 2202 9059 2209 9070
rect 2261 9100 2268 9111
rect 2602 9111 2668 9112
rect 2602 9100 2609 9111
rect 2261 9070 2609 9100
rect 2261 9059 2268 9070
rect 2202 9058 2268 9059
rect 2602 9059 2609 9070
rect 2661 9100 2668 9111
rect 3002 9111 3068 9112
rect 3002 9100 3009 9111
rect 2661 9070 3009 9100
rect 2661 9059 2668 9070
rect 2602 9058 2668 9059
rect 3002 9059 3009 9070
rect 3061 9100 3068 9111
rect 3402 9111 3468 9112
rect 3402 9100 3409 9111
rect 3061 9070 3409 9100
rect 3061 9059 3068 9070
rect 3002 9058 3068 9059
rect 3402 9059 3409 9070
rect 3461 9100 3468 9111
rect 3802 9111 3868 9112
rect 3802 9100 3809 9111
rect 3461 9070 3809 9100
rect 3461 9059 3468 9070
rect 3402 9058 3468 9059
rect 3802 9059 3809 9070
rect 3861 9100 3868 9111
rect 4202 9111 4268 9112
rect 4202 9100 4209 9111
rect 3861 9070 4209 9100
rect 3861 9059 3868 9070
rect 3802 9058 3868 9059
rect 4202 9059 4209 9070
rect 4261 9100 4268 9111
rect 4602 9111 4668 9112
rect 4602 9100 4609 9111
rect 4261 9070 4609 9100
rect 4261 9059 4268 9070
rect 4202 9058 4268 9059
rect 4602 9059 4609 9070
rect 4661 9100 4668 9111
rect 5002 9111 5068 9112
rect 5002 9100 5009 9111
rect 4661 9070 5009 9100
rect 4661 9059 4668 9070
rect 4602 9058 4668 9059
rect 5002 9059 5009 9070
rect 5061 9100 5068 9111
rect 5402 9111 5468 9112
rect 5402 9100 5409 9111
rect 5061 9070 5409 9100
rect 5061 9059 5068 9070
rect 5002 9058 5068 9059
rect 5402 9059 5409 9070
rect 5461 9100 5468 9111
rect 5802 9111 5868 9112
rect 5802 9100 5809 9111
rect 5461 9070 5809 9100
rect 5461 9059 5468 9070
rect 5402 9058 5468 9059
rect 5802 9059 5809 9070
rect 5861 9100 5868 9111
rect 6202 9111 6268 9112
rect 6202 9100 6209 9111
rect 5861 9070 6209 9100
rect 5861 9059 5868 9070
rect 5802 9058 5868 9059
rect 6202 9059 6209 9070
rect 6261 9100 6268 9111
rect 6704 9111 6770 9112
rect 6704 9100 6711 9111
rect 6261 9070 6711 9100
rect 6261 9059 6268 9070
rect 6202 9058 6268 9059
rect 6704 9059 6711 9070
rect 6763 9059 6770 9111
rect 6704 9058 6770 9059
rect 2 9041 68 9042
rect 2 9030 9 9041
rect 0 9000 9 9030
rect 2 8989 9 9000
rect 61 9030 68 9041
rect 402 9041 468 9042
rect 402 9030 409 9041
rect 61 9000 409 9030
rect 61 8989 68 9000
rect 2 8988 68 8989
rect 402 8989 409 9000
rect 461 9030 468 9041
rect 802 9041 868 9042
rect 802 9030 809 9041
rect 461 9000 809 9030
rect 461 8989 468 9000
rect 402 8988 468 8989
rect 802 8989 809 9000
rect 861 9030 868 9041
rect 1202 9041 1268 9042
rect 1202 9030 1209 9041
rect 861 9000 1209 9030
rect 861 8989 868 9000
rect 802 8988 868 8989
rect 1202 8989 1209 9000
rect 1261 9030 1268 9041
rect 1602 9041 1668 9042
rect 1602 9030 1609 9041
rect 1261 9000 1609 9030
rect 1261 8989 1268 9000
rect 1202 8988 1268 8989
rect 1602 8989 1609 9000
rect 1661 9030 1668 9041
rect 2002 9041 2068 9042
rect 2002 9030 2009 9041
rect 1661 9000 2009 9030
rect 1661 8989 1668 9000
rect 1602 8988 1668 8989
rect 2002 8989 2009 9000
rect 2061 9030 2068 9041
rect 2402 9041 2468 9042
rect 2402 9030 2409 9041
rect 2061 9000 2409 9030
rect 2061 8989 2068 9000
rect 2002 8988 2068 8989
rect 2402 8989 2409 9000
rect 2461 9030 2468 9041
rect 2802 9041 2868 9042
rect 2802 9030 2809 9041
rect 2461 9000 2809 9030
rect 2461 8989 2468 9000
rect 2402 8988 2468 8989
rect 2802 8989 2809 9000
rect 2861 9030 2868 9041
rect 3202 9041 3268 9042
rect 3202 9030 3209 9041
rect 2861 9000 3209 9030
rect 2861 8989 2868 9000
rect 2802 8988 2868 8989
rect 3202 8989 3209 9000
rect 3261 9030 3268 9041
rect 3602 9041 3668 9042
rect 3602 9030 3609 9041
rect 3261 9000 3609 9030
rect 3261 8989 3268 9000
rect 3202 8988 3268 8989
rect 3602 8989 3609 9000
rect 3661 9030 3668 9041
rect 4002 9041 4068 9042
rect 4002 9030 4009 9041
rect 3661 9000 4009 9030
rect 3661 8989 3668 9000
rect 3602 8988 3668 8989
rect 4002 8989 4009 9000
rect 4061 9030 4068 9041
rect 4402 9041 4468 9042
rect 4402 9030 4409 9041
rect 4061 9000 4409 9030
rect 4061 8989 4068 9000
rect 4002 8988 4068 8989
rect 4402 8989 4409 9000
rect 4461 9030 4468 9041
rect 4802 9041 4868 9042
rect 4802 9030 4809 9041
rect 4461 9000 4809 9030
rect 4461 8989 4468 9000
rect 4402 8988 4468 8989
rect 4802 8989 4809 9000
rect 4861 9030 4868 9041
rect 5202 9041 5268 9042
rect 5202 9030 5209 9041
rect 4861 9000 5209 9030
rect 4861 8989 4868 9000
rect 4802 8988 4868 8989
rect 5202 8989 5209 9000
rect 5261 9030 5268 9041
rect 5602 9041 5668 9042
rect 5602 9030 5609 9041
rect 5261 9000 5609 9030
rect 5261 8989 5268 9000
rect 5202 8988 5268 8989
rect 5602 8989 5609 9000
rect 5661 9030 5668 9041
rect 6002 9041 6068 9042
rect 6002 9030 6009 9041
rect 5661 9000 6009 9030
rect 5661 8989 5668 9000
rect 5602 8988 5668 8989
rect 6002 8989 6009 9000
rect 6061 9030 6068 9041
rect 6402 9041 6468 9042
rect 6402 9030 6409 9041
rect 6061 9000 6409 9030
rect 6061 8989 6068 9000
rect 6002 8988 6068 8989
rect 6402 8989 6409 9000
rect 6461 9030 6468 9041
rect 6500 9041 6566 9042
rect 6500 9030 6507 9041
rect 6461 9000 6507 9030
rect 6461 8989 6468 9000
rect 6402 8988 6468 8989
rect 6500 8989 6507 9000
rect 6559 8989 6566 9041
rect 6500 8988 6566 8989
rect 202 8971 268 8972
rect 202 8960 209 8971
rect 0 8930 209 8960
rect 202 8919 209 8930
rect 261 8960 268 8971
rect 602 8971 668 8972
rect 602 8960 609 8971
rect 261 8930 609 8960
rect 261 8919 268 8930
rect 202 8918 268 8919
rect 602 8919 609 8930
rect 661 8960 668 8971
rect 1002 8971 1068 8972
rect 1002 8960 1009 8971
rect 661 8930 1009 8960
rect 661 8919 668 8930
rect 602 8918 668 8919
rect 1002 8919 1009 8930
rect 1061 8960 1068 8971
rect 1402 8971 1468 8972
rect 1402 8960 1409 8971
rect 1061 8930 1409 8960
rect 1061 8919 1068 8930
rect 1002 8918 1068 8919
rect 1402 8919 1409 8930
rect 1461 8960 1468 8971
rect 1802 8971 1868 8972
rect 1802 8960 1809 8971
rect 1461 8930 1809 8960
rect 1461 8919 1468 8930
rect 1402 8918 1468 8919
rect 1802 8919 1809 8930
rect 1861 8960 1868 8971
rect 2202 8971 2268 8972
rect 2202 8960 2209 8971
rect 1861 8930 2209 8960
rect 1861 8919 1868 8930
rect 1802 8918 1868 8919
rect 2202 8919 2209 8930
rect 2261 8960 2268 8971
rect 2602 8971 2668 8972
rect 2602 8960 2609 8971
rect 2261 8930 2609 8960
rect 2261 8919 2268 8930
rect 2202 8918 2268 8919
rect 2602 8919 2609 8930
rect 2661 8960 2668 8971
rect 3002 8971 3068 8972
rect 3002 8960 3009 8971
rect 2661 8930 3009 8960
rect 2661 8919 2668 8930
rect 2602 8918 2668 8919
rect 3002 8919 3009 8930
rect 3061 8960 3068 8971
rect 3402 8971 3468 8972
rect 3402 8960 3409 8971
rect 3061 8930 3409 8960
rect 3061 8919 3068 8930
rect 3002 8918 3068 8919
rect 3402 8919 3409 8930
rect 3461 8960 3468 8971
rect 3802 8971 3868 8972
rect 3802 8960 3809 8971
rect 3461 8930 3809 8960
rect 3461 8919 3468 8930
rect 3402 8918 3468 8919
rect 3802 8919 3809 8930
rect 3861 8960 3868 8971
rect 4202 8971 4268 8972
rect 4202 8960 4209 8971
rect 3861 8930 4209 8960
rect 3861 8919 3868 8930
rect 3802 8918 3868 8919
rect 4202 8919 4209 8930
rect 4261 8960 4268 8971
rect 4602 8971 4668 8972
rect 4602 8960 4609 8971
rect 4261 8930 4609 8960
rect 4261 8919 4268 8930
rect 4202 8918 4268 8919
rect 4602 8919 4609 8930
rect 4661 8960 4668 8971
rect 5002 8971 5068 8972
rect 5002 8960 5009 8971
rect 4661 8930 5009 8960
rect 4661 8919 4668 8930
rect 4602 8918 4668 8919
rect 5002 8919 5009 8930
rect 5061 8960 5068 8971
rect 5402 8971 5468 8972
rect 5402 8960 5409 8971
rect 5061 8930 5409 8960
rect 5061 8919 5068 8930
rect 5002 8918 5068 8919
rect 5402 8919 5409 8930
rect 5461 8960 5468 8971
rect 5802 8971 5868 8972
rect 5802 8960 5809 8971
rect 5461 8930 5809 8960
rect 5461 8919 5468 8930
rect 5402 8918 5468 8919
rect 5802 8919 5809 8930
rect 5861 8960 5868 8971
rect 6202 8971 6268 8972
rect 6202 8960 6209 8971
rect 5861 8930 6209 8960
rect 5861 8919 5868 8930
rect 5802 8918 5868 8919
rect 6202 8919 6209 8930
rect 6261 8960 6268 8971
rect 6704 8971 6770 8972
rect 6704 8960 6711 8971
rect 6261 8930 6711 8960
rect 6261 8919 6268 8930
rect 6202 8918 6268 8919
rect 6704 8919 6711 8930
rect 6763 8919 6770 8971
rect 6704 8918 6770 8919
rect 2 8901 68 8902
rect 2 8890 9 8901
rect 0 8860 9 8890
rect 2 8849 9 8860
rect 61 8890 68 8901
rect 402 8901 468 8902
rect 402 8890 409 8901
rect 61 8860 409 8890
rect 61 8849 68 8860
rect 2 8848 68 8849
rect 402 8849 409 8860
rect 461 8890 468 8901
rect 802 8901 868 8902
rect 802 8890 809 8901
rect 461 8860 809 8890
rect 461 8849 468 8860
rect 402 8848 468 8849
rect 802 8849 809 8860
rect 861 8890 868 8901
rect 1202 8901 1268 8902
rect 1202 8890 1209 8901
rect 861 8860 1209 8890
rect 861 8849 868 8860
rect 802 8848 868 8849
rect 1202 8849 1209 8860
rect 1261 8890 1268 8901
rect 1602 8901 1668 8902
rect 1602 8890 1609 8901
rect 1261 8860 1609 8890
rect 1261 8849 1268 8860
rect 1202 8848 1268 8849
rect 1602 8849 1609 8860
rect 1661 8890 1668 8901
rect 2002 8901 2068 8902
rect 2002 8890 2009 8901
rect 1661 8860 2009 8890
rect 1661 8849 1668 8860
rect 1602 8848 1668 8849
rect 2002 8849 2009 8860
rect 2061 8890 2068 8901
rect 2402 8901 2468 8902
rect 2402 8890 2409 8901
rect 2061 8860 2409 8890
rect 2061 8849 2068 8860
rect 2002 8848 2068 8849
rect 2402 8849 2409 8860
rect 2461 8890 2468 8901
rect 2802 8901 2868 8902
rect 2802 8890 2809 8901
rect 2461 8860 2809 8890
rect 2461 8849 2468 8860
rect 2402 8848 2468 8849
rect 2802 8849 2809 8860
rect 2861 8890 2868 8901
rect 3202 8901 3268 8902
rect 3202 8890 3209 8901
rect 2861 8860 3209 8890
rect 2861 8849 2868 8860
rect 2802 8848 2868 8849
rect 3202 8849 3209 8860
rect 3261 8890 3268 8901
rect 3602 8901 3668 8902
rect 3602 8890 3609 8901
rect 3261 8860 3609 8890
rect 3261 8849 3268 8860
rect 3202 8848 3268 8849
rect 3602 8849 3609 8860
rect 3661 8890 3668 8901
rect 4002 8901 4068 8902
rect 4002 8890 4009 8901
rect 3661 8860 4009 8890
rect 3661 8849 3668 8860
rect 3602 8848 3668 8849
rect 4002 8849 4009 8860
rect 4061 8890 4068 8901
rect 4402 8901 4468 8902
rect 4402 8890 4409 8901
rect 4061 8860 4409 8890
rect 4061 8849 4068 8860
rect 4002 8848 4068 8849
rect 4402 8849 4409 8860
rect 4461 8890 4468 8901
rect 4802 8901 4868 8902
rect 4802 8890 4809 8901
rect 4461 8860 4809 8890
rect 4461 8849 4468 8860
rect 4402 8848 4468 8849
rect 4802 8849 4809 8860
rect 4861 8890 4868 8901
rect 5202 8901 5268 8902
rect 5202 8890 5209 8901
rect 4861 8860 5209 8890
rect 4861 8849 4868 8860
rect 4802 8848 4868 8849
rect 5202 8849 5209 8860
rect 5261 8890 5268 8901
rect 5602 8901 5668 8902
rect 5602 8890 5609 8901
rect 5261 8860 5609 8890
rect 5261 8849 5268 8860
rect 5202 8848 5268 8849
rect 5602 8849 5609 8860
rect 5661 8890 5668 8901
rect 6002 8901 6068 8902
rect 6002 8890 6009 8901
rect 5661 8860 6009 8890
rect 5661 8849 5668 8860
rect 5602 8848 5668 8849
rect 6002 8849 6009 8860
rect 6061 8890 6068 8901
rect 6402 8901 6468 8902
rect 6402 8890 6409 8901
rect 6061 8860 6409 8890
rect 6061 8849 6068 8860
rect 6002 8848 6068 8849
rect 6402 8849 6409 8860
rect 6461 8890 6468 8901
rect 6500 8901 6566 8902
rect 6500 8890 6507 8901
rect 6461 8860 6507 8890
rect 6461 8849 6468 8860
rect 6402 8848 6468 8849
rect 6500 8849 6507 8860
rect 6559 8849 6566 8901
rect 6500 8848 6566 8849
rect 202 8831 268 8832
rect 202 8820 209 8831
rect 0 8790 209 8820
rect 202 8779 209 8790
rect 261 8820 268 8831
rect 602 8831 668 8832
rect 602 8820 609 8831
rect 261 8790 609 8820
rect 261 8779 268 8790
rect 202 8778 268 8779
rect 602 8779 609 8790
rect 661 8820 668 8831
rect 1002 8831 1068 8832
rect 1002 8820 1009 8831
rect 661 8790 1009 8820
rect 661 8779 668 8790
rect 602 8778 668 8779
rect 1002 8779 1009 8790
rect 1061 8820 1068 8831
rect 1402 8831 1468 8832
rect 1402 8820 1409 8831
rect 1061 8790 1409 8820
rect 1061 8779 1068 8790
rect 1002 8778 1068 8779
rect 1402 8779 1409 8790
rect 1461 8820 1468 8831
rect 1802 8831 1868 8832
rect 1802 8820 1809 8831
rect 1461 8790 1809 8820
rect 1461 8779 1468 8790
rect 1402 8778 1468 8779
rect 1802 8779 1809 8790
rect 1861 8820 1868 8831
rect 2202 8831 2268 8832
rect 2202 8820 2209 8831
rect 1861 8790 2209 8820
rect 1861 8779 1868 8790
rect 1802 8778 1868 8779
rect 2202 8779 2209 8790
rect 2261 8820 2268 8831
rect 2602 8831 2668 8832
rect 2602 8820 2609 8831
rect 2261 8790 2609 8820
rect 2261 8779 2268 8790
rect 2202 8778 2268 8779
rect 2602 8779 2609 8790
rect 2661 8820 2668 8831
rect 3002 8831 3068 8832
rect 3002 8820 3009 8831
rect 2661 8790 3009 8820
rect 2661 8779 2668 8790
rect 2602 8778 2668 8779
rect 3002 8779 3009 8790
rect 3061 8820 3068 8831
rect 3402 8831 3468 8832
rect 3402 8820 3409 8831
rect 3061 8790 3409 8820
rect 3061 8779 3068 8790
rect 3002 8778 3068 8779
rect 3402 8779 3409 8790
rect 3461 8820 3468 8831
rect 3802 8831 3868 8832
rect 3802 8820 3809 8831
rect 3461 8790 3809 8820
rect 3461 8779 3468 8790
rect 3402 8778 3468 8779
rect 3802 8779 3809 8790
rect 3861 8820 3868 8831
rect 4202 8831 4268 8832
rect 4202 8820 4209 8831
rect 3861 8790 4209 8820
rect 3861 8779 3868 8790
rect 3802 8778 3868 8779
rect 4202 8779 4209 8790
rect 4261 8820 4268 8831
rect 4602 8831 4668 8832
rect 4602 8820 4609 8831
rect 4261 8790 4609 8820
rect 4261 8779 4268 8790
rect 4202 8778 4268 8779
rect 4602 8779 4609 8790
rect 4661 8820 4668 8831
rect 5002 8831 5068 8832
rect 5002 8820 5009 8831
rect 4661 8790 5009 8820
rect 4661 8779 4668 8790
rect 4602 8778 4668 8779
rect 5002 8779 5009 8790
rect 5061 8820 5068 8831
rect 5402 8831 5468 8832
rect 5402 8820 5409 8831
rect 5061 8790 5409 8820
rect 5061 8779 5068 8790
rect 5002 8778 5068 8779
rect 5402 8779 5409 8790
rect 5461 8820 5468 8831
rect 5802 8831 5868 8832
rect 5802 8820 5809 8831
rect 5461 8790 5809 8820
rect 5461 8779 5468 8790
rect 5402 8778 5468 8779
rect 5802 8779 5809 8790
rect 5861 8820 5868 8831
rect 6202 8831 6268 8832
rect 6202 8820 6209 8831
rect 5861 8790 6209 8820
rect 5861 8779 5868 8790
rect 5802 8778 5868 8779
rect 6202 8779 6209 8790
rect 6261 8820 6268 8831
rect 6704 8831 6770 8832
rect 6704 8820 6711 8831
rect 6261 8790 6711 8820
rect 6261 8779 6268 8790
rect 6202 8778 6268 8779
rect 6704 8779 6711 8790
rect 6763 8779 6770 8831
rect 6704 8778 6770 8779
rect 2 8761 68 8762
rect 2 8750 9 8761
rect 0 8720 9 8750
rect 2 8709 9 8720
rect 61 8750 68 8761
rect 402 8761 468 8762
rect 402 8750 409 8761
rect 61 8720 409 8750
rect 61 8709 68 8720
rect 2 8708 68 8709
rect 402 8709 409 8720
rect 461 8750 468 8761
rect 802 8761 868 8762
rect 802 8750 809 8761
rect 461 8720 809 8750
rect 461 8709 468 8720
rect 402 8708 468 8709
rect 802 8709 809 8720
rect 861 8750 868 8761
rect 1202 8761 1268 8762
rect 1202 8750 1209 8761
rect 861 8720 1209 8750
rect 861 8709 868 8720
rect 802 8708 868 8709
rect 1202 8709 1209 8720
rect 1261 8750 1268 8761
rect 1602 8761 1668 8762
rect 1602 8750 1609 8761
rect 1261 8720 1609 8750
rect 1261 8709 1268 8720
rect 1202 8708 1268 8709
rect 1602 8709 1609 8720
rect 1661 8750 1668 8761
rect 2002 8761 2068 8762
rect 2002 8750 2009 8761
rect 1661 8720 2009 8750
rect 1661 8709 1668 8720
rect 1602 8708 1668 8709
rect 2002 8709 2009 8720
rect 2061 8750 2068 8761
rect 2402 8761 2468 8762
rect 2402 8750 2409 8761
rect 2061 8720 2409 8750
rect 2061 8709 2068 8720
rect 2002 8708 2068 8709
rect 2402 8709 2409 8720
rect 2461 8750 2468 8761
rect 2802 8761 2868 8762
rect 2802 8750 2809 8761
rect 2461 8720 2809 8750
rect 2461 8709 2468 8720
rect 2402 8708 2468 8709
rect 2802 8709 2809 8720
rect 2861 8750 2868 8761
rect 3202 8761 3268 8762
rect 3202 8750 3209 8761
rect 2861 8720 3209 8750
rect 2861 8709 2868 8720
rect 2802 8708 2868 8709
rect 3202 8709 3209 8720
rect 3261 8750 3268 8761
rect 3602 8761 3668 8762
rect 3602 8750 3609 8761
rect 3261 8720 3609 8750
rect 3261 8709 3268 8720
rect 3202 8708 3268 8709
rect 3602 8709 3609 8720
rect 3661 8750 3668 8761
rect 4002 8761 4068 8762
rect 4002 8750 4009 8761
rect 3661 8720 4009 8750
rect 3661 8709 3668 8720
rect 3602 8708 3668 8709
rect 4002 8709 4009 8720
rect 4061 8750 4068 8761
rect 4402 8761 4468 8762
rect 4402 8750 4409 8761
rect 4061 8720 4409 8750
rect 4061 8709 4068 8720
rect 4002 8708 4068 8709
rect 4402 8709 4409 8720
rect 4461 8750 4468 8761
rect 4802 8761 4868 8762
rect 4802 8750 4809 8761
rect 4461 8720 4809 8750
rect 4461 8709 4468 8720
rect 4402 8708 4468 8709
rect 4802 8709 4809 8720
rect 4861 8750 4868 8761
rect 5202 8761 5268 8762
rect 5202 8750 5209 8761
rect 4861 8720 5209 8750
rect 4861 8709 4868 8720
rect 4802 8708 4868 8709
rect 5202 8709 5209 8720
rect 5261 8750 5268 8761
rect 5602 8761 5668 8762
rect 5602 8750 5609 8761
rect 5261 8720 5609 8750
rect 5261 8709 5268 8720
rect 5202 8708 5268 8709
rect 5602 8709 5609 8720
rect 5661 8750 5668 8761
rect 6002 8761 6068 8762
rect 6002 8750 6009 8761
rect 5661 8720 6009 8750
rect 5661 8709 5668 8720
rect 5602 8708 5668 8709
rect 6002 8709 6009 8720
rect 6061 8750 6068 8761
rect 6402 8761 6468 8762
rect 6402 8750 6409 8761
rect 6061 8720 6409 8750
rect 6061 8709 6068 8720
rect 6002 8708 6068 8709
rect 6402 8709 6409 8720
rect 6461 8750 6468 8761
rect 6500 8761 6566 8762
rect 6500 8750 6507 8761
rect 6461 8720 6507 8750
rect 6461 8709 6468 8720
rect 6402 8708 6468 8709
rect 6500 8709 6507 8720
rect 6559 8709 6566 8761
rect 6500 8708 6566 8709
rect 196 8691 274 8692
rect -4 8675 74 8676
rect -4 8619 7 8675
rect 63 8619 74 8675
rect 196 8635 207 8691
rect 263 8635 274 8691
rect 596 8691 674 8692
rect 196 8634 274 8635
rect 396 8675 474 8676
rect -4 8618 74 8619
rect 396 8619 407 8675
rect 463 8619 474 8675
rect 596 8635 607 8691
rect 663 8635 674 8691
rect 996 8691 1074 8692
rect 596 8634 674 8635
rect 796 8675 874 8676
rect 396 8618 474 8619
rect 796 8619 807 8675
rect 863 8619 874 8675
rect 996 8635 1007 8691
rect 1063 8635 1074 8691
rect 1396 8691 1474 8692
rect 996 8634 1074 8635
rect 1196 8675 1274 8676
rect 796 8618 874 8619
rect 1196 8619 1207 8675
rect 1263 8619 1274 8675
rect 1396 8635 1407 8691
rect 1463 8635 1474 8691
rect 1796 8691 1874 8692
rect 1396 8634 1474 8635
rect 1596 8675 1674 8676
rect 1196 8618 1274 8619
rect 1596 8619 1607 8675
rect 1663 8619 1674 8675
rect 1796 8635 1807 8691
rect 1863 8635 1874 8691
rect 2196 8691 2274 8692
rect 1796 8634 1874 8635
rect 1996 8675 2074 8676
rect 1596 8618 1674 8619
rect 1996 8619 2007 8675
rect 2063 8619 2074 8675
rect 2196 8635 2207 8691
rect 2263 8635 2274 8691
rect 2596 8691 2674 8692
rect 2196 8634 2274 8635
rect 2396 8675 2474 8676
rect 1996 8618 2074 8619
rect 2396 8619 2407 8675
rect 2463 8619 2474 8675
rect 2596 8635 2607 8691
rect 2663 8635 2674 8691
rect 2996 8691 3074 8692
rect 2596 8634 2674 8635
rect 2796 8675 2874 8676
rect 2396 8618 2474 8619
rect 2796 8619 2807 8675
rect 2863 8619 2874 8675
rect 2996 8635 3007 8691
rect 3063 8635 3074 8691
rect 3396 8691 3474 8692
rect 2996 8634 3074 8635
rect 3196 8675 3274 8676
rect 2796 8618 2874 8619
rect 3196 8619 3207 8675
rect 3263 8619 3274 8675
rect 3396 8635 3407 8691
rect 3463 8635 3474 8691
rect 3796 8691 3874 8692
rect 3396 8634 3474 8635
rect 3596 8675 3674 8676
rect 3196 8618 3274 8619
rect 3596 8619 3607 8675
rect 3663 8619 3674 8675
rect 3796 8635 3807 8691
rect 3863 8635 3874 8691
rect 4196 8691 4274 8692
rect 3796 8634 3874 8635
rect 3996 8675 4074 8676
rect 3596 8618 3674 8619
rect 3996 8619 4007 8675
rect 4063 8619 4074 8675
rect 4196 8635 4207 8691
rect 4263 8635 4274 8691
rect 4596 8691 4674 8692
rect 4196 8634 4274 8635
rect 4396 8675 4474 8676
rect 3996 8618 4074 8619
rect 4396 8619 4407 8675
rect 4463 8619 4474 8675
rect 4596 8635 4607 8691
rect 4663 8635 4674 8691
rect 4996 8691 5074 8692
rect 4596 8634 4674 8635
rect 4796 8675 4874 8676
rect 4396 8618 4474 8619
rect 4796 8619 4807 8675
rect 4863 8619 4874 8675
rect 4996 8635 5007 8691
rect 5063 8635 5074 8691
rect 5396 8691 5474 8692
rect 4996 8634 5074 8635
rect 5196 8675 5274 8676
rect 4796 8618 4874 8619
rect 5196 8619 5207 8675
rect 5263 8619 5274 8675
rect 5396 8635 5407 8691
rect 5463 8635 5474 8691
rect 5796 8691 5874 8692
rect 5396 8634 5474 8635
rect 5596 8675 5674 8676
rect 5196 8618 5274 8619
rect 5596 8619 5607 8675
rect 5663 8619 5674 8675
rect 5796 8635 5807 8691
rect 5863 8635 5874 8691
rect 6196 8691 6274 8692
rect 5796 8634 5874 8635
rect 5996 8675 6074 8676
rect 5596 8618 5674 8619
rect 5996 8619 6007 8675
rect 6063 8619 6074 8675
rect 6196 8635 6207 8691
rect 6263 8635 6274 8691
rect 6196 8634 6274 8635
rect 5996 8618 6074 8619
rect 202 8601 268 8602
rect 202 8590 209 8601
rect 0 8560 209 8590
rect 202 8549 209 8560
rect 261 8590 268 8601
rect 602 8601 668 8602
rect 602 8590 609 8601
rect 261 8560 609 8590
rect 261 8549 268 8560
rect 202 8548 268 8549
rect 602 8549 609 8560
rect 661 8590 668 8601
rect 1002 8601 1068 8602
rect 1002 8590 1009 8601
rect 661 8560 1009 8590
rect 661 8549 668 8560
rect 602 8548 668 8549
rect 1002 8549 1009 8560
rect 1061 8590 1068 8601
rect 1402 8601 1468 8602
rect 1402 8590 1409 8601
rect 1061 8560 1409 8590
rect 1061 8549 1068 8560
rect 1002 8548 1068 8549
rect 1402 8549 1409 8560
rect 1461 8590 1468 8601
rect 1802 8601 1868 8602
rect 1802 8590 1809 8601
rect 1461 8560 1809 8590
rect 1461 8549 1468 8560
rect 1402 8548 1468 8549
rect 1802 8549 1809 8560
rect 1861 8590 1868 8601
rect 2202 8601 2268 8602
rect 2202 8590 2209 8601
rect 1861 8560 2209 8590
rect 1861 8549 1868 8560
rect 1802 8548 1868 8549
rect 2202 8549 2209 8560
rect 2261 8590 2268 8601
rect 2602 8601 2668 8602
rect 2602 8590 2609 8601
rect 2261 8560 2609 8590
rect 2261 8549 2268 8560
rect 2202 8548 2268 8549
rect 2602 8549 2609 8560
rect 2661 8590 2668 8601
rect 3002 8601 3068 8602
rect 3002 8590 3009 8601
rect 2661 8560 3009 8590
rect 2661 8549 2668 8560
rect 2602 8548 2668 8549
rect 3002 8549 3009 8560
rect 3061 8590 3068 8601
rect 3402 8601 3468 8602
rect 3402 8590 3409 8601
rect 3061 8560 3409 8590
rect 3061 8549 3068 8560
rect 3002 8548 3068 8549
rect 3402 8549 3409 8560
rect 3461 8590 3468 8601
rect 3802 8601 3868 8602
rect 3802 8590 3809 8601
rect 3461 8560 3809 8590
rect 3461 8549 3468 8560
rect 3402 8548 3468 8549
rect 3802 8549 3809 8560
rect 3861 8590 3868 8601
rect 4202 8601 4268 8602
rect 4202 8590 4209 8601
rect 3861 8560 4209 8590
rect 3861 8549 3868 8560
rect 3802 8548 3868 8549
rect 4202 8549 4209 8560
rect 4261 8590 4268 8601
rect 4602 8601 4668 8602
rect 4602 8590 4609 8601
rect 4261 8560 4609 8590
rect 4261 8549 4268 8560
rect 4202 8548 4268 8549
rect 4602 8549 4609 8560
rect 4661 8590 4668 8601
rect 5002 8601 5068 8602
rect 5002 8590 5009 8601
rect 4661 8560 5009 8590
rect 4661 8549 4668 8560
rect 4602 8548 4668 8549
rect 5002 8549 5009 8560
rect 5061 8590 5068 8601
rect 5402 8601 5468 8602
rect 5402 8590 5409 8601
rect 5061 8560 5409 8590
rect 5061 8549 5068 8560
rect 5002 8548 5068 8549
rect 5402 8549 5409 8560
rect 5461 8590 5468 8601
rect 5802 8601 5868 8602
rect 5802 8590 5809 8601
rect 5461 8560 5809 8590
rect 5461 8549 5468 8560
rect 5402 8548 5468 8549
rect 5802 8549 5809 8560
rect 5861 8590 5868 8601
rect 6202 8601 6268 8602
rect 6202 8590 6209 8601
rect 5861 8560 6209 8590
rect 5861 8549 5868 8560
rect 5802 8548 5868 8549
rect 6202 8549 6209 8560
rect 6261 8590 6268 8601
rect 6704 8601 6770 8602
rect 6704 8590 6711 8601
rect 6261 8560 6711 8590
rect 6261 8549 6268 8560
rect 6202 8548 6268 8549
rect 6704 8549 6711 8560
rect 6763 8549 6770 8601
rect 6704 8548 6770 8549
rect 2 8531 68 8532
rect 2 8520 9 8531
rect 0 8490 9 8520
rect 2 8479 9 8490
rect 61 8520 68 8531
rect 402 8531 468 8532
rect 402 8520 409 8531
rect 61 8490 409 8520
rect 61 8479 68 8490
rect 2 8478 68 8479
rect 402 8479 409 8490
rect 461 8520 468 8531
rect 802 8531 868 8532
rect 802 8520 809 8531
rect 461 8490 809 8520
rect 461 8479 468 8490
rect 402 8478 468 8479
rect 802 8479 809 8490
rect 861 8520 868 8531
rect 1202 8531 1268 8532
rect 1202 8520 1209 8531
rect 861 8490 1209 8520
rect 861 8479 868 8490
rect 802 8478 868 8479
rect 1202 8479 1209 8490
rect 1261 8520 1268 8531
rect 1602 8531 1668 8532
rect 1602 8520 1609 8531
rect 1261 8490 1609 8520
rect 1261 8479 1268 8490
rect 1202 8478 1268 8479
rect 1602 8479 1609 8490
rect 1661 8520 1668 8531
rect 2002 8531 2068 8532
rect 2002 8520 2009 8531
rect 1661 8490 2009 8520
rect 1661 8479 1668 8490
rect 1602 8478 1668 8479
rect 2002 8479 2009 8490
rect 2061 8520 2068 8531
rect 2402 8531 2468 8532
rect 2402 8520 2409 8531
rect 2061 8490 2409 8520
rect 2061 8479 2068 8490
rect 2002 8478 2068 8479
rect 2402 8479 2409 8490
rect 2461 8520 2468 8531
rect 2802 8531 2868 8532
rect 2802 8520 2809 8531
rect 2461 8490 2809 8520
rect 2461 8479 2468 8490
rect 2402 8478 2468 8479
rect 2802 8479 2809 8490
rect 2861 8520 2868 8531
rect 3202 8531 3268 8532
rect 3202 8520 3209 8531
rect 2861 8490 3209 8520
rect 2861 8479 2868 8490
rect 2802 8478 2868 8479
rect 3202 8479 3209 8490
rect 3261 8520 3268 8531
rect 3602 8531 3668 8532
rect 3602 8520 3609 8531
rect 3261 8490 3609 8520
rect 3261 8479 3268 8490
rect 3202 8478 3268 8479
rect 3602 8479 3609 8490
rect 3661 8520 3668 8531
rect 4002 8531 4068 8532
rect 4002 8520 4009 8531
rect 3661 8490 4009 8520
rect 3661 8479 3668 8490
rect 3602 8478 3668 8479
rect 4002 8479 4009 8490
rect 4061 8520 4068 8531
rect 4402 8531 4468 8532
rect 4402 8520 4409 8531
rect 4061 8490 4409 8520
rect 4061 8479 4068 8490
rect 4002 8478 4068 8479
rect 4402 8479 4409 8490
rect 4461 8520 4468 8531
rect 4802 8531 4868 8532
rect 4802 8520 4809 8531
rect 4461 8490 4809 8520
rect 4461 8479 4468 8490
rect 4402 8478 4468 8479
rect 4802 8479 4809 8490
rect 4861 8520 4868 8531
rect 5202 8531 5268 8532
rect 5202 8520 5209 8531
rect 4861 8490 5209 8520
rect 4861 8479 4868 8490
rect 4802 8478 4868 8479
rect 5202 8479 5209 8490
rect 5261 8520 5268 8531
rect 5602 8531 5668 8532
rect 5602 8520 5609 8531
rect 5261 8490 5609 8520
rect 5261 8479 5268 8490
rect 5202 8478 5268 8479
rect 5602 8479 5609 8490
rect 5661 8520 5668 8531
rect 6002 8531 6068 8532
rect 6002 8520 6009 8531
rect 5661 8490 6009 8520
rect 5661 8479 5668 8490
rect 5602 8478 5668 8479
rect 6002 8479 6009 8490
rect 6061 8520 6068 8531
rect 6402 8531 6468 8532
rect 6402 8520 6409 8531
rect 6061 8490 6409 8520
rect 6061 8479 6068 8490
rect 6002 8478 6068 8479
rect 6402 8479 6409 8490
rect 6461 8520 6468 8531
rect 6500 8531 6566 8532
rect 6500 8520 6507 8531
rect 6461 8490 6507 8520
rect 6461 8479 6468 8490
rect 6402 8478 6468 8479
rect 6500 8479 6507 8490
rect 6559 8479 6566 8531
rect 6500 8478 6566 8479
rect 202 8461 268 8462
rect 202 8450 209 8461
rect 0 8420 209 8450
rect 202 8409 209 8420
rect 261 8450 268 8461
rect 602 8461 668 8462
rect 602 8450 609 8461
rect 261 8420 609 8450
rect 261 8409 268 8420
rect 202 8408 268 8409
rect 602 8409 609 8420
rect 661 8450 668 8461
rect 1002 8461 1068 8462
rect 1002 8450 1009 8461
rect 661 8420 1009 8450
rect 661 8409 668 8420
rect 602 8408 668 8409
rect 1002 8409 1009 8420
rect 1061 8450 1068 8461
rect 1402 8461 1468 8462
rect 1402 8450 1409 8461
rect 1061 8420 1409 8450
rect 1061 8409 1068 8420
rect 1002 8408 1068 8409
rect 1402 8409 1409 8420
rect 1461 8450 1468 8461
rect 1802 8461 1868 8462
rect 1802 8450 1809 8461
rect 1461 8420 1809 8450
rect 1461 8409 1468 8420
rect 1402 8408 1468 8409
rect 1802 8409 1809 8420
rect 1861 8450 1868 8461
rect 2202 8461 2268 8462
rect 2202 8450 2209 8461
rect 1861 8420 2209 8450
rect 1861 8409 1868 8420
rect 1802 8408 1868 8409
rect 2202 8409 2209 8420
rect 2261 8450 2268 8461
rect 2602 8461 2668 8462
rect 2602 8450 2609 8461
rect 2261 8420 2609 8450
rect 2261 8409 2268 8420
rect 2202 8408 2268 8409
rect 2602 8409 2609 8420
rect 2661 8450 2668 8461
rect 3002 8461 3068 8462
rect 3002 8450 3009 8461
rect 2661 8420 3009 8450
rect 2661 8409 2668 8420
rect 2602 8408 2668 8409
rect 3002 8409 3009 8420
rect 3061 8450 3068 8461
rect 3402 8461 3468 8462
rect 3402 8450 3409 8461
rect 3061 8420 3409 8450
rect 3061 8409 3068 8420
rect 3002 8408 3068 8409
rect 3402 8409 3409 8420
rect 3461 8450 3468 8461
rect 3802 8461 3868 8462
rect 3802 8450 3809 8461
rect 3461 8420 3809 8450
rect 3461 8409 3468 8420
rect 3402 8408 3468 8409
rect 3802 8409 3809 8420
rect 3861 8450 3868 8461
rect 4202 8461 4268 8462
rect 4202 8450 4209 8461
rect 3861 8420 4209 8450
rect 3861 8409 3868 8420
rect 3802 8408 3868 8409
rect 4202 8409 4209 8420
rect 4261 8450 4268 8461
rect 4602 8461 4668 8462
rect 4602 8450 4609 8461
rect 4261 8420 4609 8450
rect 4261 8409 4268 8420
rect 4202 8408 4268 8409
rect 4602 8409 4609 8420
rect 4661 8450 4668 8461
rect 5002 8461 5068 8462
rect 5002 8450 5009 8461
rect 4661 8420 5009 8450
rect 4661 8409 4668 8420
rect 4602 8408 4668 8409
rect 5002 8409 5009 8420
rect 5061 8450 5068 8461
rect 5402 8461 5468 8462
rect 5402 8450 5409 8461
rect 5061 8420 5409 8450
rect 5061 8409 5068 8420
rect 5002 8408 5068 8409
rect 5402 8409 5409 8420
rect 5461 8450 5468 8461
rect 5802 8461 5868 8462
rect 5802 8450 5809 8461
rect 5461 8420 5809 8450
rect 5461 8409 5468 8420
rect 5402 8408 5468 8409
rect 5802 8409 5809 8420
rect 5861 8450 5868 8461
rect 6202 8461 6268 8462
rect 6202 8450 6209 8461
rect 5861 8420 6209 8450
rect 5861 8409 5868 8420
rect 5802 8408 5868 8409
rect 6202 8409 6209 8420
rect 6261 8450 6268 8461
rect 6704 8461 6770 8462
rect 6704 8450 6711 8461
rect 6261 8420 6711 8450
rect 6261 8409 6268 8420
rect 6202 8408 6268 8409
rect 6704 8409 6711 8420
rect 6763 8409 6770 8461
rect 6704 8408 6770 8409
rect 2 8391 68 8392
rect 2 8380 9 8391
rect 0 8350 9 8380
rect 2 8339 9 8350
rect 61 8380 68 8391
rect 402 8391 468 8392
rect 402 8380 409 8391
rect 61 8350 409 8380
rect 61 8339 68 8350
rect 2 8338 68 8339
rect 402 8339 409 8350
rect 461 8380 468 8391
rect 802 8391 868 8392
rect 802 8380 809 8391
rect 461 8350 809 8380
rect 461 8339 468 8350
rect 402 8338 468 8339
rect 802 8339 809 8350
rect 861 8380 868 8391
rect 1202 8391 1268 8392
rect 1202 8380 1209 8391
rect 861 8350 1209 8380
rect 861 8339 868 8350
rect 802 8338 868 8339
rect 1202 8339 1209 8350
rect 1261 8380 1268 8391
rect 1602 8391 1668 8392
rect 1602 8380 1609 8391
rect 1261 8350 1609 8380
rect 1261 8339 1268 8350
rect 1202 8338 1268 8339
rect 1602 8339 1609 8350
rect 1661 8380 1668 8391
rect 2002 8391 2068 8392
rect 2002 8380 2009 8391
rect 1661 8350 2009 8380
rect 1661 8339 1668 8350
rect 1602 8338 1668 8339
rect 2002 8339 2009 8350
rect 2061 8380 2068 8391
rect 2402 8391 2468 8392
rect 2402 8380 2409 8391
rect 2061 8350 2409 8380
rect 2061 8339 2068 8350
rect 2002 8338 2068 8339
rect 2402 8339 2409 8350
rect 2461 8380 2468 8391
rect 2802 8391 2868 8392
rect 2802 8380 2809 8391
rect 2461 8350 2809 8380
rect 2461 8339 2468 8350
rect 2402 8338 2468 8339
rect 2802 8339 2809 8350
rect 2861 8380 2868 8391
rect 3202 8391 3268 8392
rect 3202 8380 3209 8391
rect 2861 8350 3209 8380
rect 2861 8339 2868 8350
rect 2802 8338 2868 8339
rect 3202 8339 3209 8350
rect 3261 8380 3268 8391
rect 3602 8391 3668 8392
rect 3602 8380 3609 8391
rect 3261 8350 3609 8380
rect 3261 8339 3268 8350
rect 3202 8338 3268 8339
rect 3602 8339 3609 8350
rect 3661 8380 3668 8391
rect 4002 8391 4068 8392
rect 4002 8380 4009 8391
rect 3661 8350 4009 8380
rect 3661 8339 3668 8350
rect 3602 8338 3668 8339
rect 4002 8339 4009 8350
rect 4061 8380 4068 8391
rect 4402 8391 4468 8392
rect 4402 8380 4409 8391
rect 4061 8350 4409 8380
rect 4061 8339 4068 8350
rect 4002 8338 4068 8339
rect 4402 8339 4409 8350
rect 4461 8380 4468 8391
rect 4802 8391 4868 8392
rect 4802 8380 4809 8391
rect 4461 8350 4809 8380
rect 4461 8339 4468 8350
rect 4402 8338 4468 8339
rect 4802 8339 4809 8350
rect 4861 8380 4868 8391
rect 5202 8391 5268 8392
rect 5202 8380 5209 8391
rect 4861 8350 5209 8380
rect 4861 8339 4868 8350
rect 4802 8338 4868 8339
rect 5202 8339 5209 8350
rect 5261 8380 5268 8391
rect 5602 8391 5668 8392
rect 5602 8380 5609 8391
rect 5261 8350 5609 8380
rect 5261 8339 5268 8350
rect 5202 8338 5268 8339
rect 5602 8339 5609 8350
rect 5661 8380 5668 8391
rect 6002 8391 6068 8392
rect 6002 8380 6009 8391
rect 5661 8350 6009 8380
rect 5661 8339 5668 8350
rect 5602 8338 5668 8339
rect 6002 8339 6009 8350
rect 6061 8380 6068 8391
rect 6402 8391 6468 8392
rect 6402 8380 6409 8391
rect 6061 8350 6409 8380
rect 6061 8339 6068 8350
rect 6002 8338 6068 8339
rect 6402 8339 6409 8350
rect 6461 8380 6468 8391
rect 6500 8391 6566 8392
rect 6500 8380 6507 8391
rect 6461 8350 6507 8380
rect 6461 8339 6468 8350
rect 6402 8338 6468 8339
rect 6500 8339 6507 8350
rect 6559 8339 6566 8391
rect 6500 8338 6566 8339
rect 202 8321 268 8322
rect 202 8310 209 8321
rect 0 8280 209 8310
rect 202 8269 209 8280
rect 261 8310 268 8321
rect 602 8321 668 8322
rect 602 8310 609 8321
rect 261 8280 609 8310
rect 261 8269 268 8280
rect 202 8268 268 8269
rect 602 8269 609 8280
rect 661 8310 668 8321
rect 1002 8321 1068 8322
rect 1002 8310 1009 8321
rect 661 8280 1009 8310
rect 661 8269 668 8280
rect 602 8268 668 8269
rect 1002 8269 1009 8280
rect 1061 8310 1068 8321
rect 1402 8321 1468 8322
rect 1402 8310 1409 8321
rect 1061 8280 1409 8310
rect 1061 8269 1068 8280
rect 1002 8268 1068 8269
rect 1402 8269 1409 8280
rect 1461 8310 1468 8321
rect 1802 8321 1868 8322
rect 1802 8310 1809 8321
rect 1461 8280 1809 8310
rect 1461 8269 1468 8280
rect 1402 8268 1468 8269
rect 1802 8269 1809 8280
rect 1861 8310 1868 8321
rect 2202 8321 2268 8322
rect 2202 8310 2209 8321
rect 1861 8280 2209 8310
rect 1861 8269 1868 8280
rect 1802 8268 1868 8269
rect 2202 8269 2209 8280
rect 2261 8310 2268 8321
rect 2602 8321 2668 8322
rect 2602 8310 2609 8321
rect 2261 8280 2609 8310
rect 2261 8269 2268 8280
rect 2202 8268 2268 8269
rect 2602 8269 2609 8280
rect 2661 8310 2668 8321
rect 3002 8321 3068 8322
rect 3002 8310 3009 8321
rect 2661 8280 3009 8310
rect 2661 8269 2668 8280
rect 2602 8268 2668 8269
rect 3002 8269 3009 8280
rect 3061 8310 3068 8321
rect 3402 8321 3468 8322
rect 3402 8310 3409 8321
rect 3061 8280 3409 8310
rect 3061 8269 3068 8280
rect 3002 8268 3068 8269
rect 3402 8269 3409 8280
rect 3461 8310 3468 8321
rect 3802 8321 3868 8322
rect 3802 8310 3809 8321
rect 3461 8280 3809 8310
rect 3461 8269 3468 8280
rect 3402 8268 3468 8269
rect 3802 8269 3809 8280
rect 3861 8310 3868 8321
rect 4202 8321 4268 8322
rect 4202 8310 4209 8321
rect 3861 8280 4209 8310
rect 3861 8269 3868 8280
rect 3802 8268 3868 8269
rect 4202 8269 4209 8280
rect 4261 8310 4268 8321
rect 4602 8321 4668 8322
rect 4602 8310 4609 8321
rect 4261 8280 4609 8310
rect 4261 8269 4268 8280
rect 4202 8268 4268 8269
rect 4602 8269 4609 8280
rect 4661 8310 4668 8321
rect 5002 8321 5068 8322
rect 5002 8310 5009 8321
rect 4661 8280 5009 8310
rect 4661 8269 4668 8280
rect 4602 8268 4668 8269
rect 5002 8269 5009 8280
rect 5061 8310 5068 8321
rect 5402 8321 5468 8322
rect 5402 8310 5409 8321
rect 5061 8280 5409 8310
rect 5061 8269 5068 8280
rect 5002 8268 5068 8269
rect 5402 8269 5409 8280
rect 5461 8310 5468 8321
rect 5802 8321 5868 8322
rect 5802 8310 5809 8321
rect 5461 8280 5809 8310
rect 5461 8269 5468 8280
rect 5402 8268 5468 8269
rect 5802 8269 5809 8280
rect 5861 8310 5868 8321
rect 6202 8321 6268 8322
rect 6202 8310 6209 8321
rect 5861 8280 6209 8310
rect 5861 8269 5868 8280
rect 5802 8268 5868 8269
rect 6202 8269 6209 8280
rect 6261 8310 6268 8321
rect 6704 8321 6770 8322
rect 6704 8310 6711 8321
rect 6261 8280 6711 8310
rect 6261 8269 6268 8280
rect 6202 8268 6268 8269
rect 6704 8269 6711 8280
rect 6763 8269 6770 8321
rect 6704 8268 6770 8269
rect 2 8251 68 8252
rect 2 8240 9 8251
rect 0 8210 9 8240
rect 2 8199 9 8210
rect 61 8240 68 8251
rect 402 8251 468 8252
rect 402 8240 409 8251
rect 61 8210 409 8240
rect 61 8199 68 8210
rect 2 8198 68 8199
rect 402 8199 409 8210
rect 461 8240 468 8251
rect 802 8251 868 8252
rect 802 8240 809 8251
rect 461 8210 809 8240
rect 461 8199 468 8210
rect 402 8198 468 8199
rect 802 8199 809 8210
rect 861 8240 868 8251
rect 1202 8251 1268 8252
rect 1202 8240 1209 8251
rect 861 8210 1209 8240
rect 861 8199 868 8210
rect 802 8198 868 8199
rect 1202 8199 1209 8210
rect 1261 8240 1268 8251
rect 1602 8251 1668 8252
rect 1602 8240 1609 8251
rect 1261 8210 1609 8240
rect 1261 8199 1268 8210
rect 1202 8198 1268 8199
rect 1602 8199 1609 8210
rect 1661 8240 1668 8251
rect 2002 8251 2068 8252
rect 2002 8240 2009 8251
rect 1661 8210 2009 8240
rect 1661 8199 1668 8210
rect 1602 8198 1668 8199
rect 2002 8199 2009 8210
rect 2061 8240 2068 8251
rect 2402 8251 2468 8252
rect 2402 8240 2409 8251
rect 2061 8210 2409 8240
rect 2061 8199 2068 8210
rect 2002 8198 2068 8199
rect 2402 8199 2409 8210
rect 2461 8240 2468 8251
rect 2802 8251 2868 8252
rect 2802 8240 2809 8251
rect 2461 8210 2809 8240
rect 2461 8199 2468 8210
rect 2402 8198 2468 8199
rect 2802 8199 2809 8210
rect 2861 8240 2868 8251
rect 3202 8251 3268 8252
rect 3202 8240 3209 8251
rect 2861 8210 3209 8240
rect 2861 8199 2868 8210
rect 2802 8198 2868 8199
rect 3202 8199 3209 8210
rect 3261 8240 3268 8251
rect 3602 8251 3668 8252
rect 3602 8240 3609 8251
rect 3261 8210 3609 8240
rect 3261 8199 3268 8210
rect 3202 8198 3268 8199
rect 3602 8199 3609 8210
rect 3661 8240 3668 8251
rect 4002 8251 4068 8252
rect 4002 8240 4009 8251
rect 3661 8210 4009 8240
rect 3661 8199 3668 8210
rect 3602 8198 3668 8199
rect 4002 8199 4009 8210
rect 4061 8240 4068 8251
rect 4402 8251 4468 8252
rect 4402 8240 4409 8251
rect 4061 8210 4409 8240
rect 4061 8199 4068 8210
rect 4002 8198 4068 8199
rect 4402 8199 4409 8210
rect 4461 8240 4468 8251
rect 4802 8251 4868 8252
rect 4802 8240 4809 8251
rect 4461 8210 4809 8240
rect 4461 8199 4468 8210
rect 4402 8198 4468 8199
rect 4802 8199 4809 8210
rect 4861 8240 4868 8251
rect 5202 8251 5268 8252
rect 5202 8240 5209 8251
rect 4861 8210 5209 8240
rect 4861 8199 4868 8210
rect 4802 8198 4868 8199
rect 5202 8199 5209 8210
rect 5261 8240 5268 8251
rect 5602 8251 5668 8252
rect 5602 8240 5609 8251
rect 5261 8210 5609 8240
rect 5261 8199 5268 8210
rect 5202 8198 5268 8199
rect 5602 8199 5609 8210
rect 5661 8240 5668 8251
rect 6002 8251 6068 8252
rect 6002 8240 6009 8251
rect 5661 8210 6009 8240
rect 5661 8199 5668 8210
rect 5602 8198 5668 8199
rect 6002 8199 6009 8210
rect 6061 8240 6068 8251
rect 6402 8251 6468 8252
rect 6402 8240 6409 8251
rect 6061 8210 6409 8240
rect 6061 8199 6068 8210
rect 6002 8198 6068 8199
rect 6402 8199 6409 8210
rect 6461 8240 6468 8251
rect 6500 8251 6566 8252
rect 6500 8240 6507 8251
rect 6461 8210 6507 8240
rect 6461 8199 6468 8210
rect 6402 8198 6468 8199
rect 6500 8199 6507 8210
rect 6559 8199 6566 8251
rect 6500 8198 6566 8199
rect 202 8181 268 8182
rect 202 8170 209 8181
rect 0 8140 209 8170
rect 202 8129 209 8140
rect 261 8170 268 8181
rect 602 8181 668 8182
rect 602 8170 609 8181
rect 261 8140 609 8170
rect 261 8129 268 8140
rect 202 8128 268 8129
rect 602 8129 609 8140
rect 661 8170 668 8181
rect 1002 8181 1068 8182
rect 1002 8170 1009 8181
rect 661 8140 1009 8170
rect 661 8129 668 8140
rect 602 8128 668 8129
rect 1002 8129 1009 8140
rect 1061 8170 1068 8181
rect 1402 8181 1468 8182
rect 1402 8170 1409 8181
rect 1061 8140 1409 8170
rect 1061 8129 1068 8140
rect 1002 8128 1068 8129
rect 1402 8129 1409 8140
rect 1461 8170 1468 8181
rect 1802 8181 1868 8182
rect 1802 8170 1809 8181
rect 1461 8140 1809 8170
rect 1461 8129 1468 8140
rect 1402 8128 1468 8129
rect 1802 8129 1809 8140
rect 1861 8170 1868 8181
rect 2202 8181 2268 8182
rect 2202 8170 2209 8181
rect 1861 8140 2209 8170
rect 1861 8129 1868 8140
rect 1802 8128 1868 8129
rect 2202 8129 2209 8140
rect 2261 8170 2268 8181
rect 2602 8181 2668 8182
rect 2602 8170 2609 8181
rect 2261 8140 2609 8170
rect 2261 8129 2268 8140
rect 2202 8128 2268 8129
rect 2602 8129 2609 8140
rect 2661 8170 2668 8181
rect 3002 8181 3068 8182
rect 3002 8170 3009 8181
rect 2661 8140 3009 8170
rect 2661 8129 2668 8140
rect 2602 8128 2668 8129
rect 3002 8129 3009 8140
rect 3061 8170 3068 8181
rect 3402 8181 3468 8182
rect 3402 8170 3409 8181
rect 3061 8140 3409 8170
rect 3061 8129 3068 8140
rect 3002 8128 3068 8129
rect 3402 8129 3409 8140
rect 3461 8170 3468 8181
rect 3802 8181 3868 8182
rect 3802 8170 3809 8181
rect 3461 8140 3809 8170
rect 3461 8129 3468 8140
rect 3402 8128 3468 8129
rect 3802 8129 3809 8140
rect 3861 8170 3868 8181
rect 4202 8181 4268 8182
rect 4202 8170 4209 8181
rect 3861 8140 4209 8170
rect 3861 8129 3868 8140
rect 3802 8128 3868 8129
rect 4202 8129 4209 8140
rect 4261 8170 4268 8181
rect 4602 8181 4668 8182
rect 4602 8170 4609 8181
rect 4261 8140 4609 8170
rect 4261 8129 4268 8140
rect 4202 8128 4268 8129
rect 4602 8129 4609 8140
rect 4661 8170 4668 8181
rect 5002 8181 5068 8182
rect 5002 8170 5009 8181
rect 4661 8140 5009 8170
rect 4661 8129 4668 8140
rect 4602 8128 4668 8129
rect 5002 8129 5009 8140
rect 5061 8170 5068 8181
rect 5402 8181 5468 8182
rect 5402 8170 5409 8181
rect 5061 8140 5409 8170
rect 5061 8129 5068 8140
rect 5002 8128 5068 8129
rect 5402 8129 5409 8140
rect 5461 8170 5468 8181
rect 5802 8181 5868 8182
rect 5802 8170 5809 8181
rect 5461 8140 5809 8170
rect 5461 8129 5468 8140
rect 5402 8128 5468 8129
rect 5802 8129 5809 8140
rect 5861 8170 5868 8181
rect 6202 8181 6268 8182
rect 6202 8170 6209 8181
rect 5861 8140 6209 8170
rect 5861 8129 5868 8140
rect 5802 8128 5868 8129
rect 6202 8129 6209 8140
rect 6261 8170 6268 8181
rect 6704 8181 6770 8182
rect 6704 8170 6711 8181
rect 6261 8140 6711 8170
rect 6261 8129 6268 8140
rect 6202 8128 6268 8129
rect 6704 8129 6711 8140
rect 6763 8129 6770 8181
rect 6704 8128 6770 8129
rect 2 8111 68 8112
rect 2 8100 9 8111
rect 0 8070 9 8100
rect 2 8059 9 8070
rect 61 8100 68 8111
rect 402 8111 468 8112
rect 402 8100 409 8111
rect 61 8070 409 8100
rect 61 8059 68 8070
rect 2 8058 68 8059
rect 402 8059 409 8070
rect 461 8100 468 8111
rect 802 8111 868 8112
rect 802 8100 809 8111
rect 461 8070 809 8100
rect 461 8059 468 8070
rect 402 8058 468 8059
rect 802 8059 809 8070
rect 861 8100 868 8111
rect 1202 8111 1268 8112
rect 1202 8100 1209 8111
rect 861 8070 1209 8100
rect 861 8059 868 8070
rect 802 8058 868 8059
rect 1202 8059 1209 8070
rect 1261 8100 1268 8111
rect 1602 8111 1668 8112
rect 1602 8100 1609 8111
rect 1261 8070 1609 8100
rect 1261 8059 1268 8070
rect 1202 8058 1268 8059
rect 1602 8059 1609 8070
rect 1661 8100 1668 8111
rect 2002 8111 2068 8112
rect 2002 8100 2009 8111
rect 1661 8070 2009 8100
rect 1661 8059 1668 8070
rect 1602 8058 1668 8059
rect 2002 8059 2009 8070
rect 2061 8100 2068 8111
rect 2402 8111 2468 8112
rect 2402 8100 2409 8111
rect 2061 8070 2409 8100
rect 2061 8059 2068 8070
rect 2002 8058 2068 8059
rect 2402 8059 2409 8070
rect 2461 8100 2468 8111
rect 2802 8111 2868 8112
rect 2802 8100 2809 8111
rect 2461 8070 2809 8100
rect 2461 8059 2468 8070
rect 2402 8058 2468 8059
rect 2802 8059 2809 8070
rect 2861 8100 2868 8111
rect 3202 8111 3268 8112
rect 3202 8100 3209 8111
rect 2861 8070 3209 8100
rect 2861 8059 2868 8070
rect 2802 8058 2868 8059
rect 3202 8059 3209 8070
rect 3261 8100 3268 8111
rect 3602 8111 3668 8112
rect 3602 8100 3609 8111
rect 3261 8070 3609 8100
rect 3261 8059 3268 8070
rect 3202 8058 3268 8059
rect 3602 8059 3609 8070
rect 3661 8100 3668 8111
rect 4002 8111 4068 8112
rect 4002 8100 4009 8111
rect 3661 8070 4009 8100
rect 3661 8059 3668 8070
rect 3602 8058 3668 8059
rect 4002 8059 4009 8070
rect 4061 8100 4068 8111
rect 4402 8111 4468 8112
rect 4402 8100 4409 8111
rect 4061 8070 4409 8100
rect 4061 8059 4068 8070
rect 4002 8058 4068 8059
rect 4402 8059 4409 8070
rect 4461 8100 4468 8111
rect 4802 8111 4868 8112
rect 4802 8100 4809 8111
rect 4461 8070 4809 8100
rect 4461 8059 4468 8070
rect 4402 8058 4468 8059
rect 4802 8059 4809 8070
rect 4861 8100 4868 8111
rect 5202 8111 5268 8112
rect 5202 8100 5209 8111
rect 4861 8070 5209 8100
rect 4861 8059 4868 8070
rect 4802 8058 4868 8059
rect 5202 8059 5209 8070
rect 5261 8100 5268 8111
rect 5602 8111 5668 8112
rect 5602 8100 5609 8111
rect 5261 8070 5609 8100
rect 5261 8059 5268 8070
rect 5202 8058 5268 8059
rect 5602 8059 5609 8070
rect 5661 8100 5668 8111
rect 6002 8111 6068 8112
rect 6002 8100 6009 8111
rect 5661 8070 6009 8100
rect 5661 8059 5668 8070
rect 5602 8058 5668 8059
rect 6002 8059 6009 8070
rect 6061 8100 6068 8111
rect 6402 8111 6468 8112
rect 6402 8100 6409 8111
rect 6061 8070 6409 8100
rect 6061 8059 6068 8070
rect 6002 8058 6068 8059
rect 6402 8059 6409 8070
rect 6461 8100 6468 8111
rect 6500 8111 6566 8112
rect 6500 8100 6507 8111
rect 6461 8070 6507 8100
rect 6461 8059 6468 8070
rect 6402 8058 6468 8059
rect 6500 8059 6507 8070
rect 6559 8059 6566 8111
rect 6500 8058 6566 8059
rect 202 8041 268 8042
rect 202 8030 209 8041
rect 0 8000 209 8030
rect 202 7989 209 8000
rect 261 8030 268 8041
rect 602 8041 668 8042
rect 602 8030 609 8041
rect 261 8000 609 8030
rect 261 7989 268 8000
rect 202 7988 268 7989
rect 602 7989 609 8000
rect 661 8030 668 8041
rect 1002 8041 1068 8042
rect 1002 8030 1009 8041
rect 661 8000 1009 8030
rect 661 7989 668 8000
rect 602 7988 668 7989
rect 1002 7989 1009 8000
rect 1061 8030 1068 8041
rect 1402 8041 1468 8042
rect 1402 8030 1409 8041
rect 1061 8000 1409 8030
rect 1061 7989 1068 8000
rect 1002 7988 1068 7989
rect 1402 7989 1409 8000
rect 1461 8030 1468 8041
rect 1802 8041 1868 8042
rect 1802 8030 1809 8041
rect 1461 8000 1809 8030
rect 1461 7989 1468 8000
rect 1402 7988 1468 7989
rect 1802 7989 1809 8000
rect 1861 8030 1868 8041
rect 2202 8041 2268 8042
rect 2202 8030 2209 8041
rect 1861 8000 2209 8030
rect 1861 7989 1868 8000
rect 1802 7988 1868 7989
rect 2202 7989 2209 8000
rect 2261 8030 2268 8041
rect 2602 8041 2668 8042
rect 2602 8030 2609 8041
rect 2261 8000 2609 8030
rect 2261 7989 2268 8000
rect 2202 7988 2268 7989
rect 2602 7989 2609 8000
rect 2661 8030 2668 8041
rect 3002 8041 3068 8042
rect 3002 8030 3009 8041
rect 2661 8000 3009 8030
rect 2661 7989 2668 8000
rect 2602 7988 2668 7989
rect 3002 7989 3009 8000
rect 3061 8030 3068 8041
rect 3402 8041 3468 8042
rect 3402 8030 3409 8041
rect 3061 8000 3409 8030
rect 3061 7989 3068 8000
rect 3002 7988 3068 7989
rect 3402 7989 3409 8000
rect 3461 8030 3468 8041
rect 3802 8041 3868 8042
rect 3802 8030 3809 8041
rect 3461 8000 3809 8030
rect 3461 7989 3468 8000
rect 3402 7988 3468 7989
rect 3802 7989 3809 8000
rect 3861 8030 3868 8041
rect 4202 8041 4268 8042
rect 4202 8030 4209 8041
rect 3861 8000 4209 8030
rect 3861 7989 3868 8000
rect 3802 7988 3868 7989
rect 4202 7989 4209 8000
rect 4261 8030 4268 8041
rect 4602 8041 4668 8042
rect 4602 8030 4609 8041
rect 4261 8000 4609 8030
rect 4261 7989 4268 8000
rect 4202 7988 4268 7989
rect 4602 7989 4609 8000
rect 4661 8030 4668 8041
rect 5002 8041 5068 8042
rect 5002 8030 5009 8041
rect 4661 8000 5009 8030
rect 4661 7989 4668 8000
rect 4602 7988 4668 7989
rect 5002 7989 5009 8000
rect 5061 8030 5068 8041
rect 5402 8041 5468 8042
rect 5402 8030 5409 8041
rect 5061 8000 5409 8030
rect 5061 7989 5068 8000
rect 5002 7988 5068 7989
rect 5402 7989 5409 8000
rect 5461 8030 5468 8041
rect 5802 8041 5868 8042
rect 5802 8030 5809 8041
rect 5461 8000 5809 8030
rect 5461 7989 5468 8000
rect 5402 7988 5468 7989
rect 5802 7989 5809 8000
rect 5861 8030 5868 8041
rect 6202 8041 6268 8042
rect 6202 8030 6209 8041
rect 5861 8000 6209 8030
rect 5861 7989 5868 8000
rect 5802 7988 5868 7989
rect 6202 7989 6209 8000
rect 6261 8030 6268 8041
rect 6704 8041 6770 8042
rect 6704 8030 6711 8041
rect 6261 8000 6711 8030
rect 6261 7989 6268 8000
rect 6202 7988 6268 7989
rect 6704 7989 6711 8000
rect 6763 7989 6770 8041
rect 6704 7988 6770 7989
rect 2 7971 68 7972
rect 2 7960 9 7971
rect 0 7930 9 7960
rect 2 7919 9 7930
rect 61 7960 68 7971
rect 402 7971 468 7972
rect 402 7960 409 7971
rect 61 7930 409 7960
rect 61 7919 68 7930
rect 2 7918 68 7919
rect 402 7919 409 7930
rect 461 7960 468 7971
rect 802 7971 868 7972
rect 802 7960 809 7971
rect 461 7930 809 7960
rect 461 7919 468 7930
rect 402 7918 468 7919
rect 802 7919 809 7930
rect 861 7960 868 7971
rect 1202 7971 1268 7972
rect 1202 7960 1209 7971
rect 861 7930 1209 7960
rect 861 7919 868 7930
rect 802 7918 868 7919
rect 1202 7919 1209 7930
rect 1261 7960 1268 7971
rect 1602 7971 1668 7972
rect 1602 7960 1609 7971
rect 1261 7930 1609 7960
rect 1261 7919 1268 7930
rect 1202 7918 1268 7919
rect 1602 7919 1609 7930
rect 1661 7960 1668 7971
rect 2002 7971 2068 7972
rect 2002 7960 2009 7971
rect 1661 7930 2009 7960
rect 1661 7919 1668 7930
rect 1602 7918 1668 7919
rect 2002 7919 2009 7930
rect 2061 7960 2068 7971
rect 2402 7971 2468 7972
rect 2402 7960 2409 7971
rect 2061 7930 2409 7960
rect 2061 7919 2068 7930
rect 2002 7918 2068 7919
rect 2402 7919 2409 7930
rect 2461 7960 2468 7971
rect 2802 7971 2868 7972
rect 2802 7960 2809 7971
rect 2461 7930 2809 7960
rect 2461 7919 2468 7930
rect 2402 7918 2468 7919
rect 2802 7919 2809 7930
rect 2861 7960 2868 7971
rect 3202 7971 3268 7972
rect 3202 7960 3209 7971
rect 2861 7930 3209 7960
rect 2861 7919 2868 7930
rect 2802 7918 2868 7919
rect 3202 7919 3209 7930
rect 3261 7960 3268 7971
rect 3602 7971 3668 7972
rect 3602 7960 3609 7971
rect 3261 7930 3609 7960
rect 3261 7919 3268 7930
rect 3202 7918 3268 7919
rect 3602 7919 3609 7930
rect 3661 7960 3668 7971
rect 4002 7971 4068 7972
rect 4002 7960 4009 7971
rect 3661 7930 4009 7960
rect 3661 7919 3668 7930
rect 3602 7918 3668 7919
rect 4002 7919 4009 7930
rect 4061 7960 4068 7971
rect 4402 7971 4468 7972
rect 4402 7960 4409 7971
rect 4061 7930 4409 7960
rect 4061 7919 4068 7930
rect 4002 7918 4068 7919
rect 4402 7919 4409 7930
rect 4461 7960 4468 7971
rect 4802 7971 4868 7972
rect 4802 7960 4809 7971
rect 4461 7930 4809 7960
rect 4461 7919 4468 7930
rect 4402 7918 4468 7919
rect 4802 7919 4809 7930
rect 4861 7960 4868 7971
rect 5202 7971 5268 7972
rect 5202 7960 5209 7971
rect 4861 7930 5209 7960
rect 4861 7919 4868 7930
rect 4802 7918 4868 7919
rect 5202 7919 5209 7930
rect 5261 7960 5268 7971
rect 5602 7971 5668 7972
rect 5602 7960 5609 7971
rect 5261 7930 5609 7960
rect 5261 7919 5268 7930
rect 5202 7918 5268 7919
rect 5602 7919 5609 7930
rect 5661 7960 5668 7971
rect 6002 7971 6068 7972
rect 6002 7960 6009 7971
rect 5661 7930 6009 7960
rect 5661 7919 5668 7930
rect 5602 7918 5668 7919
rect 6002 7919 6009 7930
rect 6061 7960 6068 7971
rect 6402 7971 6468 7972
rect 6402 7960 6409 7971
rect 6061 7930 6409 7960
rect 6061 7919 6068 7930
rect 6002 7918 6068 7919
rect 6402 7919 6409 7930
rect 6461 7960 6468 7971
rect 6500 7971 6566 7972
rect 6500 7960 6507 7971
rect 6461 7930 6507 7960
rect 6461 7919 6468 7930
rect 6402 7918 6468 7919
rect 6500 7919 6507 7930
rect 6559 7919 6566 7971
rect 6500 7918 6566 7919
rect 202 7901 268 7902
rect 202 7890 209 7901
rect 0 7860 209 7890
rect 202 7849 209 7860
rect 261 7890 268 7901
rect 602 7901 668 7902
rect 602 7890 609 7901
rect 261 7860 609 7890
rect 261 7849 268 7860
rect 202 7848 268 7849
rect 602 7849 609 7860
rect 661 7890 668 7901
rect 1002 7901 1068 7902
rect 1002 7890 1009 7901
rect 661 7860 1009 7890
rect 661 7849 668 7860
rect 602 7848 668 7849
rect 1002 7849 1009 7860
rect 1061 7890 1068 7901
rect 1402 7901 1468 7902
rect 1402 7890 1409 7901
rect 1061 7860 1409 7890
rect 1061 7849 1068 7860
rect 1002 7848 1068 7849
rect 1402 7849 1409 7860
rect 1461 7890 1468 7901
rect 1802 7901 1868 7902
rect 1802 7890 1809 7901
rect 1461 7860 1809 7890
rect 1461 7849 1468 7860
rect 1402 7848 1468 7849
rect 1802 7849 1809 7860
rect 1861 7890 1868 7901
rect 2202 7901 2268 7902
rect 2202 7890 2209 7901
rect 1861 7860 2209 7890
rect 1861 7849 1868 7860
rect 1802 7848 1868 7849
rect 2202 7849 2209 7860
rect 2261 7890 2268 7901
rect 2602 7901 2668 7902
rect 2602 7890 2609 7901
rect 2261 7860 2609 7890
rect 2261 7849 2268 7860
rect 2202 7848 2268 7849
rect 2602 7849 2609 7860
rect 2661 7890 2668 7901
rect 3002 7901 3068 7902
rect 3002 7890 3009 7901
rect 2661 7860 3009 7890
rect 2661 7849 2668 7860
rect 2602 7848 2668 7849
rect 3002 7849 3009 7860
rect 3061 7890 3068 7901
rect 3402 7901 3468 7902
rect 3402 7890 3409 7901
rect 3061 7860 3409 7890
rect 3061 7849 3068 7860
rect 3002 7848 3068 7849
rect 3402 7849 3409 7860
rect 3461 7890 3468 7901
rect 3802 7901 3868 7902
rect 3802 7890 3809 7901
rect 3461 7860 3809 7890
rect 3461 7849 3468 7860
rect 3402 7848 3468 7849
rect 3802 7849 3809 7860
rect 3861 7890 3868 7901
rect 4202 7901 4268 7902
rect 4202 7890 4209 7901
rect 3861 7860 4209 7890
rect 3861 7849 3868 7860
rect 3802 7848 3868 7849
rect 4202 7849 4209 7860
rect 4261 7890 4268 7901
rect 4602 7901 4668 7902
rect 4602 7890 4609 7901
rect 4261 7860 4609 7890
rect 4261 7849 4268 7860
rect 4202 7848 4268 7849
rect 4602 7849 4609 7860
rect 4661 7890 4668 7901
rect 5002 7901 5068 7902
rect 5002 7890 5009 7901
rect 4661 7860 5009 7890
rect 4661 7849 4668 7860
rect 4602 7848 4668 7849
rect 5002 7849 5009 7860
rect 5061 7890 5068 7901
rect 5402 7901 5468 7902
rect 5402 7890 5409 7901
rect 5061 7860 5409 7890
rect 5061 7849 5068 7860
rect 5002 7848 5068 7849
rect 5402 7849 5409 7860
rect 5461 7890 5468 7901
rect 5802 7901 5868 7902
rect 5802 7890 5809 7901
rect 5461 7860 5809 7890
rect 5461 7849 5468 7860
rect 5402 7848 5468 7849
rect 5802 7849 5809 7860
rect 5861 7890 5868 7901
rect 6202 7901 6268 7902
rect 6202 7890 6209 7901
rect 5861 7860 6209 7890
rect 5861 7849 5868 7860
rect 5802 7848 5868 7849
rect 6202 7849 6209 7860
rect 6261 7890 6268 7901
rect 6704 7901 6770 7902
rect 6704 7890 6711 7901
rect 6261 7860 6711 7890
rect 6261 7849 6268 7860
rect 6202 7848 6268 7849
rect 6704 7849 6711 7860
rect 6763 7849 6770 7901
rect 6704 7848 6770 7849
rect 2 7831 68 7832
rect 2 7820 9 7831
rect 0 7790 9 7820
rect 2 7779 9 7790
rect 61 7820 68 7831
rect 402 7831 468 7832
rect 402 7820 409 7831
rect 61 7790 409 7820
rect 61 7779 68 7790
rect 2 7778 68 7779
rect 402 7779 409 7790
rect 461 7820 468 7831
rect 802 7831 868 7832
rect 802 7820 809 7831
rect 461 7790 809 7820
rect 461 7779 468 7790
rect 402 7778 468 7779
rect 802 7779 809 7790
rect 861 7820 868 7831
rect 1202 7831 1268 7832
rect 1202 7820 1209 7831
rect 861 7790 1209 7820
rect 861 7779 868 7790
rect 802 7778 868 7779
rect 1202 7779 1209 7790
rect 1261 7820 1268 7831
rect 1602 7831 1668 7832
rect 1602 7820 1609 7831
rect 1261 7790 1609 7820
rect 1261 7779 1268 7790
rect 1202 7778 1268 7779
rect 1602 7779 1609 7790
rect 1661 7820 1668 7831
rect 2002 7831 2068 7832
rect 2002 7820 2009 7831
rect 1661 7790 2009 7820
rect 1661 7779 1668 7790
rect 1602 7778 1668 7779
rect 2002 7779 2009 7790
rect 2061 7820 2068 7831
rect 2402 7831 2468 7832
rect 2402 7820 2409 7831
rect 2061 7790 2409 7820
rect 2061 7779 2068 7790
rect 2002 7778 2068 7779
rect 2402 7779 2409 7790
rect 2461 7820 2468 7831
rect 2802 7831 2868 7832
rect 2802 7820 2809 7831
rect 2461 7790 2809 7820
rect 2461 7779 2468 7790
rect 2402 7778 2468 7779
rect 2802 7779 2809 7790
rect 2861 7820 2868 7831
rect 3202 7831 3268 7832
rect 3202 7820 3209 7831
rect 2861 7790 3209 7820
rect 2861 7779 2868 7790
rect 2802 7778 2868 7779
rect 3202 7779 3209 7790
rect 3261 7820 3268 7831
rect 3602 7831 3668 7832
rect 3602 7820 3609 7831
rect 3261 7790 3609 7820
rect 3261 7779 3268 7790
rect 3202 7778 3268 7779
rect 3602 7779 3609 7790
rect 3661 7820 3668 7831
rect 4002 7831 4068 7832
rect 4002 7820 4009 7831
rect 3661 7790 4009 7820
rect 3661 7779 3668 7790
rect 3602 7778 3668 7779
rect 4002 7779 4009 7790
rect 4061 7820 4068 7831
rect 4402 7831 4468 7832
rect 4402 7820 4409 7831
rect 4061 7790 4409 7820
rect 4061 7779 4068 7790
rect 4002 7778 4068 7779
rect 4402 7779 4409 7790
rect 4461 7820 4468 7831
rect 4802 7831 4868 7832
rect 4802 7820 4809 7831
rect 4461 7790 4809 7820
rect 4461 7779 4468 7790
rect 4402 7778 4468 7779
rect 4802 7779 4809 7790
rect 4861 7820 4868 7831
rect 5202 7831 5268 7832
rect 5202 7820 5209 7831
rect 4861 7790 5209 7820
rect 4861 7779 4868 7790
rect 4802 7778 4868 7779
rect 5202 7779 5209 7790
rect 5261 7820 5268 7831
rect 5602 7831 5668 7832
rect 5602 7820 5609 7831
rect 5261 7790 5609 7820
rect 5261 7779 5268 7790
rect 5202 7778 5268 7779
rect 5602 7779 5609 7790
rect 5661 7820 5668 7831
rect 6002 7831 6068 7832
rect 6002 7820 6009 7831
rect 5661 7790 6009 7820
rect 5661 7779 5668 7790
rect 5602 7778 5668 7779
rect 6002 7779 6009 7790
rect 6061 7820 6068 7831
rect 6402 7831 6468 7832
rect 6402 7820 6409 7831
rect 6061 7790 6409 7820
rect 6061 7779 6068 7790
rect 6002 7778 6068 7779
rect 6402 7779 6409 7790
rect 6461 7820 6468 7831
rect 6500 7831 6566 7832
rect 6500 7820 6507 7831
rect 6461 7790 6507 7820
rect 6461 7779 6468 7790
rect 6402 7778 6468 7779
rect 6500 7779 6507 7790
rect 6559 7779 6566 7831
rect 6500 7778 6566 7779
rect 202 7761 268 7762
rect 202 7750 209 7761
rect 0 7720 209 7750
rect 202 7709 209 7720
rect 261 7750 268 7761
rect 602 7761 668 7762
rect 602 7750 609 7761
rect 261 7720 609 7750
rect 261 7709 268 7720
rect 202 7708 268 7709
rect 602 7709 609 7720
rect 661 7750 668 7761
rect 1002 7761 1068 7762
rect 1002 7750 1009 7761
rect 661 7720 1009 7750
rect 661 7709 668 7720
rect 602 7708 668 7709
rect 1002 7709 1009 7720
rect 1061 7750 1068 7761
rect 1402 7761 1468 7762
rect 1402 7750 1409 7761
rect 1061 7720 1409 7750
rect 1061 7709 1068 7720
rect 1002 7708 1068 7709
rect 1402 7709 1409 7720
rect 1461 7750 1468 7761
rect 1802 7761 1868 7762
rect 1802 7750 1809 7761
rect 1461 7720 1809 7750
rect 1461 7709 1468 7720
rect 1402 7708 1468 7709
rect 1802 7709 1809 7720
rect 1861 7750 1868 7761
rect 2202 7761 2268 7762
rect 2202 7750 2209 7761
rect 1861 7720 2209 7750
rect 1861 7709 1868 7720
rect 1802 7708 1868 7709
rect 2202 7709 2209 7720
rect 2261 7750 2268 7761
rect 2602 7761 2668 7762
rect 2602 7750 2609 7761
rect 2261 7720 2609 7750
rect 2261 7709 2268 7720
rect 2202 7708 2268 7709
rect 2602 7709 2609 7720
rect 2661 7750 2668 7761
rect 3002 7761 3068 7762
rect 3002 7750 3009 7761
rect 2661 7720 3009 7750
rect 2661 7709 2668 7720
rect 2602 7708 2668 7709
rect 3002 7709 3009 7720
rect 3061 7750 3068 7761
rect 3402 7761 3468 7762
rect 3402 7750 3409 7761
rect 3061 7720 3409 7750
rect 3061 7709 3068 7720
rect 3002 7708 3068 7709
rect 3402 7709 3409 7720
rect 3461 7750 3468 7761
rect 3802 7761 3868 7762
rect 3802 7750 3809 7761
rect 3461 7720 3809 7750
rect 3461 7709 3468 7720
rect 3402 7708 3468 7709
rect 3802 7709 3809 7720
rect 3861 7750 3868 7761
rect 4202 7761 4268 7762
rect 4202 7750 4209 7761
rect 3861 7720 4209 7750
rect 3861 7709 3868 7720
rect 3802 7708 3868 7709
rect 4202 7709 4209 7720
rect 4261 7750 4268 7761
rect 4602 7761 4668 7762
rect 4602 7750 4609 7761
rect 4261 7720 4609 7750
rect 4261 7709 4268 7720
rect 4202 7708 4268 7709
rect 4602 7709 4609 7720
rect 4661 7750 4668 7761
rect 5002 7761 5068 7762
rect 5002 7750 5009 7761
rect 4661 7720 5009 7750
rect 4661 7709 4668 7720
rect 4602 7708 4668 7709
rect 5002 7709 5009 7720
rect 5061 7750 5068 7761
rect 5402 7761 5468 7762
rect 5402 7750 5409 7761
rect 5061 7720 5409 7750
rect 5061 7709 5068 7720
rect 5002 7708 5068 7709
rect 5402 7709 5409 7720
rect 5461 7750 5468 7761
rect 5802 7761 5868 7762
rect 5802 7750 5809 7761
rect 5461 7720 5809 7750
rect 5461 7709 5468 7720
rect 5402 7708 5468 7709
rect 5802 7709 5809 7720
rect 5861 7750 5868 7761
rect 6202 7761 6268 7762
rect 6202 7750 6209 7761
rect 5861 7720 6209 7750
rect 5861 7709 5868 7720
rect 5802 7708 5868 7709
rect 6202 7709 6209 7720
rect 6261 7750 6268 7761
rect 6704 7761 6770 7762
rect 6704 7750 6711 7761
rect 6261 7720 6711 7750
rect 6261 7709 6268 7720
rect 6202 7708 6268 7709
rect 6704 7709 6711 7720
rect 6763 7709 6770 7761
rect 6704 7708 6770 7709
rect 2 7691 68 7692
rect 2 7680 9 7691
rect 0 7650 9 7680
rect 2 7639 9 7650
rect 61 7680 68 7691
rect 402 7691 468 7692
rect 402 7680 409 7691
rect 61 7650 409 7680
rect 61 7639 68 7650
rect 2 7638 68 7639
rect 402 7639 409 7650
rect 461 7680 468 7691
rect 802 7691 868 7692
rect 802 7680 809 7691
rect 461 7650 809 7680
rect 461 7639 468 7650
rect 402 7638 468 7639
rect 802 7639 809 7650
rect 861 7680 868 7691
rect 1202 7691 1268 7692
rect 1202 7680 1209 7691
rect 861 7650 1209 7680
rect 861 7639 868 7650
rect 802 7638 868 7639
rect 1202 7639 1209 7650
rect 1261 7680 1268 7691
rect 1602 7691 1668 7692
rect 1602 7680 1609 7691
rect 1261 7650 1609 7680
rect 1261 7639 1268 7650
rect 1202 7638 1268 7639
rect 1602 7639 1609 7650
rect 1661 7680 1668 7691
rect 2002 7691 2068 7692
rect 2002 7680 2009 7691
rect 1661 7650 2009 7680
rect 1661 7639 1668 7650
rect 1602 7638 1668 7639
rect 2002 7639 2009 7650
rect 2061 7680 2068 7691
rect 2402 7691 2468 7692
rect 2402 7680 2409 7691
rect 2061 7650 2409 7680
rect 2061 7639 2068 7650
rect 2002 7638 2068 7639
rect 2402 7639 2409 7650
rect 2461 7680 2468 7691
rect 2802 7691 2868 7692
rect 2802 7680 2809 7691
rect 2461 7650 2809 7680
rect 2461 7639 2468 7650
rect 2402 7638 2468 7639
rect 2802 7639 2809 7650
rect 2861 7680 2868 7691
rect 3202 7691 3268 7692
rect 3202 7680 3209 7691
rect 2861 7650 3209 7680
rect 2861 7639 2868 7650
rect 2802 7638 2868 7639
rect 3202 7639 3209 7650
rect 3261 7680 3268 7691
rect 3602 7691 3668 7692
rect 3602 7680 3609 7691
rect 3261 7650 3609 7680
rect 3261 7639 3268 7650
rect 3202 7638 3268 7639
rect 3602 7639 3609 7650
rect 3661 7680 3668 7691
rect 4002 7691 4068 7692
rect 4002 7680 4009 7691
rect 3661 7650 4009 7680
rect 3661 7639 3668 7650
rect 3602 7638 3668 7639
rect 4002 7639 4009 7650
rect 4061 7680 4068 7691
rect 4402 7691 4468 7692
rect 4402 7680 4409 7691
rect 4061 7650 4409 7680
rect 4061 7639 4068 7650
rect 4002 7638 4068 7639
rect 4402 7639 4409 7650
rect 4461 7680 4468 7691
rect 4802 7691 4868 7692
rect 4802 7680 4809 7691
rect 4461 7650 4809 7680
rect 4461 7639 4468 7650
rect 4402 7638 4468 7639
rect 4802 7639 4809 7650
rect 4861 7680 4868 7691
rect 5202 7691 5268 7692
rect 5202 7680 5209 7691
rect 4861 7650 5209 7680
rect 4861 7639 4868 7650
rect 4802 7638 4868 7639
rect 5202 7639 5209 7650
rect 5261 7680 5268 7691
rect 5602 7691 5668 7692
rect 5602 7680 5609 7691
rect 5261 7650 5609 7680
rect 5261 7639 5268 7650
rect 5202 7638 5268 7639
rect 5602 7639 5609 7650
rect 5661 7680 5668 7691
rect 6002 7691 6068 7692
rect 6002 7680 6009 7691
rect 5661 7650 6009 7680
rect 5661 7639 5668 7650
rect 5602 7638 5668 7639
rect 6002 7639 6009 7650
rect 6061 7680 6068 7691
rect 6402 7691 6468 7692
rect 6402 7680 6409 7691
rect 6061 7650 6409 7680
rect 6061 7639 6068 7650
rect 6002 7638 6068 7639
rect 6402 7639 6409 7650
rect 6461 7680 6468 7691
rect 6500 7691 6566 7692
rect 6500 7680 6507 7691
rect 6461 7650 6507 7680
rect 6461 7639 6468 7650
rect 6402 7638 6468 7639
rect 6500 7639 6507 7650
rect 6559 7639 6566 7691
rect 6500 7638 6566 7639
rect 202 7621 268 7622
rect 202 7610 209 7621
rect 0 7580 209 7610
rect 202 7569 209 7580
rect 261 7610 268 7621
rect 602 7621 668 7622
rect 602 7610 609 7621
rect 261 7580 609 7610
rect 261 7569 268 7580
rect 202 7568 268 7569
rect 602 7569 609 7580
rect 661 7610 668 7621
rect 1002 7621 1068 7622
rect 1002 7610 1009 7621
rect 661 7580 1009 7610
rect 661 7569 668 7580
rect 602 7568 668 7569
rect 1002 7569 1009 7580
rect 1061 7610 1068 7621
rect 1402 7621 1468 7622
rect 1402 7610 1409 7621
rect 1061 7580 1409 7610
rect 1061 7569 1068 7580
rect 1002 7568 1068 7569
rect 1402 7569 1409 7580
rect 1461 7610 1468 7621
rect 1802 7621 1868 7622
rect 1802 7610 1809 7621
rect 1461 7580 1809 7610
rect 1461 7569 1468 7580
rect 1402 7568 1468 7569
rect 1802 7569 1809 7580
rect 1861 7610 1868 7621
rect 2202 7621 2268 7622
rect 2202 7610 2209 7621
rect 1861 7580 2209 7610
rect 1861 7569 1868 7580
rect 1802 7568 1868 7569
rect 2202 7569 2209 7580
rect 2261 7610 2268 7621
rect 2602 7621 2668 7622
rect 2602 7610 2609 7621
rect 2261 7580 2609 7610
rect 2261 7569 2268 7580
rect 2202 7568 2268 7569
rect 2602 7569 2609 7580
rect 2661 7610 2668 7621
rect 3002 7621 3068 7622
rect 3002 7610 3009 7621
rect 2661 7580 3009 7610
rect 2661 7569 2668 7580
rect 2602 7568 2668 7569
rect 3002 7569 3009 7580
rect 3061 7610 3068 7621
rect 3402 7621 3468 7622
rect 3402 7610 3409 7621
rect 3061 7580 3409 7610
rect 3061 7569 3068 7580
rect 3002 7568 3068 7569
rect 3402 7569 3409 7580
rect 3461 7610 3468 7621
rect 3802 7621 3868 7622
rect 3802 7610 3809 7621
rect 3461 7580 3809 7610
rect 3461 7569 3468 7580
rect 3402 7568 3468 7569
rect 3802 7569 3809 7580
rect 3861 7610 3868 7621
rect 4202 7621 4268 7622
rect 4202 7610 4209 7621
rect 3861 7580 4209 7610
rect 3861 7569 3868 7580
rect 3802 7568 3868 7569
rect 4202 7569 4209 7580
rect 4261 7610 4268 7621
rect 4602 7621 4668 7622
rect 4602 7610 4609 7621
rect 4261 7580 4609 7610
rect 4261 7569 4268 7580
rect 4202 7568 4268 7569
rect 4602 7569 4609 7580
rect 4661 7610 4668 7621
rect 5002 7621 5068 7622
rect 5002 7610 5009 7621
rect 4661 7580 5009 7610
rect 4661 7569 4668 7580
rect 4602 7568 4668 7569
rect 5002 7569 5009 7580
rect 5061 7610 5068 7621
rect 5402 7621 5468 7622
rect 5402 7610 5409 7621
rect 5061 7580 5409 7610
rect 5061 7569 5068 7580
rect 5002 7568 5068 7569
rect 5402 7569 5409 7580
rect 5461 7610 5468 7621
rect 5802 7621 5868 7622
rect 5802 7610 5809 7621
rect 5461 7580 5809 7610
rect 5461 7569 5468 7580
rect 5402 7568 5468 7569
rect 5802 7569 5809 7580
rect 5861 7610 5868 7621
rect 6202 7621 6268 7622
rect 6202 7610 6209 7621
rect 5861 7580 6209 7610
rect 5861 7569 5868 7580
rect 5802 7568 5868 7569
rect 6202 7569 6209 7580
rect 6261 7610 6268 7621
rect 6704 7621 6770 7622
rect 6704 7610 6711 7621
rect 6261 7580 6711 7610
rect 6261 7569 6268 7580
rect 6202 7568 6268 7569
rect 6704 7569 6711 7580
rect 6763 7569 6770 7621
rect 6704 7568 6770 7569
rect 2 7551 68 7552
rect 2 7540 9 7551
rect 0 7510 9 7540
rect 2 7499 9 7510
rect 61 7540 68 7551
rect 402 7551 468 7552
rect 402 7540 409 7551
rect 61 7510 409 7540
rect 61 7499 68 7510
rect 2 7498 68 7499
rect 402 7499 409 7510
rect 461 7540 468 7551
rect 802 7551 868 7552
rect 802 7540 809 7551
rect 461 7510 809 7540
rect 461 7499 468 7510
rect 402 7498 468 7499
rect 802 7499 809 7510
rect 861 7540 868 7551
rect 1202 7551 1268 7552
rect 1202 7540 1209 7551
rect 861 7510 1209 7540
rect 861 7499 868 7510
rect 802 7498 868 7499
rect 1202 7499 1209 7510
rect 1261 7540 1268 7551
rect 1602 7551 1668 7552
rect 1602 7540 1609 7551
rect 1261 7510 1609 7540
rect 1261 7499 1268 7510
rect 1202 7498 1268 7499
rect 1602 7499 1609 7510
rect 1661 7540 1668 7551
rect 2002 7551 2068 7552
rect 2002 7540 2009 7551
rect 1661 7510 2009 7540
rect 1661 7499 1668 7510
rect 1602 7498 1668 7499
rect 2002 7499 2009 7510
rect 2061 7540 2068 7551
rect 2402 7551 2468 7552
rect 2402 7540 2409 7551
rect 2061 7510 2409 7540
rect 2061 7499 2068 7510
rect 2002 7498 2068 7499
rect 2402 7499 2409 7510
rect 2461 7540 2468 7551
rect 2802 7551 2868 7552
rect 2802 7540 2809 7551
rect 2461 7510 2809 7540
rect 2461 7499 2468 7510
rect 2402 7498 2468 7499
rect 2802 7499 2809 7510
rect 2861 7540 2868 7551
rect 3202 7551 3268 7552
rect 3202 7540 3209 7551
rect 2861 7510 3209 7540
rect 2861 7499 2868 7510
rect 2802 7498 2868 7499
rect 3202 7499 3209 7510
rect 3261 7540 3268 7551
rect 3602 7551 3668 7552
rect 3602 7540 3609 7551
rect 3261 7510 3609 7540
rect 3261 7499 3268 7510
rect 3202 7498 3268 7499
rect 3602 7499 3609 7510
rect 3661 7540 3668 7551
rect 4002 7551 4068 7552
rect 4002 7540 4009 7551
rect 3661 7510 4009 7540
rect 3661 7499 3668 7510
rect 3602 7498 3668 7499
rect 4002 7499 4009 7510
rect 4061 7540 4068 7551
rect 4402 7551 4468 7552
rect 4402 7540 4409 7551
rect 4061 7510 4409 7540
rect 4061 7499 4068 7510
rect 4002 7498 4068 7499
rect 4402 7499 4409 7510
rect 4461 7540 4468 7551
rect 4802 7551 4868 7552
rect 4802 7540 4809 7551
rect 4461 7510 4809 7540
rect 4461 7499 4468 7510
rect 4402 7498 4468 7499
rect 4802 7499 4809 7510
rect 4861 7540 4868 7551
rect 5202 7551 5268 7552
rect 5202 7540 5209 7551
rect 4861 7510 5209 7540
rect 4861 7499 4868 7510
rect 4802 7498 4868 7499
rect 5202 7499 5209 7510
rect 5261 7540 5268 7551
rect 5602 7551 5668 7552
rect 5602 7540 5609 7551
rect 5261 7510 5609 7540
rect 5261 7499 5268 7510
rect 5202 7498 5268 7499
rect 5602 7499 5609 7510
rect 5661 7540 5668 7551
rect 6002 7551 6068 7552
rect 6002 7540 6009 7551
rect 5661 7510 6009 7540
rect 5661 7499 5668 7510
rect 5602 7498 5668 7499
rect 6002 7499 6009 7510
rect 6061 7540 6068 7551
rect 6402 7551 6468 7552
rect 6402 7540 6409 7551
rect 6061 7510 6409 7540
rect 6061 7499 6068 7510
rect 6002 7498 6068 7499
rect 6402 7499 6409 7510
rect 6461 7540 6468 7551
rect 6500 7551 6566 7552
rect 6500 7540 6507 7551
rect 6461 7510 6507 7540
rect 6461 7499 6468 7510
rect 6402 7498 6468 7499
rect 6500 7499 6507 7510
rect 6559 7499 6566 7551
rect 6500 7498 6566 7499
rect 196 7481 274 7482
rect -4 7465 74 7466
rect -4 7409 7 7465
rect 63 7409 74 7465
rect 196 7425 207 7481
rect 263 7425 274 7481
rect 596 7481 674 7482
rect 196 7424 274 7425
rect 396 7465 474 7466
rect -4 7408 74 7409
rect 396 7409 407 7465
rect 463 7409 474 7465
rect 596 7425 607 7481
rect 663 7425 674 7481
rect 996 7481 1074 7482
rect 596 7424 674 7425
rect 796 7465 874 7466
rect 396 7408 474 7409
rect 796 7409 807 7465
rect 863 7409 874 7465
rect 996 7425 1007 7481
rect 1063 7425 1074 7481
rect 1396 7481 1474 7482
rect 996 7424 1074 7425
rect 1196 7465 1274 7466
rect 796 7408 874 7409
rect 1196 7409 1207 7465
rect 1263 7409 1274 7465
rect 1396 7425 1407 7481
rect 1463 7425 1474 7481
rect 1796 7481 1874 7482
rect 1396 7424 1474 7425
rect 1596 7465 1674 7466
rect 1196 7408 1274 7409
rect 1596 7409 1607 7465
rect 1663 7409 1674 7465
rect 1796 7425 1807 7481
rect 1863 7425 1874 7481
rect 2196 7481 2274 7482
rect 1796 7424 1874 7425
rect 1996 7465 2074 7466
rect 1596 7408 1674 7409
rect 1996 7409 2007 7465
rect 2063 7409 2074 7465
rect 2196 7425 2207 7481
rect 2263 7425 2274 7481
rect 2596 7481 2674 7482
rect 2196 7424 2274 7425
rect 2396 7465 2474 7466
rect 1996 7408 2074 7409
rect 2396 7409 2407 7465
rect 2463 7409 2474 7465
rect 2596 7425 2607 7481
rect 2663 7425 2674 7481
rect 2996 7481 3074 7482
rect 2596 7424 2674 7425
rect 2796 7465 2874 7466
rect 2396 7408 2474 7409
rect 2796 7409 2807 7465
rect 2863 7409 2874 7465
rect 2996 7425 3007 7481
rect 3063 7425 3074 7481
rect 3396 7481 3474 7482
rect 2996 7424 3074 7425
rect 3196 7465 3274 7466
rect 2796 7408 2874 7409
rect 3196 7409 3207 7465
rect 3263 7409 3274 7465
rect 3396 7425 3407 7481
rect 3463 7425 3474 7481
rect 3796 7481 3874 7482
rect 3396 7424 3474 7425
rect 3596 7465 3674 7466
rect 3196 7408 3274 7409
rect 3596 7409 3607 7465
rect 3663 7409 3674 7465
rect 3796 7425 3807 7481
rect 3863 7425 3874 7481
rect 4196 7481 4274 7482
rect 3796 7424 3874 7425
rect 3996 7465 4074 7466
rect 3596 7408 3674 7409
rect 3996 7409 4007 7465
rect 4063 7409 4074 7465
rect 4196 7425 4207 7481
rect 4263 7425 4274 7481
rect 4596 7481 4674 7482
rect 4196 7424 4274 7425
rect 4396 7465 4474 7466
rect 3996 7408 4074 7409
rect 4396 7409 4407 7465
rect 4463 7409 4474 7465
rect 4596 7425 4607 7481
rect 4663 7425 4674 7481
rect 4996 7481 5074 7482
rect 4596 7424 4674 7425
rect 4796 7465 4874 7466
rect 4396 7408 4474 7409
rect 4796 7409 4807 7465
rect 4863 7409 4874 7465
rect 4996 7425 5007 7481
rect 5063 7425 5074 7481
rect 5396 7481 5474 7482
rect 4996 7424 5074 7425
rect 5196 7465 5274 7466
rect 4796 7408 4874 7409
rect 5196 7409 5207 7465
rect 5263 7409 5274 7465
rect 5396 7425 5407 7481
rect 5463 7425 5474 7481
rect 5796 7481 5874 7482
rect 5396 7424 5474 7425
rect 5596 7465 5674 7466
rect 5196 7408 5274 7409
rect 5596 7409 5607 7465
rect 5663 7409 5674 7465
rect 5796 7425 5807 7481
rect 5863 7425 5874 7481
rect 6196 7481 6274 7482
rect 5796 7424 5874 7425
rect 5996 7465 6074 7466
rect 5596 7408 5674 7409
rect 5996 7409 6007 7465
rect 6063 7409 6074 7465
rect 6196 7425 6207 7481
rect 6263 7425 6274 7481
rect 6196 7424 6274 7425
rect 5996 7408 6074 7409
rect 202 7391 268 7392
rect 202 7380 209 7391
rect 0 7350 209 7380
rect 202 7339 209 7350
rect 261 7380 268 7391
rect 602 7391 668 7392
rect 602 7380 609 7391
rect 261 7350 609 7380
rect 261 7339 268 7350
rect 202 7338 268 7339
rect 602 7339 609 7350
rect 661 7380 668 7391
rect 1002 7391 1068 7392
rect 1002 7380 1009 7391
rect 661 7350 1009 7380
rect 661 7339 668 7350
rect 602 7338 668 7339
rect 1002 7339 1009 7350
rect 1061 7380 1068 7391
rect 1402 7391 1468 7392
rect 1402 7380 1409 7391
rect 1061 7350 1409 7380
rect 1061 7339 1068 7350
rect 1002 7338 1068 7339
rect 1402 7339 1409 7350
rect 1461 7380 1468 7391
rect 1802 7391 1868 7392
rect 1802 7380 1809 7391
rect 1461 7350 1809 7380
rect 1461 7339 1468 7350
rect 1402 7338 1468 7339
rect 1802 7339 1809 7350
rect 1861 7380 1868 7391
rect 2202 7391 2268 7392
rect 2202 7380 2209 7391
rect 1861 7350 2209 7380
rect 1861 7339 1868 7350
rect 1802 7338 1868 7339
rect 2202 7339 2209 7350
rect 2261 7380 2268 7391
rect 2602 7391 2668 7392
rect 2602 7380 2609 7391
rect 2261 7350 2609 7380
rect 2261 7339 2268 7350
rect 2202 7338 2268 7339
rect 2602 7339 2609 7350
rect 2661 7380 2668 7391
rect 3002 7391 3068 7392
rect 3002 7380 3009 7391
rect 2661 7350 3009 7380
rect 2661 7339 2668 7350
rect 2602 7338 2668 7339
rect 3002 7339 3009 7350
rect 3061 7380 3068 7391
rect 3402 7391 3468 7392
rect 3402 7380 3409 7391
rect 3061 7350 3409 7380
rect 3061 7339 3068 7350
rect 3002 7338 3068 7339
rect 3402 7339 3409 7350
rect 3461 7380 3468 7391
rect 3802 7391 3868 7392
rect 3802 7380 3809 7391
rect 3461 7350 3809 7380
rect 3461 7339 3468 7350
rect 3402 7338 3468 7339
rect 3802 7339 3809 7350
rect 3861 7380 3868 7391
rect 4202 7391 4268 7392
rect 4202 7380 4209 7391
rect 3861 7350 4209 7380
rect 3861 7339 3868 7350
rect 3802 7338 3868 7339
rect 4202 7339 4209 7350
rect 4261 7380 4268 7391
rect 4602 7391 4668 7392
rect 4602 7380 4609 7391
rect 4261 7350 4609 7380
rect 4261 7339 4268 7350
rect 4202 7338 4268 7339
rect 4602 7339 4609 7350
rect 4661 7380 4668 7391
rect 5002 7391 5068 7392
rect 5002 7380 5009 7391
rect 4661 7350 5009 7380
rect 4661 7339 4668 7350
rect 4602 7338 4668 7339
rect 5002 7339 5009 7350
rect 5061 7380 5068 7391
rect 5402 7391 5468 7392
rect 5402 7380 5409 7391
rect 5061 7350 5409 7380
rect 5061 7339 5068 7350
rect 5002 7338 5068 7339
rect 5402 7339 5409 7350
rect 5461 7380 5468 7391
rect 5802 7391 5868 7392
rect 5802 7380 5809 7391
rect 5461 7350 5809 7380
rect 5461 7339 5468 7350
rect 5402 7338 5468 7339
rect 5802 7339 5809 7350
rect 5861 7380 5868 7391
rect 6202 7391 6268 7392
rect 6202 7380 6209 7391
rect 5861 7350 6209 7380
rect 5861 7339 5868 7350
rect 5802 7338 5868 7339
rect 6202 7339 6209 7350
rect 6261 7380 6268 7391
rect 6704 7391 6770 7392
rect 6704 7380 6711 7391
rect 6261 7350 6711 7380
rect 6261 7339 6268 7350
rect 6202 7338 6268 7339
rect 6704 7339 6711 7350
rect 6763 7339 6770 7391
rect 6704 7338 6770 7339
rect 2 7321 68 7322
rect 2 7310 9 7321
rect 0 7280 9 7310
rect 2 7269 9 7280
rect 61 7310 68 7321
rect 402 7321 468 7322
rect 402 7310 409 7321
rect 61 7280 409 7310
rect 61 7269 68 7280
rect 2 7268 68 7269
rect 402 7269 409 7280
rect 461 7310 468 7321
rect 802 7321 868 7322
rect 802 7310 809 7321
rect 461 7280 809 7310
rect 461 7269 468 7280
rect 402 7268 468 7269
rect 802 7269 809 7280
rect 861 7310 868 7321
rect 1202 7321 1268 7322
rect 1202 7310 1209 7321
rect 861 7280 1209 7310
rect 861 7269 868 7280
rect 802 7268 868 7269
rect 1202 7269 1209 7280
rect 1261 7310 1268 7321
rect 1602 7321 1668 7322
rect 1602 7310 1609 7321
rect 1261 7280 1609 7310
rect 1261 7269 1268 7280
rect 1202 7268 1268 7269
rect 1602 7269 1609 7280
rect 1661 7310 1668 7321
rect 2002 7321 2068 7322
rect 2002 7310 2009 7321
rect 1661 7280 2009 7310
rect 1661 7269 1668 7280
rect 1602 7268 1668 7269
rect 2002 7269 2009 7280
rect 2061 7310 2068 7321
rect 2402 7321 2468 7322
rect 2402 7310 2409 7321
rect 2061 7280 2409 7310
rect 2061 7269 2068 7280
rect 2002 7268 2068 7269
rect 2402 7269 2409 7280
rect 2461 7310 2468 7321
rect 2802 7321 2868 7322
rect 2802 7310 2809 7321
rect 2461 7280 2809 7310
rect 2461 7269 2468 7280
rect 2402 7268 2468 7269
rect 2802 7269 2809 7280
rect 2861 7310 2868 7321
rect 3202 7321 3268 7322
rect 3202 7310 3209 7321
rect 2861 7280 3209 7310
rect 2861 7269 2868 7280
rect 2802 7268 2868 7269
rect 3202 7269 3209 7280
rect 3261 7310 3268 7321
rect 3602 7321 3668 7322
rect 3602 7310 3609 7321
rect 3261 7280 3609 7310
rect 3261 7269 3268 7280
rect 3202 7268 3268 7269
rect 3602 7269 3609 7280
rect 3661 7310 3668 7321
rect 4002 7321 4068 7322
rect 4002 7310 4009 7321
rect 3661 7280 4009 7310
rect 3661 7269 3668 7280
rect 3602 7268 3668 7269
rect 4002 7269 4009 7280
rect 4061 7310 4068 7321
rect 4402 7321 4468 7322
rect 4402 7310 4409 7321
rect 4061 7280 4409 7310
rect 4061 7269 4068 7280
rect 4002 7268 4068 7269
rect 4402 7269 4409 7280
rect 4461 7310 4468 7321
rect 4802 7321 4868 7322
rect 4802 7310 4809 7321
rect 4461 7280 4809 7310
rect 4461 7269 4468 7280
rect 4402 7268 4468 7269
rect 4802 7269 4809 7280
rect 4861 7310 4868 7321
rect 5202 7321 5268 7322
rect 5202 7310 5209 7321
rect 4861 7280 5209 7310
rect 4861 7269 4868 7280
rect 4802 7268 4868 7269
rect 5202 7269 5209 7280
rect 5261 7310 5268 7321
rect 5602 7321 5668 7322
rect 5602 7310 5609 7321
rect 5261 7280 5609 7310
rect 5261 7269 5268 7280
rect 5202 7268 5268 7269
rect 5602 7269 5609 7280
rect 5661 7310 5668 7321
rect 6002 7321 6068 7322
rect 6002 7310 6009 7321
rect 5661 7280 6009 7310
rect 5661 7269 5668 7280
rect 5602 7268 5668 7269
rect 6002 7269 6009 7280
rect 6061 7310 6068 7321
rect 6402 7321 6468 7322
rect 6402 7310 6409 7321
rect 6061 7280 6409 7310
rect 6061 7269 6068 7280
rect 6002 7268 6068 7269
rect 6402 7269 6409 7280
rect 6461 7310 6468 7321
rect 6500 7321 6566 7322
rect 6500 7310 6507 7321
rect 6461 7280 6507 7310
rect 6461 7269 6468 7280
rect 6402 7268 6468 7269
rect 6500 7269 6507 7280
rect 6559 7269 6566 7321
rect 6500 7268 6566 7269
rect 202 7251 268 7252
rect 202 7240 209 7251
rect 0 7210 209 7240
rect 202 7199 209 7210
rect 261 7240 268 7251
rect 602 7251 668 7252
rect 602 7240 609 7251
rect 261 7210 609 7240
rect 261 7199 268 7210
rect 202 7198 268 7199
rect 602 7199 609 7210
rect 661 7240 668 7251
rect 1002 7251 1068 7252
rect 1002 7240 1009 7251
rect 661 7210 1009 7240
rect 661 7199 668 7210
rect 602 7198 668 7199
rect 1002 7199 1009 7210
rect 1061 7240 1068 7251
rect 1402 7251 1468 7252
rect 1402 7240 1409 7251
rect 1061 7210 1409 7240
rect 1061 7199 1068 7210
rect 1002 7198 1068 7199
rect 1402 7199 1409 7210
rect 1461 7240 1468 7251
rect 1802 7251 1868 7252
rect 1802 7240 1809 7251
rect 1461 7210 1809 7240
rect 1461 7199 1468 7210
rect 1402 7198 1468 7199
rect 1802 7199 1809 7210
rect 1861 7240 1868 7251
rect 2202 7251 2268 7252
rect 2202 7240 2209 7251
rect 1861 7210 2209 7240
rect 1861 7199 1868 7210
rect 1802 7198 1868 7199
rect 2202 7199 2209 7210
rect 2261 7240 2268 7251
rect 2602 7251 2668 7252
rect 2602 7240 2609 7251
rect 2261 7210 2609 7240
rect 2261 7199 2268 7210
rect 2202 7198 2268 7199
rect 2602 7199 2609 7210
rect 2661 7240 2668 7251
rect 3002 7251 3068 7252
rect 3002 7240 3009 7251
rect 2661 7210 3009 7240
rect 2661 7199 2668 7210
rect 2602 7198 2668 7199
rect 3002 7199 3009 7210
rect 3061 7240 3068 7251
rect 3402 7251 3468 7252
rect 3402 7240 3409 7251
rect 3061 7210 3409 7240
rect 3061 7199 3068 7210
rect 3002 7198 3068 7199
rect 3402 7199 3409 7210
rect 3461 7240 3468 7251
rect 3802 7251 3868 7252
rect 3802 7240 3809 7251
rect 3461 7210 3809 7240
rect 3461 7199 3468 7210
rect 3402 7198 3468 7199
rect 3802 7199 3809 7210
rect 3861 7240 3868 7251
rect 4202 7251 4268 7252
rect 4202 7240 4209 7251
rect 3861 7210 4209 7240
rect 3861 7199 3868 7210
rect 3802 7198 3868 7199
rect 4202 7199 4209 7210
rect 4261 7240 4268 7251
rect 4602 7251 4668 7252
rect 4602 7240 4609 7251
rect 4261 7210 4609 7240
rect 4261 7199 4268 7210
rect 4202 7198 4268 7199
rect 4602 7199 4609 7210
rect 4661 7240 4668 7251
rect 5002 7251 5068 7252
rect 5002 7240 5009 7251
rect 4661 7210 5009 7240
rect 4661 7199 4668 7210
rect 4602 7198 4668 7199
rect 5002 7199 5009 7210
rect 5061 7240 5068 7251
rect 5402 7251 5468 7252
rect 5402 7240 5409 7251
rect 5061 7210 5409 7240
rect 5061 7199 5068 7210
rect 5002 7198 5068 7199
rect 5402 7199 5409 7210
rect 5461 7240 5468 7251
rect 5802 7251 5868 7252
rect 5802 7240 5809 7251
rect 5461 7210 5809 7240
rect 5461 7199 5468 7210
rect 5402 7198 5468 7199
rect 5802 7199 5809 7210
rect 5861 7240 5868 7251
rect 6202 7251 6268 7252
rect 6202 7240 6209 7251
rect 5861 7210 6209 7240
rect 5861 7199 5868 7210
rect 5802 7198 5868 7199
rect 6202 7199 6209 7210
rect 6261 7240 6268 7251
rect 6704 7251 6770 7252
rect 6704 7240 6711 7251
rect 6261 7210 6711 7240
rect 6261 7199 6268 7210
rect 6202 7198 6268 7199
rect 6704 7199 6711 7210
rect 6763 7199 6770 7251
rect 6704 7198 6770 7199
rect 2 7181 68 7182
rect 2 7170 9 7181
rect 0 7140 9 7170
rect 2 7129 9 7140
rect 61 7170 68 7181
rect 402 7181 468 7182
rect 402 7170 409 7181
rect 61 7140 409 7170
rect 61 7129 68 7140
rect 2 7128 68 7129
rect 402 7129 409 7140
rect 461 7170 468 7181
rect 802 7181 868 7182
rect 802 7170 809 7181
rect 461 7140 809 7170
rect 461 7129 468 7140
rect 402 7128 468 7129
rect 802 7129 809 7140
rect 861 7170 868 7181
rect 1202 7181 1268 7182
rect 1202 7170 1209 7181
rect 861 7140 1209 7170
rect 861 7129 868 7140
rect 802 7128 868 7129
rect 1202 7129 1209 7140
rect 1261 7170 1268 7181
rect 1602 7181 1668 7182
rect 1602 7170 1609 7181
rect 1261 7140 1609 7170
rect 1261 7129 1268 7140
rect 1202 7128 1268 7129
rect 1602 7129 1609 7140
rect 1661 7170 1668 7181
rect 2002 7181 2068 7182
rect 2002 7170 2009 7181
rect 1661 7140 2009 7170
rect 1661 7129 1668 7140
rect 1602 7128 1668 7129
rect 2002 7129 2009 7140
rect 2061 7170 2068 7181
rect 2402 7181 2468 7182
rect 2402 7170 2409 7181
rect 2061 7140 2409 7170
rect 2061 7129 2068 7140
rect 2002 7128 2068 7129
rect 2402 7129 2409 7140
rect 2461 7170 2468 7181
rect 2802 7181 2868 7182
rect 2802 7170 2809 7181
rect 2461 7140 2809 7170
rect 2461 7129 2468 7140
rect 2402 7128 2468 7129
rect 2802 7129 2809 7140
rect 2861 7170 2868 7181
rect 3202 7181 3268 7182
rect 3202 7170 3209 7181
rect 2861 7140 3209 7170
rect 2861 7129 2868 7140
rect 2802 7128 2868 7129
rect 3202 7129 3209 7140
rect 3261 7170 3268 7181
rect 3602 7181 3668 7182
rect 3602 7170 3609 7181
rect 3261 7140 3609 7170
rect 3261 7129 3268 7140
rect 3202 7128 3268 7129
rect 3602 7129 3609 7140
rect 3661 7170 3668 7181
rect 4002 7181 4068 7182
rect 4002 7170 4009 7181
rect 3661 7140 4009 7170
rect 3661 7129 3668 7140
rect 3602 7128 3668 7129
rect 4002 7129 4009 7140
rect 4061 7170 4068 7181
rect 4402 7181 4468 7182
rect 4402 7170 4409 7181
rect 4061 7140 4409 7170
rect 4061 7129 4068 7140
rect 4002 7128 4068 7129
rect 4402 7129 4409 7140
rect 4461 7170 4468 7181
rect 4802 7181 4868 7182
rect 4802 7170 4809 7181
rect 4461 7140 4809 7170
rect 4461 7129 4468 7140
rect 4402 7128 4468 7129
rect 4802 7129 4809 7140
rect 4861 7170 4868 7181
rect 5202 7181 5268 7182
rect 5202 7170 5209 7181
rect 4861 7140 5209 7170
rect 4861 7129 4868 7140
rect 4802 7128 4868 7129
rect 5202 7129 5209 7140
rect 5261 7170 5268 7181
rect 5602 7181 5668 7182
rect 5602 7170 5609 7181
rect 5261 7140 5609 7170
rect 5261 7129 5268 7140
rect 5202 7128 5268 7129
rect 5602 7129 5609 7140
rect 5661 7170 5668 7181
rect 6002 7181 6068 7182
rect 6002 7170 6009 7181
rect 5661 7140 6009 7170
rect 5661 7129 5668 7140
rect 5602 7128 5668 7129
rect 6002 7129 6009 7140
rect 6061 7170 6068 7181
rect 6402 7181 6468 7182
rect 6402 7170 6409 7181
rect 6061 7140 6409 7170
rect 6061 7129 6068 7140
rect 6002 7128 6068 7129
rect 6402 7129 6409 7140
rect 6461 7170 6468 7181
rect 6500 7181 6566 7182
rect 6500 7170 6507 7181
rect 6461 7140 6507 7170
rect 6461 7129 6468 7140
rect 6402 7128 6468 7129
rect 6500 7129 6507 7140
rect 6559 7129 6566 7181
rect 6500 7128 6566 7129
rect 202 7111 268 7112
rect 202 7100 209 7111
rect 0 7070 209 7100
rect 202 7059 209 7070
rect 261 7100 268 7111
rect 602 7111 668 7112
rect 602 7100 609 7111
rect 261 7070 609 7100
rect 261 7059 268 7070
rect 202 7058 268 7059
rect 602 7059 609 7070
rect 661 7100 668 7111
rect 1002 7111 1068 7112
rect 1002 7100 1009 7111
rect 661 7070 1009 7100
rect 661 7059 668 7070
rect 602 7058 668 7059
rect 1002 7059 1009 7070
rect 1061 7100 1068 7111
rect 1402 7111 1468 7112
rect 1402 7100 1409 7111
rect 1061 7070 1409 7100
rect 1061 7059 1068 7070
rect 1002 7058 1068 7059
rect 1402 7059 1409 7070
rect 1461 7100 1468 7111
rect 1802 7111 1868 7112
rect 1802 7100 1809 7111
rect 1461 7070 1809 7100
rect 1461 7059 1468 7070
rect 1402 7058 1468 7059
rect 1802 7059 1809 7070
rect 1861 7100 1868 7111
rect 2202 7111 2268 7112
rect 2202 7100 2209 7111
rect 1861 7070 2209 7100
rect 1861 7059 1868 7070
rect 1802 7058 1868 7059
rect 2202 7059 2209 7070
rect 2261 7100 2268 7111
rect 2602 7111 2668 7112
rect 2602 7100 2609 7111
rect 2261 7070 2609 7100
rect 2261 7059 2268 7070
rect 2202 7058 2268 7059
rect 2602 7059 2609 7070
rect 2661 7100 2668 7111
rect 3002 7111 3068 7112
rect 3002 7100 3009 7111
rect 2661 7070 3009 7100
rect 2661 7059 2668 7070
rect 2602 7058 2668 7059
rect 3002 7059 3009 7070
rect 3061 7100 3068 7111
rect 3402 7111 3468 7112
rect 3402 7100 3409 7111
rect 3061 7070 3409 7100
rect 3061 7059 3068 7070
rect 3002 7058 3068 7059
rect 3402 7059 3409 7070
rect 3461 7100 3468 7111
rect 3802 7111 3868 7112
rect 3802 7100 3809 7111
rect 3461 7070 3809 7100
rect 3461 7059 3468 7070
rect 3402 7058 3468 7059
rect 3802 7059 3809 7070
rect 3861 7100 3868 7111
rect 4202 7111 4268 7112
rect 4202 7100 4209 7111
rect 3861 7070 4209 7100
rect 3861 7059 3868 7070
rect 3802 7058 3868 7059
rect 4202 7059 4209 7070
rect 4261 7100 4268 7111
rect 4602 7111 4668 7112
rect 4602 7100 4609 7111
rect 4261 7070 4609 7100
rect 4261 7059 4268 7070
rect 4202 7058 4268 7059
rect 4602 7059 4609 7070
rect 4661 7100 4668 7111
rect 5002 7111 5068 7112
rect 5002 7100 5009 7111
rect 4661 7070 5009 7100
rect 4661 7059 4668 7070
rect 4602 7058 4668 7059
rect 5002 7059 5009 7070
rect 5061 7100 5068 7111
rect 5402 7111 5468 7112
rect 5402 7100 5409 7111
rect 5061 7070 5409 7100
rect 5061 7059 5068 7070
rect 5002 7058 5068 7059
rect 5402 7059 5409 7070
rect 5461 7100 5468 7111
rect 5802 7111 5868 7112
rect 5802 7100 5809 7111
rect 5461 7070 5809 7100
rect 5461 7059 5468 7070
rect 5402 7058 5468 7059
rect 5802 7059 5809 7070
rect 5861 7100 5868 7111
rect 6202 7111 6268 7112
rect 6202 7100 6209 7111
rect 5861 7070 6209 7100
rect 5861 7059 5868 7070
rect 5802 7058 5868 7059
rect 6202 7059 6209 7070
rect 6261 7100 6268 7111
rect 6704 7111 6770 7112
rect 6704 7100 6711 7111
rect 6261 7070 6711 7100
rect 6261 7059 6268 7070
rect 6202 7058 6268 7059
rect 6704 7059 6711 7070
rect 6763 7059 6770 7111
rect 6704 7058 6770 7059
rect 2 7041 68 7042
rect 2 7030 9 7041
rect 0 7000 9 7030
rect 2 6989 9 7000
rect 61 7030 68 7041
rect 402 7041 468 7042
rect 402 7030 409 7041
rect 61 7000 409 7030
rect 61 6989 68 7000
rect 2 6988 68 6989
rect 402 6989 409 7000
rect 461 7030 468 7041
rect 802 7041 868 7042
rect 802 7030 809 7041
rect 461 7000 809 7030
rect 461 6989 468 7000
rect 402 6988 468 6989
rect 802 6989 809 7000
rect 861 7030 868 7041
rect 1202 7041 1268 7042
rect 1202 7030 1209 7041
rect 861 7000 1209 7030
rect 861 6989 868 7000
rect 802 6988 868 6989
rect 1202 6989 1209 7000
rect 1261 7030 1268 7041
rect 1602 7041 1668 7042
rect 1602 7030 1609 7041
rect 1261 7000 1609 7030
rect 1261 6989 1268 7000
rect 1202 6988 1268 6989
rect 1602 6989 1609 7000
rect 1661 7030 1668 7041
rect 2002 7041 2068 7042
rect 2002 7030 2009 7041
rect 1661 7000 2009 7030
rect 1661 6989 1668 7000
rect 1602 6988 1668 6989
rect 2002 6989 2009 7000
rect 2061 7030 2068 7041
rect 2402 7041 2468 7042
rect 2402 7030 2409 7041
rect 2061 7000 2409 7030
rect 2061 6989 2068 7000
rect 2002 6988 2068 6989
rect 2402 6989 2409 7000
rect 2461 7030 2468 7041
rect 2802 7041 2868 7042
rect 2802 7030 2809 7041
rect 2461 7000 2809 7030
rect 2461 6989 2468 7000
rect 2402 6988 2468 6989
rect 2802 6989 2809 7000
rect 2861 7030 2868 7041
rect 3202 7041 3268 7042
rect 3202 7030 3209 7041
rect 2861 7000 3209 7030
rect 2861 6989 2868 7000
rect 2802 6988 2868 6989
rect 3202 6989 3209 7000
rect 3261 7030 3268 7041
rect 3602 7041 3668 7042
rect 3602 7030 3609 7041
rect 3261 7000 3609 7030
rect 3261 6989 3268 7000
rect 3202 6988 3268 6989
rect 3602 6989 3609 7000
rect 3661 7030 3668 7041
rect 4002 7041 4068 7042
rect 4002 7030 4009 7041
rect 3661 7000 4009 7030
rect 3661 6989 3668 7000
rect 3602 6988 3668 6989
rect 4002 6989 4009 7000
rect 4061 7030 4068 7041
rect 4402 7041 4468 7042
rect 4402 7030 4409 7041
rect 4061 7000 4409 7030
rect 4061 6989 4068 7000
rect 4002 6988 4068 6989
rect 4402 6989 4409 7000
rect 4461 7030 4468 7041
rect 4802 7041 4868 7042
rect 4802 7030 4809 7041
rect 4461 7000 4809 7030
rect 4461 6989 4468 7000
rect 4402 6988 4468 6989
rect 4802 6989 4809 7000
rect 4861 7030 4868 7041
rect 5202 7041 5268 7042
rect 5202 7030 5209 7041
rect 4861 7000 5209 7030
rect 4861 6989 4868 7000
rect 4802 6988 4868 6989
rect 5202 6989 5209 7000
rect 5261 7030 5268 7041
rect 5602 7041 5668 7042
rect 5602 7030 5609 7041
rect 5261 7000 5609 7030
rect 5261 6989 5268 7000
rect 5202 6988 5268 6989
rect 5602 6989 5609 7000
rect 5661 7030 5668 7041
rect 6002 7041 6068 7042
rect 6002 7030 6009 7041
rect 5661 7000 6009 7030
rect 5661 6989 5668 7000
rect 5602 6988 5668 6989
rect 6002 6989 6009 7000
rect 6061 7030 6068 7041
rect 6402 7041 6468 7042
rect 6402 7030 6409 7041
rect 6061 7000 6409 7030
rect 6061 6989 6068 7000
rect 6002 6988 6068 6989
rect 6402 6989 6409 7000
rect 6461 7030 6468 7041
rect 6500 7041 6566 7042
rect 6500 7030 6507 7041
rect 6461 7000 6507 7030
rect 6461 6989 6468 7000
rect 6402 6988 6468 6989
rect 6500 6989 6507 7000
rect 6559 6989 6566 7041
rect 6500 6988 6566 6989
rect 202 6971 268 6972
rect 202 6960 209 6971
rect 0 6930 209 6960
rect 202 6919 209 6930
rect 261 6960 268 6971
rect 602 6971 668 6972
rect 602 6960 609 6971
rect 261 6930 609 6960
rect 261 6919 268 6930
rect 202 6918 268 6919
rect 602 6919 609 6930
rect 661 6960 668 6971
rect 1002 6971 1068 6972
rect 1002 6960 1009 6971
rect 661 6930 1009 6960
rect 661 6919 668 6930
rect 602 6918 668 6919
rect 1002 6919 1009 6930
rect 1061 6960 1068 6971
rect 1402 6971 1468 6972
rect 1402 6960 1409 6971
rect 1061 6930 1409 6960
rect 1061 6919 1068 6930
rect 1002 6918 1068 6919
rect 1402 6919 1409 6930
rect 1461 6960 1468 6971
rect 1802 6971 1868 6972
rect 1802 6960 1809 6971
rect 1461 6930 1809 6960
rect 1461 6919 1468 6930
rect 1402 6918 1468 6919
rect 1802 6919 1809 6930
rect 1861 6960 1868 6971
rect 2202 6971 2268 6972
rect 2202 6960 2209 6971
rect 1861 6930 2209 6960
rect 1861 6919 1868 6930
rect 1802 6918 1868 6919
rect 2202 6919 2209 6930
rect 2261 6960 2268 6971
rect 2602 6971 2668 6972
rect 2602 6960 2609 6971
rect 2261 6930 2609 6960
rect 2261 6919 2268 6930
rect 2202 6918 2268 6919
rect 2602 6919 2609 6930
rect 2661 6960 2668 6971
rect 3002 6971 3068 6972
rect 3002 6960 3009 6971
rect 2661 6930 3009 6960
rect 2661 6919 2668 6930
rect 2602 6918 2668 6919
rect 3002 6919 3009 6930
rect 3061 6960 3068 6971
rect 3402 6971 3468 6972
rect 3402 6960 3409 6971
rect 3061 6930 3409 6960
rect 3061 6919 3068 6930
rect 3002 6918 3068 6919
rect 3402 6919 3409 6930
rect 3461 6960 3468 6971
rect 3802 6971 3868 6972
rect 3802 6960 3809 6971
rect 3461 6930 3809 6960
rect 3461 6919 3468 6930
rect 3402 6918 3468 6919
rect 3802 6919 3809 6930
rect 3861 6960 3868 6971
rect 4202 6971 4268 6972
rect 4202 6960 4209 6971
rect 3861 6930 4209 6960
rect 3861 6919 3868 6930
rect 3802 6918 3868 6919
rect 4202 6919 4209 6930
rect 4261 6960 4268 6971
rect 4602 6971 4668 6972
rect 4602 6960 4609 6971
rect 4261 6930 4609 6960
rect 4261 6919 4268 6930
rect 4202 6918 4268 6919
rect 4602 6919 4609 6930
rect 4661 6960 4668 6971
rect 5002 6971 5068 6972
rect 5002 6960 5009 6971
rect 4661 6930 5009 6960
rect 4661 6919 4668 6930
rect 4602 6918 4668 6919
rect 5002 6919 5009 6930
rect 5061 6960 5068 6971
rect 5402 6971 5468 6972
rect 5402 6960 5409 6971
rect 5061 6930 5409 6960
rect 5061 6919 5068 6930
rect 5002 6918 5068 6919
rect 5402 6919 5409 6930
rect 5461 6960 5468 6971
rect 5802 6971 5868 6972
rect 5802 6960 5809 6971
rect 5461 6930 5809 6960
rect 5461 6919 5468 6930
rect 5402 6918 5468 6919
rect 5802 6919 5809 6930
rect 5861 6960 5868 6971
rect 6202 6971 6268 6972
rect 6202 6960 6209 6971
rect 5861 6930 6209 6960
rect 5861 6919 5868 6930
rect 5802 6918 5868 6919
rect 6202 6919 6209 6930
rect 6261 6960 6268 6971
rect 6704 6971 6770 6972
rect 6704 6960 6711 6971
rect 6261 6930 6711 6960
rect 6261 6919 6268 6930
rect 6202 6918 6268 6919
rect 6704 6919 6711 6930
rect 6763 6919 6770 6971
rect 6704 6918 6770 6919
rect 2 6901 68 6902
rect 2 6890 9 6901
rect 0 6860 9 6890
rect 2 6849 9 6860
rect 61 6890 68 6901
rect 402 6901 468 6902
rect 402 6890 409 6901
rect 61 6860 409 6890
rect 61 6849 68 6860
rect 2 6848 68 6849
rect 402 6849 409 6860
rect 461 6890 468 6901
rect 802 6901 868 6902
rect 802 6890 809 6901
rect 461 6860 809 6890
rect 461 6849 468 6860
rect 402 6848 468 6849
rect 802 6849 809 6860
rect 861 6890 868 6901
rect 1202 6901 1268 6902
rect 1202 6890 1209 6901
rect 861 6860 1209 6890
rect 861 6849 868 6860
rect 802 6848 868 6849
rect 1202 6849 1209 6860
rect 1261 6890 1268 6901
rect 1602 6901 1668 6902
rect 1602 6890 1609 6901
rect 1261 6860 1609 6890
rect 1261 6849 1268 6860
rect 1202 6848 1268 6849
rect 1602 6849 1609 6860
rect 1661 6890 1668 6901
rect 2002 6901 2068 6902
rect 2002 6890 2009 6901
rect 1661 6860 2009 6890
rect 1661 6849 1668 6860
rect 1602 6848 1668 6849
rect 2002 6849 2009 6860
rect 2061 6890 2068 6901
rect 2402 6901 2468 6902
rect 2402 6890 2409 6901
rect 2061 6860 2409 6890
rect 2061 6849 2068 6860
rect 2002 6848 2068 6849
rect 2402 6849 2409 6860
rect 2461 6890 2468 6901
rect 2802 6901 2868 6902
rect 2802 6890 2809 6901
rect 2461 6860 2809 6890
rect 2461 6849 2468 6860
rect 2402 6848 2468 6849
rect 2802 6849 2809 6860
rect 2861 6890 2868 6901
rect 3202 6901 3268 6902
rect 3202 6890 3209 6901
rect 2861 6860 3209 6890
rect 2861 6849 2868 6860
rect 2802 6848 2868 6849
rect 3202 6849 3209 6860
rect 3261 6890 3268 6901
rect 3602 6901 3668 6902
rect 3602 6890 3609 6901
rect 3261 6860 3609 6890
rect 3261 6849 3268 6860
rect 3202 6848 3268 6849
rect 3602 6849 3609 6860
rect 3661 6890 3668 6901
rect 4002 6901 4068 6902
rect 4002 6890 4009 6901
rect 3661 6860 4009 6890
rect 3661 6849 3668 6860
rect 3602 6848 3668 6849
rect 4002 6849 4009 6860
rect 4061 6890 4068 6901
rect 4402 6901 4468 6902
rect 4402 6890 4409 6901
rect 4061 6860 4409 6890
rect 4061 6849 4068 6860
rect 4002 6848 4068 6849
rect 4402 6849 4409 6860
rect 4461 6890 4468 6901
rect 4802 6901 4868 6902
rect 4802 6890 4809 6901
rect 4461 6860 4809 6890
rect 4461 6849 4468 6860
rect 4402 6848 4468 6849
rect 4802 6849 4809 6860
rect 4861 6890 4868 6901
rect 5202 6901 5268 6902
rect 5202 6890 5209 6901
rect 4861 6860 5209 6890
rect 4861 6849 4868 6860
rect 4802 6848 4868 6849
rect 5202 6849 5209 6860
rect 5261 6890 5268 6901
rect 5602 6901 5668 6902
rect 5602 6890 5609 6901
rect 5261 6860 5609 6890
rect 5261 6849 5268 6860
rect 5202 6848 5268 6849
rect 5602 6849 5609 6860
rect 5661 6890 5668 6901
rect 6002 6901 6068 6902
rect 6002 6890 6009 6901
rect 5661 6860 6009 6890
rect 5661 6849 5668 6860
rect 5602 6848 5668 6849
rect 6002 6849 6009 6860
rect 6061 6890 6068 6901
rect 6402 6901 6468 6902
rect 6402 6890 6409 6901
rect 6061 6860 6409 6890
rect 6061 6849 6068 6860
rect 6002 6848 6068 6849
rect 6402 6849 6409 6860
rect 6461 6890 6468 6901
rect 6500 6901 6566 6902
rect 6500 6890 6507 6901
rect 6461 6860 6507 6890
rect 6461 6849 6468 6860
rect 6402 6848 6468 6849
rect 6500 6849 6507 6860
rect 6559 6849 6566 6901
rect 6500 6848 6566 6849
rect 202 6831 268 6832
rect 202 6820 209 6831
rect 0 6790 209 6820
rect 202 6779 209 6790
rect 261 6820 268 6831
rect 602 6831 668 6832
rect 602 6820 609 6831
rect 261 6790 609 6820
rect 261 6779 268 6790
rect 202 6778 268 6779
rect 602 6779 609 6790
rect 661 6820 668 6831
rect 1002 6831 1068 6832
rect 1002 6820 1009 6831
rect 661 6790 1009 6820
rect 661 6779 668 6790
rect 602 6778 668 6779
rect 1002 6779 1009 6790
rect 1061 6820 1068 6831
rect 1402 6831 1468 6832
rect 1402 6820 1409 6831
rect 1061 6790 1409 6820
rect 1061 6779 1068 6790
rect 1002 6778 1068 6779
rect 1402 6779 1409 6790
rect 1461 6820 1468 6831
rect 1802 6831 1868 6832
rect 1802 6820 1809 6831
rect 1461 6790 1809 6820
rect 1461 6779 1468 6790
rect 1402 6778 1468 6779
rect 1802 6779 1809 6790
rect 1861 6820 1868 6831
rect 2202 6831 2268 6832
rect 2202 6820 2209 6831
rect 1861 6790 2209 6820
rect 1861 6779 1868 6790
rect 1802 6778 1868 6779
rect 2202 6779 2209 6790
rect 2261 6820 2268 6831
rect 2602 6831 2668 6832
rect 2602 6820 2609 6831
rect 2261 6790 2609 6820
rect 2261 6779 2268 6790
rect 2202 6778 2268 6779
rect 2602 6779 2609 6790
rect 2661 6820 2668 6831
rect 3002 6831 3068 6832
rect 3002 6820 3009 6831
rect 2661 6790 3009 6820
rect 2661 6779 2668 6790
rect 2602 6778 2668 6779
rect 3002 6779 3009 6790
rect 3061 6820 3068 6831
rect 3402 6831 3468 6832
rect 3402 6820 3409 6831
rect 3061 6790 3409 6820
rect 3061 6779 3068 6790
rect 3002 6778 3068 6779
rect 3402 6779 3409 6790
rect 3461 6820 3468 6831
rect 3802 6831 3868 6832
rect 3802 6820 3809 6831
rect 3461 6790 3809 6820
rect 3461 6779 3468 6790
rect 3402 6778 3468 6779
rect 3802 6779 3809 6790
rect 3861 6820 3868 6831
rect 4202 6831 4268 6832
rect 4202 6820 4209 6831
rect 3861 6790 4209 6820
rect 3861 6779 3868 6790
rect 3802 6778 3868 6779
rect 4202 6779 4209 6790
rect 4261 6820 4268 6831
rect 4602 6831 4668 6832
rect 4602 6820 4609 6831
rect 4261 6790 4609 6820
rect 4261 6779 4268 6790
rect 4202 6778 4268 6779
rect 4602 6779 4609 6790
rect 4661 6820 4668 6831
rect 5002 6831 5068 6832
rect 5002 6820 5009 6831
rect 4661 6790 5009 6820
rect 4661 6779 4668 6790
rect 4602 6778 4668 6779
rect 5002 6779 5009 6790
rect 5061 6820 5068 6831
rect 5402 6831 5468 6832
rect 5402 6820 5409 6831
rect 5061 6790 5409 6820
rect 5061 6779 5068 6790
rect 5002 6778 5068 6779
rect 5402 6779 5409 6790
rect 5461 6820 5468 6831
rect 5802 6831 5868 6832
rect 5802 6820 5809 6831
rect 5461 6790 5809 6820
rect 5461 6779 5468 6790
rect 5402 6778 5468 6779
rect 5802 6779 5809 6790
rect 5861 6820 5868 6831
rect 6202 6831 6268 6832
rect 6202 6820 6209 6831
rect 5861 6790 6209 6820
rect 5861 6779 5868 6790
rect 5802 6778 5868 6779
rect 6202 6779 6209 6790
rect 6261 6820 6268 6831
rect 6704 6831 6770 6832
rect 6704 6820 6711 6831
rect 6261 6790 6711 6820
rect 6261 6779 6268 6790
rect 6202 6778 6268 6779
rect 6704 6779 6711 6790
rect 6763 6779 6770 6831
rect 6704 6778 6770 6779
rect 2 6761 68 6762
rect 2 6750 9 6761
rect 0 6720 9 6750
rect 2 6709 9 6720
rect 61 6750 68 6761
rect 402 6761 468 6762
rect 402 6750 409 6761
rect 61 6720 409 6750
rect 61 6709 68 6720
rect 2 6708 68 6709
rect 402 6709 409 6720
rect 461 6750 468 6761
rect 802 6761 868 6762
rect 802 6750 809 6761
rect 461 6720 809 6750
rect 461 6709 468 6720
rect 402 6708 468 6709
rect 802 6709 809 6720
rect 861 6750 868 6761
rect 1202 6761 1268 6762
rect 1202 6750 1209 6761
rect 861 6720 1209 6750
rect 861 6709 868 6720
rect 802 6708 868 6709
rect 1202 6709 1209 6720
rect 1261 6750 1268 6761
rect 1602 6761 1668 6762
rect 1602 6750 1609 6761
rect 1261 6720 1609 6750
rect 1261 6709 1268 6720
rect 1202 6708 1268 6709
rect 1602 6709 1609 6720
rect 1661 6750 1668 6761
rect 2002 6761 2068 6762
rect 2002 6750 2009 6761
rect 1661 6720 2009 6750
rect 1661 6709 1668 6720
rect 1602 6708 1668 6709
rect 2002 6709 2009 6720
rect 2061 6750 2068 6761
rect 2402 6761 2468 6762
rect 2402 6750 2409 6761
rect 2061 6720 2409 6750
rect 2061 6709 2068 6720
rect 2002 6708 2068 6709
rect 2402 6709 2409 6720
rect 2461 6750 2468 6761
rect 2802 6761 2868 6762
rect 2802 6750 2809 6761
rect 2461 6720 2809 6750
rect 2461 6709 2468 6720
rect 2402 6708 2468 6709
rect 2802 6709 2809 6720
rect 2861 6750 2868 6761
rect 3202 6761 3268 6762
rect 3202 6750 3209 6761
rect 2861 6720 3209 6750
rect 2861 6709 2868 6720
rect 2802 6708 2868 6709
rect 3202 6709 3209 6720
rect 3261 6750 3268 6761
rect 3602 6761 3668 6762
rect 3602 6750 3609 6761
rect 3261 6720 3609 6750
rect 3261 6709 3268 6720
rect 3202 6708 3268 6709
rect 3602 6709 3609 6720
rect 3661 6750 3668 6761
rect 4002 6761 4068 6762
rect 4002 6750 4009 6761
rect 3661 6720 4009 6750
rect 3661 6709 3668 6720
rect 3602 6708 3668 6709
rect 4002 6709 4009 6720
rect 4061 6750 4068 6761
rect 4402 6761 4468 6762
rect 4402 6750 4409 6761
rect 4061 6720 4409 6750
rect 4061 6709 4068 6720
rect 4002 6708 4068 6709
rect 4402 6709 4409 6720
rect 4461 6750 4468 6761
rect 4802 6761 4868 6762
rect 4802 6750 4809 6761
rect 4461 6720 4809 6750
rect 4461 6709 4468 6720
rect 4402 6708 4468 6709
rect 4802 6709 4809 6720
rect 4861 6750 4868 6761
rect 5202 6761 5268 6762
rect 5202 6750 5209 6761
rect 4861 6720 5209 6750
rect 4861 6709 4868 6720
rect 4802 6708 4868 6709
rect 5202 6709 5209 6720
rect 5261 6750 5268 6761
rect 5602 6761 5668 6762
rect 5602 6750 5609 6761
rect 5261 6720 5609 6750
rect 5261 6709 5268 6720
rect 5202 6708 5268 6709
rect 5602 6709 5609 6720
rect 5661 6750 5668 6761
rect 6002 6761 6068 6762
rect 6002 6750 6009 6761
rect 5661 6720 6009 6750
rect 5661 6709 5668 6720
rect 5602 6708 5668 6709
rect 6002 6709 6009 6720
rect 6061 6750 6068 6761
rect 6402 6761 6468 6762
rect 6402 6750 6409 6761
rect 6061 6720 6409 6750
rect 6061 6709 6068 6720
rect 6002 6708 6068 6709
rect 6402 6709 6409 6720
rect 6461 6750 6468 6761
rect 6500 6761 6566 6762
rect 6500 6750 6507 6761
rect 6461 6720 6507 6750
rect 6461 6709 6468 6720
rect 6402 6708 6468 6709
rect 6500 6709 6507 6720
rect 6559 6709 6566 6761
rect 6500 6708 6566 6709
rect 202 6691 268 6692
rect 202 6680 209 6691
rect 0 6650 209 6680
rect 202 6639 209 6650
rect 261 6680 268 6691
rect 602 6691 668 6692
rect 602 6680 609 6691
rect 261 6650 609 6680
rect 261 6639 268 6650
rect 202 6638 268 6639
rect 602 6639 609 6650
rect 661 6680 668 6691
rect 1002 6691 1068 6692
rect 1002 6680 1009 6691
rect 661 6650 1009 6680
rect 661 6639 668 6650
rect 602 6638 668 6639
rect 1002 6639 1009 6650
rect 1061 6680 1068 6691
rect 1402 6691 1468 6692
rect 1402 6680 1409 6691
rect 1061 6650 1409 6680
rect 1061 6639 1068 6650
rect 1002 6638 1068 6639
rect 1402 6639 1409 6650
rect 1461 6680 1468 6691
rect 1802 6691 1868 6692
rect 1802 6680 1809 6691
rect 1461 6650 1809 6680
rect 1461 6639 1468 6650
rect 1402 6638 1468 6639
rect 1802 6639 1809 6650
rect 1861 6680 1868 6691
rect 2202 6691 2268 6692
rect 2202 6680 2209 6691
rect 1861 6650 2209 6680
rect 1861 6639 1868 6650
rect 1802 6638 1868 6639
rect 2202 6639 2209 6650
rect 2261 6680 2268 6691
rect 2602 6691 2668 6692
rect 2602 6680 2609 6691
rect 2261 6650 2609 6680
rect 2261 6639 2268 6650
rect 2202 6638 2268 6639
rect 2602 6639 2609 6650
rect 2661 6680 2668 6691
rect 3002 6691 3068 6692
rect 3002 6680 3009 6691
rect 2661 6650 3009 6680
rect 2661 6639 2668 6650
rect 2602 6638 2668 6639
rect 3002 6639 3009 6650
rect 3061 6680 3068 6691
rect 3402 6691 3468 6692
rect 3402 6680 3409 6691
rect 3061 6650 3409 6680
rect 3061 6639 3068 6650
rect 3002 6638 3068 6639
rect 3402 6639 3409 6650
rect 3461 6680 3468 6691
rect 3802 6691 3868 6692
rect 3802 6680 3809 6691
rect 3461 6650 3809 6680
rect 3461 6639 3468 6650
rect 3402 6638 3468 6639
rect 3802 6639 3809 6650
rect 3861 6680 3868 6691
rect 4202 6691 4268 6692
rect 4202 6680 4209 6691
rect 3861 6650 4209 6680
rect 3861 6639 3868 6650
rect 3802 6638 3868 6639
rect 4202 6639 4209 6650
rect 4261 6680 4268 6691
rect 4602 6691 4668 6692
rect 4602 6680 4609 6691
rect 4261 6650 4609 6680
rect 4261 6639 4268 6650
rect 4202 6638 4268 6639
rect 4602 6639 4609 6650
rect 4661 6680 4668 6691
rect 5002 6691 5068 6692
rect 5002 6680 5009 6691
rect 4661 6650 5009 6680
rect 4661 6639 4668 6650
rect 4602 6638 4668 6639
rect 5002 6639 5009 6650
rect 5061 6680 5068 6691
rect 5402 6691 5468 6692
rect 5402 6680 5409 6691
rect 5061 6650 5409 6680
rect 5061 6639 5068 6650
rect 5002 6638 5068 6639
rect 5402 6639 5409 6650
rect 5461 6680 5468 6691
rect 5802 6691 5868 6692
rect 5802 6680 5809 6691
rect 5461 6650 5809 6680
rect 5461 6639 5468 6650
rect 5402 6638 5468 6639
rect 5802 6639 5809 6650
rect 5861 6680 5868 6691
rect 6202 6691 6268 6692
rect 6202 6680 6209 6691
rect 5861 6650 6209 6680
rect 5861 6639 5868 6650
rect 5802 6638 5868 6639
rect 6202 6639 6209 6650
rect 6261 6680 6268 6691
rect 6704 6691 6770 6692
rect 6704 6680 6711 6691
rect 6261 6650 6711 6680
rect 6261 6639 6268 6650
rect 6202 6638 6268 6639
rect 6704 6639 6711 6650
rect 6763 6639 6770 6691
rect 6704 6638 6770 6639
rect 2 6621 68 6622
rect 2 6610 9 6621
rect 0 6580 9 6610
rect 2 6569 9 6580
rect 61 6610 68 6621
rect 402 6621 468 6622
rect 402 6610 409 6621
rect 61 6580 409 6610
rect 61 6569 68 6580
rect 2 6568 68 6569
rect 402 6569 409 6580
rect 461 6610 468 6621
rect 802 6621 868 6622
rect 802 6610 809 6621
rect 461 6580 809 6610
rect 461 6569 468 6580
rect 402 6568 468 6569
rect 802 6569 809 6580
rect 861 6610 868 6621
rect 1202 6621 1268 6622
rect 1202 6610 1209 6621
rect 861 6580 1209 6610
rect 861 6569 868 6580
rect 802 6568 868 6569
rect 1202 6569 1209 6580
rect 1261 6610 1268 6621
rect 1602 6621 1668 6622
rect 1602 6610 1609 6621
rect 1261 6580 1609 6610
rect 1261 6569 1268 6580
rect 1202 6568 1268 6569
rect 1602 6569 1609 6580
rect 1661 6610 1668 6621
rect 2002 6621 2068 6622
rect 2002 6610 2009 6621
rect 1661 6580 2009 6610
rect 1661 6569 1668 6580
rect 1602 6568 1668 6569
rect 2002 6569 2009 6580
rect 2061 6610 2068 6621
rect 2402 6621 2468 6622
rect 2402 6610 2409 6621
rect 2061 6580 2409 6610
rect 2061 6569 2068 6580
rect 2002 6568 2068 6569
rect 2402 6569 2409 6580
rect 2461 6610 2468 6621
rect 2802 6621 2868 6622
rect 2802 6610 2809 6621
rect 2461 6580 2809 6610
rect 2461 6569 2468 6580
rect 2402 6568 2468 6569
rect 2802 6569 2809 6580
rect 2861 6610 2868 6621
rect 3202 6621 3268 6622
rect 3202 6610 3209 6621
rect 2861 6580 3209 6610
rect 2861 6569 2868 6580
rect 2802 6568 2868 6569
rect 3202 6569 3209 6580
rect 3261 6610 3268 6621
rect 3602 6621 3668 6622
rect 3602 6610 3609 6621
rect 3261 6580 3609 6610
rect 3261 6569 3268 6580
rect 3202 6568 3268 6569
rect 3602 6569 3609 6580
rect 3661 6610 3668 6621
rect 4002 6621 4068 6622
rect 4002 6610 4009 6621
rect 3661 6580 4009 6610
rect 3661 6569 3668 6580
rect 3602 6568 3668 6569
rect 4002 6569 4009 6580
rect 4061 6610 4068 6621
rect 4402 6621 4468 6622
rect 4402 6610 4409 6621
rect 4061 6580 4409 6610
rect 4061 6569 4068 6580
rect 4002 6568 4068 6569
rect 4402 6569 4409 6580
rect 4461 6610 4468 6621
rect 4802 6621 4868 6622
rect 4802 6610 4809 6621
rect 4461 6580 4809 6610
rect 4461 6569 4468 6580
rect 4402 6568 4468 6569
rect 4802 6569 4809 6580
rect 4861 6610 4868 6621
rect 5202 6621 5268 6622
rect 5202 6610 5209 6621
rect 4861 6580 5209 6610
rect 4861 6569 4868 6580
rect 4802 6568 4868 6569
rect 5202 6569 5209 6580
rect 5261 6610 5268 6621
rect 5602 6621 5668 6622
rect 5602 6610 5609 6621
rect 5261 6580 5609 6610
rect 5261 6569 5268 6580
rect 5202 6568 5268 6569
rect 5602 6569 5609 6580
rect 5661 6610 5668 6621
rect 6002 6621 6068 6622
rect 6002 6610 6009 6621
rect 5661 6580 6009 6610
rect 5661 6569 5668 6580
rect 5602 6568 5668 6569
rect 6002 6569 6009 6580
rect 6061 6610 6068 6621
rect 6402 6621 6468 6622
rect 6402 6610 6409 6621
rect 6061 6580 6409 6610
rect 6061 6569 6068 6580
rect 6002 6568 6068 6569
rect 6402 6569 6409 6580
rect 6461 6610 6468 6621
rect 6500 6621 6566 6622
rect 6500 6610 6507 6621
rect 6461 6580 6507 6610
rect 6461 6569 6468 6580
rect 6402 6568 6468 6569
rect 6500 6569 6507 6580
rect 6559 6569 6566 6621
rect 6500 6568 6566 6569
rect 202 6551 268 6552
rect 202 6540 209 6551
rect 0 6510 209 6540
rect 202 6499 209 6510
rect 261 6540 268 6551
rect 602 6551 668 6552
rect 602 6540 609 6551
rect 261 6510 609 6540
rect 261 6499 268 6510
rect 202 6498 268 6499
rect 602 6499 609 6510
rect 661 6540 668 6551
rect 1002 6551 1068 6552
rect 1002 6540 1009 6551
rect 661 6510 1009 6540
rect 661 6499 668 6510
rect 602 6498 668 6499
rect 1002 6499 1009 6510
rect 1061 6540 1068 6551
rect 1402 6551 1468 6552
rect 1402 6540 1409 6551
rect 1061 6510 1409 6540
rect 1061 6499 1068 6510
rect 1002 6498 1068 6499
rect 1402 6499 1409 6510
rect 1461 6540 1468 6551
rect 1802 6551 1868 6552
rect 1802 6540 1809 6551
rect 1461 6510 1809 6540
rect 1461 6499 1468 6510
rect 1402 6498 1468 6499
rect 1802 6499 1809 6510
rect 1861 6540 1868 6551
rect 2202 6551 2268 6552
rect 2202 6540 2209 6551
rect 1861 6510 2209 6540
rect 1861 6499 1868 6510
rect 1802 6498 1868 6499
rect 2202 6499 2209 6510
rect 2261 6540 2268 6551
rect 2602 6551 2668 6552
rect 2602 6540 2609 6551
rect 2261 6510 2609 6540
rect 2261 6499 2268 6510
rect 2202 6498 2268 6499
rect 2602 6499 2609 6510
rect 2661 6540 2668 6551
rect 3002 6551 3068 6552
rect 3002 6540 3009 6551
rect 2661 6510 3009 6540
rect 2661 6499 2668 6510
rect 2602 6498 2668 6499
rect 3002 6499 3009 6510
rect 3061 6540 3068 6551
rect 3402 6551 3468 6552
rect 3402 6540 3409 6551
rect 3061 6510 3409 6540
rect 3061 6499 3068 6510
rect 3002 6498 3068 6499
rect 3402 6499 3409 6510
rect 3461 6540 3468 6551
rect 3802 6551 3868 6552
rect 3802 6540 3809 6551
rect 3461 6510 3809 6540
rect 3461 6499 3468 6510
rect 3402 6498 3468 6499
rect 3802 6499 3809 6510
rect 3861 6540 3868 6551
rect 4202 6551 4268 6552
rect 4202 6540 4209 6551
rect 3861 6510 4209 6540
rect 3861 6499 3868 6510
rect 3802 6498 3868 6499
rect 4202 6499 4209 6510
rect 4261 6540 4268 6551
rect 4602 6551 4668 6552
rect 4602 6540 4609 6551
rect 4261 6510 4609 6540
rect 4261 6499 4268 6510
rect 4202 6498 4268 6499
rect 4602 6499 4609 6510
rect 4661 6540 4668 6551
rect 5002 6551 5068 6552
rect 5002 6540 5009 6551
rect 4661 6510 5009 6540
rect 4661 6499 4668 6510
rect 4602 6498 4668 6499
rect 5002 6499 5009 6510
rect 5061 6540 5068 6551
rect 5402 6551 5468 6552
rect 5402 6540 5409 6551
rect 5061 6510 5409 6540
rect 5061 6499 5068 6510
rect 5002 6498 5068 6499
rect 5402 6499 5409 6510
rect 5461 6540 5468 6551
rect 5802 6551 5868 6552
rect 5802 6540 5809 6551
rect 5461 6510 5809 6540
rect 5461 6499 5468 6510
rect 5402 6498 5468 6499
rect 5802 6499 5809 6510
rect 5861 6540 5868 6551
rect 6202 6551 6268 6552
rect 6202 6540 6209 6551
rect 5861 6510 6209 6540
rect 5861 6499 5868 6510
rect 5802 6498 5868 6499
rect 6202 6499 6209 6510
rect 6261 6540 6268 6551
rect 6704 6551 6770 6552
rect 6704 6540 6711 6551
rect 6261 6510 6711 6540
rect 6261 6499 6268 6510
rect 6202 6498 6268 6499
rect 6704 6499 6711 6510
rect 6763 6499 6770 6551
rect 6704 6498 6770 6499
rect 2 6481 68 6482
rect 2 6470 9 6481
rect 0 6440 9 6470
rect 2 6429 9 6440
rect 61 6470 68 6481
rect 402 6481 468 6482
rect 402 6470 409 6481
rect 61 6440 409 6470
rect 61 6429 68 6440
rect 2 6428 68 6429
rect 402 6429 409 6440
rect 461 6470 468 6481
rect 802 6481 868 6482
rect 802 6470 809 6481
rect 461 6440 809 6470
rect 461 6429 468 6440
rect 402 6428 468 6429
rect 802 6429 809 6440
rect 861 6470 868 6481
rect 1202 6481 1268 6482
rect 1202 6470 1209 6481
rect 861 6440 1209 6470
rect 861 6429 868 6440
rect 802 6428 868 6429
rect 1202 6429 1209 6440
rect 1261 6470 1268 6481
rect 1602 6481 1668 6482
rect 1602 6470 1609 6481
rect 1261 6440 1609 6470
rect 1261 6429 1268 6440
rect 1202 6428 1268 6429
rect 1602 6429 1609 6440
rect 1661 6470 1668 6481
rect 2002 6481 2068 6482
rect 2002 6470 2009 6481
rect 1661 6440 2009 6470
rect 1661 6429 1668 6440
rect 1602 6428 1668 6429
rect 2002 6429 2009 6440
rect 2061 6470 2068 6481
rect 2402 6481 2468 6482
rect 2402 6470 2409 6481
rect 2061 6440 2409 6470
rect 2061 6429 2068 6440
rect 2002 6428 2068 6429
rect 2402 6429 2409 6440
rect 2461 6470 2468 6481
rect 2802 6481 2868 6482
rect 2802 6470 2809 6481
rect 2461 6440 2809 6470
rect 2461 6429 2468 6440
rect 2402 6428 2468 6429
rect 2802 6429 2809 6440
rect 2861 6470 2868 6481
rect 3202 6481 3268 6482
rect 3202 6470 3209 6481
rect 2861 6440 3209 6470
rect 2861 6429 2868 6440
rect 2802 6428 2868 6429
rect 3202 6429 3209 6440
rect 3261 6470 3268 6481
rect 3602 6481 3668 6482
rect 3602 6470 3609 6481
rect 3261 6440 3609 6470
rect 3261 6429 3268 6440
rect 3202 6428 3268 6429
rect 3602 6429 3609 6440
rect 3661 6470 3668 6481
rect 4002 6481 4068 6482
rect 4002 6470 4009 6481
rect 3661 6440 4009 6470
rect 3661 6429 3668 6440
rect 3602 6428 3668 6429
rect 4002 6429 4009 6440
rect 4061 6470 4068 6481
rect 4402 6481 4468 6482
rect 4402 6470 4409 6481
rect 4061 6440 4409 6470
rect 4061 6429 4068 6440
rect 4002 6428 4068 6429
rect 4402 6429 4409 6440
rect 4461 6470 4468 6481
rect 4802 6481 4868 6482
rect 4802 6470 4809 6481
rect 4461 6440 4809 6470
rect 4461 6429 4468 6440
rect 4402 6428 4468 6429
rect 4802 6429 4809 6440
rect 4861 6470 4868 6481
rect 5202 6481 5268 6482
rect 5202 6470 5209 6481
rect 4861 6440 5209 6470
rect 4861 6429 4868 6440
rect 4802 6428 4868 6429
rect 5202 6429 5209 6440
rect 5261 6470 5268 6481
rect 5602 6481 5668 6482
rect 5602 6470 5609 6481
rect 5261 6440 5609 6470
rect 5261 6429 5268 6440
rect 5202 6428 5268 6429
rect 5602 6429 5609 6440
rect 5661 6470 5668 6481
rect 6002 6481 6068 6482
rect 6002 6470 6009 6481
rect 5661 6440 6009 6470
rect 5661 6429 5668 6440
rect 5602 6428 5668 6429
rect 6002 6429 6009 6440
rect 6061 6470 6068 6481
rect 6402 6481 6468 6482
rect 6402 6470 6409 6481
rect 6061 6440 6409 6470
rect 6061 6429 6068 6440
rect 6002 6428 6068 6429
rect 6402 6429 6409 6440
rect 6461 6470 6468 6481
rect 6500 6481 6566 6482
rect 6500 6470 6507 6481
rect 6461 6440 6507 6470
rect 6461 6429 6468 6440
rect 6402 6428 6468 6429
rect 6500 6429 6507 6440
rect 6559 6429 6566 6481
rect 6500 6428 6566 6429
rect 202 6411 268 6412
rect 202 6400 209 6411
rect 0 6370 209 6400
rect 202 6359 209 6370
rect 261 6400 268 6411
rect 602 6411 668 6412
rect 602 6400 609 6411
rect 261 6370 609 6400
rect 261 6359 268 6370
rect 202 6358 268 6359
rect 602 6359 609 6370
rect 661 6400 668 6411
rect 1002 6411 1068 6412
rect 1002 6400 1009 6411
rect 661 6370 1009 6400
rect 661 6359 668 6370
rect 602 6358 668 6359
rect 1002 6359 1009 6370
rect 1061 6400 1068 6411
rect 1402 6411 1468 6412
rect 1402 6400 1409 6411
rect 1061 6370 1409 6400
rect 1061 6359 1068 6370
rect 1002 6358 1068 6359
rect 1402 6359 1409 6370
rect 1461 6400 1468 6411
rect 1802 6411 1868 6412
rect 1802 6400 1809 6411
rect 1461 6370 1809 6400
rect 1461 6359 1468 6370
rect 1402 6358 1468 6359
rect 1802 6359 1809 6370
rect 1861 6400 1868 6411
rect 2202 6411 2268 6412
rect 2202 6400 2209 6411
rect 1861 6370 2209 6400
rect 1861 6359 1868 6370
rect 1802 6358 1868 6359
rect 2202 6359 2209 6370
rect 2261 6400 2268 6411
rect 2602 6411 2668 6412
rect 2602 6400 2609 6411
rect 2261 6370 2609 6400
rect 2261 6359 2268 6370
rect 2202 6358 2268 6359
rect 2602 6359 2609 6370
rect 2661 6400 2668 6411
rect 3002 6411 3068 6412
rect 3002 6400 3009 6411
rect 2661 6370 3009 6400
rect 2661 6359 2668 6370
rect 2602 6358 2668 6359
rect 3002 6359 3009 6370
rect 3061 6400 3068 6411
rect 3402 6411 3468 6412
rect 3402 6400 3409 6411
rect 3061 6370 3409 6400
rect 3061 6359 3068 6370
rect 3002 6358 3068 6359
rect 3402 6359 3409 6370
rect 3461 6400 3468 6411
rect 3802 6411 3868 6412
rect 3802 6400 3809 6411
rect 3461 6370 3809 6400
rect 3461 6359 3468 6370
rect 3402 6358 3468 6359
rect 3802 6359 3809 6370
rect 3861 6400 3868 6411
rect 4202 6411 4268 6412
rect 4202 6400 4209 6411
rect 3861 6370 4209 6400
rect 3861 6359 3868 6370
rect 3802 6358 3868 6359
rect 4202 6359 4209 6370
rect 4261 6400 4268 6411
rect 4602 6411 4668 6412
rect 4602 6400 4609 6411
rect 4261 6370 4609 6400
rect 4261 6359 4268 6370
rect 4202 6358 4268 6359
rect 4602 6359 4609 6370
rect 4661 6400 4668 6411
rect 5002 6411 5068 6412
rect 5002 6400 5009 6411
rect 4661 6370 5009 6400
rect 4661 6359 4668 6370
rect 4602 6358 4668 6359
rect 5002 6359 5009 6370
rect 5061 6400 5068 6411
rect 5402 6411 5468 6412
rect 5402 6400 5409 6411
rect 5061 6370 5409 6400
rect 5061 6359 5068 6370
rect 5002 6358 5068 6359
rect 5402 6359 5409 6370
rect 5461 6400 5468 6411
rect 5802 6411 5868 6412
rect 5802 6400 5809 6411
rect 5461 6370 5809 6400
rect 5461 6359 5468 6370
rect 5402 6358 5468 6359
rect 5802 6359 5809 6370
rect 5861 6400 5868 6411
rect 6202 6411 6268 6412
rect 6202 6400 6209 6411
rect 5861 6370 6209 6400
rect 5861 6359 5868 6370
rect 5802 6358 5868 6359
rect 6202 6359 6209 6370
rect 6261 6400 6268 6411
rect 6704 6411 6770 6412
rect 6704 6400 6711 6411
rect 6261 6370 6711 6400
rect 6261 6359 6268 6370
rect 6202 6358 6268 6359
rect 6704 6359 6711 6370
rect 6763 6359 6770 6411
rect 6704 6358 6770 6359
rect 2 6341 68 6342
rect 2 6330 9 6341
rect 0 6300 9 6330
rect 2 6289 9 6300
rect 61 6330 68 6341
rect 402 6341 468 6342
rect 402 6330 409 6341
rect 61 6300 409 6330
rect 61 6289 68 6300
rect 2 6288 68 6289
rect 402 6289 409 6300
rect 461 6330 468 6341
rect 802 6341 868 6342
rect 802 6330 809 6341
rect 461 6300 809 6330
rect 461 6289 468 6300
rect 402 6288 468 6289
rect 802 6289 809 6300
rect 861 6330 868 6341
rect 1202 6341 1268 6342
rect 1202 6330 1209 6341
rect 861 6300 1209 6330
rect 861 6289 868 6300
rect 802 6288 868 6289
rect 1202 6289 1209 6300
rect 1261 6330 1268 6341
rect 1602 6341 1668 6342
rect 1602 6330 1609 6341
rect 1261 6300 1609 6330
rect 1261 6289 1268 6300
rect 1202 6288 1268 6289
rect 1602 6289 1609 6300
rect 1661 6330 1668 6341
rect 2002 6341 2068 6342
rect 2002 6330 2009 6341
rect 1661 6300 2009 6330
rect 1661 6289 1668 6300
rect 1602 6288 1668 6289
rect 2002 6289 2009 6300
rect 2061 6330 2068 6341
rect 2402 6341 2468 6342
rect 2402 6330 2409 6341
rect 2061 6300 2409 6330
rect 2061 6289 2068 6300
rect 2002 6288 2068 6289
rect 2402 6289 2409 6300
rect 2461 6330 2468 6341
rect 2802 6341 2868 6342
rect 2802 6330 2809 6341
rect 2461 6300 2809 6330
rect 2461 6289 2468 6300
rect 2402 6288 2468 6289
rect 2802 6289 2809 6300
rect 2861 6330 2868 6341
rect 3202 6341 3268 6342
rect 3202 6330 3209 6341
rect 2861 6300 3209 6330
rect 2861 6289 2868 6300
rect 2802 6288 2868 6289
rect 3202 6289 3209 6300
rect 3261 6330 3268 6341
rect 3602 6341 3668 6342
rect 3602 6330 3609 6341
rect 3261 6300 3609 6330
rect 3261 6289 3268 6300
rect 3202 6288 3268 6289
rect 3602 6289 3609 6300
rect 3661 6330 3668 6341
rect 4002 6341 4068 6342
rect 4002 6330 4009 6341
rect 3661 6300 4009 6330
rect 3661 6289 3668 6300
rect 3602 6288 3668 6289
rect 4002 6289 4009 6300
rect 4061 6330 4068 6341
rect 4402 6341 4468 6342
rect 4402 6330 4409 6341
rect 4061 6300 4409 6330
rect 4061 6289 4068 6300
rect 4002 6288 4068 6289
rect 4402 6289 4409 6300
rect 4461 6330 4468 6341
rect 4802 6341 4868 6342
rect 4802 6330 4809 6341
rect 4461 6300 4809 6330
rect 4461 6289 4468 6300
rect 4402 6288 4468 6289
rect 4802 6289 4809 6300
rect 4861 6330 4868 6341
rect 5202 6341 5268 6342
rect 5202 6330 5209 6341
rect 4861 6300 5209 6330
rect 4861 6289 4868 6300
rect 4802 6288 4868 6289
rect 5202 6289 5209 6300
rect 5261 6330 5268 6341
rect 5602 6341 5668 6342
rect 5602 6330 5609 6341
rect 5261 6300 5609 6330
rect 5261 6289 5268 6300
rect 5202 6288 5268 6289
rect 5602 6289 5609 6300
rect 5661 6330 5668 6341
rect 6002 6341 6068 6342
rect 6002 6330 6009 6341
rect 5661 6300 6009 6330
rect 5661 6289 5668 6300
rect 5602 6288 5668 6289
rect 6002 6289 6009 6300
rect 6061 6330 6068 6341
rect 6402 6341 6468 6342
rect 6402 6330 6409 6341
rect 6061 6300 6409 6330
rect 6061 6289 6068 6300
rect 6002 6288 6068 6289
rect 6402 6289 6409 6300
rect 6461 6330 6468 6341
rect 6500 6341 6566 6342
rect 6500 6330 6507 6341
rect 6461 6300 6507 6330
rect 6461 6289 6468 6300
rect 6402 6288 6468 6289
rect 6500 6289 6507 6300
rect 6559 6289 6566 6341
rect 6500 6288 6566 6289
rect 196 6271 274 6272
rect -4 6255 74 6256
rect -4 6199 7 6255
rect 63 6199 74 6255
rect 196 6215 207 6271
rect 263 6215 274 6271
rect 596 6271 674 6272
rect 196 6214 274 6215
rect 396 6255 474 6256
rect -4 6198 74 6199
rect 396 6199 407 6255
rect 463 6199 474 6255
rect 596 6215 607 6271
rect 663 6215 674 6271
rect 996 6271 1074 6272
rect 596 6214 674 6215
rect 796 6255 874 6256
rect 396 6198 474 6199
rect 796 6199 807 6255
rect 863 6199 874 6255
rect 996 6215 1007 6271
rect 1063 6215 1074 6271
rect 1396 6271 1474 6272
rect 996 6214 1074 6215
rect 1196 6255 1274 6256
rect 796 6198 874 6199
rect 1196 6199 1207 6255
rect 1263 6199 1274 6255
rect 1396 6215 1407 6271
rect 1463 6215 1474 6271
rect 1796 6271 1874 6272
rect 1396 6214 1474 6215
rect 1596 6255 1674 6256
rect 1196 6198 1274 6199
rect 1596 6199 1607 6255
rect 1663 6199 1674 6255
rect 1796 6215 1807 6271
rect 1863 6215 1874 6271
rect 2196 6271 2274 6272
rect 1796 6214 1874 6215
rect 1996 6255 2074 6256
rect 1596 6198 1674 6199
rect 1996 6199 2007 6255
rect 2063 6199 2074 6255
rect 2196 6215 2207 6271
rect 2263 6215 2274 6271
rect 2596 6271 2674 6272
rect 2196 6214 2274 6215
rect 2396 6255 2474 6256
rect 1996 6198 2074 6199
rect 2396 6199 2407 6255
rect 2463 6199 2474 6255
rect 2596 6215 2607 6271
rect 2663 6215 2674 6271
rect 2996 6271 3074 6272
rect 2596 6214 2674 6215
rect 2796 6255 2874 6256
rect 2396 6198 2474 6199
rect 2796 6199 2807 6255
rect 2863 6199 2874 6255
rect 2996 6215 3007 6271
rect 3063 6215 3074 6271
rect 3396 6271 3474 6272
rect 2996 6214 3074 6215
rect 3196 6255 3274 6256
rect 2796 6198 2874 6199
rect 3196 6199 3207 6255
rect 3263 6199 3274 6255
rect 3396 6215 3407 6271
rect 3463 6215 3474 6271
rect 3796 6271 3874 6272
rect 3396 6214 3474 6215
rect 3596 6255 3674 6256
rect 3196 6198 3274 6199
rect 3596 6199 3607 6255
rect 3663 6199 3674 6255
rect 3796 6215 3807 6271
rect 3863 6215 3874 6271
rect 4196 6271 4274 6272
rect 3796 6214 3874 6215
rect 3996 6255 4074 6256
rect 3596 6198 3674 6199
rect 3996 6199 4007 6255
rect 4063 6199 4074 6255
rect 4196 6215 4207 6271
rect 4263 6215 4274 6271
rect 4596 6271 4674 6272
rect 4196 6214 4274 6215
rect 4396 6255 4474 6256
rect 3996 6198 4074 6199
rect 4396 6199 4407 6255
rect 4463 6199 4474 6255
rect 4596 6215 4607 6271
rect 4663 6215 4674 6271
rect 4996 6271 5074 6272
rect 4596 6214 4674 6215
rect 4796 6255 4874 6256
rect 4396 6198 4474 6199
rect 4796 6199 4807 6255
rect 4863 6199 4874 6255
rect 4996 6215 5007 6271
rect 5063 6215 5074 6271
rect 5396 6271 5474 6272
rect 4996 6214 5074 6215
rect 5196 6255 5274 6256
rect 4796 6198 4874 6199
rect 5196 6199 5207 6255
rect 5263 6199 5274 6255
rect 5396 6215 5407 6271
rect 5463 6215 5474 6271
rect 5796 6271 5874 6272
rect 5396 6214 5474 6215
rect 5596 6255 5674 6256
rect 5196 6198 5274 6199
rect 5596 6199 5607 6255
rect 5663 6199 5674 6255
rect 5796 6215 5807 6271
rect 5863 6215 5874 6271
rect 6196 6271 6274 6272
rect 5796 6214 5874 6215
rect 5996 6255 6074 6256
rect 5596 6198 5674 6199
rect 5996 6199 6007 6255
rect 6063 6199 6074 6255
rect 6196 6215 6207 6271
rect 6263 6215 6274 6271
rect 6196 6214 6274 6215
rect 5996 6198 6074 6199
rect 202 6181 268 6182
rect 202 6170 209 6181
rect 0 6140 209 6170
rect 202 6129 209 6140
rect 261 6170 268 6181
rect 602 6181 668 6182
rect 602 6170 609 6181
rect 261 6140 609 6170
rect 261 6129 268 6140
rect 202 6128 268 6129
rect 602 6129 609 6140
rect 661 6170 668 6181
rect 1002 6181 1068 6182
rect 1002 6170 1009 6181
rect 661 6140 1009 6170
rect 661 6129 668 6140
rect 602 6128 668 6129
rect 1002 6129 1009 6140
rect 1061 6170 1068 6181
rect 1402 6181 1468 6182
rect 1402 6170 1409 6181
rect 1061 6140 1409 6170
rect 1061 6129 1068 6140
rect 1002 6128 1068 6129
rect 1402 6129 1409 6140
rect 1461 6170 1468 6181
rect 1802 6181 1868 6182
rect 1802 6170 1809 6181
rect 1461 6140 1809 6170
rect 1461 6129 1468 6140
rect 1402 6128 1468 6129
rect 1802 6129 1809 6140
rect 1861 6170 1868 6181
rect 2202 6181 2268 6182
rect 2202 6170 2209 6181
rect 1861 6140 2209 6170
rect 1861 6129 1868 6140
rect 1802 6128 1868 6129
rect 2202 6129 2209 6140
rect 2261 6170 2268 6181
rect 2602 6181 2668 6182
rect 2602 6170 2609 6181
rect 2261 6140 2609 6170
rect 2261 6129 2268 6140
rect 2202 6128 2268 6129
rect 2602 6129 2609 6140
rect 2661 6170 2668 6181
rect 3002 6181 3068 6182
rect 3002 6170 3009 6181
rect 2661 6140 3009 6170
rect 2661 6129 2668 6140
rect 2602 6128 2668 6129
rect 3002 6129 3009 6140
rect 3061 6170 3068 6181
rect 3402 6181 3468 6182
rect 3402 6170 3409 6181
rect 3061 6140 3409 6170
rect 3061 6129 3068 6140
rect 3002 6128 3068 6129
rect 3402 6129 3409 6140
rect 3461 6170 3468 6181
rect 3802 6181 3868 6182
rect 3802 6170 3809 6181
rect 3461 6140 3809 6170
rect 3461 6129 3468 6140
rect 3402 6128 3468 6129
rect 3802 6129 3809 6140
rect 3861 6170 3868 6181
rect 4202 6181 4268 6182
rect 4202 6170 4209 6181
rect 3861 6140 4209 6170
rect 3861 6129 3868 6140
rect 3802 6128 3868 6129
rect 4202 6129 4209 6140
rect 4261 6170 4268 6181
rect 4602 6181 4668 6182
rect 4602 6170 4609 6181
rect 4261 6140 4609 6170
rect 4261 6129 4268 6140
rect 4202 6128 4268 6129
rect 4602 6129 4609 6140
rect 4661 6170 4668 6181
rect 5002 6181 5068 6182
rect 5002 6170 5009 6181
rect 4661 6140 5009 6170
rect 4661 6129 4668 6140
rect 4602 6128 4668 6129
rect 5002 6129 5009 6140
rect 5061 6170 5068 6181
rect 5402 6181 5468 6182
rect 5402 6170 5409 6181
rect 5061 6140 5409 6170
rect 5061 6129 5068 6140
rect 5002 6128 5068 6129
rect 5402 6129 5409 6140
rect 5461 6170 5468 6181
rect 5802 6181 5868 6182
rect 5802 6170 5809 6181
rect 5461 6140 5809 6170
rect 5461 6129 5468 6140
rect 5402 6128 5468 6129
rect 5802 6129 5809 6140
rect 5861 6170 5868 6181
rect 6202 6181 6268 6182
rect 6202 6170 6209 6181
rect 5861 6140 6209 6170
rect 5861 6129 5868 6140
rect 5802 6128 5868 6129
rect 6202 6129 6209 6140
rect 6261 6170 6268 6181
rect 6704 6181 6770 6182
rect 6704 6170 6711 6181
rect 6261 6140 6711 6170
rect 6261 6129 6268 6140
rect 6202 6128 6268 6129
rect 6704 6129 6711 6140
rect 6763 6129 6770 6181
rect 6704 6128 6770 6129
rect 2 6111 68 6112
rect 2 6100 9 6111
rect 0 6070 9 6100
rect 2 6059 9 6070
rect 61 6100 68 6111
rect 402 6111 468 6112
rect 402 6100 409 6111
rect 61 6070 409 6100
rect 61 6059 68 6070
rect 2 6058 68 6059
rect 402 6059 409 6070
rect 461 6100 468 6111
rect 802 6111 868 6112
rect 802 6100 809 6111
rect 461 6070 809 6100
rect 461 6059 468 6070
rect 402 6058 468 6059
rect 802 6059 809 6070
rect 861 6100 868 6111
rect 1202 6111 1268 6112
rect 1202 6100 1209 6111
rect 861 6070 1209 6100
rect 861 6059 868 6070
rect 802 6058 868 6059
rect 1202 6059 1209 6070
rect 1261 6100 1268 6111
rect 1602 6111 1668 6112
rect 1602 6100 1609 6111
rect 1261 6070 1609 6100
rect 1261 6059 1268 6070
rect 1202 6058 1268 6059
rect 1602 6059 1609 6070
rect 1661 6100 1668 6111
rect 2002 6111 2068 6112
rect 2002 6100 2009 6111
rect 1661 6070 2009 6100
rect 1661 6059 1668 6070
rect 1602 6058 1668 6059
rect 2002 6059 2009 6070
rect 2061 6100 2068 6111
rect 2402 6111 2468 6112
rect 2402 6100 2409 6111
rect 2061 6070 2409 6100
rect 2061 6059 2068 6070
rect 2002 6058 2068 6059
rect 2402 6059 2409 6070
rect 2461 6100 2468 6111
rect 2802 6111 2868 6112
rect 2802 6100 2809 6111
rect 2461 6070 2809 6100
rect 2461 6059 2468 6070
rect 2402 6058 2468 6059
rect 2802 6059 2809 6070
rect 2861 6100 2868 6111
rect 3202 6111 3268 6112
rect 3202 6100 3209 6111
rect 2861 6070 3209 6100
rect 2861 6059 2868 6070
rect 2802 6058 2868 6059
rect 3202 6059 3209 6070
rect 3261 6100 3268 6111
rect 3602 6111 3668 6112
rect 3602 6100 3609 6111
rect 3261 6070 3609 6100
rect 3261 6059 3268 6070
rect 3202 6058 3268 6059
rect 3602 6059 3609 6070
rect 3661 6100 3668 6111
rect 4002 6111 4068 6112
rect 4002 6100 4009 6111
rect 3661 6070 4009 6100
rect 3661 6059 3668 6070
rect 3602 6058 3668 6059
rect 4002 6059 4009 6070
rect 4061 6100 4068 6111
rect 4402 6111 4468 6112
rect 4402 6100 4409 6111
rect 4061 6070 4409 6100
rect 4061 6059 4068 6070
rect 4002 6058 4068 6059
rect 4402 6059 4409 6070
rect 4461 6100 4468 6111
rect 4802 6111 4868 6112
rect 4802 6100 4809 6111
rect 4461 6070 4809 6100
rect 4461 6059 4468 6070
rect 4402 6058 4468 6059
rect 4802 6059 4809 6070
rect 4861 6100 4868 6111
rect 5202 6111 5268 6112
rect 5202 6100 5209 6111
rect 4861 6070 5209 6100
rect 4861 6059 4868 6070
rect 4802 6058 4868 6059
rect 5202 6059 5209 6070
rect 5261 6100 5268 6111
rect 5602 6111 5668 6112
rect 5602 6100 5609 6111
rect 5261 6070 5609 6100
rect 5261 6059 5268 6070
rect 5202 6058 5268 6059
rect 5602 6059 5609 6070
rect 5661 6100 5668 6111
rect 6002 6111 6068 6112
rect 6002 6100 6009 6111
rect 5661 6070 6009 6100
rect 5661 6059 5668 6070
rect 5602 6058 5668 6059
rect 6002 6059 6009 6070
rect 6061 6100 6068 6111
rect 6402 6111 6468 6112
rect 6402 6100 6409 6111
rect 6061 6070 6409 6100
rect 6061 6059 6068 6070
rect 6002 6058 6068 6059
rect 6402 6059 6409 6070
rect 6461 6100 6468 6111
rect 6500 6111 6566 6112
rect 6500 6100 6507 6111
rect 6461 6070 6507 6100
rect 6461 6059 6468 6070
rect 6402 6058 6468 6059
rect 6500 6059 6507 6070
rect 6559 6059 6566 6111
rect 6500 6058 6566 6059
rect 202 6041 268 6042
rect 202 6030 209 6041
rect 0 6000 209 6030
rect 202 5989 209 6000
rect 261 6030 268 6041
rect 602 6041 668 6042
rect 602 6030 609 6041
rect 261 6000 609 6030
rect 261 5989 268 6000
rect 202 5988 268 5989
rect 602 5989 609 6000
rect 661 6030 668 6041
rect 1002 6041 1068 6042
rect 1002 6030 1009 6041
rect 661 6000 1009 6030
rect 661 5989 668 6000
rect 602 5988 668 5989
rect 1002 5989 1009 6000
rect 1061 6030 1068 6041
rect 1402 6041 1468 6042
rect 1402 6030 1409 6041
rect 1061 6000 1409 6030
rect 1061 5989 1068 6000
rect 1002 5988 1068 5989
rect 1402 5989 1409 6000
rect 1461 6030 1468 6041
rect 1802 6041 1868 6042
rect 1802 6030 1809 6041
rect 1461 6000 1809 6030
rect 1461 5989 1468 6000
rect 1402 5988 1468 5989
rect 1802 5989 1809 6000
rect 1861 6030 1868 6041
rect 2202 6041 2268 6042
rect 2202 6030 2209 6041
rect 1861 6000 2209 6030
rect 1861 5989 1868 6000
rect 1802 5988 1868 5989
rect 2202 5989 2209 6000
rect 2261 6030 2268 6041
rect 2602 6041 2668 6042
rect 2602 6030 2609 6041
rect 2261 6000 2609 6030
rect 2261 5989 2268 6000
rect 2202 5988 2268 5989
rect 2602 5989 2609 6000
rect 2661 6030 2668 6041
rect 3002 6041 3068 6042
rect 3002 6030 3009 6041
rect 2661 6000 3009 6030
rect 2661 5989 2668 6000
rect 2602 5988 2668 5989
rect 3002 5989 3009 6000
rect 3061 6030 3068 6041
rect 3402 6041 3468 6042
rect 3402 6030 3409 6041
rect 3061 6000 3409 6030
rect 3061 5989 3068 6000
rect 3002 5988 3068 5989
rect 3402 5989 3409 6000
rect 3461 6030 3468 6041
rect 3802 6041 3868 6042
rect 3802 6030 3809 6041
rect 3461 6000 3809 6030
rect 3461 5989 3468 6000
rect 3402 5988 3468 5989
rect 3802 5989 3809 6000
rect 3861 6030 3868 6041
rect 4202 6041 4268 6042
rect 4202 6030 4209 6041
rect 3861 6000 4209 6030
rect 3861 5989 3868 6000
rect 3802 5988 3868 5989
rect 4202 5989 4209 6000
rect 4261 6030 4268 6041
rect 4602 6041 4668 6042
rect 4602 6030 4609 6041
rect 4261 6000 4609 6030
rect 4261 5989 4268 6000
rect 4202 5988 4268 5989
rect 4602 5989 4609 6000
rect 4661 6030 4668 6041
rect 5002 6041 5068 6042
rect 5002 6030 5009 6041
rect 4661 6000 5009 6030
rect 4661 5989 4668 6000
rect 4602 5988 4668 5989
rect 5002 5989 5009 6000
rect 5061 6030 5068 6041
rect 5402 6041 5468 6042
rect 5402 6030 5409 6041
rect 5061 6000 5409 6030
rect 5061 5989 5068 6000
rect 5002 5988 5068 5989
rect 5402 5989 5409 6000
rect 5461 6030 5468 6041
rect 5802 6041 5868 6042
rect 5802 6030 5809 6041
rect 5461 6000 5809 6030
rect 5461 5989 5468 6000
rect 5402 5988 5468 5989
rect 5802 5989 5809 6000
rect 5861 6030 5868 6041
rect 6202 6041 6268 6042
rect 6202 6030 6209 6041
rect 5861 6000 6209 6030
rect 5861 5989 5868 6000
rect 5802 5988 5868 5989
rect 6202 5989 6209 6000
rect 6261 6030 6268 6041
rect 6704 6041 6770 6042
rect 6704 6030 6711 6041
rect 6261 6000 6711 6030
rect 6261 5989 6268 6000
rect 6202 5988 6268 5989
rect 6704 5989 6711 6000
rect 6763 5989 6770 6041
rect 6704 5988 6770 5989
rect 2 5971 68 5972
rect 2 5960 9 5971
rect 0 5930 9 5960
rect 2 5919 9 5930
rect 61 5960 68 5971
rect 402 5971 468 5972
rect 402 5960 409 5971
rect 61 5930 409 5960
rect 61 5919 68 5930
rect 2 5918 68 5919
rect 402 5919 409 5930
rect 461 5960 468 5971
rect 802 5971 868 5972
rect 802 5960 809 5971
rect 461 5930 809 5960
rect 461 5919 468 5930
rect 402 5918 468 5919
rect 802 5919 809 5930
rect 861 5960 868 5971
rect 1202 5971 1268 5972
rect 1202 5960 1209 5971
rect 861 5930 1209 5960
rect 861 5919 868 5930
rect 802 5918 868 5919
rect 1202 5919 1209 5930
rect 1261 5960 1268 5971
rect 1602 5971 1668 5972
rect 1602 5960 1609 5971
rect 1261 5930 1609 5960
rect 1261 5919 1268 5930
rect 1202 5918 1268 5919
rect 1602 5919 1609 5930
rect 1661 5960 1668 5971
rect 2002 5971 2068 5972
rect 2002 5960 2009 5971
rect 1661 5930 2009 5960
rect 1661 5919 1668 5930
rect 1602 5918 1668 5919
rect 2002 5919 2009 5930
rect 2061 5960 2068 5971
rect 2402 5971 2468 5972
rect 2402 5960 2409 5971
rect 2061 5930 2409 5960
rect 2061 5919 2068 5930
rect 2002 5918 2068 5919
rect 2402 5919 2409 5930
rect 2461 5960 2468 5971
rect 2802 5971 2868 5972
rect 2802 5960 2809 5971
rect 2461 5930 2809 5960
rect 2461 5919 2468 5930
rect 2402 5918 2468 5919
rect 2802 5919 2809 5930
rect 2861 5960 2868 5971
rect 3202 5971 3268 5972
rect 3202 5960 3209 5971
rect 2861 5930 3209 5960
rect 2861 5919 2868 5930
rect 2802 5918 2868 5919
rect 3202 5919 3209 5930
rect 3261 5960 3268 5971
rect 3602 5971 3668 5972
rect 3602 5960 3609 5971
rect 3261 5930 3609 5960
rect 3261 5919 3268 5930
rect 3202 5918 3268 5919
rect 3602 5919 3609 5930
rect 3661 5960 3668 5971
rect 4002 5971 4068 5972
rect 4002 5960 4009 5971
rect 3661 5930 4009 5960
rect 3661 5919 3668 5930
rect 3602 5918 3668 5919
rect 4002 5919 4009 5930
rect 4061 5960 4068 5971
rect 4402 5971 4468 5972
rect 4402 5960 4409 5971
rect 4061 5930 4409 5960
rect 4061 5919 4068 5930
rect 4002 5918 4068 5919
rect 4402 5919 4409 5930
rect 4461 5960 4468 5971
rect 4802 5971 4868 5972
rect 4802 5960 4809 5971
rect 4461 5930 4809 5960
rect 4461 5919 4468 5930
rect 4402 5918 4468 5919
rect 4802 5919 4809 5930
rect 4861 5960 4868 5971
rect 5202 5971 5268 5972
rect 5202 5960 5209 5971
rect 4861 5930 5209 5960
rect 4861 5919 4868 5930
rect 4802 5918 4868 5919
rect 5202 5919 5209 5930
rect 5261 5960 5268 5971
rect 5602 5971 5668 5972
rect 5602 5960 5609 5971
rect 5261 5930 5609 5960
rect 5261 5919 5268 5930
rect 5202 5918 5268 5919
rect 5602 5919 5609 5930
rect 5661 5960 5668 5971
rect 6002 5971 6068 5972
rect 6002 5960 6009 5971
rect 5661 5930 6009 5960
rect 5661 5919 5668 5930
rect 5602 5918 5668 5919
rect 6002 5919 6009 5930
rect 6061 5960 6068 5971
rect 6402 5971 6468 5972
rect 6402 5960 6409 5971
rect 6061 5930 6409 5960
rect 6061 5919 6068 5930
rect 6002 5918 6068 5919
rect 6402 5919 6409 5930
rect 6461 5960 6468 5971
rect 6500 5971 6566 5972
rect 6500 5960 6507 5971
rect 6461 5930 6507 5960
rect 6461 5919 6468 5930
rect 6402 5918 6468 5919
rect 6500 5919 6507 5930
rect 6559 5919 6566 5971
rect 6500 5918 6566 5919
rect 202 5901 268 5902
rect 202 5890 209 5901
rect 0 5860 209 5890
rect 202 5849 209 5860
rect 261 5890 268 5901
rect 602 5901 668 5902
rect 602 5890 609 5901
rect 261 5860 609 5890
rect 261 5849 268 5860
rect 202 5848 268 5849
rect 602 5849 609 5860
rect 661 5890 668 5901
rect 1002 5901 1068 5902
rect 1002 5890 1009 5901
rect 661 5860 1009 5890
rect 661 5849 668 5860
rect 602 5848 668 5849
rect 1002 5849 1009 5860
rect 1061 5890 1068 5901
rect 1402 5901 1468 5902
rect 1402 5890 1409 5901
rect 1061 5860 1409 5890
rect 1061 5849 1068 5860
rect 1002 5848 1068 5849
rect 1402 5849 1409 5860
rect 1461 5890 1468 5901
rect 1802 5901 1868 5902
rect 1802 5890 1809 5901
rect 1461 5860 1809 5890
rect 1461 5849 1468 5860
rect 1402 5848 1468 5849
rect 1802 5849 1809 5860
rect 1861 5890 1868 5901
rect 2202 5901 2268 5902
rect 2202 5890 2209 5901
rect 1861 5860 2209 5890
rect 1861 5849 1868 5860
rect 1802 5848 1868 5849
rect 2202 5849 2209 5860
rect 2261 5890 2268 5901
rect 2602 5901 2668 5902
rect 2602 5890 2609 5901
rect 2261 5860 2609 5890
rect 2261 5849 2268 5860
rect 2202 5848 2268 5849
rect 2602 5849 2609 5860
rect 2661 5890 2668 5901
rect 3002 5901 3068 5902
rect 3002 5890 3009 5901
rect 2661 5860 3009 5890
rect 2661 5849 2668 5860
rect 2602 5848 2668 5849
rect 3002 5849 3009 5860
rect 3061 5890 3068 5901
rect 3402 5901 3468 5902
rect 3402 5890 3409 5901
rect 3061 5860 3409 5890
rect 3061 5849 3068 5860
rect 3002 5848 3068 5849
rect 3402 5849 3409 5860
rect 3461 5890 3468 5901
rect 3802 5901 3868 5902
rect 3802 5890 3809 5901
rect 3461 5860 3809 5890
rect 3461 5849 3468 5860
rect 3402 5848 3468 5849
rect 3802 5849 3809 5860
rect 3861 5890 3868 5901
rect 4202 5901 4268 5902
rect 4202 5890 4209 5901
rect 3861 5860 4209 5890
rect 3861 5849 3868 5860
rect 3802 5848 3868 5849
rect 4202 5849 4209 5860
rect 4261 5890 4268 5901
rect 4602 5901 4668 5902
rect 4602 5890 4609 5901
rect 4261 5860 4609 5890
rect 4261 5849 4268 5860
rect 4202 5848 4268 5849
rect 4602 5849 4609 5860
rect 4661 5890 4668 5901
rect 5002 5901 5068 5902
rect 5002 5890 5009 5901
rect 4661 5860 5009 5890
rect 4661 5849 4668 5860
rect 4602 5848 4668 5849
rect 5002 5849 5009 5860
rect 5061 5890 5068 5901
rect 5402 5901 5468 5902
rect 5402 5890 5409 5901
rect 5061 5860 5409 5890
rect 5061 5849 5068 5860
rect 5002 5848 5068 5849
rect 5402 5849 5409 5860
rect 5461 5890 5468 5901
rect 5802 5901 5868 5902
rect 5802 5890 5809 5901
rect 5461 5860 5809 5890
rect 5461 5849 5468 5860
rect 5402 5848 5468 5849
rect 5802 5849 5809 5860
rect 5861 5890 5868 5901
rect 6202 5901 6268 5902
rect 6202 5890 6209 5901
rect 5861 5860 6209 5890
rect 5861 5849 5868 5860
rect 5802 5848 5868 5849
rect 6202 5849 6209 5860
rect 6261 5890 6268 5901
rect 6704 5901 6770 5902
rect 6704 5890 6711 5901
rect 6261 5860 6711 5890
rect 6261 5849 6268 5860
rect 6202 5848 6268 5849
rect 6704 5849 6711 5860
rect 6763 5849 6770 5901
rect 6704 5848 6770 5849
rect 2 5831 68 5832
rect 2 5820 9 5831
rect 0 5790 9 5820
rect 2 5779 9 5790
rect 61 5820 68 5831
rect 402 5831 468 5832
rect 402 5820 409 5831
rect 61 5790 409 5820
rect 61 5779 68 5790
rect 2 5778 68 5779
rect 402 5779 409 5790
rect 461 5820 468 5831
rect 802 5831 868 5832
rect 802 5820 809 5831
rect 461 5790 809 5820
rect 461 5779 468 5790
rect 402 5778 468 5779
rect 802 5779 809 5790
rect 861 5820 868 5831
rect 1202 5831 1268 5832
rect 1202 5820 1209 5831
rect 861 5790 1209 5820
rect 861 5779 868 5790
rect 802 5778 868 5779
rect 1202 5779 1209 5790
rect 1261 5820 1268 5831
rect 1602 5831 1668 5832
rect 1602 5820 1609 5831
rect 1261 5790 1609 5820
rect 1261 5779 1268 5790
rect 1202 5778 1268 5779
rect 1602 5779 1609 5790
rect 1661 5820 1668 5831
rect 2002 5831 2068 5832
rect 2002 5820 2009 5831
rect 1661 5790 2009 5820
rect 1661 5779 1668 5790
rect 1602 5778 1668 5779
rect 2002 5779 2009 5790
rect 2061 5820 2068 5831
rect 2402 5831 2468 5832
rect 2402 5820 2409 5831
rect 2061 5790 2409 5820
rect 2061 5779 2068 5790
rect 2002 5778 2068 5779
rect 2402 5779 2409 5790
rect 2461 5820 2468 5831
rect 2802 5831 2868 5832
rect 2802 5820 2809 5831
rect 2461 5790 2809 5820
rect 2461 5779 2468 5790
rect 2402 5778 2468 5779
rect 2802 5779 2809 5790
rect 2861 5820 2868 5831
rect 3202 5831 3268 5832
rect 3202 5820 3209 5831
rect 2861 5790 3209 5820
rect 2861 5779 2868 5790
rect 2802 5778 2868 5779
rect 3202 5779 3209 5790
rect 3261 5820 3268 5831
rect 3602 5831 3668 5832
rect 3602 5820 3609 5831
rect 3261 5790 3609 5820
rect 3261 5779 3268 5790
rect 3202 5778 3268 5779
rect 3602 5779 3609 5790
rect 3661 5820 3668 5831
rect 4002 5831 4068 5832
rect 4002 5820 4009 5831
rect 3661 5790 4009 5820
rect 3661 5779 3668 5790
rect 3602 5778 3668 5779
rect 4002 5779 4009 5790
rect 4061 5820 4068 5831
rect 4402 5831 4468 5832
rect 4402 5820 4409 5831
rect 4061 5790 4409 5820
rect 4061 5779 4068 5790
rect 4002 5778 4068 5779
rect 4402 5779 4409 5790
rect 4461 5820 4468 5831
rect 4802 5831 4868 5832
rect 4802 5820 4809 5831
rect 4461 5790 4809 5820
rect 4461 5779 4468 5790
rect 4402 5778 4468 5779
rect 4802 5779 4809 5790
rect 4861 5820 4868 5831
rect 5202 5831 5268 5832
rect 5202 5820 5209 5831
rect 4861 5790 5209 5820
rect 4861 5779 4868 5790
rect 4802 5778 4868 5779
rect 5202 5779 5209 5790
rect 5261 5820 5268 5831
rect 5602 5831 5668 5832
rect 5602 5820 5609 5831
rect 5261 5790 5609 5820
rect 5261 5779 5268 5790
rect 5202 5778 5268 5779
rect 5602 5779 5609 5790
rect 5661 5820 5668 5831
rect 6002 5831 6068 5832
rect 6002 5820 6009 5831
rect 5661 5790 6009 5820
rect 5661 5779 5668 5790
rect 5602 5778 5668 5779
rect 6002 5779 6009 5790
rect 6061 5820 6068 5831
rect 6402 5831 6468 5832
rect 6402 5820 6409 5831
rect 6061 5790 6409 5820
rect 6061 5779 6068 5790
rect 6002 5778 6068 5779
rect 6402 5779 6409 5790
rect 6461 5820 6468 5831
rect 6500 5831 6566 5832
rect 6500 5820 6507 5831
rect 6461 5790 6507 5820
rect 6461 5779 6468 5790
rect 6402 5778 6468 5779
rect 6500 5779 6507 5790
rect 6559 5779 6566 5831
rect 6500 5778 6566 5779
rect 202 5761 268 5762
rect 202 5750 209 5761
rect 0 5720 209 5750
rect 202 5709 209 5720
rect 261 5750 268 5761
rect 602 5761 668 5762
rect 602 5750 609 5761
rect 261 5720 609 5750
rect 261 5709 268 5720
rect 202 5708 268 5709
rect 602 5709 609 5720
rect 661 5750 668 5761
rect 1002 5761 1068 5762
rect 1002 5750 1009 5761
rect 661 5720 1009 5750
rect 661 5709 668 5720
rect 602 5708 668 5709
rect 1002 5709 1009 5720
rect 1061 5750 1068 5761
rect 1402 5761 1468 5762
rect 1402 5750 1409 5761
rect 1061 5720 1409 5750
rect 1061 5709 1068 5720
rect 1002 5708 1068 5709
rect 1402 5709 1409 5720
rect 1461 5750 1468 5761
rect 1802 5761 1868 5762
rect 1802 5750 1809 5761
rect 1461 5720 1809 5750
rect 1461 5709 1468 5720
rect 1402 5708 1468 5709
rect 1802 5709 1809 5720
rect 1861 5750 1868 5761
rect 2202 5761 2268 5762
rect 2202 5750 2209 5761
rect 1861 5720 2209 5750
rect 1861 5709 1868 5720
rect 1802 5708 1868 5709
rect 2202 5709 2209 5720
rect 2261 5750 2268 5761
rect 2602 5761 2668 5762
rect 2602 5750 2609 5761
rect 2261 5720 2609 5750
rect 2261 5709 2268 5720
rect 2202 5708 2268 5709
rect 2602 5709 2609 5720
rect 2661 5750 2668 5761
rect 3002 5761 3068 5762
rect 3002 5750 3009 5761
rect 2661 5720 3009 5750
rect 2661 5709 2668 5720
rect 2602 5708 2668 5709
rect 3002 5709 3009 5720
rect 3061 5750 3068 5761
rect 3402 5761 3468 5762
rect 3402 5750 3409 5761
rect 3061 5720 3409 5750
rect 3061 5709 3068 5720
rect 3002 5708 3068 5709
rect 3402 5709 3409 5720
rect 3461 5750 3468 5761
rect 3802 5761 3868 5762
rect 3802 5750 3809 5761
rect 3461 5720 3809 5750
rect 3461 5709 3468 5720
rect 3402 5708 3468 5709
rect 3802 5709 3809 5720
rect 3861 5750 3868 5761
rect 4202 5761 4268 5762
rect 4202 5750 4209 5761
rect 3861 5720 4209 5750
rect 3861 5709 3868 5720
rect 3802 5708 3868 5709
rect 4202 5709 4209 5720
rect 4261 5750 4268 5761
rect 4602 5761 4668 5762
rect 4602 5750 4609 5761
rect 4261 5720 4609 5750
rect 4261 5709 4268 5720
rect 4202 5708 4268 5709
rect 4602 5709 4609 5720
rect 4661 5750 4668 5761
rect 5002 5761 5068 5762
rect 5002 5750 5009 5761
rect 4661 5720 5009 5750
rect 4661 5709 4668 5720
rect 4602 5708 4668 5709
rect 5002 5709 5009 5720
rect 5061 5750 5068 5761
rect 5402 5761 5468 5762
rect 5402 5750 5409 5761
rect 5061 5720 5409 5750
rect 5061 5709 5068 5720
rect 5002 5708 5068 5709
rect 5402 5709 5409 5720
rect 5461 5750 5468 5761
rect 5802 5761 5868 5762
rect 5802 5750 5809 5761
rect 5461 5720 5809 5750
rect 5461 5709 5468 5720
rect 5402 5708 5468 5709
rect 5802 5709 5809 5720
rect 5861 5750 5868 5761
rect 6202 5761 6268 5762
rect 6202 5750 6209 5761
rect 5861 5720 6209 5750
rect 5861 5709 5868 5720
rect 5802 5708 5868 5709
rect 6202 5709 6209 5720
rect 6261 5750 6268 5761
rect 6704 5761 6770 5762
rect 6704 5750 6711 5761
rect 6261 5720 6711 5750
rect 6261 5709 6268 5720
rect 6202 5708 6268 5709
rect 6704 5709 6711 5720
rect 6763 5709 6770 5761
rect 6704 5708 6770 5709
rect 2 5691 68 5692
rect 2 5680 9 5691
rect 0 5650 9 5680
rect 2 5639 9 5650
rect 61 5680 68 5691
rect 402 5691 468 5692
rect 402 5680 409 5691
rect 61 5650 409 5680
rect 61 5639 68 5650
rect 2 5638 68 5639
rect 402 5639 409 5650
rect 461 5680 468 5691
rect 802 5691 868 5692
rect 802 5680 809 5691
rect 461 5650 809 5680
rect 461 5639 468 5650
rect 402 5638 468 5639
rect 802 5639 809 5650
rect 861 5680 868 5691
rect 1202 5691 1268 5692
rect 1202 5680 1209 5691
rect 861 5650 1209 5680
rect 861 5639 868 5650
rect 802 5638 868 5639
rect 1202 5639 1209 5650
rect 1261 5680 1268 5691
rect 1602 5691 1668 5692
rect 1602 5680 1609 5691
rect 1261 5650 1609 5680
rect 1261 5639 1268 5650
rect 1202 5638 1268 5639
rect 1602 5639 1609 5650
rect 1661 5680 1668 5691
rect 2002 5691 2068 5692
rect 2002 5680 2009 5691
rect 1661 5650 2009 5680
rect 1661 5639 1668 5650
rect 1602 5638 1668 5639
rect 2002 5639 2009 5650
rect 2061 5680 2068 5691
rect 2402 5691 2468 5692
rect 2402 5680 2409 5691
rect 2061 5650 2409 5680
rect 2061 5639 2068 5650
rect 2002 5638 2068 5639
rect 2402 5639 2409 5650
rect 2461 5680 2468 5691
rect 2802 5691 2868 5692
rect 2802 5680 2809 5691
rect 2461 5650 2809 5680
rect 2461 5639 2468 5650
rect 2402 5638 2468 5639
rect 2802 5639 2809 5650
rect 2861 5680 2868 5691
rect 3202 5691 3268 5692
rect 3202 5680 3209 5691
rect 2861 5650 3209 5680
rect 2861 5639 2868 5650
rect 2802 5638 2868 5639
rect 3202 5639 3209 5650
rect 3261 5680 3268 5691
rect 3602 5691 3668 5692
rect 3602 5680 3609 5691
rect 3261 5650 3609 5680
rect 3261 5639 3268 5650
rect 3202 5638 3268 5639
rect 3602 5639 3609 5650
rect 3661 5680 3668 5691
rect 4002 5691 4068 5692
rect 4002 5680 4009 5691
rect 3661 5650 4009 5680
rect 3661 5639 3668 5650
rect 3602 5638 3668 5639
rect 4002 5639 4009 5650
rect 4061 5680 4068 5691
rect 4402 5691 4468 5692
rect 4402 5680 4409 5691
rect 4061 5650 4409 5680
rect 4061 5639 4068 5650
rect 4002 5638 4068 5639
rect 4402 5639 4409 5650
rect 4461 5680 4468 5691
rect 4802 5691 4868 5692
rect 4802 5680 4809 5691
rect 4461 5650 4809 5680
rect 4461 5639 4468 5650
rect 4402 5638 4468 5639
rect 4802 5639 4809 5650
rect 4861 5680 4868 5691
rect 5202 5691 5268 5692
rect 5202 5680 5209 5691
rect 4861 5650 5209 5680
rect 4861 5639 4868 5650
rect 4802 5638 4868 5639
rect 5202 5639 5209 5650
rect 5261 5680 5268 5691
rect 5602 5691 5668 5692
rect 5602 5680 5609 5691
rect 5261 5650 5609 5680
rect 5261 5639 5268 5650
rect 5202 5638 5268 5639
rect 5602 5639 5609 5650
rect 5661 5680 5668 5691
rect 6002 5691 6068 5692
rect 6002 5680 6009 5691
rect 5661 5650 6009 5680
rect 5661 5639 5668 5650
rect 5602 5638 5668 5639
rect 6002 5639 6009 5650
rect 6061 5680 6068 5691
rect 6402 5691 6468 5692
rect 6402 5680 6409 5691
rect 6061 5650 6409 5680
rect 6061 5639 6068 5650
rect 6002 5638 6068 5639
rect 6402 5639 6409 5650
rect 6461 5680 6468 5691
rect 6500 5691 6566 5692
rect 6500 5680 6507 5691
rect 6461 5650 6507 5680
rect 6461 5639 6468 5650
rect 6402 5638 6468 5639
rect 6500 5639 6507 5650
rect 6559 5639 6566 5691
rect 6500 5638 6566 5639
rect 202 5621 268 5622
rect 202 5610 209 5621
rect 0 5580 209 5610
rect 202 5569 209 5580
rect 261 5610 268 5621
rect 602 5621 668 5622
rect 602 5610 609 5621
rect 261 5580 609 5610
rect 261 5569 268 5580
rect 202 5568 268 5569
rect 602 5569 609 5580
rect 661 5610 668 5621
rect 1002 5621 1068 5622
rect 1002 5610 1009 5621
rect 661 5580 1009 5610
rect 661 5569 668 5580
rect 602 5568 668 5569
rect 1002 5569 1009 5580
rect 1061 5610 1068 5621
rect 1402 5621 1468 5622
rect 1402 5610 1409 5621
rect 1061 5580 1409 5610
rect 1061 5569 1068 5580
rect 1002 5568 1068 5569
rect 1402 5569 1409 5580
rect 1461 5610 1468 5621
rect 1802 5621 1868 5622
rect 1802 5610 1809 5621
rect 1461 5580 1809 5610
rect 1461 5569 1468 5580
rect 1402 5568 1468 5569
rect 1802 5569 1809 5580
rect 1861 5610 1868 5621
rect 2202 5621 2268 5622
rect 2202 5610 2209 5621
rect 1861 5580 2209 5610
rect 1861 5569 1868 5580
rect 1802 5568 1868 5569
rect 2202 5569 2209 5580
rect 2261 5610 2268 5621
rect 2602 5621 2668 5622
rect 2602 5610 2609 5621
rect 2261 5580 2609 5610
rect 2261 5569 2268 5580
rect 2202 5568 2268 5569
rect 2602 5569 2609 5580
rect 2661 5610 2668 5621
rect 3002 5621 3068 5622
rect 3002 5610 3009 5621
rect 2661 5580 3009 5610
rect 2661 5569 2668 5580
rect 2602 5568 2668 5569
rect 3002 5569 3009 5580
rect 3061 5610 3068 5621
rect 3402 5621 3468 5622
rect 3402 5610 3409 5621
rect 3061 5580 3409 5610
rect 3061 5569 3068 5580
rect 3002 5568 3068 5569
rect 3402 5569 3409 5580
rect 3461 5610 3468 5621
rect 3802 5621 3868 5622
rect 3802 5610 3809 5621
rect 3461 5580 3809 5610
rect 3461 5569 3468 5580
rect 3402 5568 3468 5569
rect 3802 5569 3809 5580
rect 3861 5610 3868 5621
rect 4202 5621 4268 5622
rect 4202 5610 4209 5621
rect 3861 5580 4209 5610
rect 3861 5569 3868 5580
rect 3802 5568 3868 5569
rect 4202 5569 4209 5580
rect 4261 5610 4268 5621
rect 4602 5621 4668 5622
rect 4602 5610 4609 5621
rect 4261 5580 4609 5610
rect 4261 5569 4268 5580
rect 4202 5568 4268 5569
rect 4602 5569 4609 5580
rect 4661 5610 4668 5621
rect 5002 5621 5068 5622
rect 5002 5610 5009 5621
rect 4661 5580 5009 5610
rect 4661 5569 4668 5580
rect 4602 5568 4668 5569
rect 5002 5569 5009 5580
rect 5061 5610 5068 5621
rect 5402 5621 5468 5622
rect 5402 5610 5409 5621
rect 5061 5580 5409 5610
rect 5061 5569 5068 5580
rect 5002 5568 5068 5569
rect 5402 5569 5409 5580
rect 5461 5610 5468 5621
rect 5802 5621 5868 5622
rect 5802 5610 5809 5621
rect 5461 5580 5809 5610
rect 5461 5569 5468 5580
rect 5402 5568 5468 5569
rect 5802 5569 5809 5580
rect 5861 5610 5868 5621
rect 6202 5621 6268 5622
rect 6202 5610 6209 5621
rect 5861 5580 6209 5610
rect 5861 5569 5868 5580
rect 5802 5568 5868 5569
rect 6202 5569 6209 5580
rect 6261 5610 6268 5621
rect 6704 5621 6770 5622
rect 6704 5610 6711 5621
rect 6261 5580 6711 5610
rect 6261 5569 6268 5580
rect 6202 5568 6268 5569
rect 6704 5569 6711 5580
rect 6763 5569 6770 5621
rect 6704 5568 6770 5569
rect 2 5551 68 5552
rect 2 5540 9 5551
rect 0 5510 9 5540
rect 2 5499 9 5510
rect 61 5540 68 5551
rect 402 5551 468 5552
rect 402 5540 409 5551
rect 61 5510 409 5540
rect 61 5499 68 5510
rect 2 5498 68 5499
rect 402 5499 409 5510
rect 461 5540 468 5551
rect 802 5551 868 5552
rect 802 5540 809 5551
rect 461 5510 809 5540
rect 461 5499 468 5510
rect 402 5498 468 5499
rect 802 5499 809 5510
rect 861 5540 868 5551
rect 1202 5551 1268 5552
rect 1202 5540 1209 5551
rect 861 5510 1209 5540
rect 861 5499 868 5510
rect 802 5498 868 5499
rect 1202 5499 1209 5510
rect 1261 5540 1268 5551
rect 1602 5551 1668 5552
rect 1602 5540 1609 5551
rect 1261 5510 1609 5540
rect 1261 5499 1268 5510
rect 1202 5498 1268 5499
rect 1602 5499 1609 5510
rect 1661 5540 1668 5551
rect 2002 5551 2068 5552
rect 2002 5540 2009 5551
rect 1661 5510 2009 5540
rect 1661 5499 1668 5510
rect 1602 5498 1668 5499
rect 2002 5499 2009 5510
rect 2061 5540 2068 5551
rect 2402 5551 2468 5552
rect 2402 5540 2409 5551
rect 2061 5510 2409 5540
rect 2061 5499 2068 5510
rect 2002 5498 2068 5499
rect 2402 5499 2409 5510
rect 2461 5540 2468 5551
rect 2802 5551 2868 5552
rect 2802 5540 2809 5551
rect 2461 5510 2809 5540
rect 2461 5499 2468 5510
rect 2402 5498 2468 5499
rect 2802 5499 2809 5510
rect 2861 5540 2868 5551
rect 3202 5551 3268 5552
rect 3202 5540 3209 5551
rect 2861 5510 3209 5540
rect 2861 5499 2868 5510
rect 2802 5498 2868 5499
rect 3202 5499 3209 5510
rect 3261 5540 3268 5551
rect 3602 5551 3668 5552
rect 3602 5540 3609 5551
rect 3261 5510 3609 5540
rect 3261 5499 3268 5510
rect 3202 5498 3268 5499
rect 3602 5499 3609 5510
rect 3661 5540 3668 5551
rect 4002 5551 4068 5552
rect 4002 5540 4009 5551
rect 3661 5510 4009 5540
rect 3661 5499 3668 5510
rect 3602 5498 3668 5499
rect 4002 5499 4009 5510
rect 4061 5540 4068 5551
rect 4402 5551 4468 5552
rect 4402 5540 4409 5551
rect 4061 5510 4409 5540
rect 4061 5499 4068 5510
rect 4002 5498 4068 5499
rect 4402 5499 4409 5510
rect 4461 5540 4468 5551
rect 4802 5551 4868 5552
rect 4802 5540 4809 5551
rect 4461 5510 4809 5540
rect 4461 5499 4468 5510
rect 4402 5498 4468 5499
rect 4802 5499 4809 5510
rect 4861 5540 4868 5551
rect 5202 5551 5268 5552
rect 5202 5540 5209 5551
rect 4861 5510 5209 5540
rect 4861 5499 4868 5510
rect 4802 5498 4868 5499
rect 5202 5499 5209 5510
rect 5261 5540 5268 5551
rect 5602 5551 5668 5552
rect 5602 5540 5609 5551
rect 5261 5510 5609 5540
rect 5261 5499 5268 5510
rect 5202 5498 5268 5499
rect 5602 5499 5609 5510
rect 5661 5540 5668 5551
rect 6002 5551 6068 5552
rect 6002 5540 6009 5551
rect 5661 5510 6009 5540
rect 5661 5499 5668 5510
rect 5602 5498 5668 5499
rect 6002 5499 6009 5510
rect 6061 5540 6068 5551
rect 6402 5551 6468 5552
rect 6402 5540 6409 5551
rect 6061 5510 6409 5540
rect 6061 5499 6068 5510
rect 6002 5498 6068 5499
rect 6402 5499 6409 5510
rect 6461 5540 6468 5551
rect 6500 5551 6566 5552
rect 6500 5540 6507 5551
rect 6461 5510 6507 5540
rect 6461 5499 6468 5510
rect 6402 5498 6468 5499
rect 6500 5499 6507 5510
rect 6559 5499 6566 5551
rect 6500 5498 6566 5499
rect 202 5481 268 5482
rect 202 5470 209 5481
rect 0 5440 209 5470
rect 202 5429 209 5440
rect 261 5470 268 5481
rect 602 5481 668 5482
rect 602 5470 609 5481
rect 261 5440 609 5470
rect 261 5429 268 5440
rect 202 5428 268 5429
rect 602 5429 609 5440
rect 661 5470 668 5481
rect 1002 5481 1068 5482
rect 1002 5470 1009 5481
rect 661 5440 1009 5470
rect 661 5429 668 5440
rect 602 5428 668 5429
rect 1002 5429 1009 5440
rect 1061 5470 1068 5481
rect 1402 5481 1468 5482
rect 1402 5470 1409 5481
rect 1061 5440 1409 5470
rect 1061 5429 1068 5440
rect 1002 5428 1068 5429
rect 1402 5429 1409 5440
rect 1461 5470 1468 5481
rect 1802 5481 1868 5482
rect 1802 5470 1809 5481
rect 1461 5440 1809 5470
rect 1461 5429 1468 5440
rect 1402 5428 1468 5429
rect 1802 5429 1809 5440
rect 1861 5470 1868 5481
rect 2202 5481 2268 5482
rect 2202 5470 2209 5481
rect 1861 5440 2209 5470
rect 1861 5429 1868 5440
rect 1802 5428 1868 5429
rect 2202 5429 2209 5440
rect 2261 5470 2268 5481
rect 2602 5481 2668 5482
rect 2602 5470 2609 5481
rect 2261 5440 2609 5470
rect 2261 5429 2268 5440
rect 2202 5428 2268 5429
rect 2602 5429 2609 5440
rect 2661 5470 2668 5481
rect 3002 5481 3068 5482
rect 3002 5470 3009 5481
rect 2661 5440 3009 5470
rect 2661 5429 2668 5440
rect 2602 5428 2668 5429
rect 3002 5429 3009 5440
rect 3061 5470 3068 5481
rect 3402 5481 3468 5482
rect 3402 5470 3409 5481
rect 3061 5440 3409 5470
rect 3061 5429 3068 5440
rect 3002 5428 3068 5429
rect 3402 5429 3409 5440
rect 3461 5470 3468 5481
rect 3802 5481 3868 5482
rect 3802 5470 3809 5481
rect 3461 5440 3809 5470
rect 3461 5429 3468 5440
rect 3402 5428 3468 5429
rect 3802 5429 3809 5440
rect 3861 5470 3868 5481
rect 4202 5481 4268 5482
rect 4202 5470 4209 5481
rect 3861 5440 4209 5470
rect 3861 5429 3868 5440
rect 3802 5428 3868 5429
rect 4202 5429 4209 5440
rect 4261 5470 4268 5481
rect 4602 5481 4668 5482
rect 4602 5470 4609 5481
rect 4261 5440 4609 5470
rect 4261 5429 4268 5440
rect 4202 5428 4268 5429
rect 4602 5429 4609 5440
rect 4661 5470 4668 5481
rect 5002 5481 5068 5482
rect 5002 5470 5009 5481
rect 4661 5440 5009 5470
rect 4661 5429 4668 5440
rect 4602 5428 4668 5429
rect 5002 5429 5009 5440
rect 5061 5470 5068 5481
rect 5402 5481 5468 5482
rect 5402 5470 5409 5481
rect 5061 5440 5409 5470
rect 5061 5429 5068 5440
rect 5002 5428 5068 5429
rect 5402 5429 5409 5440
rect 5461 5470 5468 5481
rect 5802 5481 5868 5482
rect 5802 5470 5809 5481
rect 5461 5440 5809 5470
rect 5461 5429 5468 5440
rect 5402 5428 5468 5429
rect 5802 5429 5809 5440
rect 5861 5470 5868 5481
rect 6202 5481 6268 5482
rect 6202 5470 6209 5481
rect 5861 5440 6209 5470
rect 5861 5429 5868 5440
rect 5802 5428 5868 5429
rect 6202 5429 6209 5440
rect 6261 5470 6268 5481
rect 6704 5481 6770 5482
rect 6704 5470 6711 5481
rect 6261 5440 6711 5470
rect 6261 5429 6268 5440
rect 6202 5428 6268 5429
rect 6704 5429 6711 5440
rect 6763 5429 6770 5481
rect 6704 5428 6770 5429
rect 2 5411 68 5412
rect 2 5400 9 5411
rect 0 5370 9 5400
rect 2 5359 9 5370
rect 61 5400 68 5411
rect 402 5411 468 5412
rect 402 5400 409 5411
rect 61 5370 409 5400
rect 61 5359 68 5370
rect 2 5358 68 5359
rect 402 5359 409 5370
rect 461 5400 468 5411
rect 802 5411 868 5412
rect 802 5400 809 5411
rect 461 5370 809 5400
rect 461 5359 468 5370
rect 402 5358 468 5359
rect 802 5359 809 5370
rect 861 5400 868 5411
rect 1202 5411 1268 5412
rect 1202 5400 1209 5411
rect 861 5370 1209 5400
rect 861 5359 868 5370
rect 802 5358 868 5359
rect 1202 5359 1209 5370
rect 1261 5400 1268 5411
rect 1602 5411 1668 5412
rect 1602 5400 1609 5411
rect 1261 5370 1609 5400
rect 1261 5359 1268 5370
rect 1202 5358 1268 5359
rect 1602 5359 1609 5370
rect 1661 5400 1668 5411
rect 2002 5411 2068 5412
rect 2002 5400 2009 5411
rect 1661 5370 2009 5400
rect 1661 5359 1668 5370
rect 1602 5358 1668 5359
rect 2002 5359 2009 5370
rect 2061 5400 2068 5411
rect 2402 5411 2468 5412
rect 2402 5400 2409 5411
rect 2061 5370 2409 5400
rect 2061 5359 2068 5370
rect 2002 5358 2068 5359
rect 2402 5359 2409 5370
rect 2461 5400 2468 5411
rect 2802 5411 2868 5412
rect 2802 5400 2809 5411
rect 2461 5370 2809 5400
rect 2461 5359 2468 5370
rect 2402 5358 2468 5359
rect 2802 5359 2809 5370
rect 2861 5400 2868 5411
rect 3202 5411 3268 5412
rect 3202 5400 3209 5411
rect 2861 5370 3209 5400
rect 2861 5359 2868 5370
rect 2802 5358 2868 5359
rect 3202 5359 3209 5370
rect 3261 5400 3268 5411
rect 3602 5411 3668 5412
rect 3602 5400 3609 5411
rect 3261 5370 3609 5400
rect 3261 5359 3268 5370
rect 3202 5358 3268 5359
rect 3602 5359 3609 5370
rect 3661 5400 3668 5411
rect 4002 5411 4068 5412
rect 4002 5400 4009 5411
rect 3661 5370 4009 5400
rect 3661 5359 3668 5370
rect 3602 5358 3668 5359
rect 4002 5359 4009 5370
rect 4061 5400 4068 5411
rect 4402 5411 4468 5412
rect 4402 5400 4409 5411
rect 4061 5370 4409 5400
rect 4061 5359 4068 5370
rect 4002 5358 4068 5359
rect 4402 5359 4409 5370
rect 4461 5400 4468 5411
rect 4802 5411 4868 5412
rect 4802 5400 4809 5411
rect 4461 5370 4809 5400
rect 4461 5359 4468 5370
rect 4402 5358 4468 5359
rect 4802 5359 4809 5370
rect 4861 5400 4868 5411
rect 5202 5411 5268 5412
rect 5202 5400 5209 5411
rect 4861 5370 5209 5400
rect 4861 5359 4868 5370
rect 4802 5358 4868 5359
rect 5202 5359 5209 5370
rect 5261 5400 5268 5411
rect 5602 5411 5668 5412
rect 5602 5400 5609 5411
rect 5261 5370 5609 5400
rect 5261 5359 5268 5370
rect 5202 5358 5268 5359
rect 5602 5359 5609 5370
rect 5661 5400 5668 5411
rect 6002 5411 6068 5412
rect 6002 5400 6009 5411
rect 5661 5370 6009 5400
rect 5661 5359 5668 5370
rect 5602 5358 5668 5359
rect 6002 5359 6009 5370
rect 6061 5400 6068 5411
rect 6402 5411 6468 5412
rect 6402 5400 6409 5411
rect 6061 5370 6409 5400
rect 6061 5359 6068 5370
rect 6002 5358 6068 5359
rect 6402 5359 6409 5370
rect 6461 5400 6468 5411
rect 6500 5411 6566 5412
rect 6500 5400 6507 5411
rect 6461 5370 6507 5400
rect 6461 5359 6468 5370
rect 6402 5358 6468 5359
rect 6500 5359 6507 5370
rect 6559 5359 6566 5411
rect 6500 5358 6566 5359
rect 202 5341 268 5342
rect 202 5330 209 5341
rect 0 5300 209 5330
rect 202 5289 209 5300
rect 261 5330 268 5341
rect 602 5341 668 5342
rect 602 5330 609 5341
rect 261 5300 609 5330
rect 261 5289 268 5300
rect 202 5288 268 5289
rect 602 5289 609 5300
rect 661 5330 668 5341
rect 1002 5341 1068 5342
rect 1002 5330 1009 5341
rect 661 5300 1009 5330
rect 661 5289 668 5300
rect 602 5288 668 5289
rect 1002 5289 1009 5300
rect 1061 5330 1068 5341
rect 1402 5341 1468 5342
rect 1402 5330 1409 5341
rect 1061 5300 1409 5330
rect 1061 5289 1068 5300
rect 1002 5288 1068 5289
rect 1402 5289 1409 5300
rect 1461 5330 1468 5341
rect 1802 5341 1868 5342
rect 1802 5330 1809 5341
rect 1461 5300 1809 5330
rect 1461 5289 1468 5300
rect 1402 5288 1468 5289
rect 1802 5289 1809 5300
rect 1861 5330 1868 5341
rect 2202 5341 2268 5342
rect 2202 5330 2209 5341
rect 1861 5300 2209 5330
rect 1861 5289 1868 5300
rect 1802 5288 1868 5289
rect 2202 5289 2209 5300
rect 2261 5330 2268 5341
rect 2602 5341 2668 5342
rect 2602 5330 2609 5341
rect 2261 5300 2609 5330
rect 2261 5289 2268 5300
rect 2202 5288 2268 5289
rect 2602 5289 2609 5300
rect 2661 5330 2668 5341
rect 3002 5341 3068 5342
rect 3002 5330 3009 5341
rect 2661 5300 3009 5330
rect 2661 5289 2668 5300
rect 2602 5288 2668 5289
rect 3002 5289 3009 5300
rect 3061 5330 3068 5341
rect 3402 5341 3468 5342
rect 3402 5330 3409 5341
rect 3061 5300 3409 5330
rect 3061 5289 3068 5300
rect 3002 5288 3068 5289
rect 3402 5289 3409 5300
rect 3461 5330 3468 5341
rect 3802 5341 3868 5342
rect 3802 5330 3809 5341
rect 3461 5300 3809 5330
rect 3461 5289 3468 5300
rect 3402 5288 3468 5289
rect 3802 5289 3809 5300
rect 3861 5330 3868 5341
rect 4202 5341 4268 5342
rect 4202 5330 4209 5341
rect 3861 5300 4209 5330
rect 3861 5289 3868 5300
rect 3802 5288 3868 5289
rect 4202 5289 4209 5300
rect 4261 5330 4268 5341
rect 4602 5341 4668 5342
rect 4602 5330 4609 5341
rect 4261 5300 4609 5330
rect 4261 5289 4268 5300
rect 4202 5288 4268 5289
rect 4602 5289 4609 5300
rect 4661 5330 4668 5341
rect 5002 5341 5068 5342
rect 5002 5330 5009 5341
rect 4661 5300 5009 5330
rect 4661 5289 4668 5300
rect 4602 5288 4668 5289
rect 5002 5289 5009 5300
rect 5061 5330 5068 5341
rect 5402 5341 5468 5342
rect 5402 5330 5409 5341
rect 5061 5300 5409 5330
rect 5061 5289 5068 5300
rect 5002 5288 5068 5289
rect 5402 5289 5409 5300
rect 5461 5330 5468 5341
rect 5802 5341 5868 5342
rect 5802 5330 5809 5341
rect 5461 5300 5809 5330
rect 5461 5289 5468 5300
rect 5402 5288 5468 5289
rect 5802 5289 5809 5300
rect 5861 5330 5868 5341
rect 6202 5341 6268 5342
rect 6202 5330 6209 5341
rect 5861 5300 6209 5330
rect 5861 5289 5868 5300
rect 5802 5288 5868 5289
rect 6202 5289 6209 5300
rect 6261 5330 6268 5341
rect 6704 5341 6770 5342
rect 6704 5330 6711 5341
rect 6261 5300 6711 5330
rect 6261 5289 6268 5300
rect 6202 5288 6268 5289
rect 6704 5289 6711 5300
rect 6763 5289 6770 5341
rect 6704 5288 6770 5289
rect 2 5271 68 5272
rect 2 5260 9 5271
rect 0 5230 9 5260
rect 2 5219 9 5230
rect 61 5260 68 5271
rect 402 5271 468 5272
rect 402 5260 409 5271
rect 61 5230 409 5260
rect 61 5219 68 5230
rect 2 5218 68 5219
rect 402 5219 409 5230
rect 461 5260 468 5271
rect 802 5271 868 5272
rect 802 5260 809 5271
rect 461 5230 809 5260
rect 461 5219 468 5230
rect 402 5218 468 5219
rect 802 5219 809 5230
rect 861 5260 868 5271
rect 1202 5271 1268 5272
rect 1202 5260 1209 5271
rect 861 5230 1209 5260
rect 861 5219 868 5230
rect 802 5218 868 5219
rect 1202 5219 1209 5230
rect 1261 5260 1268 5271
rect 1602 5271 1668 5272
rect 1602 5260 1609 5271
rect 1261 5230 1609 5260
rect 1261 5219 1268 5230
rect 1202 5218 1268 5219
rect 1602 5219 1609 5230
rect 1661 5260 1668 5271
rect 2002 5271 2068 5272
rect 2002 5260 2009 5271
rect 1661 5230 2009 5260
rect 1661 5219 1668 5230
rect 1602 5218 1668 5219
rect 2002 5219 2009 5230
rect 2061 5260 2068 5271
rect 2402 5271 2468 5272
rect 2402 5260 2409 5271
rect 2061 5230 2409 5260
rect 2061 5219 2068 5230
rect 2002 5218 2068 5219
rect 2402 5219 2409 5230
rect 2461 5260 2468 5271
rect 2802 5271 2868 5272
rect 2802 5260 2809 5271
rect 2461 5230 2809 5260
rect 2461 5219 2468 5230
rect 2402 5218 2468 5219
rect 2802 5219 2809 5230
rect 2861 5260 2868 5271
rect 3202 5271 3268 5272
rect 3202 5260 3209 5271
rect 2861 5230 3209 5260
rect 2861 5219 2868 5230
rect 2802 5218 2868 5219
rect 3202 5219 3209 5230
rect 3261 5260 3268 5271
rect 3602 5271 3668 5272
rect 3602 5260 3609 5271
rect 3261 5230 3609 5260
rect 3261 5219 3268 5230
rect 3202 5218 3268 5219
rect 3602 5219 3609 5230
rect 3661 5260 3668 5271
rect 4002 5271 4068 5272
rect 4002 5260 4009 5271
rect 3661 5230 4009 5260
rect 3661 5219 3668 5230
rect 3602 5218 3668 5219
rect 4002 5219 4009 5230
rect 4061 5260 4068 5271
rect 4402 5271 4468 5272
rect 4402 5260 4409 5271
rect 4061 5230 4409 5260
rect 4061 5219 4068 5230
rect 4002 5218 4068 5219
rect 4402 5219 4409 5230
rect 4461 5260 4468 5271
rect 4802 5271 4868 5272
rect 4802 5260 4809 5271
rect 4461 5230 4809 5260
rect 4461 5219 4468 5230
rect 4402 5218 4468 5219
rect 4802 5219 4809 5230
rect 4861 5260 4868 5271
rect 5202 5271 5268 5272
rect 5202 5260 5209 5271
rect 4861 5230 5209 5260
rect 4861 5219 4868 5230
rect 4802 5218 4868 5219
rect 5202 5219 5209 5230
rect 5261 5260 5268 5271
rect 5602 5271 5668 5272
rect 5602 5260 5609 5271
rect 5261 5230 5609 5260
rect 5261 5219 5268 5230
rect 5202 5218 5268 5219
rect 5602 5219 5609 5230
rect 5661 5260 5668 5271
rect 6002 5271 6068 5272
rect 6002 5260 6009 5271
rect 5661 5230 6009 5260
rect 5661 5219 5668 5230
rect 5602 5218 5668 5219
rect 6002 5219 6009 5230
rect 6061 5260 6068 5271
rect 6402 5271 6468 5272
rect 6402 5260 6409 5271
rect 6061 5230 6409 5260
rect 6061 5219 6068 5230
rect 6002 5218 6068 5219
rect 6402 5219 6409 5230
rect 6461 5260 6468 5271
rect 6500 5271 6566 5272
rect 6500 5260 6507 5271
rect 6461 5230 6507 5260
rect 6461 5219 6468 5230
rect 6402 5218 6468 5219
rect 6500 5219 6507 5230
rect 6559 5219 6566 5271
rect 6500 5218 6566 5219
rect 202 5201 268 5202
rect 202 5190 209 5201
rect 0 5160 209 5190
rect 202 5149 209 5160
rect 261 5190 268 5201
rect 602 5201 668 5202
rect 602 5190 609 5201
rect 261 5160 609 5190
rect 261 5149 268 5160
rect 202 5148 268 5149
rect 602 5149 609 5160
rect 661 5190 668 5201
rect 1002 5201 1068 5202
rect 1002 5190 1009 5201
rect 661 5160 1009 5190
rect 661 5149 668 5160
rect 602 5148 668 5149
rect 1002 5149 1009 5160
rect 1061 5190 1068 5201
rect 1402 5201 1468 5202
rect 1402 5190 1409 5201
rect 1061 5160 1409 5190
rect 1061 5149 1068 5160
rect 1002 5148 1068 5149
rect 1402 5149 1409 5160
rect 1461 5190 1468 5201
rect 1802 5201 1868 5202
rect 1802 5190 1809 5201
rect 1461 5160 1809 5190
rect 1461 5149 1468 5160
rect 1402 5148 1468 5149
rect 1802 5149 1809 5160
rect 1861 5190 1868 5201
rect 2202 5201 2268 5202
rect 2202 5190 2209 5201
rect 1861 5160 2209 5190
rect 1861 5149 1868 5160
rect 1802 5148 1868 5149
rect 2202 5149 2209 5160
rect 2261 5190 2268 5201
rect 2602 5201 2668 5202
rect 2602 5190 2609 5201
rect 2261 5160 2609 5190
rect 2261 5149 2268 5160
rect 2202 5148 2268 5149
rect 2602 5149 2609 5160
rect 2661 5190 2668 5201
rect 3002 5201 3068 5202
rect 3002 5190 3009 5201
rect 2661 5160 3009 5190
rect 2661 5149 2668 5160
rect 2602 5148 2668 5149
rect 3002 5149 3009 5160
rect 3061 5190 3068 5201
rect 3402 5201 3468 5202
rect 3402 5190 3409 5201
rect 3061 5160 3409 5190
rect 3061 5149 3068 5160
rect 3002 5148 3068 5149
rect 3402 5149 3409 5160
rect 3461 5190 3468 5201
rect 3802 5201 3868 5202
rect 3802 5190 3809 5201
rect 3461 5160 3809 5190
rect 3461 5149 3468 5160
rect 3402 5148 3468 5149
rect 3802 5149 3809 5160
rect 3861 5190 3868 5201
rect 4202 5201 4268 5202
rect 4202 5190 4209 5201
rect 3861 5160 4209 5190
rect 3861 5149 3868 5160
rect 3802 5148 3868 5149
rect 4202 5149 4209 5160
rect 4261 5190 4268 5201
rect 4602 5201 4668 5202
rect 4602 5190 4609 5201
rect 4261 5160 4609 5190
rect 4261 5149 4268 5160
rect 4202 5148 4268 5149
rect 4602 5149 4609 5160
rect 4661 5190 4668 5201
rect 5002 5201 5068 5202
rect 5002 5190 5009 5201
rect 4661 5160 5009 5190
rect 4661 5149 4668 5160
rect 4602 5148 4668 5149
rect 5002 5149 5009 5160
rect 5061 5190 5068 5201
rect 5402 5201 5468 5202
rect 5402 5190 5409 5201
rect 5061 5160 5409 5190
rect 5061 5149 5068 5160
rect 5002 5148 5068 5149
rect 5402 5149 5409 5160
rect 5461 5190 5468 5201
rect 5802 5201 5868 5202
rect 5802 5190 5809 5201
rect 5461 5160 5809 5190
rect 5461 5149 5468 5160
rect 5402 5148 5468 5149
rect 5802 5149 5809 5160
rect 5861 5190 5868 5201
rect 6202 5201 6268 5202
rect 6202 5190 6209 5201
rect 5861 5160 6209 5190
rect 5861 5149 5868 5160
rect 5802 5148 5868 5149
rect 6202 5149 6209 5160
rect 6261 5190 6268 5201
rect 6704 5201 6770 5202
rect 6704 5190 6711 5201
rect 6261 5160 6711 5190
rect 6261 5149 6268 5160
rect 6202 5148 6268 5149
rect 6704 5149 6711 5160
rect 6763 5149 6770 5201
rect 6704 5148 6770 5149
rect 2 5131 68 5132
rect 2 5120 9 5131
rect 0 5090 9 5120
rect 2 5079 9 5090
rect 61 5120 68 5131
rect 402 5131 468 5132
rect 402 5120 409 5131
rect 61 5090 409 5120
rect 61 5079 68 5090
rect 2 5078 68 5079
rect 402 5079 409 5090
rect 461 5120 468 5131
rect 802 5131 868 5132
rect 802 5120 809 5131
rect 461 5090 809 5120
rect 461 5079 468 5090
rect 402 5078 468 5079
rect 802 5079 809 5090
rect 861 5120 868 5131
rect 1202 5131 1268 5132
rect 1202 5120 1209 5131
rect 861 5090 1209 5120
rect 861 5079 868 5090
rect 802 5078 868 5079
rect 1202 5079 1209 5090
rect 1261 5120 1268 5131
rect 1602 5131 1668 5132
rect 1602 5120 1609 5131
rect 1261 5090 1609 5120
rect 1261 5079 1268 5090
rect 1202 5078 1268 5079
rect 1602 5079 1609 5090
rect 1661 5120 1668 5131
rect 2002 5131 2068 5132
rect 2002 5120 2009 5131
rect 1661 5090 2009 5120
rect 1661 5079 1668 5090
rect 1602 5078 1668 5079
rect 2002 5079 2009 5090
rect 2061 5120 2068 5131
rect 2402 5131 2468 5132
rect 2402 5120 2409 5131
rect 2061 5090 2409 5120
rect 2061 5079 2068 5090
rect 2002 5078 2068 5079
rect 2402 5079 2409 5090
rect 2461 5120 2468 5131
rect 2802 5131 2868 5132
rect 2802 5120 2809 5131
rect 2461 5090 2809 5120
rect 2461 5079 2468 5090
rect 2402 5078 2468 5079
rect 2802 5079 2809 5090
rect 2861 5120 2868 5131
rect 3202 5131 3268 5132
rect 3202 5120 3209 5131
rect 2861 5090 3209 5120
rect 2861 5079 2868 5090
rect 2802 5078 2868 5079
rect 3202 5079 3209 5090
rect 3261 5120 3268 5131
rect 3602 5131 3668 5132
rect 3602 5120 3609 5131
rect 3261 5090 3609 5120
rect 3261 5079 3268 5090
rect 3202 5078 3268 5079
rect 3602 5079 3609 5090
rect 3661 5120 3668 5131
rect 4002 5131 4068 5132
rect 4002 5120 4009 5131
rect 3661 5090 4009 5120
rect 3661 5079 3668 5090
rect 3602 5078 3668 5079
rect 4002 5079 4009 5090
rect 4061 5120 4068 5131
rect 4402 5131 4468 5132
rect 4402 5120 4409 5131
rect 4061 5090 4409 5120
rect 4061 5079 4068 5090
rect 4002 5078 4068 5079
rect 4402 5079 4409 5090
rect 4461 5120 4468 5131
rect 4802 5131 4868 5132
rect 4802 5120 4809 5131
rect 4461 5090 4809 5120
rect 4461 5079 4468 5090
rect 4402 5078 4468 5079
rect 4802 5079 4809 5090
rect 4861 5120 4868 5131
rect 5202 5131 5268 5132
rect 5202 5120 5209 5131
rect 4861 5090 5209 5120
rect 4861 5079 4868 5090
rect 4802 5078 4868 5079
rect 5202 5079 5209 5090
rect 5261 5120 5268 5131
rect 5602 5131 5668 5132
rect 5602 5120 5609 5131
rect 5261 5090 5609 5120
rect 5261 5079 5268 5090
rect 5202 5078 5268 5079
rect 5602 5079 5609 5090
rect 5661 5120 5668 5131
rect 6002 5131 6068 5132
rect 6002 5120 6009 5131
rect 5661 5090 6009 5120
rect 5661 5079 5668 5090
rect 5602 5078 5668 5079
rect 6002 5079 6009 5090
rect 6061 5120 6068 5131
rect 6402 5131 6468 5132
rect 6402 5120 6409 5131
rect 6061 5090 6409 5120
rect 6061 5079 6068 5090
rect 6002 5078 6068 5079
rect 6402 5079 6409 5090
rect 6461 5120 6468 5131
rect 6500 5131 6566 5132
rect 6500 5120 6507 5131
rect 6461 5090 6507 5120
rect 6461 5079 6468 5090
rect 6402 5078 6468 5079
rect 6500 5079 6507 5090
rect 6559 5079 6566 5131
rect 6500 5078 6566 5079
rect 196 4921 274 4922
rect -4 4905 74 4906
rect -4 4849 7 4905
rect 63 4849 74 4905
rect 196 4865 207 4921
rect 263 4865 274 4921
rect 596 4921 674 4922
rect 196 4864 274 4865
rect 396 4905 474 4906
rect -4 4848 74 4849
rect 396 4849 407 4905
rect 463 4849 474 4905
rect 596 4865 607 4921
rect 663 4865 674 4921
rect 996 4921 1074 4922
rect 596 4864 674 4865
rect 796 4905 874 4906
rect 396 4848 474 4849
rect 796 4849 807 4905
rect 863 4849 874 4905
rect 996 4865 1007 4921
rect 1063 4865 1074 4921
rect 1396 4921 1474 4922
rect 996 4864 1074 4865
rect 1196 4905 1274 4906
rect 796 4848 874 4849
rect 1196 4849 1207 4905
rect 1263 4849 1274 4905
rect 1396 4865 1407 4921
rect 1463 4865 1474 4921
rect 1796 4921 1874 4922
rect 1396 4864 1474 4865
rect 1596 4905 1674 4906
rect 1196 4848 1274 4849
rect 1596 4849 1607 4905
rect 1663 4849 1674 4905
rect 1796 4865 1807 4921
rect 1863 4865 1874 4921
rect 2196 4921 2274 4922
rect 1796 4864 1874 4865
rect 1996 4905 2074 4906
rect 1596 4848 1674 4849
rect 1996 4849 2007 4905
rect 2063 4849 2074 4905
rect 2196 4865 2207 4921
rect 2263 4865 2274 4921
rect 2596 4921 2674 4922
rect 2196 4864 2274 4865
rect 2396 4905 2474 4906
rect 1996 4848 2074 4849
rect 2396 4849 2407 4905
rect 2463 4849 2474 4905
rect 2596 4865 2607 4921
rect 2663 4865 2674 4921
rect 2996 4921 3074 4922
rect 2596 4864 2674 4865
rect 2796 4905 2874 4906
rect 2396 4848 2474 4849
rect 2796 4849 2807 4905
rect 2863 4849 2874 4905
rect 2996 4865 3007 4921
rect 3063 4865 3074 4921
rect 3396 4921 3474 4922
rect 2996 4864 3074 4865
rect 3196 4905 3274 4906
rect 2796 4848 2874 4849
rect 3196 4849 3207 4905
rect 3263 4849 3274 4905
rect 3396 4865 3407 4921
rect 3463 4865 3474 4921
rect 3796 4921 3874 4922
rect 3396 4864 3474 4865
rect 3596 4905 3674 4906
rect 3196 4848 3274 4849
rect 3596 4849 3607 4905
rect 3663 4849 3674 4905
rect 3796 4865 3807 4921
rect 3863 4865 3874 4921
rect 4196 4921 4274 4922
rect 3796 4864 3874 4865
rect 3996 4905 4074 4906
rect 3596 4848 3674 4849
rect 3996 4849 4007 4905
rect 4063 4849 4074 4905
rect 4196 4865 4207 4921
rect 4263 4865 4274 4921
rect 4596 4921 4674 4922
rect 4196 4864 4274 4865
rect 4396 4905 4474 4906
rect 3996 4848 4074 4849
rect 4396 4849 4407 4905
rect 4463 4849 4474 4905
rect 4596 4865 4607 4921
rect 4663 4865 4674 4921
rect 4996 4921 5074 4922
rect 4596 4864 4674 4865
rect 4796 4905 4874 4906
rect 4396 4848 4474 4849
rect 4796 4849 4807 4905
rect 4863 4849 4874 4905
rect 4996 4865 5007 4921
rect 5063 4865 5074 4921
rect 5396 4921 5474 4922
rect 4996 4864 5074 4865
rect 5196 4905 5274 4906
rect 4796 4848 4874 4849
rect 5196 4849 5207 4905
rect 5263 4849 5274 4905
rect 5396 4865 5407 4921
rect 5463 4865 5474 4921
rect 5796 4921 5874 4922
rect 5396 4864 5474 4865
rect 5596 4905 5674 4906
rect 5196 4848 5274 4849
rect 5596 4849 5607 4905
rect 5663 4849 5674 4905
rect 5796 4865 5807 4921
rect 5863 4865 5874 4921
rect 6196 4921 6274 4922
rect 5796 4864 5874 4865
rect 5996 4905 6074 4906
rect 5596 4848 5674 4849
rect 5996 4849 6007 4905
rect 6063 4849 6074 4905
rect 6196 4865 6207 4921
rect 6263 4865 6274 4921
rect 6196 4864 6274 4865
rect 5996 4848 6074 4849
rect 202 4831 268 4832
rect 202 4820 209 4831
rect 0 4790 209 4820
rect 202 4779 209 4790
rect 261 4820 268 4831
rect 602 4831 668 4832
rect 602 4820 609 4831
rect 261 4790 609 4820
rect 261 4779 268 4790
rect 202 4778 268 4779
rect 602 4779 609 4790
rect 661 4820 668 4831
rect 1002 4831 1068 4832
rect 1002 4820 1009 4831
rect 661 4790 1009 4820
rect 661 4779 668 4790
rect 602 4778 668 4779
rect 1002 4779 1009 4790
rect 1061 4820 1068 4831
rect 1402 4831 1468 4832
rect 1402 4820 1409 4831
rect 1061 4790 1409 4820
rect 1061 4779 1068 4790
rect 1002 4778 1068 4779
rect 1402 4779 1409 4790
rect 1461 4820 1468 4831
rect 1802 4831 1868 4832
rect 1802 4820 1809 4831
rect 1461 4790 1809 4820
rect 1461 4779 1468 4790
rect 1402 4778 1468 4779
rect 1802 4779 1809 4790
rect 1861 4820 1868 4831
rect 2202 4831 2268 4832
rect 2202 4820 2209 4831
rect 1861 4790 2209 4820
rect 1861 4779 1868 4790
rect 1802 4778 1868 4779
rect 2202 4779 2209 4790
rect 2261 4820 2268 4831
rect 2602 4831 2668 4832
rect 2602 4820 2609 4831
rect 2261 4790 2609 4820
rect 2261 4779 2268 4790
rect 2202 4778 2268 4779
rect 2602 4779 2609 4790
rect 2661 4820 2668 4831
rect 3002 4831 3068 4832
rect 3002 4820 3009 4831
rect 2661 4790 3009 4820
rect 2661 4779 2668 4790
rect 2602 4778 2668 4779
rect 3002 4779 3009 4790
rect 3061 4820 3068 4831
rect 3402 4831 3468 4832
rect 3402 4820 3409 4831
rect 3061 4790 3409 4820
rect 3061 4779 3068 4790
rect 3002 4778 3068 4779
rect 3402 4779 3409 4790
rect 3461 4820 3468 4831
rect 3802 4831 3868 4832
rect 3802 4820 3809 4831
rect 3461 4790 3809 4820
rect 3461 4779 3468 4790
rect 3402 4778 3468 4779
rect 3802 4779 3809 4790
rect 3861 4820 3868 4831
rect 4202 4831 4268 4832
rect 4202 4820 4209 4831
rect 3861 4790 4209 4820
rect 3861 4779 3868 4790
rect 3802 4778 3868 4779
rect 4202 4779 4209 4790
rect 4261 4820 4268 4831
rect 4602 4831 4668 4832
rect 4602 4820 4609 4831
rect 4261 4790 4609 4820
rect 4261 4779 4268 4790
rect 4202 4778 4268 4779
rect 4602 4779 4609 4790
rect 4661 4820 4668 4831
rect 5002 4831 5068 4832
rect 5002 4820 5009 4831
rect 4661 4790 5009 4820
rect 4661 4779 4668 4790
rect 4602 4778 4668 4779
rect 5002 4779 5009 4790
rect 5061 4820 5068 4831
rect 5402 4831 5468 4832
rect 5402 4820 5409 4831
rect 5061 4790 5409 4820
rect 5061 4779 5068 4790
rect 5002 4778 5068 4779
rect 5402 4779 5409 4790
rect 5461 4820 5468 4831
rect 5802 4831 5868 4832
rect 5802 4820 5809 4831
rect 5461 4790 5809 4820
rect 5461 4779 5468 4790
rect 5402 4778 5468 4779
rect 5802 4779 5809 4790
rect 5861 4820 5868 4831
rect 6202 4831 6268 4832
rect 6202 4820 6209 4831
rect 5861 4790 6209 4820
rect 5861 4779 5868 4790
rect 5802 4778 5868 4779
rect 6202 4779 6209 4790
rect 6261 4820 6268 4831
rect 6704 4831 6770 4832
rect 6704 4820 6711 4831
rect 6261 4790 6711 4820
rect 6261 4779 6268 4790
rect 6202 4778 6268 4779
rect 6704 4779 6711 4790
rect 6763 4779 6770 4831
rect 6704 4778 6770 4779
rect 2 4761 68 4762
rect 2 4750 9 4761
rect 0 4720 9 4750
rect 2 4709 9 4720
rect 61 4750 68 4761
rect 402 4761 468 4762
rect 402 4750 409 4761
rect 61 4720 409 4750
rect 61 4709 68 4720
rect 2 4708 68 4709
rect 402 4709 409 4720
rect 461 4750 468 4761
rect 802 4761 868 4762
rect 802 4750 809 4761
rect 461 4720 809 4750
rect 461 4709 468 4720
rect 402 4708 468 4709
rect 802 4709 809 4720
rect 861 4750 868 4761
rect 1202 4761 1268 4762
rect 1202 4750 1209 4761
rect 861 4720 1209 4750
rect 861 4709 868 4720
rect 802 4708 868 4709
rect 1202 4709 1209 4720
rect 1261 4750 1268 4761
rect 1602 4761 1668 4762
rect 1602 4750 1609 4761
rect 1261 4720 1609 4750
rect 1261 4709 1268 4720
rect 1202 4708 1268 4709
rect 1602 4709 1609 4720
rect 1661 4750 1668 4761
rect 2002 4761 2068 4762
rect 2002 4750 2009 4761
rect 1661 4720 2009 4750
rect 1661 4709 1668 4720
rect 1602 4708 1668 4709
rect 2002 4709 2009 4720
rect 2061 4750 2068 4761
rect 2402 4761 2468 4762
rect 2402 4750 2409 4761
rect 2061 4720 2409 4750
rect 2061 4709 2068 4720
rect 2002 4708 2068 4709
rect 2402 4709 2409 4720
rect 2461 4750 2468 4761
rect 2802 4761 2868 4762
rect 2802 4750 2809 4761
rect 2461 4720 2809 4750
rect 2461 4709 2468 4720
rect 2402 4708 2468 4709
rect 2802 4709 2809 4720
rect 2861 4750 2868 4761
rect 3202 4761 3268 4762
rect 3202 4750 3209 4761
rect 2861 4720 3209 4750
rect 2861 4709 2868 4720
rect 2802 4708 2868 4709
rect 3202 4709 3209 4720
rect 3261 4750 3268 4761
rect 3602 4761 3668 4762
rect 3602 4750 3609 4761
rect 3261 4720 3609 4750
rect 3261 4709 3268 4720
rect 3202 4708 3268 4709
rect 3602 4709 3609 4720
rect 3661 4750 3668 4761
rect 4002 4761 4068 4762
rect 4002 4750 4009 4761
rect 3661 4720 4009 4750
rect 3661 4709 3668 4720
rect 3602 4708 3668 4709
rect 4002 4709 4009 4720
rect 4061 4750 4068 4761
rect 4402 4761 4468 4762
rect 4402 4750 4409 4761
rect 4061 4720 4409 4750
rect 4061 4709 4068 4720
rect 4002 4708 4068 4709
rect 4402 4709 4409 4720
rect 4461 4750 4468 4761
rect 4802 4761 4868 4762
rect 4802 4750 4809 4761
rect 4461 4720 4809 4750
rect 4461 4709 4468 4720
rect 4402 4708 4468 4709
rect 4802 4709 4809 4720
rect 4861 4750 4868 4761
rect 5202 4761 5268 4762
rect 5202 4750 5209 4761
rect 4861 4720 5209 4750
rect 4861 4709 4868 4720
rect 4802 4708 4868 4709
rect 5202 4709 5209 4720
rect 5261 4750 5268 4761
rect 5602 4761 5668 4762
rect 5602 4750 5609 4761
rect 5261 4720 5609 4750
rect 5261 4709 5268 4720
rect 5202 4708 5268 4709
rect 5602 4709 5609 4720
rect 5661 4750 5668 4761
rect 6002 4761 6068 4762
rect 6002 4750 6009 4761
rect 5661 4720 6009 4750
rect 5661 4709 5668 4720
rect 5602 4708 5668 4709
rect 6002 4709 6009 4720
rect 6061 4750 6068 4761
rect 6402 4761 6468 4762
rect 6402 4750 6409 4761
rect 6061 4720 6409 4750
rect 6061 4709 6068 4720
rect 6002 4708 6068 4709
rect 6402 4709 6409 4720
rect 6461 4750 6468 4761
rect 6500 4761 6566 4762
rect 6500 4750 6507 4761
rect 6461 4720 6507 4750
rect 6461 4709 6468 4720
rect 6402 4708 6468 4709
rect 6500 4709 6507 4720
rect 6559 4709 6566 4761
rect 6500 4708 6566 4709
rect 202 4691 268 4692
rect 202 4680 209 4691
rect 0 4650 209 4680
rect 202 4639 209 4650
rect 261 4680 268 4691
rect 602 4691 668 4692
rect 602 4680 609 4691
rect 261 4650 609 4680
rect 261 4639 268 4650
rect 202 4638 268 4639
rect 602 4639 609 4650
rect 661 4680 668 4691
rect 1002 4691 1068 4692
rect 1002 4680 1009 4691
rect 661 4650 1009 4680
rect 661 4639 668 4650
rect 602 4638 668 4639
rect 1002 4639 1009 4650
rect 1061 4680 1068 4691
rect 1402 4691 1468 4692
rect 1402 4680 1409 4691
rect 1061 4650 1409 4680
rect 1061 4639 1068 4650
rect 1002 4638 1068 4639
rect 1402 4639 1409 4650
rect 1461 4680 1468 4691
rect 1802 4691 1868 4692
rect 1802 4680 1809 4691
rect 1461 4650 1809 4680
rect 1461 4639 1468 4650
rect 1402 4638 1468 4639
rect 1802 4639 1809 4650
rect 1861 4680 1868 4691
rect 2202 4691 2268 4692
rect 2202 4680 2209 4691
rect 1861 4650 2209 4680
rect 1861 4639 1868 4650
rect 1802 4638 1868 4639
rect 2202 4639 2209 4650
rect 2261 4680 2268 4691
rect 2602 4691 2668 4692
rect 2602 4680 2609 4691
rect 2261 4650 2609 4680
rect 2261 4639 2268 4650
rect 2202 4638 2268 4639
rect 2602 4639 2609 4650
rect 2661 4680 2668 4691
rect 3002 4691 3068 4692
rect 3002 4680 3009 4691
rect 2661 4650 3009 4680
rect 2661 4639 2668 4650
rect 2602 4638 2668 4639
rect 3002 4639 3009 4650
rect 3061 4680 3068 4691
rect 3402 4691 3468 4692
rect 3402 4680 3409 4691
rect 3061 4650 3409 4680
rect 3061 4639 3068 4650
rect 3002 4638 3068 4639
rect 3402 4639 3409 4650
rect 3461 4680 3468 4691
rect 3802 4691 3868 4692
rect 3802 4680 3809 4691
rect 3461 4650 3809 4680
rect 3461 4639 3468 4650
rect 3402 4638 3468 4639
rect 3802 4639 3809 4650
rect 3861 4680 3868 4691
rect 4202 4691 4268 4692
rect 4202 4680 4209 4691
rect 3861 4650 4209 4680
rect 3861 4639 3868 4650
rect 3802 4638 3868 4639
rect 4202 4639 4209 4650
rect 4261 4680 4268 4691
rect 4602 4691 4668 4692
rect 4602 4680 4609 4691
rect 4261 4650 4609 4680
rect 4261 4639 4268 4650
rect 4202 4638 4268 4639
rect 4602 4639 4609 4650
rect 4661 4680 4668 4691
rect 5002 4691 5068 4692
rect 5002 4680 5009 4691
rect 4661 4650 5009 4680
rect 4661 4639 4668 4650
rect 4602 4638 4668 4639
rect 5002 4639 5009 4650
rect 5061 4680 5068 4691
rect 5402 4691 5468 4692
rect 5402 4680 5409 4691
rect 5061 4650 5409 4680
rect 5061 4639 5068 4650
rect 5002 4638 5068 4639
rect 5402 4639 5409 4650
rect 5461 4680 5468 4691
rect 5802 4691 5868 4692
rect 5802 4680 5809 4691
rect 5461 4650 5809 4680
rect 5461 4639 5468 4650
rect 5402 4638 5468 4639
rect 5802 4639 5809 4650
rect 5861 4680 5868 4691
rect 6202 4691 6268 4692
rect 6202 4680 6209 4691
rect 5861 4650 6209 4680
rect 5861 4639 5868 4650
rect 5802 4638 5868 4639
rect 6202 4639 6209 4650
rect 6261 4680 6268 4691
rect 6704 4691 6770 4692
rect 6704 4680 6711 4691
rect 6261 4650 6711 4680
rect 6261 4639 6268 4650
rect 6202 4638 6268 4639
rect 6704 4639 6711 4650
rect 6763 4639 6770 4691
rect 6704 4638 6770 4639
rect 2 4621 68 4622
rect 2 4610 9 4621
rect 0 4580 9 4610
rect 2 4569 9 4580
rect 61 4610 68 4621
rect 402 4621 468 4622
rect 402 4610 409 4621
rect 61 4580 409 4610
rect 61 4569 68 4580
rect 2 4568 68 4569
rect 402 4569 409 4580
rect 461 4610 468 4621
rect 802 4621 868 4622
rect 802 4610 809 4621
rect 461 4580 809 4610
rect 461 4569 468 4580
rect 402 4568 468 4569
rect 802 4569 809 4580
rect 861 4610 868 4621
rect 1202 4621 1268 4622
rect 1202 4610 1209 4621
rect 861 4580 1209 4610
rect 861 4569 868 4580
rect 802 4568 868 4569
rect 1202 4569 1209 4580
rect 1261 4610 1268 4621
rect 1602 4621 1668 4622
rect 1602 4610 1609 4621
rect 1261 4580 1609 4610
rect 1261 4569 1268 4580
rect 1202 4568 1268 4569
rect 1602 4569 1609 4580
rect 1661 4610 1668 4621
rect 2002 4621 2068 4622
rect 2002 4610 2009 4621
rect 1661 4580 2009 4610
rect 1661 4569 1668 4580
rect 1602 4568 1668 4569
rect 2002 4569 2009 4580
rect 2061 4610 2068 4621
rect 2402 4621 2468 4622
rect 2402 4610 2409 4621
rect 2061 4580 2409 4610
rect 2061 4569 2068 4580
rect 2002 4568 2068 4569
rect 2402 4569 2409 4580
rect 2461 4610 2468 4621
rect 2802 4621 2868 4622
rect 2802 4610 2809 4621
rect 2461 4580 2809 4610
rect 2461 4569 2468 4580
rect 2402 4568 2468 4569
rect 2802 4569 2809 4580
rect 2861 4610 2868 4621
rect 3202 4621 3268 4622
rect 3202 4610 3209 4621
rect 2861 4580 3209 4610
rect 2861 4569 2868 4580
rect 2802 4568 2868 4569
rect 3202 4569 3209 4580
rect 3261 4610 3268 4621
rect 3602 4621 3668 4622
rect 3602 4610 3609 4621
rect 3261 4580 3609 4610
rect 3261 4569 3268 4580
rect 3202 4568 3268 4569
rect 3602 4569 3609 4580
rect 3661 4610 3668 4621
rect 4002 4621 4068 4622
rect 4002 4610 4009 4621
rect 3661 4580 4009 4610
rect 3661 4569 3668 4580
rect 3602 4568 3668 4569
rect 4002 4569 4009 4580
rect 4061 4610 4068 4621
rect 4402 4621 4468 4622
rect 4402 4610 4409 4621
rect 4061 4580 4409 4610
rect 4061 4569 4068 4580
rect 4002 4568 4068 4569
rect 4402 4569 4409 4580
rect 4461 4610 4468 4621
rect 4802 4621 4868 4622
rect 4802 4610 4809 4621
rect 4461 4580 4809 4610
rect 4461 4569 4468 4580
rect 4402 4568 4468 4569
rect 4802 4569 4809 4580
rect 4861 4610 4868 4621
rect 5202 4621 5268 4622
rect 5202 4610 5209 4621
rect 4861 4580 5209 4610
rect 4861 4569 4868 4580
rect 4802 4568 4868 4569
rect 5202 4569 5209 4580
rect 5261 4610 5268 4621
rect 5602 4621 5668 4622
rect 5602 4610 5609 4621
rect 5261 4580 5609 4610
rect 5261 4569 5268 4580
rect 5202 4568 5268 4569
rect 5602 4569 5609 4580
rect 5661 4610 5668 4621
rect 6002 4621 6068 4622
rect 6002 4610 6009 4621
rect 5661 4580 6009 4610
rect 5661 4569 5668 4580
rect 5602 4568 5668 4569
rect 6002 4569 6009 4580
rect 6061 4610 6068 4621
rect 6402 4621 6468 4622
rect 6402 4610 6409 4621
rect 6061 4580 6409 4610
rect 6061 4569 6068 4580
rect 6002 4568 6068 4569
rect 6402 4569 6409 4580
rect 6461 4610 6468 4621
rect 6500 4621 6566 4622
rect 6500 4610 6507 4621
rect 6461 4580 6507 4610
rect 6461 4569 6468 4580
rect 6402 4568 6468 4569
rect 6500 4569 6507 4580
rect 6559 4569 6566 4621
rect 6500 4568 6566 4569
rect 202 4551 268 4552
rect 202 4540 209 4551
rect 0 4510 209 4540
rect 202 4499 209 4510
rect 261 4540 268 4551
rect 602 4551 668 4552
rect 602 4540 609 4551
rect 261 4510 609 4540
rect 261 4499 268 4510
rect 202 4498 268 4499
rect 602 4499 609 4510
rect 661 4540 668 4551
rect 1002 4551 1068 4552
rect 1002 4540 1009 4551
rect 661 4510 1009 4540
rect 661 4499 668 4510
rect 602 4498 668 4499
rect 1002 4499 1009 4510
rect 1061 4540 1068 4551
rect 1402 4551 1468 4552
rect 1402 4540 1409 4551
rect 1061 4510 1409 4540
rect 1061 4499 1068 4510
rect 1002 4498 1068 4499
rect 1402 4499 1409 4510
rect 1461 4540 1468 4551
rect 1802 4551 1868 4552
rect 1802 4540 1809 4551
rect 1461 4510 1809 4540
rect 1461 4499 1468 4510
rect 1402 4498 1468 4499
rect 1802 4499 1809 4510
rect 1861 4540 1868 4551
rect 2202 4551 2268 4552
rect 2202 4540 2209 4551
rect 1861 4510 2209 4540
rect 1861 4499 1868 4510
rect 1802 4498 1868 4499
rect 2202 4499 2209 4510
rect 2261 4540 2268 4551
rect 2602 4551 2668 4552
rect 2602 4540 2609 4551
rect 2261 4510 2609 4540
rect 2261 4499 2268 4510
rect 2202 4498 2268 4499
rect 2602 4499 2609 4510
rect 2661 4540 2668 4551
rect 3002 4551 3068 4552
rect 3002 4540 3009 4551
rect 2661 4510 3009 4540
rect 2661 4499 2668 4510
rect 2602 4498 2668 4499
rect 3002 4499 3009 4510
rect 3061 4540 3068 4551
rect 3402 4551 3468 4552
rect 3402 4540 3409 4551
rect 3061 4510 3409 4540
rect 3061 4499 3068 4510
rect 3002 4498 3068 4499
rect 3402 4499 3409 4510
rect 3461 4540 3468 4551
rect 3802 4551 3868 4552
rect 3802 4540 3809 4551
rect 3461 4510 3809 4540
rect 3461 4499 3468 4510
rect 3402 4498 3468 4499
rect 3802 4499 3809 4510
rect 3861 4540 3868 4551
rect 4202 4551 4268 4552
rect 4202 4540 4209 4551
rect 3861 4510 4209 4540
rect 3861 4499 3868 4510
rect 3802 4498 3868 4499
rect 4202 4499 4209 4510
rect 4261 4540 4268 4551
rect 4602 4551 4668 4552
rect 4602 4540 4609 4551
rect 4261 4510 4609 4540
rect 4261 4499 4268 4510
rect 4202 4498 4268 4499
rect 4602 4499 4609 4510
rect 4661 4540 4668 4551
rect 5002 4551 5068 4552
rect 5002 4540 5009 4551
rect 4661 4510 5009 4540
rect 4661 4499 4668 4510
rect 4602 4498 4668 4499
rect 5002 4499 5009 4510
rect 5061 4540 5068 4551
rect 5402 4551 5468 4552
rect 5402 4540 5409 4551
rect 5061 4510 5409 4540
rect 5061 4499 5068 4510
rect 5002 4498 5068 4499
rect 5402 4499 5409 4510
rect 5461 4540 5468 4551
rect 5802 4551 5868 4552
rect 5802 4540 5809 4551
rect 5461 4510 5809 4540
rect 5461 4499 5468 4510
rect 5402 4498 5468 4499
rect 5802 4499 5809 4510
rect 5861 4540 5868 4551
rect 6202 4551 6268 4552
rect 6202 4540 6209 4551
rect 5861 4510 6209 4540
rect 5861 4499 5868 4510
rect 5802 4498 5868 4499
rect 6202 4499 6209 4510
rect 6261 4540 6268 4551
rect 6704 4551 6770 4552
rect 6704 4540 6711 4551
rect 6261 4510 6711 4540
rect 6261 4499 6268 4510
rect 6202 4498 6268 4499
rect 6704 4499 6711 4510
rect 6763 4499 6770 4551
rect 6704 4498 6770 4499
rect 2 4481 68 4482
rect 2 4470 9 4481
rect 0 4440 9 4470
rect 2 4429 9 4440
rect 61 4470 68 4481
rect 402 4481 468 4482
rect 402 4470 409 4481
rect 61 4440 409 4470
rect 61 4429 68 4440
rect 2 4428 68 4429
rect 402 4429 409 4440
rect 461 4470 468 4481
rect 802 4481 868 4482
rect 802 4470 809 4481
rect 461 4440 809 4470
rect 461 4429 468 4440
rect 402 4428 468 4429
rect 802 4429 809 4440
rect 861 4470 868 4481
rect 1202 4481 1268 4482
rect 1202 4470 1209 4481
rect 861 4440 1209 4470
rect 861 4429 868 4440
rect 802 4428 868 4429
rect 1202 4429 1209 4440
rect 1261 4470 1268 4481
rect 1602 4481 1668 4482
rect 1602 4470 1609 4481
rect 1261 4440 1609 4470
rect 1261 4429 1268 4440
rect 1202 4428 1268 4429
rect 1602 4429 1609 4440
rect 1661 4470 1668 4481
rect 2002 4481 2068 4482
rect 2002 4470 2009 4481
rect 1661 4440 2009 4470
rect 1661 4429 1668 4440
rect 1602 4428 1668 4429
rect 2002 4429 2009 4440
rect 2061 4470 2068 4481
rect 2402 4481 2468 4482
rect 2402 4470 2409 4481
rect 2061 4440 2409 4470
rect 2061 4429 2068 4440
rect 2002 4428 2068 4429
rect 2402 4429 2409 4440
rect 2461 4470 2468 4481
rect 2802 4481 2868 4482
rect 2802 4470 2809 4481
rect 2461 4440 2809 4470
rect 2461 4429 2468 4440
rect 2402 4428 2468 4429
rect 2802 4429 2809 4440
rect 2861 4470 2868 4481
rect 3202 4481 3268 4482
rect 3202 4470 3209 4481
rect 2861 4440 3209 4470
rect 2861 4429 2868 4440
rect 2802 4428 2868 4429
rect 3202 4429 3209 4440
rect 3261 4470 3268 4481
rect 3602 4481 3668 4482
rect 3602 4470 3609 4481
rect 3261 4440 3609 4470
rect 3261 4429 3268 4440
rect 3202 4428 3268 4429
rect 3602 4429 3609 4440
rect 3661 4470 3668 4481
rect 4002 4481 4068 4482
rect 4002 4470 4009 4481
rect 3661 4440 4009 4470
rect 3661 4429 3668 4440
rect 3602 4428 3668 4429
rect 4002 4429 4009 4440
rect 4061 4470 4068 4481
rect 4402 4481 4468 4482
rect 4402 4470 4409 4481
rect 4061 4440 4409 4470
rect 4061 4429 4068 4440
rect 4002 4428 4068 4429
rect 4402 4429 4409 4440
rect 4461 4470 4468 4481
rect 4802 4481 4868 4482
rect 4802 4470 4809 4481
rect 4461 4440 4809 4470
rect 4461 4429 4468 4440
rect 4402 4428 4468 4429
rect 4802 4429 4809 4440
rect 4861 4470 4868 4481
rect 5202 4481 5268 4482
rect 5202 4470 5209 4481
rect 4861 4440 5209 4470
rect 4861 4429 4868 4440
rect 4802 4428 4868 4429
rect 5202 4429 5209 4440
rect 5261 4470 5268 4481
rect 5602 4481 5668 4482
rect 5602 4470 5609 4481
rect 5261 4440 5609 4470
rect 5261 4429 5268 4440
rect 5202 4428 5268 4429
rect 5602 4429 5609 4440
rect 5661 4470 5668 4481
rect 6002 4481 6068 4482
rect 6002 4470 6009 4481
rect 5661 4440 6009 4470
rect 5661 4429 5668 4440
rect 5602 4428 5668 4429
rect 6002 4429 6009 4440
rect 6061 4470 6068 4481
rect 6402 4481 6468 4482
rect 6402 4470 6409 4481
rect 6061 4440 6409 4470
rect 6061 4429 6068 4440
rect 6002 4428 6068 4429
rect 6402 4429 6409 4440
rect 6461 4470 6468 4481
rect 6500 4481 6566 4482
rect 6500 4470 6507 4481
rect 6461 4440 6507 4470
rect 6461 4429 6468 4440
rect 6402 4428 6468 4429
rect 6500 4429 6507 4440
rect 6559 4429 6566 4481
rect 6500 4428 6566 4429
rect 202 4411 268 4412
rect 202 4400 209 4411
rect 0 4370 209 4400
rect 202 4359 209 4370
rect 261 4400 268 4411
rect 602 4411 668 4412
rect 602 4400 609 4411
rect 261 4370 609 4400
rect 261 4359 268 4370
rect 202 4358 268 4359
rect 602 4359 609 4370
rect 661 4400 668 4411
rect 1002 4411 1068 4412
rect 1002 4400 1009 4411
rect 661 4370 1009 4400
rect 661 4359 668 4370
rect 602 4358 668 4359
rect 1002 4359 1009 4370
rect 1061 4400 1068 4411
rect 1402 4411 1468 4412
rect 1402 4400 1409 4411
rect 1061 4370 1409 4400
rect 1061 4359 1068 4370
rect 1002 4358 1068 4359
rect 1402 4359 1409 4370
rect 1461 4400 1468 4411
rect 1802 4411 1868 4412
rect 1802 4400 1809 4411
rect 1461 4370 1809 4400
rect 1461 4359 1468 4370
rect 1402 4358 1468 4359
rect 1802 4359 1809 4370
rect 1861 4400 1868 4411
rect 2202 4411 2268 4412
rect 2202 4400 2209 4411
rect 1861 4370 2209 4400
rect 1861 4359 1868 4370
rect 1802 4358 1868 4359
rect 2202 4359 2209 4370
rect 2261 4400 2268 4411
rect 2602 4411 2668 4412
rect 2602 4400 2609 4411
rect 2261 4370 2609 4400
rect 2261 4359 2268 4370
rect 2202 4358 2268 4359
rect 2602 4359 2609 4370
rect 2661 4400 2668 4411
rect 3002 4411 3068 4412
rect 3002 4400 3009 4411
rect 2661 4370 3009 4400
rect 2661 4359 2668 4370
rect 2602 4358 2668 4359
rect 3002 4359 3009 4370
rect 3061 4400 3068 4411
rect 3402 4411 3468 4412
rect 3402 4400 3409 4411
rect 3061 4370 3409 4400
rect 3061 4359 3068 4370
rect 3002 4358 3068 4359
rect 3402 4359 3409 4370
rect 3461 4400 3468 4411
rect 3802 4411 3868 4412
rect 3802 4400 3809 4411
rect 3461 4370 3809 4400
rect 3461 4359 3468 4370
rect 3402 4358 3468 4359
rect 3802 4359 3809 4370
rect 3861 4400 3868 4411
rect 4202 4411 4268 4412
rect 4202 4400 4209 4411
rect 3861 4370 4209 4400
rect 3861 4359 3868 4370
rect 3802 4358 3868 4359
rect 4202 4359 4209 4370
rect 4261 4400 4268 4411
rect 4602 4411 4668 4412
rect 4602 4400 4609 4411
rect 4261 4370 4609 4400
rect 4261 4359 4268 4370
rect 4202 4358 4268 4359
rect 4602 4359 4609 4370
rect 4661 4400 4668 4411
rect 5002 4411 5068 4412
rect 5002 4400 5009 4411
rect 4661 4370 5009 4400
rect 4661 4359 4668 4370
rect 4602 4358 4668 4359
rect 5002 4359 5009 4370
rect 5061 4400 5068 4411
rect 5402 4411 5468 4412
rect 5402 4400 5409 4411
rect 5061 4370 5409 4400
rect 5061 4359 5068 4370
rect 5002 4358 5068 4359
rect 5402 4359 5409 4370
rect 5461 4400 5468 4411
rect 5802 4411 5868 4412
rect 5802 4400 5809 4411
rect 5461 4370 5809 4400
rect 5461 4359 5468 4370
rect 5402 4358 5468 4359
rect 5802 4359 5809 4370
rect 5861 4400 5868 4411
rect 6202 4411 6268 4412
rect 6202 4400 6209 4411
rect 5861 4370 6209 4400
rect 5861 4359 5868 4370
rect 5802 4358 5868 4359
rect 6202 4359 6209 4370
rect 6261 4400 6268 4411
rect 6704 4411 6770 4412
rect 6704 4400 6711 4411
rect 6261 4370 6711 4400
rect 6261 4359 6268 4370
rect 6202 4358 6268 4359
rect 6704 4359 6711 4370
rect 6763 4359 6770 4411
rect 6704 4358 6770 4359
rect 2 4341 68 4342
rect 2 4330 9 4341
rect 0 4300 9 4330
rect 2 4289 9 4300
rect 61 4330 68 4341
rect 402 4341 468 4342
rect 402 4330 409 4341
rect 61 4300 409 4330
rect 61 4289 68 4300
rect 2 4288 68 4289
rect 402 4289 409 4300
rect 461 4330 468 4341
rect 802 4341 868 4342
rect 802 4330 809 4341
rect 461 4300 809 4330
rect 461 4289 468 4300
rect 402 4288 468 4289
rect 802 4289 809 4300
rect 861 4330 868 4341
rect 1202 4341 1268 4342
rect 1202 4330 1209 4341
rect 861 4300 1209 4330
rect 861 4289 868 4300
rect 802 4288 868 4289
rect 1202 4289 1209 4300
rect 1261 4330 1268 4341
rect 1602 4341 1668 4342
rect 1602 4330 1609 4341
rect 1261 4300 1609 4330
rect 1261 4289 1268 4300
rect 1202 4288 1268 4289
rect 1602 4289 1609 4300
rect 1661 4330 1668 4341
rect 2002 4341 2068 4342
rect 2002 4330 2009 4341
rect 1661 4300 2009 4330
rect 1661 4289 1668 4300
rect 1602 4288 1668 4289
rect 2002 4289 2009 4300
rect 2061 4330 2068 4341
rect 2402 4341 2468 4342
rect 2402 4330 2409 4341
rect 2061 4300 2409 4330
rect 2061 4289 2068 4300
rect 2002 4288 2068 4289
rect 2402 4289 2409 4300
rect 2461 4330 2468 4341
rect 2802 4341 2868 4342
rect 2802 4330 2809 4341
rect 2461 4300 2809 4330
rect 2461 4289 2468 4300
rect 2402 4288 2468 4289
rect 2802 4289 2809 4300
rect 2861 4330 2868 4341
rect 3202 4341 3268 4342
rect 3202 4330 3209 4341
rect 2861 4300 3209 4330
rect 2861 4289 2868 4300
rect 2802 4288 2868 4289
rect 3202 4289 3209 4300
rect 3261 4330 3268 4341
rect 3602 4341 3668 4342
rect 3602 4330 3609 4341
rect 3261 4300 3609 4330
rect 3261 4289 3268 4300
rect 3202 4288 3268 4289
rect 3602 4289 3609 4300
rect 3661 4330 3668 4341
rect 4002 4341 4068 4342
rect 4002 4330 4009 4341
rect 3661 4300 4009 4330
rect 3661 4289 3668 4300
rect 3602 4288 3668 4289
rect 4002 4289 4009 4300
rect 4061 4330 4068 4341
rect 4402 4341 4468 4342
rect 4402 4330 4409 4341
rect 4061 4300 4409 4330
rect 4061 4289 4068 4300
rect 4002 4288 4068 4289
rect 4402 4289 4409 4300
rect 4461 4330 4468 4341
rect 4802 4341 4868 4342
rect 4802 4330 4809 4341
rect 4461 4300 4809 4330
rect 4461 4289 4468 4300
rect 4402 4288 4468 4289
rect 4802 4289 4809 4300
rect 4861 4330 4868 4341
rect 5202 4341 5268 4342
rect 5202 4330 5209 4341
rect 4861 4300 5209 4330
rect 4861 4289 4868 4300
rect 4802 4288 4868 4289
rect 5202 4289 5209 4300
rect 5261 4330 5268 4341
rect 5602 4341 5668 4342
rect 5602 4330 5609 4341
rect 5261 4300 5609 4330
rect 5261 4289 5268 4300
rect 5202 4288 5268 4289
rect 5602 4289 5609 4300
rect 5661 4330 5668 4341
rect 6002 4341 6068 4342
rect 6002 4330 6009 4341
rect 5661 4300 6009 4330
rect 5661 4289 5668 4300
rect 5602 4288 5668 4289
rect 6002 4289 6009 4300
rect 6061 4330 6068 4341
rect 6402 4341 6468 4342
rect 6402 4330 6409 4341
rect 6061 4300 6409 4330
rect 6061 4289 6068 4300
rect 6002 4288 6068 4289
rect 6402 4289 6409 4300
rect 6461 4330 6468 4341
rect 6500 4341 6566 4342
rect 6500 4330 6507 4341
rect 6461 4300 6507 4330
rect 6461 4289 6468 4300
rect 6402 4288 6468 4289
rect 6500 4289 6507 4300
rect 6559 4289 6566 4341
rect 6500 4288 6566 4289
rect 202 4271 268 4272
rect 202 4260 209 4271
rect 0 4230 209 4260
rect 202 4219 209 4230
rect 261 4260 268 4271
rect 602 4271 668 4272
rect 602 4260 609 4271
rect 261 4230 609 4260
rect 261 4219 268 4230
rect 202 4218 268 4219
rect 602 4219 609 4230
rect 661 4260 668 4271
rect 1002 4271 1068 4272
rect 1002 4260 1009 4271
rect 661 4230 1009 4260
rect 661 4219 668 4230
rect 602 4218 668 4219
rect 1002 4219 1009 4230
rect 1061 4260 1068 4271
rect 1402 4271 1468 4272
rect 1402 4260 1409 4271
rect 1061 4230 1409 4260
rect 1061 4219 1068 4230
rect 1002 4218 1068 4219
rect 1402 4219 1409 4230
rect 1461 4260 1468 4271
rect 1802 4271 1868 4272
rect 1802 4260 1809 4271
rect 1461 4230 1809 4260
rect 1461 4219 1468 4230
rect 1402 4218 1468 4219
rect 1802 4219 1809 4230
rect 1861 4260 1868 4271
rect 2202 4271 2268 4272
rect 2202 4260 2209 4271
rect 1861 4230 2209 4260
rect 1861 4219 1868 4230
rect 1802 4218 1868 4219
rect 2202 4219 2209 4230
rect 2261 4260 2268 4271
rect 2602 4271 2668 4272
rect 2602 4260 2609 4271
rect 2261 4230 2609 4260
rect 2261 4219 2268 4230
rect 2202 4218 2268 4219
rect 2602 4219 2609 4230
rect 2661 4260 2668 4271
rect 3002 4271 3068 4272
rect 3002 4260 3009 4271
rect 2661 4230 3009 4260
rect 2661 4219 2668 4230
rect 2602 4218 2668 4219
rect 3002 4219 3009 4230
rect 3061 4260 3068 4271
rect 3402 4271 3468 4272
rect 3402 4260 3409 4271
rect 3061 4230 3409 4260
rect 3061 4219 3068 4230
rect 3002 4218 3068 4219
rect 3402 4219 3409 4230
rect 3461 4260 3468 4271
rect 3802 4271 3868 4272
rect 3802 4260 3809 4271
rect 3461 4230 3809 4260
rect 3461 4219 3468 4230
rect 3402 4218 3468 4219
rect 3802 4219 3809 4230
rect 3861 4260 3868 4271
rect 4202 4271 4268 4272
rect 4202 4260 4209 4271
rect 3861 4230 4209 4260
rect 3861 4219 3868 4230
rect 3802 4218 3868 4219
rect 4202 4219 4209 4230
rect 4261 4260 4268 4271
rect 4602 4271 4668 4272
rect 4602 4260 4609 4271
rect 4261 4230 4609 4260
rect 4261 4219 4268 4230
rect 4202 4218 4268 4219
rect 4602 4219 4609 4230
rect 4661 4260 4668 4271
rect 5002 4271 5068 4272
rect 5002 4260 5009 4271
rect 4661 4230 5009 4260
rect 4661 4219 4668 4230
rect 4602 4218 4668 4219
rect 5002 4219 5009 4230
rect 5061 4260 5068 4271
rect 5402 4271 5468 4272
rect 5402 4260 5409 4271
rect 5061 4230 5409 4260
rect 5061 4219 5068 4230
rect 5002 4218 5068 4219
rect 5402 4219 5409 4230
rect 5461 4260 5468 4271
rect 5802 4271 5868 4272
rect 5802 4260 5809 4271
rect 5461 4230 5809 4260
rect 5461 4219 5468 4230
rect 5402 4218 5468 4219
rect 5802 4219 5809 4230
rect 5861 4260 5868 4271
rect 6202 4271 6268 4272
rect 6202 4260 6209 4271
rect 5861 4230 6209 4260
rect 5861 4219 5868 4230
rect 5802 4218 5868 4219
rect 6202 4219 6209 4230
rect 6261 4260 6268 4271
rect 6704 4271 6770 4272
rect 6704 4260 6711 4271
rect 6261 4230 6711 4260
rect 6261 4219 6268 4230
rect 6202 4218 6268 4219
rect 6704 4219 6711 4230
rect 6763 4219 6770 4271
rect 6704 4218 6770 4219
rect 2 4201 68 4202
rect 2 4190 9 4201
rect 0 4160 9 4190
rect 2 4149 9 4160
rect 61 4190 68 4201
rect 402 4201 468 4202
rect 402 4190 409 4201
rect 61 4160 409 4190
rect 61 4149 68 4160
rect 2 4148 68 4149
rect 402 4149 409 4160
rect 461 4190 468 4201
rect 802 4201 868 4202
rect 802 4190 809 4201
rect 461 4160 809 4190
rect 461 4149 468 4160
rect 402 4148 468 4149
rect 802 4149 809 4160
rect 861 4190 868 4201
rect 1202 4201 1268 4202
rect 1202 4190 1209 4201
rect 861 4160 1209 4190
rect 861 4149 868 4160
rect 802 4148 868 4149
rect 1202 4149 1209 4160
rect 1261 4190 1268 4201
rect 1602 4201 1668 4202
rect 1602 4190 1609 4201
rect 1261 4160 1609 4190
rect 1261 4149 1268 4160
rect 1202 4148 1268 4149
rect 1602 4149 1609 4160
rect 1661 4190 1668 4201
rect 2002 4201 2068 4202
rect 2002 4190 2009 4201
rect 1661 4160 2009 4190
rect 1661 4149 1668 4160
rect 1602 4148 1668 4149
rect 2002 4149 2009 4160
rect 2061 4190 2068 4201
rect 2402 4201 2468 4202
rect 2402 4190 2409 4201
rect 2061 4160 2409 4190
rect 2061 4149 2068 4160
rect 2002 4148 2068 4149
rect 2402 4149 2409 4160
rect 2461 4190 2468 4201
rect 2802 4201 2868 4202
rect 2802 4190 2809 4201
rect 2461 4160 2809 4190
rect 2461 4149 2468 4160
rect 2402 4148 2468 4149
rect 2802 4149 2809 4160
rect 2861 4190 2868 4201
rect 3202 4201 3268 4202
rect 3202 4190 3209 4201
rect 2861 4160 3209 4190
rect 2861 4149 2868 4160
rect 2802 4148 2868 4149
rect 3202 4149 3209 4160
rect 3261 4190 3268 4201
rect 3602 4201 3668 4202
rect 3602 4190 3609 4201
rect 3261 4160 3609 4190
rect 3261 4149 3268 4160
rect 3202 4148 3268 4149
rect 3602 4149 3609 4160
rect 3661 4190 3668 4201
rect 4002 4201 4068 4202
rect 4002 4190 4009 4201
rect 3661 4160 4009 4190
rect 3661 4149 3668 4160
rect 3602 4148 3668 4149
rect 4002 4149 4009 4160
rect 4061 4190 4068 4201
rect 4402 4201 4468 4202
rect 4402 4190 4409 4201
rect 4061 4160 4409 4190
rect 4061 4149 4068 4160
rect 4002 4148 4068 4149
rect 4402 4149 4409 4160
rect 4461 4190 4468 4201
rect 4802 4201 4868 4202
rect 4802 4190 4809 4201
rect 4461 4160 4809 4190
rect 4461 4149 4468 4160
rect 4402 4148 4468 4149
rect 4802 4149 4809 4160
rect 4861 4190 4868 4201
rect 5202 4201 5268 4202
rect 5202 4190 5209 4201
rect 4861 4160 5209 4190
rect 4861 4149 4868 4160
rect 4802 4148 4868 4149
rect 5202 4149 5209 4160
rect 5261 4190 5268 4201
rect 5602 4201 5668 4202
rect 5602 4190 5609 4201
rect 5261 4160 5609 4190
rect 5261 4149 5268 4160
rect 5202 4148 5268 4149
rect 5602 4149 5609 4160
rect 5661 4190 5668 4201
rect 6002 4201 6068 4202
rect 6002 4190 6009 4201
rect 5661 4160 6009 4190
rect 5661 4149 5668 4160
rect 5602 4148 5668 4149
rect 6002 4149 6009 4160
rect 6061 4190 6068 4201
rect 6402 4201 6468 4202
rect 6402 4190 6409 4201
rect 6061 4160 6409 4190
rect 6061 4149 6068 4160
rect 6002 4148 6068 4149
rect 6402 4149 6409 4160
rect 6461 4190 6468 4201
rect 6500 4201 6566 4202
rect 6500 4190 6507 4201
rect 6461 4160 6507 4190
rect 6461 4149 6468 4160
rect 6402 4148 6468 4149
rect 6500 4149 6507 4160
rect 6559 4149 6566 4201
rect 6500 4148 6566 4149
rect 202 4131 268 4132
rect 202 4120 209 4131
rect 0 4090 209 4120
rect 202 4079 209 4090
rect 261 4120 268 4131
rect 602 4131 668 4132
rect 602 4120 609 4131
rect 261 4090 609 4120
rect 261 4079 268 4090
rect 202 4078 268 4079
rect 602 4079 609 4090
rect 661 4120 668 4131
rect 1002 4131 1068 4132
rect 1002 4120 1009 4131
rect 661 4090 1009 4120
rect 661 4079 668 4090
rect 602 4078 668 4079
rect 1002 4079 1009 4090
rect 1061 4120 1068 4131
rect 1402 4131 1468 4132
rect 1402 4120 1409 4131
rect 1061 4090 1409 4120
rect 1061 4079 1068 4090
rect 1002 4078 1068 4079
rect 1402 4079 1409 4090
rect 1461 4120 1468 4131
rect 1802 4131 1868 4132
rect 1802 4120 1809 4131
rect 1461 4090 1809 4120
rect 1461 4079 1468 4090
rect 1402 4078 1468 4079
rect 1802 4079 1809 4090
rect 1861 4120 1868 4131
rect 2202 4131 2268 4132
rect 2202 4120 2209 4131
rect 1861 4090 2209 4120
rect 1861 4079 1868 4090
rect 1802 4078 1868 4079
rect 2202 4079 2209 4090
rect 2261 4120 2268 4131
rect 2602 4131 2668 4132
rect 2602 4120 2609 4131
rect 2261 4090 2609 4120
rect 2261 4079 2268 4090
rect 2202 4078 2268 4079
rect 2602 4079 2609 4090
rect 2661 4120 2668 4131
rect 3002 4131 3068 4132
rect 3002 4120 3009 4131
rect 2661 4090 3009 4120
rect 2661 4079 2668 4090
rect 2602 4078 2668 4079
rect 3002 4079 3009 4090
rect 3061 4120 3068 4131
rect 3402 4131 3468 4132
rect 3402 4120 3409 4131
rect 3061 4090 3409 4120
rect 3061 4079 3068 4090
rect 3002 4078 3068 4079
rect 3402 4079 3409 4090
rect 3461 4120 3468 4131
rect 3802 4131 3868 4132
rect 3802 4120 3809 4131
rect 3461 4090 3809 4120
rect 3461 4079 3468 4090
rect 3402 4078 3468 4079
rect 3802 4079 3809 4090
rect 3861 4120 3868 4131
rect 4202 4131 4268 4132
rect 4202 4120 4209 4131
rect 3861 4090 4209 4120
rect 3861 4079 3868 4090
rect 3802 4078 3868 4079
rect 4202 4079 4209 4090
rect 4261 4120 4268 4131
rect 4602 4131 4668 4132
rect 4602 4120 4609 4131
rect 4261 4090 4609 4120
rect 4261 4079 4268 4090
rect 4202 4078 4268 4079
rect 4602 4079 4609 4090
rect 4661 4120 4668 4131
rect 5002 4131 5068 4132
rect 5002 4120 5009 4131
rect 4661 4090 5009 4120
rect 4661 4079 4668 4090
rect 4602 4078 4668 4079
rect 5002 4079 5009 4090
rect 5061 4120 5068 4131
rect 5402 4131 5468 4132
rect 5402 4120 5409 4131
rect 5061 4090 5409 4120
rect 5061 4079 5068 4090
rect 5002 4078 5068 4079
rect 5402 4079 5409 4090
rect 5461 4120 5468 4131
rect 5802 4131 5868 4132
rect 5802 4120 5809 4131
rect 5461 4090 5809 4120
rect 5461 4079 5468 4090
rect 5402 4078 5468 4079
rect 5802 4079 5809 4090
rect 5861 4120 5868 4131
rect 6202 4131 6268 4132
rect 6202 4120 6209 4131
rect 5861 4090 6209 4120
rect 5861 4079 5868 4090
rect 5802 4078 5868 4079
rect 6202 4079 6209 4090
rect 6261 4120 6268 4131
rect 6704 4131 6770 4132
rect 6704 4120 6711 4131
rect 6261 4090 6711 4120
rect 6261 4079 6268 4090
rect 6202 4078 6268 4079
rect 6704 4079 6711 4090
rect 6763 4079 6770 4131
rect 6704 4078 6770 4079
rect 2 4061 68 4062
rect 2 4050 9 4061
rect 0 4020 9 4050
rect 2 4009 9 4020
rect 61 4050 68 4061
rect 402 4061 468 4062
rect 402 4050 409 4061
rect 61 4020 409 4050
rect 61 4009 68 4020
rect 2 4008 68 4009
rect 402 4009 409 4020
rect 461 4050 468 4061
rect 802 4061 868 4062
rect 802 4050 809 4061
rect 461 4020 809 4050
rect 461 4009 468 4020
rect 402 4008 468 4009
rect 802 4009 809 4020
rect 861 4050 868 4061
rect 1202 4061 1268 4062
rect 1202 4050 1209 4061
rect 861 4020 1209 4050
rect 861 4009 868 4020
rect 802 4008 868 4009
rect 1202 4009 1209 4020
rect 1261 4050 1268 4061
rect 1602 4061 1668 4062
rect 1602 4050 1609 4061
rect 1261 4020 1609 4050
rect 1261 4009 1268 4020
rect 1202 4008 1268 4009
rect 1602 4009 1609 4020
rect 1661 4050 1668 4061
rect 2002 4061 2068 4062
rect 2002 4050 2009 4061
rect 1661 4020 2009 4050
rect 1661 4009 1668 4020
rect 1602 4008 1668 4009
rect 2002 4009 2009 4020
rect 2061 4050 2068 4061
rect 2402 4061 2468 4062
rect 2402 4050 2409 4061
rect 2061 4020 2409 4050
rect 2061 4009 2068 4020
rect 2002 4008 2068 4009
rect 2402 4009 2409 4020
rect 2461 4050 2468 4061
rect 2802 4061 2868 4062
rect 2802 4050 2809 4061
rect 2461 4020 2809 4050
rect 2461 4009 2468 4020
rect 2402 4008 2468 4009
rect 2802 4009 2809 4020
rect 2861 4050 2868 4061
rect 3202 4061 3268 4062
rect 3202 4050 3209 4061
rect 2861 4020 3209 4050
rect 2861 4009 2868 4020
rect 2802 4008 2868 4009
rect 3202 4009 3209 4020
rect 3261 4050 3268 4061
rect 3602 4061 3668 4062
rect 3602 4050 3609 4061
rect 3261 4020 3609 4050
rect 3261 4009 3268 4020
rect 3202 4008 3268 4009
rect 3602 4009 3609 4020
rect 3661 4050 3668 4061
rect 4002 4061 4068 4062
rect 4002 4050 4009 4061
rect 3661 4020 4009 4050
rect 3661 4009 3668 4020
rect 3602 4008 3668 4009
rect 4002 4009 4009 4020
rect 4061 4050 4068 4061
rect 4402 4061 4468 4062
rect 4402 4050 4409 4061
rect 4061 4020 4409 4050
rect 4061 4009 4068 4020
rect 4002 4008 4068 4009
rect 4402 4009 4409 4020
rect 4461 4050 4468 4061
rect 4802 4061 4868 4062
rect 4802 4050 4809 4061
rect 4461 4020 4809 4050
rect 4461 4009 4468 4020
rect 4402 4008 4468 4009
rect 4802 4009 4809 4020
rect 4861 4050 4868 4061
rect 5202 4061 5268 4062
rect 5202 4050 5209 4061
rect 4861 4020 5209 4050
rect 4861 4009 4868 4020
rect 4802 4008 4868 4009
rect 5202 4009 5209 4020
rect 5261 4050 5268 4061
rect 5602 4061 5668 4062
rect 5602 4050 5609 4061
rect 5261 4020 5609 4050
rect 5261 4009 5268 4020
rect 5202 4008 5268 4009
rect 5602 4009 5609 4020
rect 5661 4050 5668 4061
rect 6002 4061 6068 4062
rect 6002 4050 6009 4061
rect 5661 4020 6009 4050
rect 5661 4009 5668 4020
rect 5602 4008 5668 4009
rect 6002 4009 6009 4020
rect 6061 4050 6068 4061
rect 6402 4061 6468 4062
rect 6402 4050 6409 4061
rect 6061 4020 6409 4050
rect 6061 4009 6068 4020
rect 6002 4008 6068 4009
rect 6402 4009 6409 4020
rect 6461 4050 6468 4061
rect 6500 4061 6566 4062
rect 6500 4050 6507 4061
rect 6461 4020 6507 4050
rect 6461 4009 6468 4020
rect 6402 4008 6468 4009
rect 6500 4009 6507 4020
rect 6559 4009 6566 4061
rect 6500 4008 6566 4009
rect 202 3991 268 3992
rect 202 3980 209 3991
rect 0 3950 209 3980
rect 202 3939 209 3950
rect 261 3980 268 3991
rect 602 3991 668 3992
rect 602 3980 609 3991
rect 261 3950 609 3980
rect 261 3939 268 3950
rect 202 3938 268 3939
rect 602 3939 609 3950
rect 661 3980 668 3991
rect 1002 3991 1068 3992
rect 1002 3980 1009 3991
rect 661 3950 1009 3980
rect 661 3939 668 3950
rect 602 3938 668 3939
rect 1002 3939 1009 3950
rect 1061 3980 1068 3991
rect 1402 3991 1468 3992
rect 1402 3980 1409 3991
rect 1061 3950 1409 3980
rect 1061 3939 1068 3950
rect 1002 3938 1068 3939
rect 1402 3939 1409 3950
rect 1461 3980 1468 3991
rect 1802 3991 1868 3992
rect 1802 3980 1809 3991
rect 1461 3950 1809 3980
rect 1461 3939 1468 3950
rect 1402 3938 1468 3939
rect 1802 3939 1809 3950
rect 1861 3980 1868 3991
rect 2202 3991 2268 3992
rect 2202 3980 2209 3991
rect 1861 3950 2209 3980
rect 1861 3939 1868 3950
rect 1802 3938 1868 3939
rect 2202 3939 2209 3950
rect 2261 3980 2268 3991
rect 2602 3991 2668 3992
rect 2602 3980 2609 3991
rect 2261 3950 2609 3980
rect 2261 3939 2268 3950
rect 2202 3938 2268 3939
rect 2602 3939 2609 3950
rect 2661 3980 2668 3991
rect 3002 3991 3068 3992
rect 3002 3980 3009 3991
rect 2661 3950 3009 3980
rect 2661 3939 2668 3950
rect 2602 3938 2668 3939
rect 3002 3939 3009 3950
rect 3061 3980 3068 3991
rect 3402 3991 3468 3992
rect 3402 3980 3409 3991
rect 3061 3950 3409 3980
rect 3061 3939 3068 3950
rect 3002 3938 3068 3939
rect 3402 3939 3409 3950
rect 3461 3980 3468 3991
rect 3802 3991 3868 3992
rect 3802 3980 3809 3991
rect 3461 3950 3809 3980
rect 3461 3939 3468 3950
rect 3402 3938 3468 3939
rect 3802 3939 3809 3950
rect 3861 3980 3868 3991
rect 4202 3991 4268 3992
rect 4202 3980 4209 3991
rect 3861 3950 4209 3980
rect 3861 3939 3868 3950
rect 3802 3938 3868 3939
rect 4202 3939 4209 3950
rect 4261 3980 4268 3991
rect 4602 3991 4668 3992
rect 4602 3980 4609 3991
rect 4261 3950 4609 3980
rect 4261 3939 4268 3950
rect 4202 3938 4268 3939
rect 4602 3939 4609 3950
rect 4661 3980 4668 3991
rect 5002 3991 5068 3992
rect 5002 3980 5009 3991
rect 4661 3950 5009 3980
rect 4661 3939 4668 3950
rect 4602 3938 4668 3939
rect 5002 3939 5009 3950
rect 5061 3980 5068 3991
rect 5402 3991 5468 3992
rect 5402 3980 5409 3991
rect 5061 3950 5409 3980
rect 5061 3939 5068 3950
rect 5002 3938 5068 3939
rect 5402 3939 5409 3950
rect 5461 3980 5468 3991
rect 5802 3991 5868 3992
rect 5802 3980 5809 3991
rect 5461 3950 5809 3980
rect 5461 3939 5468 3950
rect 5402 3938 5468 3939
rect 5802 3939 5809 3950
rect 5861 3980 5868 3991
rect 6202 3991 6268 3992
rect 6202 3980 6209 3991
rect 5861 3950 6209 3980
rect 5861 3939 5868 3950
rect 5802 3938 5868 3939
rect 6202 3939 6209 3950
rect 6261 3980 6268 3991
rect 6704 3991 6770 3992
rect 6704 3980 6711 3991
rect 6261 3950 6711 3980
rect 6261 3939 6268 3950
rect 6202 3938 6268 3939
rect 6704 3939 6711 3950
rect 6763 3939 6770 3991
rect 6704 3938 6770 3939
rect 2 3921 68 3922
rect 2 3910 9 3921
rect 0 3880 9 3910
rect 2 3869 9 3880
rect 61 3910 68 3921
rect 402 3921 468 3922
rect 402 3910 409 3921
rect 61 3880 409 3910
rect 61 3869 68 3880
rect 2 3868 68 3869
rect 402 3869 409 3880
rect 461 3910 468 3921
rect 802 3921 868 3922
rect 802 3910 809 3921
rect 461 3880 809 3910
rect 461 3869 468 3880
rect 402 3868 468 3869
rect 802 3869 809 3880
rect 861 3910 868 3921
rect 1202 3921 1268 3922
rect 1202 3910 1209 3921
rect 861 3880 1209 3910
rect 861 3869 868 3880
rect 802 3868 868 3869
rect 1202 3869 1209 3880
rect 1261 3910 1268 3921
rect 1602 3921 1668 3922
rect 1602 3910 1609 3921
rect 1261 3880 1609 3910
rect 1261 3869 1268 3880
rect 1202 3868 1268 3869
rect 1602 3869 1609 3880
rect 1661 3910 1668 3921
rect 2002 3921 2068 3922
rect 2002 3910 2009 3921
rect 1661 3880 2009 3910
rect 1661 3869 1668 3880
rect 1602 3868 1668 3869
rect 2002 3869 2009 3880
rect 2061 3910 2068 3921
rect 2402 3921 2468 3922
rect 2402 3910 2409 3921
rect 2061 3880 2409 3910
rect 2061 3869 2068 3880
rect 2002 3868 2068 3869
rect 2402 3869 2409 3880
rect 2461 3910 2468 3921
rect 2802 3921 2868 3922
rect 2802 3910 2809 3921
rect 2461 3880 2809 3910
rect 2461 3869 2468 3880
rect 2402 3868 2468 3869
rect 2802 3869 2809 3880
rect 2861 3910 2868 3921
rect 3202 3921 3268 3922
rect 3202 3910 3209 3921
rect 2861 3880 3209 3910
rect 2861 3869 2868 3880
rect 2802 3868 2868 3869
rect 3202 3869 3209 3880
rect 3261 3910 3268 3921
rect 3602 3921 3668 3922
rect 3602 3910 3609 3921
rect 3261 3880 3609 3910
rect 3261 3869 3268 3880
rect 3202 3868 3268 3869
rect 3602 3869 3609 3880
rect 3661 3910 3668 3921
rect 4002 3921 4068 3922
rect 4002 3910 4009 3921
rect 3661 3880 4009 3910
rect 3661 3869 3668 3880
rect 3602 3868 3668 3869
rect 4002 3869 4009 3880
rect 4061 3910 4068 3921
rect 4402 3921 4468 3922
rect 4402 3910 4409 3921
rect 4061 3880 4409 3910
rect 4061 3869 4068 3880
rect 4002 3868 4068 3869
rect 4402 3869 4409 3880
rect 4461 3910 4468 3921
rect 4802 3921 4868 3922
rect 4802 3910 4809 3921
rect 4461 3880 4809 3910
rect 4461 3869 4468 3880
rect 4402 3868 4468 3869
rect 4802 3869 4809 3880
rect 4861 3910 4868 3921
rect 5202 3921 5268 3922
rect 5202 3910 5209 3921
rect 4861 3880 5209 3910
rect 4861 3869 4868 3880
rect 4802 3868 4868 3869
rect 5202 3869 5209 3880
rect 5261 3910 5268 3921
rect 5602 3921 5668 3922
rect 5602 3910 5609 3921
rect 5261 3880 5609 3910
rect 5261 3869 5268 3880
rect 5202 3868 5268 3869
rect 5602 3869 5609 3880
rect 5661 3910 5668 3921
rect 6002 3921 6068 3922
rect 6002 3910 6009 3921
rect 5661 3880 6009 3910
rect 5661 3869 5668 3880
rect 5602 3868 5668 3869
rect 6002 3869 6009 3880
rect 6061 3910 6068 3921
rect 6402 3921 6468 3922
rect 6402 3910 6409 3921
rect 6061 3880 6409 3910
rect 6061 3869 6068 3880
rect 6002 3868 6068 3869
rect 6402 3869 6409 3880
rect 6461 3910 6468 3921
rect 6500 3921 6566 3922
rect 6500 3910 6507 3921
rect 6461 3880 6507 3910
rect 6461 3869 6468 3880
rect 6402 3868 6468 3869
rect 6500 3869 6507 3880
rect 6559 3869 6566 3921
rect 6500 3868 6566 3869
rect 202 3851 268 3852
rect 202 3840 209 3851
rect 0 3810 209 3840
rect 202 3799 209 3810
rect 261 3840 268 3851
rect 602 3851 668 3852
rect 602 3840 609 3851
rect 261 3810 609 3840
rect 261 3799 268 3810
rect 202 3798 268 3799
rect 602 3799 609 3810
rect 661 3840 668 3851
rect 1002 3851 1068 3852
rect 1002 3840 1009 3851
rect 661 3810 1009 3840
rect 661 3799 668 3810
rect 602 3798 668 3799
rect 1002 3799 1009 3810
rect 1061 3840 1068 3851
rect 1402 3851 1468 3852
rect 1402 3840 1409 3851
rect 1061 3810 1409 3840
rect 1061 3799 1068 3810
rect 1002 3798 1068 3799
rect 1402 3799 1409 3810
rect 1461 3840 1468 3851
rect 1802 3851 1868 3852
rect 1802 3840 1809 3851
rect 1461 3810 1809 3840
rect 1461 3799 1468 3810
rect 1402 3798 1468 3799
rect 1802 3799 1809 3810
rect 1861 3840 1868 3851
rect 2202 3851 2268 3852
rect 2202 3840 2209 3851
rect 1861 3810 2209 3840
rect 1861 3799 1868 3810
rect 1802 3798 1868 3799
rect 2202 3799 2209 3810
rect 2261 3840 2268 3851
rect 2602 3851 2668 3852
rect 2602 3840 2609 3851
rect 2261 3810 2609 3840
rect 2261 3799 2268 3810
rect 2202 3798 2268 3799
rect 2602 3799 2609 3810
rect 2661 3840 2668 3851
rect 3002 3851 3068 3852
rect 3002 3840 3009 3851
rect 2661 3810 3009 3840
rect 2661 3799 2668 3810
rect 2602 3798 2668 3799
rect 3002 3799 3009 3810
rect 3061 3840 3068 3851
rect 3402 3851 3468 3852
rect 3402 3840 3409 3851
rect 3061 3810 3409 3840
rect 3061 3799 3068 3810
rect 3002 3798 3068 3799
rect 3402 3799 3409 3810
rect 3461 3840 3468 3851
rect 3802 3851 3868 3852
rect 3802 3840 3809 3851
rect 3461 3810 3809 3840
rect 3461 3799 3468 3810
rect 3402 3798 3468 3799
rect 3802 3799 3809 3810
rect 3861 3840 3868 3851
rect 4202 3851 4268 3852
rect 4202 3840 4209 3851
rect 3861 3810 4209 3840
rect 3861 3799 3868 3810
rect 3802 3798 3868 3799
rect 4202 3799 4209 3810
rect 4261 3840 4268 3851
rect 4602 3851 4668 3852
rect 4602 3840 4609 3851
rect 4261 3810 4609 3840
rect 4261 3799 4268 3810
rect 4202 3798 4268 3799
rect 4602 3799 4609 3810
rect 4661 3840 4668 3851
rect 5002 3851 5068 3852
rect 5002 3840 5009 3851
rect 4661 3810 5009 3840
rect 4661 3799 4668 3810
rect 4602 3798 4668 3799
rect 5002 3799 5009 3810
rect 5061 3840 5068 3851
rect 5402 3851 5468 3852
rect 5402 3840 5409 3851
rect 5061 3810 5409 3840
rect 5061 3799 5068 3810
rect 5002 3798 5068 3799
rect 5402 3799 5409 3810
rect 5461 3840 5468 3851
rect 5802 3851 5868 3852
rect 5802 3840 5809 3851
rect 5461 3810 5809 3840
rect 5461 3799 5468 3810
rect 5402 3798 5468 3799
rect 5802 3799 5809 3810
rect 5861 3840 5868 3851
rect 6202 3851 6268 3852
rect 6202 3840 6209 3851
rect 5861 3810 6209 3840
rect 5861 3799 5868 3810
rect 5802 3798 5868 3799
rect 6202 3799 6209 3810
rect 6261 3840 6268 3851
rect 6704 3851 6770 3852
rect 6704 3840 6711 3851
rect 6261 3810 6711 3840
rect 6261 3799 6268 3810
rect 6202 3798 6268 3799
rect 6704 3799 6711 3810
rect 6763 3799 6770 3851
rect 6704 3798 6770 3799
rect 2 3781 68 3782
rect 2 3770 9 3781
rect 0 3740 9 3770
rect 2 3729 9 3740
rect 61 3770 68 3781
rect 402 3781 468 3782
rect 402 3770 409 3781
rect 61 3740 409 3770
rect 61 3729 68 3740
rect 2 3728 68 3729
rect 402 3729 409 3740
rect 461 3770 468 3781
rect 802 3781 868 3782
rect 802 3770 809 3781
rect 461 3740 809 3770
rect 461 3729 468 3740
rect 402 3728 468 3729
rect 802 3729 809 3740
rect 861 3770 868 3781
rect 1202 3781 1268 3782
rect 1202 3770 1209 3781
rect 861 3740 1209 3770
rect 861 3729 868 3740
rect 802 3728 868 3729
rect 1202 3729 1209 3740
rect 1261 3770 1268 3781
rect 1602 3781 1668 3782
rect 1602 3770 1609 3781
rect 1261 3740 1609 3770
rect 1261 3729 1268 3740
rect 1202 3728 1268 3729
rect 1602 3729 1609 3740
rect 1661 3770 1668 3781
rect 2002 3781 2068 3782
rect 2002 3770 2009 3781
rect 1661 3740 2009 3770
rect 1661 3729 1668 3740
rect 1602 3728 1668 3729
rect 2002 3729 2009 3740
rect 2061 3770 2068 3781
rect 2402 3781 2468 3782
rect 2402 3770 2409 3781
rect 2061 3740 2409 3770
rect 2061 3729 2068 3740
rect 2002 3728 2068 3729
rect 2402 3729 2409 3740
rect 2461 3770 2468 3781
rect 2802 3781 2868 3782
rect 2802 3770 2809 3781
rect 2461 3740 2809 3770
rect 2461 3729 2468 3740
rect 2402 3728 2468 3729
rect 2802 3729 2809 3740
rect 2861 3770 2868 3781
rect 3202 3781 3268 3782
rect 3202 3770 3209 3781
rect 2861 3740 3209 3770
rect 2861 3729 2868 3740
rect 2802 3728 2868 3729
rect 3202 3729 3209 3740
rect 3261 3770 3268 3781
rect 3602 3781 3668 3782
rect 3602 3770 3609 3781
rect 3261 3740 3609 3770
rect 3261 3729 3268 3740
rect 3202 3728 3268 3729
rect 3602 3729 3609 3740
rect 3661 3770 3668 3781
rect 4002 3781 4068 3782
rect 4002 3770 4009 3781
rect 3661 3740 4009 3770
rect 3661 3729 3668 3740
rect 3602 3728 3668 3729
rect 4002 3729 4009 3740
rect 4061 3770 4068 3781
rect 4402 3781 4468 3782
rect 4402 3770 4409 3781
rect 4061 3740 4409 3770
rect 4061 3729 4068 3740
rect 4002 3728 4068 3729
rect 4402 3729 4409 3740
rect 4461 3770 4468 3781
rect 4802 3781 4868 3782
rect 4802 3770 4809 3781
rect 4461 3740 4809 3770
rect 4461 3729 4468 3740
rect 4402 3728 4468 3729
rect 4802 3729 4809 3740
rect 4861 3770 4868 3781
rect 5202 3781 5268 3782
rect 5202 3770 5209 3781
rect 4861 3740 5209 3770
rect 4861 3729 4868 3740
rect 4802 3728 4868 3729
rect 5202 3729 5209 3740
rect 5261 3770 5268 3781
rect 5602 3781 5668 3782
rect 5602 3770 5609 3781
rect 5261 3740 5609 3770
rect 5261 3729 5268 3740
rect 5202 3728 5268 3729
rect 5602 3729 5609 3740
rect 5661 3770 5668 3781
rect 6002 3781 6068 3782
rect 6002 3770 6009 3781
rect 5661 3740 6009 3770
rect 5661 3729 5668 3740
rect 5602 3728 5668 3729
rect 6002 3729 6009 3740
rect 6061 3770 6068 3781
rect 6402 3781 6468 3782
rect 6402 3770 6409 3781
rect 6061 3740 6409 3770
rect 6061 3729 6068 3740
rect 6002 3728 6068 3729
rect 6402 3729 6409 3740
rect 6461 3770 6468 3781
rect 6500 3781 6566 3782
rect 6500 3770 6507 3781
rect 6461 3740 6507 3770
rect 6461 3729 6468 3740
rect 6402 3728 6468 3729
rect 6500 3729 6507 3740
rect 6559 3729 6566 3781
rect 6500 3728 6566 3729
rect 196 3711 274 3712
rect -4 3695 74 3696
rect -4 3639 7 3695
rect 63 3639 74 3695
rect 196 3655 207 3711
rect 263 3655 274 3711
rect 596 3711 674 3712
rect 196 3654 274 3655
rect 396 3695 474 3696
rect -4 3638 74 3639
rect 396 3639 407 3695
rect 463 3639 474 3695
rect 596 3655 607 3711
rect 663 3655 674 3711
rect 996 3711 1074 3712
rect 596 3654 674 3655
rect 796 3695 874 3696
rect 396 3638 474 3639
rect 796 3639 807 3695
rect 863 3639 874 3695
rect 996 3655 1007 3711
rect 1063 3655 1074 3711
rect 1396 3711 1474 3712
rect 996 3654 1074 3655
rect 1196 3695 1274 3696
rect 796 3638 874 3639
rect 1196 3639 1207 3695
rect 1263 3639 1274 3695
rect 1396 3655 1407 3711
rect 1463 3655 1474 3711
rect 1796 3711 1874 3712
rect 1396 3654 1474 3655
rect 1596 3695 1674 3696
rect 1196 3638 1274 3639
rect 1596 3639 1607 3695
rect 1663 3639 1674 3695
rect 1796 3655 1807 3711
rect 1863 3655 1874 3711
rect 2196 3711 2274 3712
rect 1796 3654 1874 3655
rect 1996 3695 2074 3696
rect 1596 3638 1674 3639
rect 1996 3639 2007 3695
rect 2063 3639 2074 3695
rect 2196 3655 2207 3711
rect 2263 3655 2274 3711
rect 2596 3711 2674 3712
rect 2196 3654 2274 3655
rect 2396 3695 2474 3696
rect 1996 3638 2074 3639
rect 2396 3639 2407 3695
rect 2463 3639 2474 3695
rect 2596 3655 2607 3711
rect 2663 3655 2674 3711
rect 2996 3711 3074 3712
rect 2596 3654 2674 3655
rect 2796 3695 2874 3696
rect 2396 3638 2474 3639
rect 2796 3639 2807 3695
rect 2863 3639 2874 3695
rect 2996 3655 3007 3711
rect 3063 3655 3074 3711
rect 3396 3711 3474 3712
rect 2996 3654 3074 3655
rect 3196 3695 3274 3696
rect 2796 3638 2874 3639
rect 3196 3639 3207 3695
rect 3263 3639 3274 3695
rect 3396 3655 3407 3711
rect 3463 3655 3474 3711
rect 3796 3711 3874 3712
rect 3396 3654 3474 3655
rect 3596 3695 3674 3696
rect 3196 3638 3274 3639
rect 3596 3639 3607 3695
rect 3663 3639 3674 3695
rect 3796 3655 3807 3711
rect 3863 3655 3874 3711
rect 4196 3711 4274 3712
rect 3796 3654 3874 3655
rect 3996 3695 4074 3696
rect 3596 3638 3674 3639
rect 3996 3639 4007 3695
rect 4063 3639 4074 3695
rect 4196 3655 4207 3711
rect 4263 3655 4274 3711
rect 4596 3711 4674 3712
rect 4196 3654 4274 3655
rect 4396 3695 4474 3696
rect 3996 3638 4074 3639
rect 4396 3639 4407 3695
rect 4463 3639 4474 3695
rect 4596 3655 4607 3711
rect 4663 3655 4674 3711
rect 4996 3711 5074 3712
rect 4596 3654 4674 3655
rect 4796 3695 4874 3696
rect 4396 3638 4474 3639
rect 4796 3639 4807 3695
rect 4863 3639 4874 3695
rect 4996 3655 5007 3711
rect 5063 3655 5074 3711
rect 5396 3711 5474 3712
rect 4996 3654 5074 3655
rect 5196 3695 5274 3696
rect 4796 3638 4874 3639
rect 5196 3639 5207 3695
rect 5263 3639 5274 3695
rect 5396 3655 5407 3711
rect 5463 3655 5474 3711
rect 5796 3711 5874 3712
rect 5396 3654 5474 3655
rect 5596 3695 5674 3696
rect 5196 3638 5274 3639
rect 5596 3639 5607 3695
rect 5663 3639 5674 3695
rect 5796 3655 5807 3711
rect 5863 3655 5874 3711
rect 6196 3711 6274 3712
rect 5796 3654 5874 3655
rect 5996 3695 6074 3696
rect 5596 3638 5674 3639
rect 5996 3639 6007 3695
rect 6063 3639 6074 3695
rect 6196 3655 6207 3711
rect 6263 3655 6274 3711
rect 6196 3654 6274 3655
rect 5996 3638 6074 3639
rect 202 3621 268 3622
rect 202 3610 209 3621
rect 0 3580 209 3610
rect 202 3569 209 3580
rect 261 3610 268 3621
rect 602 3621 668 3622
rect 602 3610 609 3621
rect 261 3580 609 3610
rect 261 3569 268 3580
rect 202 3568 268 3569
rect 602 3569 609 3580
rect 661 3610 668 3621
rect 1002 3621 1068 3622
rect 1002 3610 1009 3621
rect 661 3580 1009 3610
rect 661 3569 668 3580
rect 602 3568 668 3569
rect 1002 3569 1009 3580
rect 1061 3610 1068 3621
rect 1402 3621 1468 3622
rect 1402 3610 1409 3621
rect 1061 3580 1409 3610
rect 1061 3569 1068 3580
rect 1002 3568 1068 3569
rect 1402 3569 1409 3580
rect 1461 3610 1468 3621
rect 1802 3621 1868 3622
rect 1802 3610 1809 3621
rect 1461 3580 1809 3610
rect 1461 3569 1468 3580
rect 1402 3568 1468 3569
rect 1802 3569 1809 3580
rect 1861 3610 1868 3621
rect 2202 3621 2268 3622
rect 2202 3610 2209 3621
rect 1861 3580 2209 3610
rect 1861 3569 1868 3580
rect 1802 3568 1868 3569
rect 2202 3569 2209 3580
rect 2261 3610 2268 3621
rect 2602 3621 2668 3622
rect 2602 3610 2609 3621
rect 2261 3580 2609 3610
rect 2261 3569 2268 3580
rect 2202 3568 2268 3569
rect 2602 3569 2609 3580
rect 2661 3610 2668 3621
rect 3002 3621 3068 3622
rect 3002 3610 3009 3621
rect 2661 3580 3009 3610
rect 2661 3569 2668 3580
rect 2602 3568 2668 3569
rect 3002 3569 3009 3580
rect 3061 3610 3068 3621
rect 3402 3621 3468 3622
rect 3402 3610 3409 3621
rect 3061 3580 3409 3610
rect 3061 3569 3068 3580
rect 3002 3568 3068 3569
rect 3402 3569 3409 3580
rect 3461 3610 3468 3621
rect 3802 3621 3868 3622
rect 3802 3610 3809 3621
rect 3461 3580 3809 3610
rect 3461 3569 3468 3580
rect 3402 3568 3468 3569
rect 3802 3569 3809 3580
rect 3861 3610 3868 3621
rect 4202 3621 4268 3622
rect 4202 3610 4209 3621
rect 3861 3580 4209 3610
rect 3861 3569 3868 3580
rect 3802 3568 3868 3569
rect 4202 3569 4209 3580
rect 4261 3610 4268 3621
rect 4602 3621 4668 3622
rect 4602 3610 4609 3621
rect 4261 3580 4609 3610
rect 4261 3569 4268 3580
rect 4202 3568 4268 3569
rect 4602 3569 4609 3580
rect 4661 3610 4668 3621
rect 5002 3621 5068 3622
rect 5002 3610 5009 3621
rect 4661 3580 5009 3610
rect 4661 3569 4668 3580
rect 4602 3568 4668 3569
rect 5002 3569 5009 3580
rect 5061 3610 5068 3621
rect 5402 3621 5468 3622
rect 5402 3610 5409 3621
rect 5061 3580 5409 3610
rect 5061 3569 5068 3580
rect 5002 3568 5068 3569
rect 5402 3569 5409 3580
rect 5461 3610 5468 3621
rect 5802 3621 5868 3622
rect 5802 3610 5809 3621
rect 5461 3580 5809 3610
rect 5461 3569 5468 3580
rect 5402 3568 5468 3569
rect 5802 3569 5809 3580
rect 5861 3610 5868 3621
rect 6202 3621 6268 3622
rect 6202 3610 6209 3621
rect 5861 3580 6209 3610
rect 5861 3569 5868 3580
rect 5802 3568 5868 3569
rect 6202 3569 6209 3580
rect 6261 3610 6268 3621
rect 6704 3621 6770 3622
rect 6704 3610 6711 3621
rect 6261 3580 6711 3610
rect 6261 3569 6268 3580
rect 6202 3568 6268 3569
rect 6704 3569 6711 3580
rect 6763 3569 6770 3621
rect 6704 3568 6770 3569
rect 2 3551 68 3552
rect 2 3540 9 3551
rect 0 3510 9 3540
rect 2 3499 9 3510
rect 61 3540 68 3551
rect 402 3551 468 3552
rect 402 3540 409 3551
rect 61 3510 409 3540
rect 61 3499 68 3510
rect 2 3498 68 3499
rect 402 3499 409 3510
rect 461 3540 468 3551
rect 802 3551 868 3552
rect 802 3540 809 3551
rect 461 3510 809 3540
rect 461 3499 468 3510
rect 402 3498 468 3499
rect 802 3499 809 3510
rect 861 3540 868 3551
rect 1202 3551 1268 3552
rect 1202 3540 1209 3551
rect 861 3510 1209 3540
rect 861 3499 868 3510
rect 802 3498 868 3499
rect 1202 3499 1209 3510
rect 1261 3540 1268 3551
rect 1602 3551 1668 3552
rect 1602 3540 1609 3551
rect 1261 3510 1609 3540
rect 1261 3499 1268 3510
rect 1202 3498 1268 3499
rect 1602 3499 1609 3510
rect 1661 3540 1668 3551
rect 2002 3551 2068 3552
rect 2002 3540 2009 3551
rect 1661 3510 2009 3540
rect 1661 3499 1668 3510
rect 1602 3498 1668 3499
rect 2002 3499 2009 3510
rect 2061 3540 2068 3551
rect 2402 3551 2468 3552
rect 2402 3540 2409 3551
rect 2061 3510 2409 3540
rect 2061 3499 2068 3510
rect 2002 3498 2068 3499
rect 2402 3499 2409 3510
rect 2461 3540 2468 3551
rect 2802 3551 2868 3552
rect 2802 3540 2809 3551
rect 2461 3510 2809 3540
rect 2461 3499 2468 3510
rect 2402 3498 2468 3499
rect 2802 3499 2809 3510
rect 2861 3540 2868 3551
rect 3202 3551 3268 3552
rect 3202 3540 3209 3551
rect 2861 3510 3209 3540
rect 2861 3499 2868 3510
rect 2802 3498 2868 3499
rect 3202 3499 3209 3510
rect 3261 3540 3268 3551
rect 3602 3551 3668 3552
rect 3602 3540 3609 3551
rect 3261 3510 3609 3540
rect 3261 3499 3268 3510
rect 3202 3498 3268 3499
rect 3602 3499 3609 3510
rect 3661 3540 3668 3551
rect 4002 3551 4068 3552
rect 4002 3540 4009 3551
rect 3661 3510 4009 3540
rect 3661 3499 3668 3510
rect 3602 3498 3668 3499
rect 4002 3499 4009 3510
rect 4061 3540 4068 3551
rect 4402 3551 4468 3552
rect 4402 3540 4409 3551
rect 4061 3510 4409 3540
rect 4061 3499 4068 3510
rect 4002 3498 4068 3499
rect 4402 3499 4409 3510
rect 4461 3540 4468 3551
rect 4802 3551 4868 3552
rect 4802 3540 4809 3551
rect 4461 3510 4809 3540
rect 4461 3499 4468 3510
rect 4402 3498 4468 3499
rect 4802 3499 4809 3510
rect 4861 3540 4868 3551
rect 5202 3551 5268 3552
rect 5202 3540 5209 3551
rect 4861 3510 5209 3540
rect 4861 3499 4868 3510
rect 4802 3498 4868 3499
rect 5202 3499 5209 3510
rect 5261 3540 5268 3551
rect 5602 3551 5668 3552
rect 5602 3540 5609 3551
rect 5261 3510 5609 3540
rect 5261 3499 5268 3510
rect 5202 3498 5268 3499
rect 5602 3499 5609 3510
rect 5661 3540 5668 3551
rect 6002 3551 6068 3552
rect 6002 3540 6009 3551
rect 5661 3510 6009 3540
rect 5661 3499 5668 3510
rect 5602 3498 5668 3499
rect 6002 3499 6009 3510
rect 6061 3540 6068 3551
rect 6402 3551 6468 3552
rect 6402 3540 6409 3551
rect 6061 3510 6409 3540
rect 6061 3499 6068 3510
rect 6002 3498 6068 3499
rect 6402 3499 6409 3510
rect 6461 3540 6468 3551
rect 6500 3551 6566 3552
rect 6500 3540 6507 3551
rect 6461 3510 6507 3540
rect 6461 3499 6468 3510
rect 6402 3498 6468 3499
rect 6500 3499 6507 3510
rect 6559 3499 6566 3551
rect 6500 3498 6566 3499
rect 202 3481 268 3482
rect 202 3470 209 3481
rect 0 3440 209 3470
rect 202 3429 209 3440
rect 261 3470 268 3481
rect 602 3481 668 3482
rect 602 3470 609 3481
rect 261 3440 609 3470
rect 261 3429 268 3440
rect 202 3428 268 3429
rect 602 3429 609 3440
rect 661 3470 668 3481
rect 1002 3481 1068 3482
rect 1002 3470 1009 3481
rect 661 3440 1009 3470
rect 661 3429 668 3440
rect 602 3428 668 3429
rect 1002 3429 1009 3440
rect 1061 3470 1068 3481
rect 1402 3481 1468 3482
rect 1402 3470 1409 3481
rect 1061 3440 1409 3470
rect 1061 3429 1068 3440
rect 1002 3428 1068 3429
rect 1402 3429 1409 3440
rect 1461 3470 1468 3481
rect 1802 3481 1868 3482
rect 1802 3470 1809 3481
rect 1461 3440 1809 3470
rect 1461 3429 1468 3440
rect 1402 3428 1468 3429
rect 1802 3429 1809 3440
rect 1861 3470 1868 3481
rect 2202 3481 2268 3482
rect 2202 3470 2209 3481
rect 1861 3440 2209 3470
rect 1861 3429 1868 3440
rect 1802 3428 1868 3429
rect 2202 3429 2209 3440
rect 2261 3470 2268 3481
rect 2602 3481 2668 3482
rect 2602 3470 2609 3481
rect 2261 3440 2609 3470
rect 2261 3429 2268 3440
rect 2202 3428 2268 3429
rect 2602 3429 2609 3440
rect 2661 3470 2668 3481
rect 3002 3481 3068 3482
rect 3002 3470 3009 3481
rect 2661 3440 3009 3470
rect 2661 3429 2668 3440
rect 2602 3428 2668 3429
rect 3002 3429 3009 3440
rect 3061 3470 3068 3481
rect 3402 3481 3468 3482
rect 3402 3470 3409 3481
rect 3061 3440 3409 3470
rect 3061 3429 3068 3440
rect 3002 3428 3068 3429
rect 3402 3429 3409 3440
rect 3461 3470 3468 3481
rect 3802 3481 3868 3482
rect 3802 3470 3809 3481
rect 3461 3440 3809 3470
rect 3461 3429 3468 3440
rect 3402 3428 3468 3429
rect 3802 3429 3809 3440
rect 3861 3470 3868 3481
rect 4202 3481 4268 3482
rect 4202 3470 4209 3481
rect 3861 3440 4209 3470
rect 3861 3429 3868 3440
rect 3802 3428 3868 3429
rect 4202 3429 4209 3440
rect 4261 3470 4268 3481
rect 4602 3481 4668 3482
rect 4602 3470 4609 3481
rect 4261 3440 4609 3470
rect 4261 3429 4268 3440
rect 4202 3428 4268 3429
rect 4602 3429 4609 3440
rect 4661 3470 4668 3481
rect 5002 3481 5068 3482
rect 5002 3470 5009 3481
rect 4661 3440 5009 3470
rect 4661 3429 4668 3440
rect 4602 3428 4668 3429
rect 5002 3429 5009 3440
rect 5061 3470 5068 3481
rect 5402 3481 5468 3482
rect 5402 3470 5409 3481
rect 5061 3440 5409 3470
rect 5061 3429 5068 3440
rect 5002 3428 5068 3429
rect 5402 3429 5409 3440
rect 5461 3470 5468 3481
rect 5802 3481 5868 3482
rect 5802 3470 5809 3481
rect 5461 3440 5809 3470
rect 5461 3429 5468 3440
rect 5402 3428 5468 3429
rect 5802 3429 5809 3440
rect 5861 3470 5868 3481
rect 6202 3481 6268 3482
rect 6202 3470 6209 3481
rect 5861 3440 6209 3470
rect 5861 3429 5868 3440
rect 5802 3428 5868 3429
rect 6202 3429 6209 3440
rect 6261 3470 6268 3481
rect 6704 3481 6770 3482
rect 6704 3470 6711 3481
rect 6261 3440 6711 3470
rect 6261 3429 6268 3440
rect 6202 3428 6268 3429
rect 6704 3429 6711 3440
rect 6763 3429 6770 3481
rect 6704 3428 6770 3429
rect 2 3411 68 3412
rect 2 3400 9 3411
rect 0 3370 9 3400
rect 2 3359 9 3370
rect 61 3400 68 3411
rect 402 3411 468 3412
rect 402 3400 409 3411
rect 61 3370 409 3400
rect 61 3359 68 3370
rect 2 3358 68 3359
rect 402 3359 409 3370
rect 461 3400 468 3411
rect 802 3411 868 3412
rect 802 3400 809 3411
rect 461 3370 809 3400
rect 461 3359 468 3370
rect 402 3358 468 3359
rect 802 3359 809 3370
rect 861 3400 868 3411
rect 1202 3411 1268 3412
rect 1202 3400 1209 3411
rect 861 3370 1209 3400
rect 861 3359 868 3370
rect 802 3358 868 3359
rect 1202 3359 1209 3370
rect 1261 3400 1268 3411
rect 1602 3411 1668 3412
rect 1602 3400 1609 3411
rect 1261 3370 1609 3400
rect 1261 3359 1268 3370
rect 1202 3358 1268 3359
rect 1602 3359 1609 3370
rect 1661 3400 1668 3411
rect 2002 3411 2068 3412
rect 2002 3400 2009 3411
rect 1661 3370 2009 3400
rect 1661 3359 1668 3370
rect 1602 3358 1668 3359
rect 2002 3359 2009 3370
rect 2061 3400 2068 3411
rect 2402 3411 2468 3412
rect 2402 3400 2409 3411
rect 2061 3370 2409 3400
rect 2061 3359 2068 3370
rect 2002 3358 2068 3359
rect 2402 3359 2409 3370
rect 2461 3400 2468 3411
rect 2802 3411 2868 3412
rect 2802 3400 2809 3411
rect 2461 3370 2809 3400
rect 2461 3359 2468 3370
rect 2402 3358 2468 3359
rect 2802 3359 2809 3370
rect 2861 3400 2868 3411
rect 3202 3411 3268 3412
rect 3202 3400 3209 3411
rect 2861 3370 3209 3400
rect 2861 3359 2868 3370
rect 2802 3358 2868 3359
rect 3202 3359 3209 3370
rect 3261 3400 3268 3411
rect 3602 3411 3668 3412
rect 3602 3400 3609 3411
rect 3261 3370 3609 3400
rect 3261 3359 3268 3370
rect 3202 3358 3268 3359
rect 3602 3359 3609 3370
rect 3661 3400 3668 3411
rect 4002 3411 4068 3412
rect 4002 3400 4009 3411
rect 3661 3370 4009 3400
rect 3661 3359 3668 3370
rect 3602 3358 3668 3359
rect 4002 3359 4009 3370
rect 4061 3400 4068 3411
rect 4402 3411 4468 3412
rect 4402 3400 4409 3411
rect 4061 3370 4409 3400
rect 4061 3359 4068 3370
rect 4002 3358 4068 3359
rect 4402 3359 4409 3370
rect 4461 3400 4468 3411
rect 4802 3411 4868 3412
rect 4802 3400 4809 3411
rect 4461 3370 4809 3400
rect 4461 3359 4468 3370
rect 4402 3358 4468 3359
rect 4802 3359 4809 3370
rect 4861 3400 4868 3411
rect 5202 3411 5268 3412
rect 5202 3400 5209 3411
rect 4861 3370 5209 3400
rect 4861 3359 4868 3370
rect 4802 3358 4868 3359
rect 5202 3359 5209 3370
rect 5261 3400 5268 3411
rect 5602 3411 5668 3412
rect 5602 3400 5609 3411
rect 5261 3370 5609 3400
rect 5261 3359 5268 3370
rect 5202 3358 5268 3359
rect 5602 3359 5609 3370
rect 5661 3400 5668 3411
rect 6002 3411 6068 3412
rect 6002 3400 6009 3411
rect 5661 3370 6009 3400
rect 5661 3359 5668 3370
rect 5602 3358 5668 3359
rect 6002 3359 6009 3370
rect 6061 3400 6068 3411
rect 6402 3411 6468 3412
rect 6402 3400 6409 3411
rect 6061 3370 6409 3400
rect 6061 3359 6068 3370
rect 6002 3358 6068 3359
rect 6402 3359 6409 3370
rect 6461 3400 6468 3411
rect 6500 3411 6566 3412
rect 6500 3400 6507 3411
rect 6461 3370 6507 3400
rect 6461 3359 6468 3370
rect 6402 3358 6468 3359
rect 6500 3359 6507 3370
rect 6559 3359 6566 3411
rect 6500 3358 6566 3359
rect 202 3341 268 3342
rect 202 3330 209 3341
rect 0 3300 209 3330
rect 202 3289 209 3300
rect 261 3330 268 3341
rect 602 3341 668 3342
rect 602 3330 609 3341
rect 261 3300 609 3330
rect 261 3289 268 3300
rect 202 3288 268 3289
rect 602 3289 609 3300
rect 661 3330 668 3341
rect 1002 3341 1068 3342
rect 1002 3330 1009 3341
rect 661 3300 1009 3330
rect 661 3289 668 3300
rect 602 3288 668 3289
rect 1002 3289 1009 3300
rect 1061 3330 1068 3341
rect 1402 3341 1468 3342
rect 1402 3330 1409 3341
rect 1061 3300 1409 3330
rect 1061 3289 1068 3300
rect 1002 3288 1068 3289
rect 1402 3289 1409 3300
rect 1461 3330 1468 3341
rect 1802 3341 1868 3342
rect 1802 3330 1809 3341
rect 1461 3300 1809 3330
rect 1461 3289 1468 3300
rect 1402 3288 1468 3289
rect 1802 3289 1809 3300
rect 1861 3330 1868 3341
rect 2202 3341 2268 3342
rect 2202 3330 2209 3341
rect 1861 3300 2209 3330
rect 1861 3289 1868 3300
rect 1802 3288 1868 3289
rect 2202 3289 2209 3300
rect 2261 3330 2268 3341
rect 2602 3341 2668 3342
rect 2602 3330 2609 3341
rect 2261 3300 2609 3330
rect 2261 3289 2268 3300
rect 2202 3288 2268 3289
rect 2602 3289 2609 3300
rect 2661 3330 2668 3341
rect 3002 3341 3068 3342
rect 3002 3330 3009 3341
rect 2661 3300 3009 3330
rect 2661 3289 2668 3300
rect 2602 3288 2668 3289
rect 3002 3289 3009 3300
rect 3061 3330 3068 3341
rect 3402 3341 3468 3342
rect 3402 3330 3409 3341
rect 3061 3300 3409 3330
rect 3061 3289 3068 3300
rect 3002 3288 3068 3289
rect 3402 3289 3409 3300
rect 3461 3330 3468 3341
rect 3802 3341 3868 3342
rect 3802 3330 3809 3341
rect 3461 3300 3809 3330
rect 3461 3289 3468 3300
rect 3402 3288 3468 3289
rect 3802 3289 3809 3300
rect 3861 3330 3868 3341
rect 4202 3341 4268 3342
rect 4202 3330 4209 3341
rect 3861 3300 4209 3330
rect 3861 3289 3868 3300
rect 3802 3288 3868 3289
rect 4202 3289 4209 3300
rect 4261 3330 4268 3341
rect 4602 3341 4668 3342
rect 4602 3330 4609 3341
rect 4261 3300 4609 3330
rect 4261 3289 4268 3300
rect 4202 3288 4268 3289
rect 4602 3289 4609 3300
rect 4661 3330 4668 3341
rect 5002 3341 5068 3342
rect 5002 3330 5009 3341
rect 4661 3300 5009 3330
rect 4661 3289 4668 3300
rect 4602 3288 4668 3289
rect 5002 3289 5009 3300
rect 5061 3330 5068 3341
rect 5402 3341 5468 3342
rect 5402 3330 5409 3341
rect 5061 3300 5409 3330
rect 5061 3289 5068 3300
rect 5002 3288 5068 3289
rect 5402 3289 5409 3300
rect 5461 3330 5468 3341
rect 5802 3341 5868 3342
rect 5802 3330 5809 3341
rect 5461 3300 5809 3330
rect 5461 3289 5468 3300
rect 5402 3288 5468 3289
rect 5802 3289 5809 3300
rect 5861 3330 5868 3341
rect 6202 3341 6268 3342
rect 6202 3330 6209 3341
rect 5861 3300 6209 3330
rect 5861 3289 5868 3300
rect 5802 3288 5868 3289
rect 6202 3289 6209 3300
rect 6261 3330 6268 3341
rect 6704 3341 6770 3342
rect 6704 3330 6711 3341
rect 6261 3300 6711 3330
rect 6261 3289 6268 3300
rect 6202 3288 6268 3289
rect 6704 3289 6711 3300
rect 6763 3289 6770 3341
rect 6704 3288 6770 3289
rect 2 3271 68 3272
rect 2 3260 9 3271
rect 0 3230 9 3260
rect 2 3219 9 3230
rect 61 3260 68 3271
rect 402 3271 468 3272
rect 402 3260 409 3271
rect 61 3230 409 3260
rect 61 3219 68 3230
rect 2 3218 68 3219
rect 402 3219 409 3230
rect 461 3260 468 3271
rect 802 3271 868 3272
rect 802 3260 809 3271
rect 461 3230 809 3260
rect 461 3219 468 3230
rect 402 3218 468 3219
rect 802 3219 809 3230
rect 861 3260 868 3271
rect 1202 3271 1268 3272
rect 1202 3260 1209 3271
rect 861 3230 1209 3260
rect 861 3219 868 3230
rect 802 3218 868 3219
rect 1202 3219 1209 3230
rect 1261 3260 1268 3271
rect 1602 3271 1668 3272
rect 1602 3260 1609 3271
rect 1261 3230 1609 3260
rect 1261 3219 1268 3230
rect 1202 3218 1268 3219
rect 1602 3219 1609 3230
rect 1661 3260 1668 3271
rect 2002 3271 2068 3272
rect 2002 3260 2009 3271
rect 1661 3230 2009 3260
rect 1661 3219 1668 3230
rect 1602 3218 1668 3219
rect 2002 3219 2009 3230
rect 2061 3260 2068 3271
rect 2402 3271 2468 3272
rect 2402 3260 2409 3271
rect 2061 3230 2409 3260
rect 2061 3219 2068 3230
rect 2002 3218 2068 3219
rect 2402 3219 2409 3230
rect 2461 3260 2468 3271
rect 2802 3271 2868 3272
rect 2802 3260 2809 3271
rect 2461 3230 2809 3260
rect 2461 3219 2468 3230
rect 2402 3218 2468 3219
rect 2802 3219 2809 3230
rect 2861 3260 2868 3271
rect 3202 3271 3268 3272
rect 3202 3260 3209 3271
rect 2861 3230 3209 3260
rect 2861 3219 2868 3230
rect 2802 3218 2868 3219
rect 3202 3219 3209 3230
rect 3261 3260 3268 3271
rect 3602 3271 3668 3272
rect 3602 3260 3609 3271
rect 3261 3230 3609 3260
rect 3261 3219 3268 3230
rect 3202 3218 3268 3219
rect 3602 3219 3609 3230
rect 3661 3260 3668 3271
rect 4002 3271 4068 3272
rect 4002 3260 4009 3271
rect 3661 3230 4009 3260
rect 3661 3219 3668 3230
rect 3602 3218 3668 3219
rect 4002 3219 4009 3230
rect 4061 3260 4068 3271
rect 4402 3271 4468 3272
rect 4402 3260 4409 3271
rect 4061 3230 4409 3260
rect 4061 3219 4068 3230
rect 4002 3218 4068 3219
rect 4402 3219 4409 3230
rect 4461 3260 4468 3271
rect 4802 3271 4868 3272
rect 4802 3260 4809 3271
rect 4461 3230 4809 3260
rect 4461 3219 4468 3230
rect 4402 3218 4468 3219
rect 4802 3219 4809 3230
rect 4861 3260 4868 3271
rect 5202 3271 5268 3272
rect 5202 3260 5209 3271
rect 4861 3230 5209 3260
rect 4861 3219 4868 3230
rect 4802 3218 4868 3219
rect 5202 3219 5209 3230
rect 5261 3260 5268 3271
rect 5602 3271 5668 3272
rect 5602 3260 5609 3271
rect 5261 3230 5609 3260
rect 5261 3219 5268 3230
rect 5202 3218 5268 3219
rect 5602 3219 5609 3230
rect 5661 3260 5668 3271
rect 6002 3271 6068 3272
rect 6002 3260 6009 3271
rect 5661 3230 6009 3260
rect 5661 3219 5668 3230
rect 5602 3218 5668 3219
rect 6002 3219 6009 3230
rect 6061 3260 6068 3271
rect 6402 3271 6468 3272
rect 6402 3260 6409 3271
rect 6061 3230 6409 3260
rect 6061 3219 6068 3230
rect 6002 3218 6068 3219
rect 6402 3219 6409 3230
rect 6461 3260 6468 3271
rect 6500 3271 6566 3272
rect 6500 3260 6507 3271
rect 6461 3230 6507 3260
rect 6461 3219 6468 3230
rect 6402 3218 6468 3219
rect 6500 3219 6507 3230
rect 6559 3219 6566 3271
rect 6500 3218 6566 3219
rect 202 3201 268 3202
rect 202 3190 209 3201
rect 0 3160 209 3190
rect 202 3149 209 3160
rect 261 3190 268 3201
rect 602 3201 668 3202
rect 602 3190 609 3201
rect 261 3160 609 3190
rect 261 3149 268 3160
rect 202 3148 268 3149
rect 602 3149 609 3160
rect 661 3190 668 3201
rect 1002 3201 1068 3202
rect 1002 3190 1009 3201
rect 661 3160 1009 3190
rect 661 3149 668 3160
rect 602 3148 668 3149
rect 1002 3149 1009 3160
rect 1061 3190 1068 3201
rect 1402 3201 1468 3202
rect 1402 3190 1409 3201
rect 1061 3160 1409 3190
rect 1061 3149 1068 3160
rect 1002 3148 1068 3149
rect 1402 3149 1409 3160
rect 1461 3190 1468 3201
rect 1802 3201 1868 3202
rect 1802 3190 1809 3201
rect 1461 3160 1809 3190
rect 1461 3149 1468 3160
rect 1402 3148 1468 3149
rect 1802 3149 1809 3160
rect 1861 3190 1868 3201
rect 2202 3201 2268 3202
rect 2202 3190 2209 3201
rect 1861 3160 2209 3190
rect 1861 3149 1868 3160
rect 1802 3148 1868 3149
rect 2202 3149 2209 3160
rect 2261 3190 2268 3201
rect 2602 3201 2668 3202
rect 2602 3190 2609 3201
rect 2261 3160 2609 3190
rect 2261 3149 2268 3160
rect 2202 3148 2268 3149
rect 2602 3149 2609 3160
rect 2661 3190 2668 3201
rect 3002 3201 3068 3202
rect 3002 3190 3009 3201
rect 2661 3160 3009 3190
rect 2661 3149 2668 3160
rect 2602 3148 2668 3149
rect 3002 3149 3009 3160
rect 3061 3190 3068 3201
rect 3402 3201 3468 3202
rect 3402 3190 3409 3201
rect 3061 3160 3409 3190
rect 3061 3149 3068 3160
rect 3002 3148 3068 3149
rect 3402 3149 3409 3160
rect 3461 3190 3468 3201
rect 3802 3201 3868 3202
rect 3802 3190 3809 3201
rect 3461 3160 3809 3190
rect 3461 3149 3468 3160
rect 3402 3148 3468 3149
rect 3802 3149 3809 3160
rect 3861 3190 3868 3201
rect 4202 3201 4268 3202
rect 4202 3190 4209 3201
rect 3861 3160 4209 3190
rect 3861 3149 3868 3160
rect 3802 3148 3868 3149
rect 4202 3149 4209 3160
rect 4261 3190 4268 3201
rect 4602 3201 4668 3202
rect 4602 3190 4609 3201
rect 4261 3160 4609 3190
rect 4261 3149 4268 3160
rect 4202 3148 4268 3149
rect 4602 3149 4609 3160
rect 4661 3190 4668 3201
rect 5002 3201 5068 3202
rect 5002 3190 5009 3201
rect 4661 3160 5009 3190
rect 4661 3149 4668 3160
rect 4602 3148 4668 3149
rect 5002 3149 5009 3160
rect 5061 3190 5068 3201
rect 5402 3201 5468 3202
rect 5402 3190 5409 3201
rect 5061 3160 5409 3190
rect 5061 3149 5068 3160
rect 5002 3148 5068 3149
rect 5402 3149 5409 3160
rect 5461 3190 5468 3201
rect 5802 3201 5868 3202
rect 5802 3190 5809 3201
rect 5461 3160 5809 3190
rect 5461 3149 5468 3160
rect 5402 3148 5468 3149
rect 5802 3149 5809 3160
rect 5861 3190 5868 3201
rect 6202 3201 6268 3202
rect 6202 3190 6209 3201
rect 5861 3160 6209 3190
rect 5861 3149 5868 3160
rect 5802 3148 5868 3149
rect 6202 3149 6209 3160
rect 6261 3190 6268 3201
rect 6704 3201 6770 3202
rect 6704 3190 6711 3201
rect 6261 3160 6711 3190
rect 6261 3149 6268 3160
rect 6202 3148 6268 3149
rect 6704 3149 6711 3160
rect 6763 3149 6770 3201
rect 6704 3148 6770 3149
rect 2 3131 68 3132
rect 2 3120 9 3131
rect 0 3090 9 3120
rect 2 3079 9 3090
rect 61 3120 68 3131
rect 402 3131 468 3132
rect 402 3120 409 3131
rect 61 3090 409 3120
rect 61 3079 68 3090
rect 2 3078 68 3079
rect 402 3079 409 3090
rect 461 3120 468 3131
rect 802 3131 868 3132
rect 802 3120 809 3131
rect 461 3090 809 3120
rect 461 3079 468 3090
rect 402 3078 468 3079
rect 802 3079 809 3090
rect 861 3120 868 3131
rect 1202 3131 1268 3132
rect 1202 3120 1209 3131
rect 861 3090 1209 3120
rect 861 3079 868 3090
rect 802 3078 868 3079
rect 1202 3079 1209 3090
rect 1261 3120 1268 3131
rect 1602 3131 1668 3132
rect 1602 3120 1609 3131
rect 1261 3090 1609 3120
rect 1261 3079 1268 3090
rect 1202 3078 1268 3079
rect 1602 3079 1609 3090
rect 1661 3120 1668 3131
rect 2002 3131 2068 3132
rect 2002 3120 2009 3131
rect 1661 3090 2009 3120
rect 1661 3079 1668 3090
rect 1602 3078 1668 3079
rect 2002 3079 2009 3090
rect 2061 3120 2068 3131
rect 2402 3131 2468 3132
rect 2402 3120 2409 3131
rect 2061 3090 2409 3120
rect 2061 3079 2068 3090
rect 2002 3078 2068 3079
rect 2402 3079 2409 3090
rect 2461 3120 2468 3131
rect 2802 3131 2868 3132
rect 2802 3120 2809 3131
rect 2461 3090 2809 3120
rect 2461 3079 2468 3090
rect 2402 3078 2468 3079
rect 2802 3079 2809 3090
rect 2861 3120 2868 3131
rect 3202 3131 3268 3132
rect 3202 3120 3209 3131
rect 2861 3090 3209 3120
rect 2861 3079 2868 3090
rect 2802 3078 2868 3079
rect 3202 3079 3209 3090
rect 3261 3120 3268 3131
rect 3602 3131 3668 3132
rect 3602 3120 3609 3131
rect 3261 3090 3609 3120
rect 3261 3079 3268 3090
rect 3202 3078 3268 3079
rect 3602 3079 3609 3090
rect 3661 3120 3668 3131
rect 4002 3131 4068 3132
rect 4002 3120 4009 3131
rect 3661 3090 4009 3120
rect 3661 3079 3668 3090
rect 3602 3078 3668 3079
rect 4002 3079 4009 3090
rect 4061 3120 4068 3131
rect 4402 3131 4468 3132
rect 4402 3120 4409 3131
rect 4061 3090 4409 3120
rect 4061 3079 4068 3090
rect 4002 3078 4068 3079
rect 4402 3079 4409 3090
rect 4461 3120 4468 3131
rect 4802 3131 4868 3132
rect 4802 3120 4809 3131
rect 4461 3090 4809 3120
rect 4461 3079 4468 3090
rect 4402 3078 4468 3079
rect 4802 3079 4809 3090
rect 4861 3120 4868 3131
rect 5202 3131 5268 3132
rect 5202 3120 5209 3131
rect 4861 3090 5209 3120
rect 4861 3079 4868 3090
rect 4802 3078 4868 3079
rect 5202 3079 5209 3090
rect 5261 3120 5268 3131
rect 5602 3131 5668 3132
rect 5602 3120 5609 3131
rect 5261 3090 5609 3120
rect 5261 3079 5268 3090
rect 5202 3078 5268 3079
rect 5602 3079 5609 3090
rect 5661 3120 5668 3131
rect 6002 3131 6068 3132
rect 6002 3120 6009 3131
rect 5661 3090 6009 3120
rect 5661 3079 5668 3090
rect 5602 3078 5668 3079
rect 6002 3079 6009 3090
rect 6061 3120 6068 3131
rect 6402 3131 6468 3132
rect 6402 3120 6409 3131
rect 6061 3090 6409 3120
rect 6061 3079 6068 3090
rect 6002 3078 6068 3079
rect 6402 3079 6409 3090
rect 6461 3120 6468 3131
rect 6500 3131 6566 3132
rect 6500 3120 6507 3131
rect 6461 3090 6507 3120
rect 6461 3079 6468 3090
rect 6402 3078 6468 3079
rect 6500 3079 6507 3090
rect 6559 3079 6566 3131
rect 6500 3078 6566 3079
rect 202 3061 268 3062
rect 202 3050 209 3061
rect 0 3020 209 3050
rect 202 3009 209 3020
rect 261 3050 268 3061
rect 602 3061 668 3062
rect 602 3050 609 3061
rect 261 3020 609 3050
rect 261 3009 268 3020
rect 202 3008 268 3009
rect 602 3009 609 3020
rect 661 3050 668 3061
rect 1002 3061 1068 3062
rect 1002 3050 1009 3061
rect 661 3020 1009 3050
rect 661 3009 668 3020
rect 602 3008 668 3009
rect 1002 3009 1009 3020
rect 1061 3050 1068 3061
rect 1402 3061 1468 3062
rect 1402 3050 1409 3061
rect 1061 3020 1409 3050
rect 1061 3009 1068 3020
rect 1002 3008 1068 3009
rect 1402 3009 1409 3020
rect 1461 3050 1468 3061
rect 1802 3061 1868 3062
rect 1802 3050 1809 3061
rect 1461 3020 1809 3050
rect 1461 3009 1468 3020
rect 1402 3008 1468 3009
rect 1802 3009 1809 3020
rect 1861 3050 1868 3061
rect 2202 3061 2268 3062
rect 2202 3050 2209 3061
rect 1861 3020 2209 3050
rect 1861 3009 1868 3020
rect 1802 3008 1868 3009
rect 2202 3009 2209 3020
rect 2261 3050 2268 3061
rect 2602 3061 2668 3062
rect 2602 3050 2609 3061
rect 2261 3020 2609 3050
rect 2261 3009 2268 3020
rect 2202 3008 2268 3009
rect 2602 3009 2609 3020
rect 2661 3050 2668 3061
rect 3002 3061 3068 3062
rect 3002 3050 3009 3061
rect 2661 3020 3009 3050
rect 2661 3009 2668 3020
rect 2602 3008 2668 3009
rect 3002 3009 3009 3020
rect 3061 3050 3068 3061
rect 3402 3061 3468 3062
rect 3402 3050 3409 3061
rect 3061 3020 3409 3050
rect 3061 3009 3068 3020
rect 3002 3008 3068 3009
rect 3402 3009 3409 3020
rect 3461 3050 3468 3061
rect 3802 3061 3868 3062
rect 3802 3050 3809 3061
rect 3461 3020 3809 3050
rect 3461 3009 3468 3020
rect 3402 3008 3468 3009
rect 3802 3009 3809 3020
rect 3861 3050 3868 3061
rect 4202 3061 4268 3062
rect 4202 3050 4209 3061
rect 3861 3020 4209 3050
rect 3861 3009 3868 3020
rect 3802 3008 3868 3009
rect 4202 3009 4209 3020
rect 4261 3050 4268 3061
rect 4602 3061 4668 3062
rect 4602 3050 4609 3061
rect 4261 3020 4609 3050
rect 4261 3009 4268 3020
rect 4202 3008 4268 3009
rect 4602 3009 4609 3020
rect 4661 3050 4668 3061
rect 5002 3061 5068 3062
rect 5002 3050 5009 3061
rect 4661 3020 5009 3050
rect 4661 3009 4668 3020
rect 4602 3008 4668 3009
rect 5002 3009 5009 3020
rect 5061 3050 5068 3061
rect 5402 3061 5468 3062
rect 5402 3050 5409 3061
rect 5061 3020 5409 3050
rect 5061 3009 5068 3020
rect 5002 3008 5068 3009
rect 5402 3009 5409 3020
rect 5461 3050 5468 3061
rect 5802 3061 5868 3062
rect 5802 3050 5809 3061
rect 5461 3020 5809 3050
rect 5461 3009 5468 3020
rect 5402 3008 5468 3009
rect 5802 3009 5809 3020
rect 5861 3050 5868 3061
rect 6202 3061 6268 3062
rect 6202 3050 6209 3061
rect 5861 3020 6209 3050
rect 5861 3009 5868 3020
rect 5802 3008 5868 3009
rect 6202 3009 6209 3020
rect 6261 3050 6268 3061
rect 6704 3061 6770 3062
rect 6704 3050 6711 3061
rect 6261 3020 6711 3050
rect 6261 3009 6268 3020
rect 6202 3008 6268 3009
rect 6704 3009 6711 3020
rect 6763 3009 6770 3061
rect 6704 3008 6770 3009
rect 2 2991 68 2992
rect 2 2980 9 2991
rect 0 2950 9 2980
rect 2 2939 9 2950
rect 61 2980 68 2991
rect 402 2991 468 2992
rect 402 2980 409 2991
rect 61 2950 409 2980
rect 61 2939 68 2950
rect 2 2938 68 2939
rect 402 2939 409 2950
rect 461 2980 468 2991
rect 802 2991 868 2992
rect 802 2980 809 2991
rect 461 2950 809 2980
rect 461 2939 468 2950
rect 402 2938 468 2939
rect 802 2939 809 2950
rect 861 2980 868 2991
rect 1202 2991 1268 2992
rect 1202 2980 1209 2991
rect 861 2950 1209 2980
rect 861 2939 868 2950
rect 802 2938 868 2939
rect 1202 2939 1209 2950
rect 1261 2980 1268 2991
rect 1602 2991 1668 2992
rect 1602 2980 1609 2991
rect 1261 2950 1609 2980
rect 1261 2939 1268 2950
rect 1202 2938 1268 2939
rect 1602 2939 1609 2950
rect 1661 2980 1668 2991
rect 2002 2991 2068 2992
rect 2002 2980 2009 2991
rect 1661 2950 2009 2980
rect 1661 2939 1668 2950
rect 1602 2938 1668 2939
rect 2002 2939 2009 2950
rect 2061 2980 2068 2991
rect 2402 2991 2468 2992
rect 2402 2980 2409 2991
rect 2061 2950 2409 2980
rect 2061 2939 2068 2950
rect 2002 2938 2068 2939
rect 2402 2939 2409 2950
rect 2461 2980 2468 2991
rect 2802 2991 2868 2992
rect 2802 2980 2809 2991
rect 2461 2950 2809 2980
rect 2461 2939 2468 2950
rect 2402 2938 2468 2939
rect 2802 2939 2809 2950
rect 2861 2980 2868 2991
rect 3202 2991 3268 2992
rect 3202 2980 3209 2991
rect 2861 2950 3209 2980
rect 2861 2939 2868 2950
rect 2802 2938 2868 2939
rect 3202 2939 3209 2950
rect 3261 2980 3268 2991
rect 3602 2991 3668 2992
rect 3602 2980 3609 2991
rect 3261 2950 3609 2980
rect 3261 2939 3268 2950
rect 3202 2938 3268 2939
rect 3602 2939 3609 2950
rect 3661 2980 3668 2991
rect 4002 2991 4068 2992
rect 4002 2980 4009 2991
rect 3661 2950 4009 2980
rect 3661 2939 3668 2950
rect 3602 2938 3668 2939
rect 4002 2939 4009 2950
rect 4061 2980 4068 2991
rect 4402 2991 4468 2992
rect 4402 2980 4409 2991
rect 4061 2950 4409 2980
rect 4061 2939 4068 2950
rect 4002 2938 4068 2939
rect 4402 2939 4409 2950
rect 4461 2980 4468 2991
rect 4802 2991 4868 2992
rect 4802 2980 4809 2991
rect 4461 2950 4809 2980
rect 4461 2939 4468 2950
rect 4402 2938 4468 2939
rect 4802 2939 4809 2950
rect 4861 2980 4868 2991
rect 5202 2991 5268 2992
rect 5202 2980 5209 2991
rect 4861 2950 5209 2980
rect 4861 2939 4868 2950
rect 4802 2938 4868 2939
rect 5202 2939 5209 2950
rect 5261 2980 5268 2991
rect 5602 2991 5668 2992
rect 5602 2980 5609 2991
rect 5261 2950 5609 2980
rect 5261 2939 5268 2950
rect 5202 2938 5268 2939
rect 5602 2939 5609 2950
rect 5661 2980 5668 2991
rect 6002 2991 6068 2992
rect 6002 2980 6009 2991
rect 5661 2950 6009 2980
rect 5661 2939 5668 2950
rect 5602 2938 5668 2939
rect 6002 2939 6009 2950
rect 6061 2980 6068 2991
rect 6402 2991 6468 2992
rect 6402 2980 6409 2991
rect 6061 2950 6409 2980
rect 6061 2939 6068 2950
rect 6002 2938 6068 2939
rect 6402 2939 6409 2950
rect 6461 2980 6468 2991
rect 6500 2991 6566 2992
rect 6500 2980 6507 2991
rect 6461 2950 6507 2980
rect 6461 2939 6468 2950
rect 6402 2938 6468 2939
rect 6500 2939 6507 2950
rect 6559 2939 6566 2991
rect 6500 2938 6566 2939
rect 202 2921 268 2922
rect 202 2910 209 2921
rect 0 2880 209 2910
rect 202 2869 209 2880
rect 261 2910 268 2921
rect 602 2921 668 2922
rect 602 2910 609 2921
rect 261 2880 609 2910
rect 261 2869 268 2880
rect 202 2868 268 2869
rect 602 2869 609 2880
rect 661 2910 668 2921
rect 1002 2921 1068 2922
rect 1002 2910 1009 2921
rect 661 2880 1009 2910
rect 661 2869 668 2880
rect 602 2868 668 2869
rect 1002 2869 1009 2880
rect 1061 2910 1068 2921
rect 1402 2921 1468 2922
rect 1402 2910 1409 2921
rect 1061 2880 1409 2910
rect 1061 2869 1068 2880
rect 1002 2868 1068 2869
rect 1402 2869 1409 2880
rect 1461 2910 1468 2921
rect 1802 2921 1868 2922
rect 1802 2910 1809 2921
rect 1461 2880 1809 2910
rect 1461 2869 1468 2880
rect 1402 2868 1468 2869
rect 1802 2869 1809 2880
rect 1861 2910 1868 2921
rect 2202 2921 2268 2922
rect 2202 2910 2209 2921
rect 1861 2880 2209 2910
rect 1861 2869 1868 2880
rect 1802 2868 1868 2869
rect 2202 2869 2209 2880
rect 2261 2910 2268 2921
rect 2602 2921 2668 2922
rect 2602 2910 2609 2921
rect 2261 2880 2609 2910
rect 2261 2869 2268 2880
rect 2202 2868 2268 2869
rect 2602 2869 2609 2880
rect 2661 2910 2668 2921
rect 3002 2921 3068 2922
rect 3002 2910 3009 2921
rect 2661 2880 3009 2910
rect 2661 2869 2668 2880
rect 2602 2868 2668 2869
rect 3002 2869 3009 2880
rect 3061 2910 3068 2921
rect 3402 2921 3468 2922
rect 3402 2910 3409 2921
rect 3061 2880 3409 2910
rect 3061 2869 3068 2880
rect 3002 2868 3068 2869
rect 3402 2869 3409 2880
rect 3461 2910 3468 2921
rect 3802 2921 3868 2922
rect 3802 2910 3809 2921
rect 3461 2880 3809 2910
rect 3461 2869 3468 2880
rect 3402 2868 3468 2869
rect 3802 2869 3809 2880
rect 3861 2910 3868 2921
rect 4202 2921 4268 2922
rect 4202 2910 4209 2921
rect 3861 2880 4209 2910
rect 3861 2869 3868 2880
rect 3802 2868 3868 2869
rect 4202 2869 4209 2880
rect 4261 2910 4268 2921
rect 4602 2921 4668 2922
rect 4602 2910 4609 2921
rect 4261 2880 4609 2910
rect 4261 2869 4268 2880
rect 4202 2868 4268 2869
rect 4602 2869 4609 2880
rect 4661 2910 4668 2921
rect 5002 2921 5068 2922
rect 5002 2910 5009 2921
rect 4661 2880 5009 2910
rect 4661 2869 4668 2880
rect 4602 2868 4668 2869
rect 5002 2869 5009 2880
rect 5061 2910 5068 2921
rect 5402 2921 5468 2922
rect 5402 2910 5409 2921
rect 5061 2880 5409 2910
rect 5061 2869 5068 2880
rect 5002 2868 5068 2869
rect 5402 2869 5409 2880
rect 5461 2910 5468 2921
rect 5802 2921 5868 2922
rect 5802 2910 5809 2921
rect 5461 2880 5809 2910
rect 5461 2869 5468 2880
rect 5402 2868 5468 2869
rect 5802 2869 5809 2880
rect 5861 2910 5868 2921
rect 6202 2921 6268 2922
rect 6202 2910 6209 2921
rect 5861 2880 6209 2910
rect 5861 2869 5868 2880
rect 5802 2868 5868 2869
rect 6202 2869 6209 2880
rect 6261 2910 6268 2921
rect 6704 2921 6770 2922
rect 6704 2910 6711 2921
rect 6261 2880 6711 2910
rect 6261 2869 6268 2880
rect 6202 2868 6268 2869
rect 6704 2869 6711 2880
rect 6763 2869 6770 2921
rect 6704 2868 6770 2869
rect 2 2851 68 2852
rect 2 2840 9 2851
rect 0 2810 9 2840
rect 2 2799 9 2810
rect 61 2840 68 2851
rect 402 2851 468 2852
rect 402 2840 409 2851
rect 61 2810 409 2840
rect 61 2799 68 2810
rect 2 2798 68 2799
rect 402 2799 409 2810
rect 461 2840 468 2851
rect 802 2851 868 2852
rect 802 2840 809 2851
rect 461 2810 809 2840
rect 461 2799 468 2810
rect 402 2798 468 2799
rect 802 2799 809 2810
rect 861 2840 868 2851
rect 1202 2851 1268 2852
rect 1202 2840 1209 2851
rect 861 2810 1209 2840
rect 861 2799 868 2810
rect 802 2798 868 2799
rect 1202 2799 1209 2810
rect 1261 2840 1268 2851
rect 1602 2851 1668 2852
rect 1602 2840 1609 2851
rect 1261 2810 1609 2840
rect 1261 2799 1268 2810
rect 1202 2798 1268 2799
rect 1602 2799 1609 2810
rect 1661 2840 1668 2851
rect 2002 2851 2068 2852
rect 2002 2840 2009 2851
rect 1661 2810 2009 2840
rect 1661 2799 1668 2810
rect 1602 2798 1668 2799
rect 2002 2799 2009 2810
rect 2061 2840 2068 2851
rect 2402 2851 2468 2852
rect 2402 2840 2409 2851
rect 2061 2810 2409 2840
rect 2061 2799 2068 2810
rect 2002 2798 2068 2799
rect 2402 2799 2409 2810
rect 2461 2840 2468 2851
rect 2802 2851 2868 2852
rect 2802 2840 2809 2851
rect 2461 2810 2809 2840
rect 2461 2799 2468 2810
rect 2402 2798 2468 2799
rect 2802 2799 2809 2810
rect 2861 2840 2868 2851
rect 3202 2851 3268 2852
rect 3202 2840 3209 2851
rect 2861 2810 3209 2840
rect 2861 2799 2868 2810
rect 2802 2798 2868 2799
rect 3202 2799 3209 2810
rect 3261 2840 3268 2851
rect 3602 2851 3668 2852
rect 3602 2840 3609 2851
rect 3261 2810 3609 2840
rect 3261 2799 3268 2810
rect 3202 2798 3268 2799
rect 3602 2799 3609 2810
rect 3661 2840 3668 2851
rect 4002 2851 4068 2852
rect 4002 2840 4009 2851
rect 3661 2810 4009 2840
rect 3661 2799 3668 2810
rect 3602 2798 3668 2799
rect 4002 2799 4009 2810
rect 4061 2840 4068 2851
rect 4402 2851 4468 2852
rect 4402 2840 4409 2851
rect 4061 2810 4409 2840
rect 4061 2799 4068 2810
rect 4002 2798 4068 2799
rect 4402 2799 4409 2810
rect 4461 2840 4468 2851
rect 4802 2851 4868 2852
rect 4802 2840 4809 2851
rect 4461 2810 4809 2840
rect 4461 2799 4468 2810
rect 4402 2798 4468 2799
rect 4802 2799 4809 2810
rect 4861 2840 4868 2851
rect 5202 2851 5268 2852
rect 5202 2840 5209 2851
rect 4861 2810 5209 2840
rect 4861 2799 4868 2810
rect 4802 2798 4868 2799
rect 5202 2799 5209 2810
rect 5261 2840 5268 2851
rect 5602 2851 5668 2852
rect 5602 2840 5609 2851
rect 5261 2810 5609 2840
rect 5261 2799 5268 2810
rect 5202 2798 5268 2799
rect 5602 2799 5609 2810
rect 5661 2840 5668 2851
rect 6002 2851 6068 2852
rect 6002 2840 6009 2851
rect 5661 2810 6009 2840
rect 5661 2799 5668 2810
rect 5602 2798 5668 2799
rect 6002 2799 6009 2810
rect 6061 2840 6068 2851
rect 6402 2851 6468 2852
rect 6402 2840 6409 2851
rect 6061 2810 6409 2840
rect 6061 2799 6068 2810
rect 6002 2798 6068 2799
rect 6402 2799 6409 2810
rect 6461 2840 6468 2851
rect 6500 2851 6566 2852
rect 6500 2840 6507 2851
rect 6461 2810 6507 2840
rect 6461 2799 6468 2810
rect 6402 2798 6468 2799
rect 6500 2799 6507 2810
rect 6559 2799 6566 2851
rect 6500 2798 6566 2799
rect 202 2781 268 2782
rect 202 2770 209 2781
rect 0 2740 209 2770
rect 202 2729 209 2740
rect 261 2770 268 2781
rect 602 2781 668 2782
rect 602 2770 609 2781
rect 261 2740 609 2770
rect 261 2729 268 2740
rect 202 2728 268 2729
rect 602 2729 609 2740
rect 661 2770 668 2781
rect 1002 2781 1068 2782
rect 1002 2770 1009 2781
rect 661 2740 1009 2770
rect 661 2729 668 2740
rect 602 2728 668 2729
rect 1002 2729 1009 2740
rect 1061 2770 1068 2781
rect 1402 2781 1468 2782
rect 1402 2770 1409 2781
rect 1061 2740 1409 2770
rect 1061 2729 1068 2740
rect 1002 2728 1068 2729
rect 1402 2729 1409 2740
rect 1461 2770 1468 2781
rect 1802 2781 1868 2782
rect 1802 2770 1809 2781
rect 1461 2740 1809 2770
rect 1461 2729 1468 2740
rect 1402 2728 1468 2729
rect 1802 2729 1809 2740
rect 1861 2770 1868 2781
rect 2202 2781 2268 2782
rect 2202 2770 2209 2781
rect 1861 2740 2209 2770
rect 1861 2729 1868 2740
rect 1802 2728 1868 2729
rect 2202 2729 2209 2740
rect 2261 2770 2268 2781
rect 2602 2781 2668 2782
rect 2602 2770 2609 2781
rect 2261 2740 2609 2770
rect 2261 2729 2268 2740
rect 2202 2728 2268 2729
rect 2602 2729 2609 2740
rect 2661 2770 2668 2781
rect 3002 2781 3068 2782
rect 3002 2770 3009 2781
rect 2661 2740 3009 2770
rect 2661 2729 2668 2740
rect 2602 2728 2668 2729
rect 3002 2729 3009 2740
rect 3061 2770 3068 2781
rect 3402 2781 3468 2782
rect 3402 2770 3409 2781
rect 3061 2740 3409 2770
rect 3061 2729 3068 2740
rect 3002 2728 3068 2729
rect 3402 2729 3409 2740
rect 3461 2770 3468 2781
rect 3802 2781 3868 2782
rect 3802 2770 3809 2781
rect 3461 2740 3809 2770
rect 3461 2729 3468 2740
rect 3402 2728 3468 2729
rect 3802 2729 3809 2740
rect 3861 2770 3868 2781
rect 4202 2781 4268 2782
rect 4202 2770 4209 2781
rect 3861 2740 4209 2770
rect 3861 2729 3868 2740
rect 3802 2728 3868 2729
rect 4202 2729 4209 2740
rect 4261 2770 4268 2781
rect 4602 2781 4668 2782
rect 4602 2770 4609 2781
rect 4261 2740 4609 2770
rect 4261 2729 4268 2740
rect 4202 2728 4268 2729
rect 4602 2729 4609 2740
rect 4661 2770 4668 2781
rect 5002 2781 5068 2782
rect 5002 2770 5009 2781
rect 4661 2740 5009 2770
rect 4661 2729 4668 2740
rect 4602 2728 4668 2729
rect 5002 2729 5009 2740
rect 5061 2770 5068 2781
rect 5402 2781 5468 2782
rect 5402 2770 5409 2781
rect 5061 2740 5409 2770
rect 5061 2729 5068 2740
rect 5002 2728 5068 2729
rect 5402 2729 5409 2740
rect 5461 2770 5468 2781
rect 5802 2781 5868 2782
rect 5802 2770 5809 2781
rect 5461 2740 5809 2770
rect 5461 2729 5468 2740
rect 5402 2728 5468 2729
rect 5802 2729 5809 2740
rect 5861 2770 5868 2781
rect 6202 2781 6268 2782
rect 6202 2770 6209 2781
rect 5861 2740 6209 2770
rect 5861 2729 5868 2740
rect 5802 2728 5868 2729
rect 6202 2729 6209 2740
rect 6261 2770 6268 2781
rect 6704 2781 6770 2782
rect 6704 2770 6711 2781
rect 6261 2740 6711 2770
rect 6261 2729 6268 2740
rect 6202 2728 6268 2729
rect 6704 2729 6711 2740
rect 6763 2729 6770 2781
rect 6704 2728 6770 2729
rect 2 2711 68 2712
rect 2 2700 9 2711
rect 0 2670 9 2700
rect 2 2659 9 2670
rect 61 2700 68 2711
rect 402 2711 468 2712
rect 402 2700 409 2711
rect 61 2670 409 2700
rect 61 2659 68 2670
rect 2 2658 68 2659
rect 402 2659 409 2670
rect 461 2700 468 2711
rect 802 2711 868 2712
rect 802 2700 809 2711
rect 461 2670 809 2700
rect 461 2659 468 2670
rect 402 2658 468 2659
rect 802 2659 809 2670
rect 861 2700 868 2711
rect 1202 2711 1268 2712
rect 1202 2700 1209 2711
rect 861 2670 1209 2700
rect 861 2659 868 2670
rect 802 2658 868 2659
rect 1202 2659 1209 2670
rect 1261 2700 1268 2711
rect 1602 2711 1668 2712
rect 1602 2700 1609 2711
rect 1261 2670 1609 2700
rect 1261 2659 1268 2670
rect 1202 2658 1268 2659
rect 1602 2659 1609 2670
rect 1661 2700 1668 2711
rect 2002 2711 2068 2712
rect 2002 2700 2009 2711
rect 1661 2670 2009 2700
rect 1661 2659 1668 2670
rect 1602 2658 1668 2659
rect 2002 2659 2009 2670
rect 2061 2700 2068 2711
rect 2402 2711 2468 2712
rect 2402 2700 2409 2711
rect 2061 2670 2409 2700
rect 2061 2659 2068 2670
rect 2002 2658 2068 2659
rect 2402 2659 2409 2670
rect 2461 2700 2468 2711
rect 2802 2711 2868 2712
rect 2802 2700 2809 2711
rect 2461 2670 2809 2700
rect 2461 2659 2468 2670
rect 2402 2658 2468 2659
rect 2802 2659 2809 2670
rect 2861 2700 2868 2711
rect 3202 2711 3268 2712
rect 3202 2700 3209 2711
rect 2861 2670 3209 2700
rect 2861 2659 2868 2670
rect 2802 2658 2868 2659
rect 3202 2659 3209 2670
rect 3261 2700 3268 2711
rect 3602 2711 3668 2712
rect 3602 2700 3609 2711
rect 3261 2670 3609 2700
rect 3261 2659 3268 2670
rect 3202 2658 3268 2659
rect 3602 2659 3609 2670
rect 3661 2700 3668 2711
rect 4002 2711 4068 2712
rect 4002 2700 4009 2711
rect 3661 2670 4009 2700
rect 3661 2659 3668 2670
rect 3602 2658 3668 2659
rect 4002 2659 4009 2670
rect 4061 2700 4068 2711
rect 4402 2711 4468 2712
rect 4402 2700 4409 2711
rect 4061 2670 4409 2700
rect 4061 2659 4068 2670
rect 4002 2658 4068 2659
rect 4402 2659 4409 2670
rect 4461 2700 4468 2711
rect 4802 2711 4868 2712
rect 4802 2700 4809 2711
rect 4461 2670 4809 2700
rect 4461 2659 4468 2670
rect 4402 2658 4468 2659
rect 4802 2659 4809 2670
rect 4861 2700 4868 2711
rect 5202 2711 5268 2712
rect 5202 2700 5209 2711
rect 4861 2670 5209 2700
rect 4861 2659 4868 2670
rect 4802 2658 4868 2659
rect 5202 2659 5209 2670
rect 5261 2700 5268 2711
rect 5602 2711 5668 2712
rect 5602 2700 5609 2711
rect 5261 2670 5609 2700
rect 5261 2659 5268 2670
rect 5202 2658 5268 2659
rect 5602 2659 5609 2670
rect 5661 2700 5668 2711
rect 6002 2711 6068 2712
rect 6002 2700 6009 2711
rect 5661 2670 6009 2700
rect 5661 2659 5668 2670
rect 5602 2658 5668 2659
rect 6002 2659 6009 2670
rect 6061 2700 6068 2711
rect 6402 2711 6468 2712
rect 6402 2700 6409 2711
rect 6061 2670 6409 2700
rect 6061 2659 6068 2670
rect 6002 2658 6068 2659
rect 6402 2659 6409 2670
rect 6461 2700 6468 2711
rect 6500 2711 6566 2712
rect 6500 2700 6507 2711
rect 6461 2670 6507 2700
rect 6461 2659 6468 2670
rect 6402 2658 6468 2659
rect 6500 2659 6507 2670
rect 6559 2659 6566 2711
rect 6500 2658 6566 2659
rect 202 2641 268 2642
rect 202 2630 209 2641
rect 0 2600 209 2630
rect 202 2589 209 2600
rect 261 2630 268 2641
rect 602 2641 668 2642
rect 602 2630 609 2641
rect 261 2600 609 2630
rect 261 2589 268 2600
rect 202 2588 268 2589
rect 602 2589 609 2600
rect 661 2630 668 2641
rect 1002 2641 1068 2642
rect 1002 2630 1009 2641
rect 661 2600 1009 2630
rect 661 2589 668 2600
rect 602 2588 668 2589
rect 1002 2589 1009 2600
rect 1061 2630 1068 2641
rect 1402 2641 1468 2642
rect 1402 2630 1409 2641
rect 1061 2600 1409 2630
rect 1061 2589 1068 2600
rect 1002 2588 1068 2589
rect 1402 2589 1409 2600
rect 1461 2630 1468 2641
rect 1802 2641 1868 2642
rect 1802 2630 1809 2641
rect 1461 2600 1809 2630
rect 1461 2589 1468 2600
rect 1402 2588 1468 2589
rect 1802 2589 1809 2600
rect 1861 2630 1868 2641
rect 2202 2641 2268 2642
rect 2202 2630 2209 2641
rect 1861 2600 2209 2630
rect 1861 2589 1868 2600
rect 1802 2588 1868 2589
rect 2202 2589 2209 2600
rect 2261 2630 2268 2641
rect 2602 2641 2668 2642
rect 2602 2630 2609 2641
rect 2261 2600 2609 2630
rect 2261 2589 2268 2600
rect 2202 2588 2268 2589
rect 2602 2589 2609 2600
rect 2661 2630 2668 2641
rect 3002 2641 3068 2642
rect 3002 2630 3009 2641
rect 2661 2600 3009 2630
rect 2661 2589 2668 2600
rect 2602 2588 2668 2589
rect 3002 2589 3009 2600
rect 3061 2630 3068 2641
rect 3402 2641 3468 2642
rect 3402 2630 3409 2641
rect 3061 2600 3409 2630
rect 3061 2589 3068 2600
rect 3002 2588 3068 2589
rect 3402 2589 3409 2600
rect 3461 2630 3468 2641
rect 3802 2641 3868 2642
rect 3802 2630 3809 2641
rect 3461 2600 3809 2630
rect 3461 2589 3468 2600
rect 3402 2588 3468 2589
rect 3802 2589 3809 2600
rect 3861 2630 3868 2641
rect 4202 2641 4268 2642
rect 4202 2630 4209 2641
rect 3861 2600 4209 2630
rect 3861 2589 3868 2600
rect 3802 2588 3868 2589
rect 4202 2589 4209 2600
rect 4261 2630 4268 2641
rect 4602 2641 4668 2642
rect 4602 2630 4609 2641
rect 4261 2600 4609 2630
rect 4261 2589 4268 2600
rect 4202 2588 4268 2589
rect 4602 2589 4609 2600
rect 4661 2630 4668 2641
rect 5002 2641 5068 2642
rect 5002 2630 5009 2641
rect 4661 2600 5009 2630
rect 4661 2589 4668 2600
rect 4602 2588 4668 2589
rect 5002 2589 5009 2600
rect 5061 2630 5068 2641
rect 5402 2641 5468 2642
rect 5402 2630 5409 2641
rect 5061 2600 5409 2630
rect 5061 2589 5068 2600
rect 5002 2588 5068 2589
rect 5402 2589 5409 2600
rect 5461 2630 5468 2641
rect 5802 2641 5868 2642
rect 5802 2630 5809 2641
rect 5461 2600 5809 2630
rect 5461 2589 5468 2600
rect 5402 2588 5468 2589
rect 5802 2589 5809 2600
rect 5861 2630 5868 2641
rect 6202 2641 6268 2642
rect 6202 2630 6209 2641
rect 5861 2600 6209 2630
rect 5861 2589 5868 2600
rect 5802 2588 5868 2589
rect 6202 2589 6209 2600
rect 6261 2630 6268 2641
rect 6704 2641 6770 2642
rect 6704 2630 6711 2641
rect 6261 2600 6711 2630
rect 6261 2589 6268 2600
rect 6202 2588 6268 2589
rect 6704 2589 6711 2600
rect 6763 2589 6770 2641
rect 6704 2588 6770 2589
rect 2 2571 68 2572
rect 2 2560 9 2571
rect 0 2530 9 2560
rect 2 2519 9 2530
rect 61 2560 68 2571
rect 402 2571 468 2572
rect 402 2560 409 2571
rect 61 2530 409 2560
rect 61 2519 68 2530
rect 2 2518 68 2519
rect 402 2519 409 2530
rect 461 2560 468 2571
rect 802 2571 868 2572
rect 802 2560 809 2571
rect 461 2530 809 2560
rect 461 2519 468 2530
rect 402 2518 468 2519
rect 802 2519 809 2530
rect 861 2560 868 2571
rect 1202 2571 1268 2572
rect 1202 2560 1209 2571
rect 861 2530 1209 2560
rect 861 2519 868 2530
rect 802 2518 868 2519
rect 1202 2519 1209 2530
rect 1261 2560 1268 2571
rect 1602 2571 1668 2572
rect 1602 2560 1609 2571
rect 1261 2530 1609 2560
rect 1261 2519 1268 2530
rect 1202 2518 1268 2519
rect 1602 2519 1609 2530
rect 1661 2560 1668 2571
rect 2002 2571 2068 2572
rect 2002 2560 2009 2571
rect 1661 2530 2009 2560
rect 1661 2519 1668 2530
rect 1602 2518 1668 2519
rect 2002 2519 2009 2530
rect 2061 2560 2068 2571
rect 2402 2571 2468 2572
rect 2402 2560 2409 2571
rect 2061 2530 2409 2560
rect 2061 2519 2068 2530
rect 2002 2518 2068 2519
rect 2402 2519 2409 2530
rect 2461 2560 2468 2571
rect 2802 2571 2868 2572
rect 2802 2560 2809 2571
rect 2461 2530 2809 2560
rect 2461 2519 2468 2530
rect 2402 2518 2468 2519
rect 2802 2519 2809 2530
rect 2861 2560 2868 2571
rect 3202 2571 3268 2572
rect 3202 2560 3209 2571
rect 2861 2530 3209 2560
rect 2861 2519 2868 2530
rect 2802 2518 2868 2519
rect 3202 2519 3209 2530
rect 3261 2560 3268 2571
rect 3602 2571 3668 2572
rect 3602 2560 3609 2571
rect 3261 2530 3609 2560
rect 3261 2519 3268 2530
rect 3202 2518 3268 2519
rect 3602 2519 3609 2530
rect 3661 2560 3668 2571
rect 4002 2571 4068 2572
rect 4002 2560 4009 2571
rect 3661 2530 4009 2560
rect 3661 2519 3668 2530
rect 3602 2518 3668 2519
rect 4002 2519 4009 2530
rect 4061 2560 4068 2571
rect 4402 2571 4468 2572
rect 4402 2560 4409 2571
rect 4061 2530 4409 2560
rect 4061 2519 4068 2530
rect 4002 2518 4068 2519
rect 4402 2519 4409 2530
rect 4461 2560 4468 2571
rect 4802 2571 4868 2572
rect 4802 2560 4809 2571
rect 4461 2530 4809 2560
rect 4461 2519 4468 2530
rect 4402 2518 4468 2519
rect 4802 2519 4809 2530
rect 4861 2560 4868 2571
rect 5202 2571 5268 2572
rect 5202 2560 5209 2571
rect 4861 2530 5209 2560
rect 4861 2519 4868 2530
rect 4802 2518 4868 2519
rect 5202 2519 5209 2530
rect 5261 2560 5268 2571
rect 5602 2571 5668 2572
rect 5602 2560 5609 2571
rect 5261 2530 5609 2560
rect 5261 2519 5268 2530
rect 5202 2518 5268 2519
rect 5602 2519 5609 2530
rect 5661 2560 5668 2571
rect 6002 2571 6068 2572
rect 6002 2560 6009 2571
rect 5661 2530 6009 2560
rect 5661 2519 5668 2530
rect 5602 2518 5668 2519
rect 6002 2519 6009 2530
rect 6061 2560 6068 2571
rect 6402 2571 6468 2572
rect 6402 2560 6409 2571
rect 6061 2530 6409 2560
rect 6061 2519 6068 2530
rect 6002 2518 6068 2519
rect 6402 2519 6409 2530
rect 6461 2560 6468 2571
rect 6500 2571 6566 2572
rect 6500 2560 6507 2571
rect 6461 2530 6507 2560
rect 6461 2519 6468 2530
rect 6402 2518 6468 2519
rect 6500 2519 6507 2530
rect 6559 2519 6566 2571
rect 6500 2518 6566 2519
rect 196 2501 274 2502
rect -4 2485 74 2486
rect -4 2429 7 2485
rect 63 2429 74 2485
rect 196 2445 207 2501
rect 263 2445 274 2501
rect 596 2501 674 2502
rect 196 2444 274 2445
rect 396 2485 474 2486
rect -4 2428 74 2429
rect 396 2429 407 2485
rect 463 2429 474 2485
rect 596 2445 607 2501
rect 663 2445 674 2501
rect 996 2501 1074 2502
rect 596 2444 674 2445
rect 796 2485 874 2486
rect 396 2428 474 2429
rect 796 2429 807 2485
rect 863 2429 874 2485
rect 996 2445 1007 2501
rect 1063 2445 1074 2501
rect 1396 2501 1474 2502
rect 996 2444 1074 2445
rect 1196 2485 1274 2486
rect 796 2428 874 2429
rect 1196 2429 1207 2485
rect 1263 2429 1274 2485
rect 1396 2445 1407 2501
rect 1463 2445 1474 2501
rect 1796 2501 1874 2502
rect 1396 2444 1474 2445
rect 1596 2485 1674 2486
rect 1196 2428 1274 2429
rect 1596 2429 1607 2485
rect 1663 2429 1674 2485
rect 1796 2445 1807 2501
rect 1863 2445 1874 2501
rect 2196 2501 2274 2502
rect 1796 2444 1874 2445
rect 1996 2485 2074 2486
rect 1596 2428 1674 2429
rect 1996 2429 2007 2485
rect 2063 2429 2074 2485
rect 2196 2445 2207 2501
rect 2263 2445 2274 2501
rect 2596 2501 2674 2502
rect 2196 2444 2274 2445
rect 2396 2485 2474 2486
rect 1996 2428 2074 2429
rect 2396 2429 2407 2485
rect 2463 2429 2474 2485
rect 2596 2445 2607 2501
rect 2663 2445 2674 2501
rect 2996 2501 3074 2502
rect 2596 2444 2674 2445
rect 2796 2485 2874 2486
rect 2396 2428 2474 2429
rect 2796 2429 2807 2485
rect 2863 2429 2874 2485
rect 2996 2445 3007 2501
rect 3063 2445 3074 2501
rect 3396 2501 3474 2502
rect 2996 2444 3074 2445
rect 3196 2485 3274 2486
rect 2796 2428 2874 2429
rect 3196 2429 3207 2485
rect 3263 2429 3274 2485
rect 3396 2445 3407 2501
rect 3463 2445 3474 2501
rect 3796 2501 3874 2502
rect 3396 2444 3474 2445
rect 3596 2485 3674 2486
rect 3196 2428 3274 2429
rect 3596 2429 3607 2485
rect 3663 2429 3674 2485
rect 3796 2445 3807 2501
rect 3863 2445 3874 2501
rect 4196 2501 4274 2502
rect 3796 2444 3874 2445
rect 3996 2485 4074 2486
rect 3596 2428 3674 2429
rect 3996 2429 4007 2485
rect 4063 2429 4074 2485
rect 4196 2445 4207 2501
rect 4263 2445 4274 2501
rect 4596 2501 4674 2502
rect 4196 2444 4274 2445
rect 4396 2485 4474 2486
rect 3996 2428 4074 2429
rect 4396 2429 4407 2485
rect 4463 2429 4474 2485
rect 4596 2445 4607 2501
rect 4663 2445 4674 2501
rect 4996 2501 5074 2502
rect 4596 2444 4674 2445
rect 4796 2485 4874 2486
rect 4396 2428 4474 2429
rect 4796 2429 4807 2485
rect 4863 2429 4874 2485
rect 4996 2445 5007 2501
rect 5063 2445 5074 2501
rect 5396 2501 5474 2502
rect 4996 2444 5074 2445
rect 5196 2485 5274 2486
rect 4796 2428 4874 2429
rect 5196 2429 5207 2485
rect 5263 2429 5274 2485
rect 5396 2445 5407 2501
rect 5463 2445 5474 2501
rect 5796 2501 5874 2502
rect 5396 2444 5474 2445
rect 5596 2485 5674 2486
rect 5196 2428 5274 2429
rect 5596 2429 5607 2485
rect 5663 2429 5674 2485
rect 5796 2445 5807 2501
rect 5863 2445 5874 2501
rect 6196 2501 6274 2502
rect 5796 2444 5874 2445
rect 5996 2485 6074 2486
rect 5596 2428 5674 2429
rect 5996 2429 6007 2485
rect 6063 2429 6074 2485
rect 6196 2445 6207 2501
rect 6263 2445 6274 2501
rect 6196 2444 6274 2445
rect 5996 2428 6074 2429
rect 202 2411 268 2412
rect 202 2400 209 2411
rect 0 2370 209 2400
rect 202 2359 209 2370
rect 261 2400 268 2411
rect 602 2411 668 2412
rect 602 2400 609 2411
rect 261 2370 609 2400
rect 261 2359 268 2370
rect 202 2358 268 2359
rect 602 2359 609 2370
rect 661 2400 668 2411
rect 1002 2411 1068 2412
rect 1002 2400 1009 2411
rect 661 2370 1009 2400
rect 661 2359 668 2370
rect 602 2358 668 2359
rect 1002 2359 1009 2370
rect 1061 2400 1068 2411
rect 1402 2411 1468 2412
rect 1402 2400 1409 2411
rect 1061 2370 1409 2400
rect 1061 2359 1068 2370
rect 1002 2358 1068 2359
rect 1402 2359 1409 2370
rect 1461 2400 1468 2411
rect 1802 2411 1868 2412
rect 1802 2400 1809 2411
rect 1461 2370 1809 2400
rect 1461 2359 1468 2370
rect 1402 2358 1468 2359
rect 1802 2359 1809 2370
rect 1861 2400 1868 2411
rect 2202 2411 2268 2412
rect 2202 2400 2209 2411
rect 1861 2370 2209 2400
rect 1861 2359 1868 2370
rect 1802 2358 1868 2359
rect 2202 2359 2209 2370
rect 2261 2400 2268 2411
rect 2602 2411 2668 2412
rect 2602 2400 2609 2411
rect 2261 2370 2609 2400
rect 2261 2359 2268 2370
rect 2202 2358 2268 2359
rect 2602 2359 2609 2370
rect 2661 2400 2668 2411
rect 3002 2411 3068 2412
rect 3002 2400 3009 2411
rect 2661 2370 3009 2400
rect 2661 2359 2668 2370
rect 2602 2358 2668 2359
rect 3002 2359 3009 2370
rect 3061 2400 3068 2411
rect 3402 2411 3468 2412
rect 3402 2400 3409 2411
rect 3061 2370 3409 2400
rect 3061 2359 3068 2370
rect 3002 2358 3068 2359
rect 3402 2359 3409 2370
rect 3461 2400 3468 2411
rect 3802 2411 3868 2412
rect 3802 2400 3809 2411
rect 3461 2370 3809 2400
rect 3461 2359 3468 2370
rect 3402 2358 3468 2359
rect 3802 2359 3809 2370
rect 3861 2400 3868 2411
rect 4202 2411 4268 2412
rect 4202 2400 4209 2411
rect 3861 2370 4209 2400
rect 3861 2359 3868 2370
rect 3802 2358 3868 2359
rect 4202 2359 4209 2370
rect 4261 2400 4268 2411
rect 4602 2411 4668 2412
rect 4602 2400 4609 2411
rect 4261 2370 4609 2400
rect 4261 2359 4268 2370
rect 4202 2358 4268 2359
rect 4602 2359 4609 2370
rect 4661 2400 4668 2411
rect 5002 2411 5068 2412
rect 5002 2400 5009 2411
rect 4661 2370 5009 2400
rect 4661 2359 4668 2370
rect 4602 2358 4668 2359
rect 5002 2359 5009 2370
rect 5061 2400 5068 2411
rect 5402 2411 5468 2412
rect 5402 2400 5409 2411
rect 5061 2370 5409 2400
rect 5061 2359 5068 2370
rect 5002 2358 5068 2359
rect 5402 2359 5409 2370
rect 5461 2400 5468 2411
rect 5802 2411 5868 2412
rect 5802 2400 5809 2411
rect 5461 2370 5809 2400
rect 5461 2359 5468 2370
rect 5402 2358 5468 2359
rect 5802 2359 5809 2370
rect 5861 2400 5868 2411
rect 6202 2411 6268 2412
rect 6202 2400 6209 2411
rect 5861 2370 6209 2400
rect 5861 2359 5868 2370
rect 5802 2358 5868 2359
rect 6202 2359 6209 2370
rect 6261 2400 6268 2411
rect 6704 2411 6770 2412
rect 6704 2400 6711 2411
rect 6261 2370 6711 2400
rect 6261 2359 6268 2370
rect 6202 2358 6268 2359
rect 6704 2359 6711 2370
rect 6763 2359 6770 2411
rect 6704 2358 6770 2359
rect 2 2341 68 2342
rect 2 2330 9 2341
rect 0 2300 9 2330
rect 2 2289 9 2300
rect 61 2330 68 2341
rect 402 2341 468 2342
rect 402 2330 409 2341
rect 61 2300 409 2330
rect 61 2289 68 2300
rect 2 2288 68 2289
rect 402 2289 409 2300
rect 461 2330 468 2341
rect 802 2341 868 2342
rect 802 2330 809 2341
rect 461 2300 809 2330
rect 461 2289 468 2300
rect 402 2288 468 2289
rect 802 2289 809 2300
rect 861 2330 868 2341
rect 1202 2341 1268 2342
rect 1202 2330 1209 2341
rect 861 2300 1209 2330
rect 861 2289 868 2300
rect 802 2288 868 2289
rect 1202 2289 1209 2300
rect 1261 2330 1268 2341
rect 1602 2341 1668 2342
rect 1602 2330 1609 2341
rect 1261 2300 1609 2330
rect 1261 2289 1268 2300
rect 1202 2288 1268 2289
rect 1602 2289 1609 2300
rect 1661 2330 1668 2341
rect 2002 2341 2068 2342
rect 2002 2330 2009 2341
rect 1661 2300 2009 2330
rect 1661 2289 1668 2300
rect 1602 2288 1668 2289
rect 2002 2289 2009 2300
rect 2061 2330 2068 2341
rect 2402 2341 2468 2342
rect 2402 2330 2409 2341
rect 2061 2300 2409 2330
rect 2061 2289 2068 2300
rect 2002 2288 2068 2289
rect 2402 2289 2409 2300
rect 2461 2330 2468 2341
rect 2802 2341 2868 2342
rect 2802 2330 2809 2341
rect 2461 2300 2809 2330
rect 2461 2289 2468 2300
rect 2402 2288 2468 2289
rect 2802 2289 2809 2300
rect 2861 2330 2868 2341
rect 3202 2341 3268 2342
rect 3202 2330 3209 2341
rect 2861 2300 3209 2330
rect 2861 2289 2868 2300
rect 2802 2288 2868 2289
rect 3202 2289 3209 2300
rect 3261 2330 3268 2341
rect 3602 2341 3668 2342
rect 3602 2330 3609 2341
rect 3261 2300 3609 2330
rect 3261 2289 3268 2300
rect 3202 2288 3268 2289
rect 3602 2289 3609 2300
rect 3661 2330 3668 2341
rect 4002 2341 4068 2342
rect 4002 2330 4009 2341
rect 3661 2300 4009 2330
rect 3661 2289 3668 2300
rect 3602 2288 3668 2289
rect 4002 2289 4009 2300
rect 4061 2330 4068 2341
rect 4402 2341 4468 2342
rect 4402 2330 4409 2341
rect 4061 2300 4409 2330
rect 4061 2289 4068 2300
rect 4002 2288 4068 2289
rect 4402 2289 4409 2300
rect 4461 2330 4468 2341
rect 4802 2341 4868 2342
rect 4802 2330 4809 2341
rect 4461 2300 4809 2330
rect 4461 2289 4468 2300
rect 4402 2288 4468 2289
rect 4802 2289 4809 2300
rect 4861 2330 4868 2341
rect 5202 2341 5268 2342
rect 5202 2330 5209 2341
rect 4861 2300 5209 2330
rect 4861 2289 4868 2300
rect 4802 2288 4868 2289
rect 5202 2289 5209 2300
rect 5261 2330 5268 2341
rect 5602 2341 5668 2342
rect 5602 2330 5609 2341
rect 5261 2300 5609 2330
rect 5261 2289 5268 2300
rect 5202 2288 5268 2289
rect 5602 2289 5609 2300
rect 5661 2330 5668 2341
rect 6002 2341 6068 2342
rect 6002 2330 6009 2341
rect 5661 2300 6009 2330
rect 5661 2289 5668 2300
rect 5602 2288 5668 2289
rect 6002 2289 6009 2300
rect 6061 2330 6068 2341
rect 6402 2341 6468 2342
rect 6402 2330 6409 2341
rect 6061 2300 6409 2330
rect 6061 2289 6068 2300
rect 6002 2288 6068 2289
rect 6402 2289 6409 2300
rect 6461 2330 6468 2341
rect 6500 2341 6566 2342
rect 6500 2330 6507 2341
rect 6461 2300 6507 2330
rect 6461 2289 6468 2300
rect 6402 2288 6468 2289
rect 6500 2289 6507 2300
rect 6559 2289 6566 2341
rect 6500 2288 6566 2289
rect 202 2271 268 2272
rect 202 2260 209 2271
rect 0 2230 209 2260
rect 202 2219 209 2230
rect 261 2260 268 2271
rect 602 2271 668 2272
rect 602 2260 609 2271
rect 261 2230 609 2260
rect 261 2219 268 2230
rect 202 2218 268 2219
rect 602 2219 609 2230
rect 661 2260 668 2271
rect 1002 2271 1068 2272
rect 1002 2260 1009 2271
rect 661 2230 1009 2260
rect 661 2219 668 2230
rect 602 2218 668 2219
rect 1002 2219 1009 2230
rect 1061 2260 1068 2271
rect 1402 2271 1468 2272
rect 1402 2260 1409 2271
rect 1061 2230 1409 2260
rect 1061 2219 1068 2230
rect 1002 2218 1068 2219
rect 1402 2219 1409 2230
rect 1461 2260 1468 2271
rect 1802 2271 1868 2272
rect 1802 2260 1809 2271
rect 1461 2230 1809 2260
rect 1461 2219 1468 2230
rect 1402 2218 1468 2219
rect 1802 2219 1809 2230
rect 1861 2260 1868 2271
rect 2202 2271 2268 2272
rect 2202 2260 2209 2271
rect 1861 2230 2209 2260
rect 1861 2219 1868 2230
rect 1802 2218 1868 2219
rect 2202 2219 2209 2230
rect 2261 2260 2268 2271
rect 2602 2271 2668 2272
rect 2602 2260 2609 2271
rect 2261 2230 2609 2260
rect 2261 2219 2268 2230
rect 2202 2218 2268 2219
rect 2602 2219 2609 2230
rect 2661 2260 2668 2271
rect 3002 2271 3068 2272
rect 3002 2260 3009 2271
rect 2661 2230 3009 2260
rect 2661 2219 2668 2230
rect 2602 2218 2668 2219
rect 3002 2219 3009 2230
rect 3061 2260 3068 2271
rect 3402 2271 3468 2272
rect 3402 2260 3409 2271
rect 3061 2230 3409 2260
rect 3061 2219 3068 2230
rect 3002 2218 3068 2219
rect 3402 2219 3409 2230
rect 3461 2260 3468 2271
rect 3802 2271 3868 2272
rect 3802 2260 3809 2271
rect 3461 2230 3809 2260
rect 3461 2219 3468 2230
rect 3402 2218 3468 2219
rect 3802 2219 3809 2230
rect 3861 2260 3868 2271
rect 4202 2271 4268 2272
rect 4202 2260 4209 2271
rect 3861 2230 4209 2260
rect 3861 2219 3868 2230
rect 3802 2218 3868 2219
rect 4202 2219 4209 2230
rect 4261 2260 4268 2271
rect 4602 2271 4668 2272
rect 4602 2260 4609 2271
rect 4261 2230 4609 2260
rect 4261 2219 4268 2230
rect 4202 2218 4268 2219
rect 4602 2219 4609 2230
rect 4661 2260 4668 2271
rect 5002 2271 5068 2272
rect 5002 2260 5009 2271
rect 4661 2230 5009 2260
rect 4661 2219 4668 2230
rect 4602 2218 4668 2219
rect 5002 2219 5009 2230
rect 5061 2260 5068 2271
rect 5402 2271 5468 2272
rect 5402 2260 5409 2271
rect 5061 2230 5409 2260
rect 5061 2219 5068 2230
rect 5002 2218 5068 2219
rect 5402 2219 5409 2230
rect 5461 2260 5468 2271
rect 5802 2271 5868 2272
rect 5802 2260 5809 2271
rect 5461 2230 5809 2260
rect 5461 2219 5468 2230
rect 5402 2218 5468 2219
rect 5802 2219 5809 2230
rect 5861 2260 5868 2271
rect 6202 2271 6268 2272
rect 6202 2260 6209 2271
rect 5861 2230 6209 2260
rect 5861 2219 5868 2230
rect 5802 2218 5868 2219
rect 6202 2219 6209 2230
rect 6261 2260 6268 2271
rect 6704 2271 6770 2272
rect 6704 2260 6711 2271
rect 6261 2230 6711 2260
rect 6261 2219 6268 2230
rect 6202 2218 6268 2219
rect 6704 2219 6711 2230
rect 6763 2219 6770 2271
rect 6704 2218 6770 2219
rect 2 2201 68 2202
rect 2 2190 9 2201
rect 0 2160 9 2190
rect 2 2149 9 2160
rect 61 2190 68 2201
rect 402 2201 468 2202
rect 402 2190 409 2201
rect 61 2160 409 2190
rect 61 2149 68 2160
rect 2 2148 68 2149
rect 402 2149 409 2160
rect 461 2190 468 2201
rect 802 2201 868 2202
rect 802 2190 809 2201
rect 461 2160 809 2190
rect 461 2149 468 2160
rect 402 2148 468 2149
rect 802 2149 809 2160
rect 861 2190 868 2201
rect 1202 2201 1268 2202
rect 1202 2190 1209 2201
rect 861 2160 1209 2190
rect 861 2149 868 2160
rect 802 2148 868 2149
rect 1202 2149 1209 2160
rect 1261 2190 1268 2201
rect 1602 2201 1668 2202
rect 1602 2190 1609 2201
rect 1261 2160 1609 2190
rect 1261 2149 1268 2160
rect 1202 2148 1268 2149
rect 1602 2149 1609 2160
rect 1661 2190 1668 2201
rect 2002 2201 2068 2202
rect 2002 2190 2009 2201
rect 1661 2160 2009 2190
rect 1661 2149 1668 2160
rect 1602 2148 1668 2149
rect 2002 2149 2009 2160
rect 2061 2190 2068 2201
rect 2402 2201 2468 2202
rect 2402 2190 2409 2201
rect 2061 2160 2409 2190
rect 2061 2149 2068 2160
rect 2002 2148 2068 2149
rect 2402 2149 2409 2160
rect 2461 2190 2468 2201
rect 2802 2201 2868 2202
rect 2802 2190 2809 2201
rect 2461 2160 2809 2190
rect 2461 2149 2468 2160
rect 2402 2148 2468 2149
rect 2802 2149 2809 2160
rect 2861 2190 2868 2201
rect 3202 2201 3268 2202
rect 3202 2190 3209 2201
rect 2861 2160 3209 2190
rect 2861 2149 2868 2160
rect 2802 2148 2868 2149
rect 3202 2149 3209 2160
rect 3261 2190 3268 2201
rect 3602 2201 3668 2202
rect 3602 2190 3609 2201
rect 3261 2160 3609 2190
rect 3261 2149 3268 2160
rect 3202 2148 3268 2149
rect 3602 2149 3609 2160
rect 3661 2190 3668 2201
rect 4002 2201 4068 2202
rect 4002 2190 4009 2201
rect 3661 2160 4009 2190
rect 3661 2149 3668 2160
rect 3602 2148 3668 2149
rect 4002 2149 4009 2160
rect 4061 2190 4068 2201
rect 4402 2201 4468 2202
rect 4402 2190 4409 2201
rect 4061 2160 4409 2190
rect 4061 2149 4068 2160
rect 4002 2148 4068 2149
rect 4402 2149 4409 2160
rect 4461 2190 4468 2201
rect 4802 2201 4868 2202
rect 4802 2190 4809 2201
rect 4461 2160 4809 2190
rect 4461 2149 4468 2160
rect 4402 2148 4468 2149
rect 4802 2149 4809 2160
rect 4861 2190 4868 2201
rect 5202 2201 5268 2202
rect 5202 2190 5209 2201
rect 4861 2160 5209 2190
rect 4861 2149 4868 2160
rect 4802 2148 4868 2149
rect 5202 2149 5209 2160
rect 5261 2190 5268 2201
rect 5602 2201 5668 2202
rect 5602 2190 5609 2201
rect 5261 2160 5609 2190
rect 5261 2149 5268 2160
rect 5202 2148 5268 2149
rect 5602 2149 5609 2160
rect 5661 2190 5668 2201
rect 6002 2201 6068 2202
rect 6002 2190 6009 2201
rect 5661 2160 6009 2190
rect 5661 2149 5668 2160
rect 5602 2148 5668 2149
rect 6002 2149 6009 2160
rect 6061 2190 6068 2201
rect 6402 2201 6468 2202
rect 6402 2190 6409 2201
rect 6061 2160 6409 2190
rect 6061 2149 6068 2160
rect 6002 2148 6068 2149
rect 6402 2149 6409 2160
rect 6461 2190 6468 2201
rect 6500 2201 6566 2202
rect 6500 2190 6507 2201
rect 6461 2160 6507 2190
rect 6461 2149 6468 2160
rect 6402 2148 6468 2149
rect 6500 2149 6507 2160
rect 6559 2149 6566 2201
rect 6500 2148 6566 2149
rect 202 2131 268 2132
rect 202 2120 209 2131
rect 0 2090 209 2120
rect 202 2079 209 2090
rect 261 2120 268 2131
rect 602 2131 668 2132
rect 602 2120 609 2131
rect 261 2090 609 2120
rect 261 2079 268 2090
rect 202 2078 268 2079
rect 602 2079 609 2090
rect 661 2120 668 2131
rect 1002 2131 1068 2132
rect 1002 2120 1009 2131
rect 661 2090 1009 2120
rect 661 2079 668 2090
rect 602 2078 668 2079
rect 1002 2079 1009 2090
rect 1061 2120 1068 2131
rect 1402 2131 1468 2132
rect 1402 2120 1409 2131
rect 1061 2090 1409 2120
rect 1061 2079 1068 2090
rect 1002 2078 1068 2079
rect 1402 2079 1409 2090
rect 1461 2120 1468 2131
rect 1802 2131 1868 2132
rect 1802 2120 1809 2131
rect 1461 2090 1809 2120
rect 1461 2079 1468 2090
rect 1402 2078 1468 2079
rect 1802 2079 1809 2090
rect 1861 2120 1868 2131
rect 2202 2131 2268 2132
rect 2202 2120 2209 2131
rect 1861 2090 2209 2120
rect 1861 2079 1868 2090
rect 1802 2078 1868 2079
rect 2202 2079 2209 2090
rect 2261 2120 2268 2131
rect 2602 2131 2668 2132
rect 2602 2120 2609 2131
rect 2261 2090 2609 2120
rect 2261 2079 2268 2090
rect 2202 2078 2268 2079
rect 2602 2079 2609 2090
rect 2661 2120 2668 2131
rect 3002 2131 3068 2132
rect 3002 2120 3009 2131
rect 2661 2090 3009 2120
rect 2661 2079 2668 2090
rect 2602 2078 2668 2079
rect 3002 2079 3009 2090
rect 3061 2120 3068 2131
rect 3402 2131 3468 2132
rect 3402 2120 3409 2131
rect 3061 2090 3409 2120
rect 3061 2079 3068 2090
rect 3002 2078 3068 2079
rect 3402 2079 3409 2090
rect 3461 2120 3468 2131
rect 3802 2131 3868 2132
rect 3802 2120 3809 2131
rect 3461 2090 3809 2120
rect 3461 2079 3468 2090
rect 3402 2078 3468 2079
rect 3802 2079 3809 2090
rect 3861 2120 3868 2131
rect 4202 2131 4268 2132
rect 4202 2120 4209 2131
rect 3861 2090 4209 2120
rect 3861 2079 3868 2090
rect 3802 2078 3868 2079
rect 4202 2079 4209 2090
rect 4261 2120 4268 2131
rect 4602 2131 4668 2132
rect 4602 2120 4609 2131
rect 4261 2090 4609 2120
rect 4261 2079 4268 2090
rect 4202 2078 4268 2079
rect 4602 2079 4609 2090
rect 4661 2120 4668 2131
rect 5002 2131 5068 2132
rect 5002 2120 5009 2131
rect 4661 2090 5009 2120
rect 4661 2079 4668 2090
rect 4602 2078 4668 2079
rect 5002 2079 5009 2090
rect 5061 2120 5068 2131
rect 5402 2131 5468 2132
rect 5402 2120 5409 2131
rect 5061 2090 5409 2120
rect 5061 2079 5068 2090
rect 5002 2078 5068 2079
rect 5402 2079 5409 2090
rect 5461 2120 5468 2131
rect 5802 2131 5868 2132
rect 5802 2120 5809 2131
rect 5461 2090 5809 2120
rect 5461 2079 5468 2090
rect 5402 2078 5468 2079
rect 5802 2079 5809 2090
rect 5861 2120 5868 2131
rect 6202 2131 6268 2132
rect 6202 2120 6209 2131
rect 5861 2090 6209 2120
rect 5861 2079 5868 2090
rect 5802 2078 5868 2079
rect 6202 2079 6209 2090
rect 6261 2120 6268 2131
rect 6704 2131 6770 2132
rect 6704 2120 6711 2131
rect 6261 2090 6711 2120
rect 6261 2079 6268 2090
rect 6202 2078 6268 2079
rect 6704 2079 6711 2090
rect 6763 2079 6770 2131
rect 6704 2078 6770 2079
rect 2 2061 68 2062
rect 2 2050 9 2061
rect 0 2020 9 2050
rect 2 2009 9 2020
rect 61 2050 68 2061
rect 402 2061 468 2062
rect 402 2050 409 2061
rect 61 2020 409 2050
rect 61 2009 68 2020
rect 2 2008 68 2009
rect 402 2009 409 2020
rect 461 2050 468 2061
rect 802 2061 868 2062
rect 802 2050 809 2061
rect 461 2020 809 2050
rect 461 2009 468 2020
rect 402 2008 468 2009
rect 802 2009 809 2020
rect 861 2050 868 2061
rect 1202 2061 1268 2062
rect 1202 2050 1209 2061
rect 861 2020 1209 2050
rect 861 2009 868 2020
rect 802 2008 868 2009
rect 1202 2009 1209 2020
rect 1261 2050 1268 2061
rect 1602 2061 1668 2062
rect 1602 2050 1609 2061
rect 1261 2020 1609 2050
rect 1261 2009 1268 2020
rect 1202 2008 1268 2009
rect 1602 2009 1609 2020
rect 1661 2050 1668 2061
rect 2002 2061 2068 2062
rect 2002 2050 2009 2061
rect 1661 2020 2009 2050
rect 1661 2009 1668 2020
rect 1602 2008 1668 2009
rect 2002 2009 2009 2020
rect 2061 2050 2068 2061
rect 2402 2061 2468 2062
rect 2402 2050 2409 2061
rect 2061 2020 2409 2050
rect 2061 2009 2068 2020
rect 2002 2008 2068 2009
rect 2402 2009 2409 2020
rect 2461 2050 2468 2061
rect 2802 2061 2868 2062
rect 2802 2050 2809 2061
rect 2461 2020 2809 2050
rect 2461 2009 2468 2020
rect 2402 2008 2468 2009
rect 2802 2009 2809 2020
rect 2861 2050 2868 2061
rect 3202 2061 3268 2062
rect 3202 2050 3209 2061
rect 2861 2020 3209 2050
rect 2861 2009 2868 2020
rect 2802 2008 2868 2009
rect 3202 2009 3209 2020
rect 3261 2050 3268 2061
rect 3602 2061 3668 2062
rect 3602 2050 3609 2061
rect 3261 2020 3609 2050
rect 3261 2009 3268 2020
rect 3202 2008 3268 2009
rect 3602 2009 3609 2020
rect 3661 2050 3668 2061
rect 4002 2061 4068 2062
rect 4002 2050 4009 2061
rect 3661 2020 4009 2050
rect 3661 2009 3668 2020
rect 3602 2008 3668 2009
rect 4002 2009 4009 2020
rect 4061 2050 4068 2061
rect 4402 2061 4468 2062
rect 4402 2050 4409 2061
rect 4061 2020 4409 2050
rect 4061 2009 4068 2020
rect 4002 2008 4068 2009
rect 4402 2009 4409 2020
rect 4461 2050 4468 2061
rect 4802 2061 4868 2062
rect 4802 2050 4809 2061
rect 4461 2020 4809 2050
rect 4461 2009 4468 2020
rect 4402 2008 4468 2009
rect 4802 2009 4809 2020
rect 4861 2050 4868 2061
rect 5202 2061 5268 2062
rect 5202 2050 5209 2061
rect 4861 2020 5209 2050
rect 4861 2009 4868 2020
rect 4802 2008 4868 2009
rect 5202 2009 5209 2020
rect 5261 2050 5268 2061
rect 5602 2061 5668 2062
rect 5602 2050 5609 2061
rect 5261 2020 5609 2050
rect 5261 2009 5268 2020
rect 5202 2008 5268 2009
rect 5602 2009 5609 2020
rect 5661 2050 5668 2061
rect 6002 2061 6068 2062
rect 6002 2050 6009 2061
rect 5661 2020 6009 2050
rect 5661 2009 5668 2020
rect 5602 2008 5668 2009
rect 6002 2009 6009 2020
rect 6061 2050 6068 2061
rect 6402 2061 6468 2062
rect 6402 2050 6409 2061
rect 6061 2020 6409 2050
rect 6061 2009 6068 2020
rect 6002 2008 6068 2009
rect 6402 2009 6409 2020
rect 6461 2050 6468 2061
rect 6500 2061 6566 2062
rect 6500 2050 6507 2061
rect 6461 2020 6507 2050
rect 6461 2009 6468 2020
rect 6402 2008 6468 2009
rect 6500 2009 6507 2020
rect 6559 2009 6566 2061
rect 6500 2008 6566 2009
rect 202 1991 268 1992
rect 202 1980 209 1991
rect 0 1950 209 1980
rect 202 1939 209 1950
rect 261 1980 268 1991
rect 602 1991 668 1992
rect 602 1980 609 1991
rect 261 1950 609 1980
rect 261 1939 268 1950
rect 202 1938 268 1939
rect 602 1939 609 1950
rect 661 1980 668 1991
rect 1002 1991 1068 1992
rect 1002 1980 1009 1991
rect 661 1950 1009 1980
rect 661 1939 668 1950
rect 602 1938 668 1939
rect 1002 1939 1009 1950
rect 1061 1980 1068 1991
rect 1402 1991 1468 1992
rect 1402 1980 1409 1991
rect 1061 1950 1409 1980
rect 1061 1939 1068 1950
rect 1002 1938 1068 1939
rect 1402 1939 1409 1950
rect 1461 1980 1468 1991
rect 1802 1991 1868 1992
rect 1802 1980 1809 1991
rect 1461 1950 1809 1980
rect 1461 1939 1468 1950
rect 1402 1938 1468 1939
rect 1802 1939 1809 1950
rect 1861 1980 1868 1991
rect 2202 1991 2268 1992
rect 2202 1980 2209 1991
rect 1861 1950 2209 1980
rect 1861 1939 1868 1950
rect 1802 1938 1868 1939
rect 2202 1939 2209 1950
rect 2261 1980 2268 1991
rect 2602 1991 2668 1992
rect 2602 1980 2609 1991
rect 2261 1950 2609 1980
rect 2261 1939 2268 1950
rect 2202 1938 2268 1939
rect 2602 1939 2609 1950
rect 2661 1980 2668 1991
rect 3002 1991 3068 1992
rect 3002 1980 3009 1991
rect 2661 1950 3009 1980
rect 2661 1939 2668 1950
rect 2602 1938 2668 1939
rect 3002 1939 3009 1950
rect 3061 1980 3068 1991
rect 3402 1991 3468 1992
rect 3402 1980 3409 1991
rect 3061 1950 3409 1980
rect 3061 1939 3068 1950
rect 3002 1938 3068 1939
rect 3402 1939 3409 1950
rect 3461 1980 3468 1991
rect 3802 1991 3868 1992
rect 3802 1980 3809 1991
rect 3461 1950 3809 1980
rect 3461 1939 3468 1950
rect 3402 1938 3468 1939
rect 3802 1939 3809 1950
rect 3861 1980 3868 1991
rect 4202 1991 4268 1992
rect 4202 1980 4209 1991
rect 3861 1950 4209 1980
rect 3861 1939 3868 1950
rect 3802 1938 3868 1939
rect 4202 1939 4209 1950
rect 4261 1980 4268 1991
rect 4602 1991 4668 1992
rect 4602 1980 4609 1991
rect 4261 1950 4609 1980
rect 4261 1939 4268 1950
rect 4202 1938 4268 1939
rect 4602 1939 4609 1950
rect 4661 1980 4668 1991
rect 5002 1991 5068 1992
rect 5002 1980 5009 1991
rect 4661 1950 5009 1980
rect 4661 1939 4668 1950
rect 4602 1938 4668 1939
rect 5002 1939 5009 1950
rect 5061 1980 5068 1991
rect 5402 1991 5468 1992
rect 5402 1980 5409 1991
rect 5061 1950 5409 1980
rect 5061 1939 5068 1950
rect 5002 1938 5068 1939
rect 5402 1939 5409 1950
rect 5461 1980 5468 1991
rect 5802 1991 5868 1992
rect 5802 1980 5809 1991
rect 5461 1950 5809 1980
rect 5461 1939 5468 1950
rect 5402 1938 5468 1939
rect 5802 1939 5809 1950
rect 5861 1980 5868 1991
rect 6202 1991 6268 1992
rect 6202 1980 6209 1991
rect 5861 1950 6209 1980
rect 5861 1939 5868 1950
rect 5802 1938 5868 1939
rect 6202 1939 6209 1950
rect 6261 1980 6268 1991
rect 6704 1991 6770 1992
rect 6704 1980 6711 1991
rect 6261 1950 6711 1980
rect 6261 1939 6268 1950
rect 6202 1938 6268 1939
rect 6704 1939 6711 1950
rect 6763 1939 6770 1991
rect 6704 1938 6770 1939
rect 2 1921 68 1922
rect 2 1910 9 1921
rect 0 1880 9 1910
rect 2 1869 9 1880
rect 61 1910 68 1921
rect 402 1921 468 1922
rect 402 1910 409 1921
rect 61 1880 409 1910
rect 61 1869 68 1880
rect 2 1868 68 1869
rect 402 1869 409 1880
rect 461 1910 468 1921
rect 802 1921 868 1922
rect 802 1910 809 1921
rect 461 1880 809 1910
rect 461 1869 468 1880
rect 402 1868 468 1869
rect 802 1869 809 1880
rect 861 1910 868 1921
rect 1202 1921 1268 1922
rect 1202 1910 1209 1921
rect 861 1880 1209 1910
rect 861 1869 868 1880
rect 802 1868 868 1869
rect 1202 1869 1209 1880
rect 1261 1910 1268 1921
rect 1602 1921 1668 1922
rect 1602 1910 1609 1921
rect 1261 1880 1609 1910
rect 1261 1869 1268 1880
rect 1202 1868 1268 1869
rect 1602 1869 1609 1880
rect 1661 1910 1668 1921
rect 2002 1921 2068 1922
rect 2002 1910 2009 1921
rect 1661 1880 2009 1910
rect 1661 1869 1668 1880
rect 1602 1868 1668 1869
rect 2002 1869 2009 1880
rect 2061 1910 2068 1921
rect 2402 1921 2468 1922
rect 2402 1910 2409 1921
rect 2061 1880 2409 1910
rect 2061 1869 2068 1880
rect 2002 1868 2068 1869
rect 2402 1869 2409 1880
rect 2461 1910 2468 1921
rect 2802 1921 2868 1922
rect 2802 1910 2809 1921
rect 2461 1880 2809 1910
rect 2461 1869 2468 1880
rect 2402 1868 2468 1869
rect 2802 1869 2809 1880
rect 2861 1910 2868 1921
rect 3202 1921 3268 1922
rect 3202 1910 3209 1921
rect 2861 1880 3209 1910
rect 2861 1869 2868 1880
rect 2802 1868 2868 1869
rect 3202 1869 3209 1880
rect 3261 1910 3268 1921
rect 3602 1921 3668 1922
rect 3602 1910 3609 1921
rect 3261 1880 3609 1910
rect 3261 1869 3268 1880
rect 3202 1868 3268 1869
rect 3602 1869 3609 1880
rect 3661 1910 3668 1921
rect 4002 1921 4068 1922
rect 4002 1910 4009 1921
rect 3661 1880 4009 1910
rect 3661 1869 3668 1880
rect 3602 1868 3668 1869
rect 4002 1869 4009 1880
rect 4061 1910 4068 1921
rect 4402 1921 4468 1922
rect 4402 1910 4409 1921
rect 4061 1880 4409 1910
rect 4061 1869 4068 1880
rect 4002 1868 4068 1869
rect 4402 1869 4409 1880
rect 4461 1910 4468 1921
rect 4802 1921 4868 1922
rect 4802 1910 4809 1921
rect 4461 1880 4809 1910
rect 4461 1869 4468 1880
rect 4402 1868 4468 1869
rect 4802 1869 4809 1880
rect 4861 1910 4868 1921
rect 5202 1921 5268 1922
rect 5202 1910 5209 1921
rect 4861 1880 5209 1910
rect 4861 1869 4868 1880
rect 4802 1868 4868 1869
rect 5202 1869 5209 1880
rect 5261 1910 5268 1921
rect 5602 1921 5668 1922
rect 5602 1910 5609 1921
rect 5261 1880 5609 1910
rect 5261 1869 5268 1880
rect 5202 1868 5268 1869
rect 5602 1869 5609 1880
rect 5661 1910 5668 1921
rect 6002 1921 6068 1922
rect 6002 1910 6009 1921
rect 5661 1880 6009 1910
rect 5661 1869 5668 1880
rect 5602 1868 5668 1869
rect 6002 1869 6009 1880
rect 6061 1910 6068 1921
rect 6402 1921 6468 1922
rect 6402 1910 6409 1921
rect 6061 1880 6409 1910
rect 6061 1869 6068 1880
rect 6002 1868 6068 1869
rect 6402 1869 6409 1880
rect 6461 1910 6468 1921
rect 6500 1921 6566 1922
rect 6500 1910 6507 1921
rect 6461 1880 6507 1910
rect 6461 1869 6468 1880
rect 6402 1868 6468 1869
rect 6500 1869 6507 1880
rect 6559 1869 6566 1921
rect 6500 1868 6566 1869
rect 202 1851 268 1852
rect 202 1840 209 1851
rect 0 1810 209 1840
rect 202 1799 209 1810
rect 261 1840 268 1851
rect 602 1851 668 1852
rect 602 1840 609 1851
rect 261 1810 609 1840
rect 261 1799 268 1810
rect 202 1798 268 1799
rect 602 1799 609 1810
rect 661 1840 668 1851
rect 1002 1851 1068 1852
rect 1002 1840 1009 1851
rect 661 1810 1009 1840
rect 661 1799 668 1810
rect 602 1798 668 1799
rect 1002 1799 1009 1810
rect 1061 1840 1068 1851
rect 1402 1851 1468 1852
rect 1402 1840 1409 1851
rect 1061 1810 1409 1840
rect 1061 1799 1068 1810
rect 1002 1798 1068 1799
rect 1402 1799 1409 1810
rect 1461 1840 1468 1851
rect 1802 1851 1868 1852
rect 1802 1840 1809 1851
rect 1461 1810 1809 1840
rect 1461 1799 1468 1810
rect 1402 1798 1468 1799
rect 1802 1799 1809 1810
rect 1861 1840 1868 1851
rect 2202 1851 2268 1852
rect 2202 1840 2209 1851
rect 1861 1810 2209 1840
rect 1861 1799 1868 1810
rect 1802 1798 1868 1799
rect 2202 1799 2209 1810
rect 2261 1840 2268 1851
rect 2602 1851 2668 1852
rect 2602 1840 2609 1851
rect 2261 1810 2609 1840
rect 2261 1799 2268 1810
rect 2202 1798 2268 1799
rect 2602 1799 2609 1810
rect 2661 1840 2668 1851
rect 3002 1851 3068 1852
rect 3002 1840 3009 1851
rect 2661 1810 3009 1840
rect 2661 1799 2668 1810
rect 2602 1798 2668 1799
rect 3002 1799 3009 1810
rect 3061 1840 3068 1851
rect 3402 1851 3468 1852
rect 3402 1840 3409 1851
rect 3061 1810 3409 1840
rect 3061 1799 3068 1810
rect 3002 1798 3068 1799
rect 3402 1799 3409 1810
rect 3461 1840 3468 1851
rect 3802 1851 3868 1852
rect 3802 1840 3809 1851
rect 3461 1810 3809 1840
rect 3461 1799 3468 1810
rect 3402 1798 3468 1799
rect 3802 1799 3809 1810
rect 3861 1840 3868 1851
rect 4202 1851 4268 1852
rect 4202 1840 4209 1851
rect 3861 1810 4209 1840
rect 3861 1799 3868 1810
rect 3802 1798 3868 1799
rect 4202 1799 4209 1810
rect 4261 1840 4268 1851
rect 4602 1851 4668 1852
rect 4602 1840 4609 1851
rect 4261 1810 4609 1840
rect 4261 1799 4268 1810
rect 4202 1798 4268 1799
rect 4602 1799 4609 1810
rect 4661 1840 4668 1851
rect 5002 1851 5068 1852
rect 5002 1840 5009 1851
rect 4661 1810 5009 1840
rect 4661 1799 4668 1810
rect 4602 1798 4668 1799
rect 5002 1799 5009 1810
rect 5061 1840 5068 1851
rect 5402 1851 5468 1852
rect 5402 1840 5409 1851
rect 5061 1810 5409 1840
rect 5061 1799 5068 1810
rect 5002 1798 5068 1799
rect 5402 1799 5409 1810
rect 5461 1840 5468 1851
rect 5802 1851 5868 1852
rect 5802 1840 5809 1851
rect 5461 1810 5809 1840
rect 5461 1799 5468 1810
rect 5402 1798 5468 1799
rect 5802 1799 5809 1810
rect 5861 1840 5868 1851
rect 6202 1851 6268 1852
rect 6202 1840 6209 1851
rect 5861 1810 6209 1840
rect 5861 1799 5868 1810
rect 5802 1798 5868 1799
rect 6202 1799 6209 1810
rect 6261 1840 6268 1851
rect 6704 1851 6770 1852
rect 6704 1840 6711 1851
rect 6261 1810 6711 1840
rect 6261 1799 6268 1810
rect 6202 1798 6268 1799
rect 6704 1799 6711 1810
rect 6763 1799 6770 1851
rect 6704 1798 6770 1799
rect 2 1781 68 1782
rect 2 1770 9 1781
rect 0 1740 9 1770
rect 2 1729 9 1740
rect 61 1770 68 1781
rect 402 1781 468 1782
rect 402 1770 409 1781
rect 61 1740 409 1770
rect 61 1729 68 1740
rect 2 1728 68 1729
rect 402 1729 409 1740
rect 461 1770 468 1781
rect 802 1781 868 1782
rect 802 1770 809 1781
rect 461 1740 809 1770
rect 461 1729 468 1740
rect 402 1728 468 1729
rect 802 1729 809 1740
rect 861 1770 868 1781
rect 1202 1781 1268 1782
rect 1202 1770 1209 1781
rect 861 1740 1209 1770
rect 861 1729 868 1740
rect 802 1728 868 1729
rect 1202 1729 1209 1740
rect 1261 1770 1268 1781
rect 1602 1781 1668 1782
rect 1602 1770 1609 1781
rect 1261 1740 1609 1770
rect 1261 1729 1268 1740
rect 1202 1728 1268 1729
rect 1602 1729 1609 1740
rect 1661 1770 1668 1781
rect 2002 1781 2068 1782
rect 2002 1770 2009 1781
rect 1661 1740 2009 1770
rect 1661 1729 1668 1740
rect 1602 1728 1668 1729
rect 2002 1729 2009 1740
rect 2061 1770 2068 1781
rect 2402 1781 2468 1782
rect 2402 1770 2409 1781
rect 2061 1740 2409 1770
rect 2061 1729 2068 1740
rect 2002 1728 2068 1729
rect 2402 1729 2409 1740
rect 2461 1770 2468 1781
rect 2802 1781 2868 1782
rect 2802 1770 2809 1781
rect 2461 1740 2809 1770
rect 2461 1729 2468 1740
rect 2402 1728 2468 1729
rect 2802 1729 2809 1740
rect 2861 1770 2868 1781
rect 3202 1781 3268 1782
rect 3202 1770 3209 1781
rect 2861 1740 3209 1770
rect 2861 1729 2868 1740
rect 2802 1728 2868 1729
rect 3202 1729 3209 1740
rect 3261 1770 3268 1781
rect 3602 1781 3668 1782
rect 3602 1770 3609 1781
rect 3261 1740 3609 1770
rect 3261 1729 3268 1740
rect 3202 1728 3268 1729
rect 3602 1729 3609 1740
rect 3661 1770 3668 1781
rect 4002 1781 4068 1782
rect 4002 1770 4009 1781
rect 3661 1740 4009 1770
rect 3661 1729 3668 1740
rect 3602 1728 3668 1729
rect 4002 1729 4009 1740
rect 4061 1770 4068 1781
rect 4402 1781 4468 1782
rect 4402 1770 4409 1781
rect 4061 1740 4409 1770
rect 4061 1729 4068 1740
rect 4002 1728 4068 1729
rect 4402 1729 4409 1740
rect 4461 1770 4468 1781
rect 4802 1781 4868 1782
rect 4802 1770 4809 1781
rect 4461 1740 4809 1770
rect 4461 1729 4468 1740
rect 4402 1728 4468 1729
rect 4802 1729 4809 1740
rect 4861 1770 4868 1781
rect 5202 1781 5268 1782
rect 5202 1770 5209 1781
rect 4861 1740 5209 1770
rect 4861 1729 4868 1740
rect 4802 1728 4868 1729
rect 5202 1729 5209 1740
rect 5261 1770 5268 1781
rect 5602 1781 5668 1782
rect 5602 1770 5609 1781
rect 5261 1740 5609 1770
rect 5261 1729 5268 1740
rect 5202 1728 5268 1729
rect 5602 1729 5609 1740
rect 5661 1770 5668 1781
rect 6002 1781 6068 1782
rect 6002 1770 6009 1781
rect 5661 1740 6009 1770
rect 5661 1729 5668 1740
rect 5602 1728 5668 1729
rect 6002 1729 6009 1740
rect 6061 1770 6068 1781
rect 6402 1781 6468 1782
rect 6402 1770 6409 1781
rect 6061 1740 6409 1770
rect 6061 1729 6068 1740
rect 6002 1728 6068 1729
rect 6402 1729 6409 1740
rect 6461 1770 6468 1781
rect 6500 1781 6566 1782
rect 6500 1770 6507 1781
rect 6461 1740 6507 1770
rect 6461 1729 6468 1740
rect 6402 1728 6468 1729
rect 6500 1729 6507 1740
rect 6559 1729 6566 1781
rect 6500 1728 6566 1729
rect 202 1711 268 1712
rect 202 1700 209 1711
rect 0 1670 209 1700
rect 202 1659 209 1670
rect 261 1700 268 1711
rect 602 1711 668 1712
rect 602 1700 609 1711
rect 261 1670 609 1700
rect 261 1659 268 1670
rect 202 1658 268 1659
rect 602 1659 609 1670
rect 661 1700 668 1711
rect 1002 1711 1068 1712
rect 1002 1700 1009 1711
rect 661 1670 1009 1700
rect 661 1659 668 1670
rect 602 1658 668 1659
rect 1002 1659 1009 1670
rect 1061 1700 1068 1711
rect 1402 1711 1468 1712
rect 1402 1700 1409 1711
rect 1061 1670 1409 1700
rect 1061 1659 1068 1670
rect 1002 1658 1068 1659
rect 1402 1659 1409 1670
rect 1461 1700 1468 1711
rect 1802 1711 1868 1712
rect 1802 1700 1809 1711
rect 1461 1670 1809 1700
rect 1461 1659 1468 1670
rect 1402 1658 1468 1659
rect 1802 1659 1809 1670
rect 1861 1700 1868 1711
rect 2202 1711 2268 1712
rect 2202 1700 2209 1711
rect 1861 1670 2209 1700
rect 1861 1659 1868 1670
rect 1802 1658 1868 1659
rect 2202 1659 2209 1670
rect 2261 1700 2268 1711
rect 2602 1711 2668 1712
rect 2602 1700 2609 1711
rect 2261 1670 2609 1700
rect 2261 1659 2268 1670
rect 2202 1658 2268 1659
rect 2602 1659 2609 1670
rect 2661 1700 2668 1711
rect 3002 1711 3068 1712
rect 3002 1700 3009 1711
rect 2661 1670 3009 1700
rect 2661 1659 2668 1670
rect 2602 1658 2668 1659
rect 3002 1659 3009 1670
rect 3061 1700 3068 1711
rect 3402 1711 3468 1712
rect 3402 1700 3409 1711
rect 3061 1670 3409 1700
rect 3061 1659 3068 1670
rect 3002 1658 3068 1659
rect 3402 1659 3409 1670
rect 3461 1700 3468 1711
rect 3802 1711 3868 1712
rect 3802 1700 3809 1711
rect 3461 1670 3809 1700
rect 3461 1659 3468 1670
rect 3402 1658 3468 1659
rect 3802 1659 3809 1670
rect 3861 1700 3868 1711
rect 4202 1711 4268 1712
rect 4202 1700 4209 1711
rect 3861 1670 4209 1700
rect 3861 1659 3868 1670
rect 3802 1658 3868 1659
rect 4202 1659 4209 1670
rect 4261 1700 4268 1711
rect 4602 1711 4668 1712
rect 4602 1700 4609 1711
rect 4261 1670 4609 1700
rect 4261 1659 4268 1670
rect 4202 1658 4268 1659
rect 4602 1659 4609 1670
rect 4661 1700 4668 1711
rect 5002 1711 5068 1712
rect 5002 1700 5009 1711
rect 4661 1670 5009 1700
rect 4661 1659 4668 1670
rect 4602 1658 4668 1659
rect 5002 1659 5009 1670
rect 5061 1700 5068 1711
rect 5402 1711 5468 1712
rect 5402 1700 5409 1711
rect 5061 1670 5409 1700
rect 5061 1659 5068 1670
rect 5002 1658 5068 1659
rect 5402 1659 5409 1670
rect 5461 1700 5468 1711
rect 5802 1711 5868 1712
rect 5802 1700 5809 1711
rect 5461 1670 5809 1700
rect 5461 1659 5468 1670
rect 5402 1658 5468 1659
rect 5802 1659 5809 1670
rect 5861 1700 5868 1711
rect 6202 1711 6268 1712
rect 6202 1700 6209 1711
rect 5861 1670 6209 1700
rect 5861 1659 5868 1670
rect 5802 1658 5868 1659
rect 6202 1659 6209 1670
rect 6261 1700 6268 1711
rect 6704 1711 6770 1712
rect 6704 1700 6711 1711
rect 6261 1670 6711 1700
rect 6261 1659 6268 1670
rect 6202 1658 6268 1659
rect 6704 1659 6711 1670
rect 6763 1659 6770 1711
rect 6704 1658 6770 1659
rect 2 1641 68 1642
rect 2 1630 9 1641
rect 0 1600 9 1630
rect 2 1589 9 1600
rect 61 1630 68 1641
rect 402 1641 468 1642
rect 402 1630 409 1641
rect 61 1600 409 1630
rect 61 1589 68 1600
rect 2 1588 68 1589
rect 402 1589 409 1600
rect 461 1630 468 1641
rect 802 1641 868 1642
rect 802 1630 809 1641
rect 461 1600 809 1630
rect 461 1589 468 1600
rect 402 1588 468 1589
rect 802 1589 809 1600
rect 861 1630 868 1641
rect 1202 1641 1268 1642
rect 1202 1630 1209 1641
rect 861 1600 1209 1630
rect 861 1589 868 1600
rect 802 1588 868 1589
rect 1202 1589 1209 1600
rect 1261 1630 1268 1641
rect 1602 1641 1668 1642
rect 1602 1630 1609 1641
rect 1261 1600 1609 1630
rect 1261 1589 1268 1600
rect 1202 1588 1268 1589
rect 1602 1589 1609 1600
rect 1661 1630 1668 1641
rect 2002 1641 2068 1642
rect 2002 1630 2009 1641
rect 1661 1600 2009 1630
rect 1661 1589 1668 1600
rect 1602 1588 1668 1589
rect 2002 1589 2009 1600
rect 2061 1630 2068 1641
rect 2402 1641 2468 1642
rect 2402 1630 2409 1641
rect 2061 1600 2409 1630
rect 2061 1589 2068 1600
rect 2002 1588 2068 1589
rect 2402 1589 2409 1600
rect 2461 1630 2468 1641
rect 2802 1641 2868 1642
rect 2802 1630 2809 1641
rect 2461 1600 2809 1630
rect 2461 1589 2468 1600
rect 2402 1588 2468 1589
rect 2802 1589 2809 1600
rect 2861 1630 2868 1641
rect 3202 1641 3268 1642
rect 3202 1630 3209 1641
rect 2861 1600 3209 1630
rect 2861 1589 2868 1600
rect 2802 1588 2868 1589
rect 3202 1589 3209 1600
rect 3261 1630 3268 1641
rect 3602 1641 3668 1642
rect 3602 1630 3609 1641
rect 3261 1600 3609 1630
rect 3261 1589 3268 1600
rect 3202 1588 3268 1589
rect 3602 1589 3609 1600
rect 3661 1630 3668 1641
rect 4002 1641 4068 1642
rect 4002 1630 4009 1641
rect 3661 1600 4009 1630
rect 3661 1589 3668 1600
rect 3602 1588 3668 1589
rect 4002 1589 4009 1600
rect 4061 1630 4068 1641
rect 4402 1641 4468 1642
rect 4402 1630 4409 1641
rect 4061 1600 4409 1630
rect 4061 1589 4068 1600
rect 4002 1588 4068 1589
rect 4402 1589 4409 1600
rect 4461 1630 4468 1641
rect 4802 1641 4868 1642
rect 4802 1630 4809 1641
rect 4461 1600 4809 1630
rect 4461 1589 4468 1600
rect 4402 1588 4468 1589
rect 4802 1589 4809 1600
rect 4861 1630 4868 1641
rect 5202 1641 5268 1642
rect 5202 1630 5209 1641
rect 4861 1600 5209 1630
rect 4861 1589 4868 1600
rect 4802 1588 4868 1589
rect 5202 1589 5209 1600
rect 5261 1630 5268 1641
rect 5602 1641 5668 1642
rect 5602 1630 5609 1641
rect 5261 1600 5609 1630
rect 5261 1589 5268 1600
rect 5202 1588 5268 1589
rect 5602 1589 5609 1600
rect 5661 1630 5668 1641
rect 6002 1641 6068 1642
rect 6002 1630 6009 1641
rect 5661 1600 6009 1630
rect 5661 1589 5668 1600
rect 5602 1588 5668 1589
rect 6002 1589 6009 1600
rect 6061 1630 6068 1641
rect 6402 1641 6468 1642
rect 6402 1630 6409 1641
rect 6061 1600 6409 1630
rect 6061 1589 6068 1600
rect 6002 1588 6068 1589
rect 6402 1589 6409 1600
rect 6461 1630 6468 1641
rect 6500 1641 6566 1642
rect 6500 1630 6507 1641
rect 6461 1600 6507 1630
rect 6461 1589 6468 1600
rect 6402 1588 6468 1589
rect 6500 1589 6507 1600
rect 6559 1589 6566 1641
rect 6500 1588 6566 1589
rect 202 1571 268 1572
rect 202 1560 209 1571
rect 0 1530 209 1560
rect 202 1519 209 1530
rect 261 1560 268 1571
rect 602 1571 668 1572
rect 602 1560 609 1571
rect 261 1530 609 1560
rect 261 1519 268 1530
rect 202 1518 268 1519
rect 602 1519 609 1530
rect 661 1560 668 1571
rect 1002 1571 1068 1572
rect 1002 1560 1009 1571
rect 661 1530 1009 1560
rect 661 1519 668 1530
rect 602 1518 668 1519
rect 1002 1519 1009 1530
rect 1061 1560 1068 1571
rect 1402 1571 1468 1572
rect 1402 1560 1409 1571
rect 1061 1530 1409 1560
rect 1061 1519 1068 1530
rect 1002 1518 1068 1519
rect 1402 1519 1409 1530
rect 1461 1560 1468 1571
rect 1802 1571 1868 1572
rect 1802 1560 1809 1571
rect 1461 1530 1809 1560
rect 1461 1519 1468 1530
rect 1402 1518 1468 1519
rect 1802 1519 1809 1530
rect 1861 1560 1868 1571
rect 2202 1571 2268 1572
rect 2202 1560 2209 1571
rect 1861 1530 2209 1560
rect 1861 1519 1868 1530
rect 1802 1518 1868 1519
rect 2202 1519 2209 1530
rect 2261 1560 2268 1571
rect 2602 1571 2668 1572
rect 2602 1560 2609 1571
rect 2261 1530 2609 1560
rect 2261 1519 2268 1530
rect 2202 1518 2268 1519
rect 2602 1519 2609 1530
rect 2661 1560 2668 1571
rect 3002 1571 3068 1572
rect 3002 1560 3009 1571
rect 2661 1530 3009 1560
rect 2661 1519 2668 1530
rect 2602 1518 2668 1519
rect 3002 1519 3009 1530
rect 3061 1560 3068 1571
rect 3402 1571 3468 1572
rect 3402 1560 3409 1571
rect 3061 1530 3409 1560
rect 3061 1519 3068 1530
rect 3002 1518 3068 1519
rect 3402 1519 3409 1530
rect 3461 1560 3468 1571
rect 3802 1571 3868 1572
rect 3802 1560 3809 1571
rect 3461 1530 3809 1560
rect 3461 1519 3468 1530
rect 3402 1518 3468 1519
rect 3802 1519 3809 1530
rect 3861 1560 3868 1571
rect 4202 1571 4268 1572
rect 4202 1560 4209 1571
rect 3861 1530 4209 1560
rect 3861 1519 3868 1530
rect 3802 1518 3868 1519
rect 4202 1519 4209 1530
rect 4261 1560 4268 1571
rect 4602 1571 4668 1572
rect 4602 1560 4609 1571
rect 4261 1530 4609 1560
rect 4261 1519 4268 1530
rect 4202 1518 4268 1519
rect 4602 1519 4609 1530
rect 4661 1560 4668 1571
rect 5002 1571 5068 1572
rect 5002 1560 5009 1571
rect 4661 1530 5009 1560
rect 4661 1519 4668 1530
rect 4602 1518 4668 1519
rect 5002 1519 5009 1530
rect 5061 1560 5068 1571
rect 5402 1571 5468 1572
rect 5402 1560 5409 1571
rect 5061 1530 5409 1560
rect 5061 1519 5068 1530
rect 5002 1518 5068 1519
rect 5402 1519 5409 1530
rect 5461 1560 5468 1571
rect 5802 1571 5868 1572
rect 5802 1560 5809 1571
rect 5461 1530 5809 1560
rect 5461 1519 5468 1530
rect 5402 1518 5468 1519
rect 5802 1519 5809 1530
rect 5861 1560 5868 1571
rect 6202 1571 6268 1572
rect 6202 1560 6209 1571
rect 5861 1530 6209 1560
rect 5861 1519 5868 1530
rect 5802 1518 5868 1519
rect 6202 1519 6209 1530
rect 6261 1560 6268 1571
rect 6704 1571 6770 1572
rect 6704 1560 6711 1571
rect 6261 1530 6711 1560
rect 6261 1519 6268 1530
rect 6202 1518 6268 1519
rect 6704 1519 6711 1530
rect 6763 1519 6770 1571
rect 6704 1518 6770 1519
rect 2 1501 68 1502
rect 2 1490 9 1501
rect 0 1460 9 1490
rect 2 1449 9 1460
rect 61 1490 68 1501
rect 402 1501 468 1502
rect 402 1490 409 1501
rect 61 1460 409 1490
rect 61 1449 68 1460
rect 2 1448 68 1449
rect 402 1449 409 1460
rect 461 1490 468 1501
rect 802 1501 868 1502
rect 802 1490 809 1501
rect 461 1460 809 1490
rect 461 1449 468 1460
rect 402 1448 468 1449
rect 802 1449 809 1460
rect 861 1490 868 1501
rect 1202 1501 1268 1502
rect 1202 1490 1209 1501
rect 861 1460 1209 1490
rect 861 1449 868 1460
rect 802 1448 868 1449
rect 1202 1449 1209 1460
rect 1261 1490 1268 1501
rect 1602 1501 1668 1502
rect 1602 1490 1609 1501
rect 1261 1460 1609 1490
rect 1261 1449 1268 1460
rect 1202 1448 1268 1449
rect 1602 1449 1609 1460
rect 1661 1490 1668 1501
rect 2002 1501 2068 1502
rect 2002 1490 2009 1501
rect 1661 1460 2009 1490
rect 1661 1449 1668 1460
rect 1602 1448 1668 1449
rect 2002 1449 2009 1460
rect 2061 1490 2068 1501
rect 2402 1501 2468 1502
rect 2402 1490 2409 1501
rect 2061 1460 2409 1490
rect 2061 1449 2068 1460
rect 2002 1448 2068 1449
rect 2402 1449 2409 1460
rect 2461 1490 2468 1501
rect 2802 1501 2868 1502
rect 2802 1490 2809 1501
rect 2461 1460 2809 1490
rect 2461 1449 2468 1460
rect 2402 1448 2468 1449
rect 2802 1449 2809 1460
rect 2861 1490 2868 1501
rect 3202 1501 3268 1502
rect 3202 1490 3209 1501
rect 2861 1460 3209 1490
rect 2861 1449 2868 1460
rect 2802 1448 2868 1449
rect 3202 1449 3209 1460
rect 3261 1490 3268 1501
rect 3602 1501 3668 1502
rect 3602 1490 3609 1501
rect 3261 1460 3609 1490
rect 3261 1449 3268 1460
rect 3202 1448 3268 1449
rect 3602 1449 3609 1460
rect 3661 1490 3668 1501
rect 4002 1501 4068 1502
rect 4002 1490 4009 1501
rect 3661 1460 4009 1490
rect 3661 1449 3668 1460
rect 3602 1448 3668 1449
rect 4002 1449 4009 1460
rect 4061 1490 4068 1501
rect 4402 1501 4468 1502
rect 4402 1490 4409 1501
rect 4061 1460 4409 1490
rect 4061 1449 4068 1460
rect 4002 1448 4068 1449
rect 4402 1449 4409 1460
rect 4461 1490 4468 1501
rect 4802 1501 4868 1502
rect 4802 1490 4809 1501
rect 4461 1460 4809 1490
rect 4461 1449 4468 1460
rect 4402 1448 4468 1449
rect 4802 1449 4809 1460
rect 4861 1490 4868 1501
rect 5202 1501 5268 1502
rect 5202 1490 5209 1501
rect 4861 1460 5209 1490
rect 4861 1449 4868 1460
rect 4802 1448 4868 1449
rect 5202 1449 5209 1460
rect 5261 1490 5268 1501
rect 5602 1501 5668 1502
rect 5602 1490 5609 1501
rect 5261 1460 5609 1490
rect 5261 1449 5268 1460
rect 5202 1448 5268 1449
rect 5602 1449 5609 1460
rect 5661 1490 5668 1501
rect 6002 1501 6068 1502
rect 6002 1490 6009 1501
rect 5661 1460 6009 1490
rect 5661 1449 5668 1460
rect 5602 1448 5668 1449
rect 6002 1449 6009 1460
rect 6061 1490 6068 1501
rect 6402 1501 6468 1502
rect 6402 1490 6409 1501
rect 6061 1460 6409 1490
rect 6061 1449 6068 1460
rect 6002 1448 6068 1449
rect 6402 1449 6409 1460
rect 6461 1490 6468 1501
rect 6500 1501 6566 1502
rect 6500 1490 6507 1501
rect 6461 1460 6507 1490
rect 6461 1449 6468 1460
rect 6402 1448 6468 1449
rect 6500 1449 6507 1460
rect 6559 1449 6566 1501
rect 6500 1448 6566 1449
rect 202 1431 268 1432
rect 202 1420 209 1431
rect 0 1390 209 1420
rect 202 1379 209 1390
rect 261 1420 268 1431
rect 602 1431 668 1432
rect 602 1420 609 1431
rect 261 1390 609 1420
rect 261 1379 268 1390
rect 202 1378 268 1379
rect 602 1379 609 1390
rect 661 1420 668 1431
rect 1002 1431 1068 1432
rect 1002 1420 1009 1431
rect 661 1390 1009 1420
rect 661 1379 668 1390
rect 602 1378 668 1379
rect 1002 1379 1009 1390
rect 1061 1420 1068 1431
rect 1402 1431 1468 1432
rect 1402 1420 1409 1431
rect 1061 1390 1409 1420
rect 1061 1379 1068 1390
rect 1002 1378 1068 1379
rect 1402 1379 1409 1390
rect 1461 1420 1468 1431
rect 1802 1431 1868 1432
rect 1802 1420 1809 1431
rect 1461 1390 1809 1420
rect 1461 1379 1468 1390
rect 1402 1378 1468 1379
rect 1802 1379 1809 1390
rect 1861 1420 1868 1431
rect 2202 1431 2268 1432
rect 2202 1420 2209 1431
rect 1861 1390 2209 1420
rect 1861 1379 1868 1390
rect 1802 1378 1868 1379
rect 2202 1379 2209 1390
rect 2261 1420 2268 1431
rect 2602 1431 2668 1432
rect 2602 1420 2609 1431
rect 2261 1390 2609 1420
rect 2261 1379 2268 1390
rect 2202 1378 2268 1379
rect 2602 1379 2609 1390
rect 2661 1420 2668 1431
rect 3002 1431 3068 1432
rect 3002 1420 3009 1431
rect 2661 1390 3009 1420
rect 2661 1379 2668 1390
rect 2602 1378 2668 1379
rect 3002 1379 3009 1390
rect 3061 1420 3068 1431
rect 3402 1431 3468 1432
rect 3402 1420 3409 1431
rect 3061 1390 3409 1420
rect 3061 1379 3068 1390
rect 3002 1378 3068 1379
rect 3402 1379 3409 1390
rect 3461 1420 3468 1431
rect 3802 1431 3868 1432
rect 3802 1420 3809 1431
rect 3461 1390 3809 1420
rect 3461 1379 3468 1390
rect 3402 1378 3468 1379
rect 3802 1379 3809 1390
rect 3861 1420 3868 1431
rect 4202 1431 4268 1432
rect 4202 1420 4209 1431
rect 3861 1390 4209 1420
rect 3861 1379 3868 1390
rect 3802 1378 3868 1379
rect 4202 1379 4209 1390
rect 4261 1420 4268 1431
rect 4602 1431 4668 1432
rect 4602 1420 4609 1431
rect 4261 1390 4609 1420
rect 4261 1379 4268 1390
rect 4202 1378 4268 1379
rect 4602 1379 4609 1390
rect 4661 1420 4668 1431
rect 5002 1431 5068 1432
rect 5002 1420 5009 1431
rect 4661 1390 5009 1420
rect 4661 1379 4668 1390
rect 4602 1378 4668 1379
rect 5002 1379 5009 1390
rect 5061 1420 5068 1431
rect 5402 1431 5468 1432
rect 5402 1420 5409 1431
rect 5061 1390 5409 1420
rect 5061 1379 5068 1390
rect 5002 1378 5068 1379
rect 5402 1379 5409 1390
rect 5461 1420 5468 1431
rect 5802 1431 5868 1432
rect 5802 1420 5809 1431
rect 5461 1390 5809 1420
rect 5461 1379 5468 1390
rect 5402 1378 5468 1379
rect 5802 1379 5809 1390
rect 5861 1420 5868 1431
rect 6202 1431 6268 1432
rect 6202 1420 6209 1431
rect 5861 1390 6209 1420
rect 5861 1379 5868 1390
rect 5802 1378 5868 1379
rect 6202 1379 6209 1390
rect 6261 1420 6268 1431
rect 6704 1431 6770 1432
rect 6704 1420 6711 1431
rect 6261 1390 6711 1420
rect 6261 1379 6268 1390
rect 6202 1378 6268 1379
rect 6704 1379 6711 1390
rect 6763 1379 6770 1431
rect 6704 1378 6770 1379
rect 2 1361 68 1362
rect 2 1350 9 1361
rect 0 1320 9 1350
rect 2 1309 9 1320
rect 61 1350 68 1361
rect 402 1361 468 1362
rect 402 1350 409 1361
rect 61 1320 409 1350
rect 61 1309 68 1320
rect 2 1308 68 1309
rect 402 1309 409 1320
rect 461 1350 468 1361
rect 802 1361 868 1362
rect 802 1350 809 1361
rect 461 1320 809 1350
rect 461 1309 468 1320
rect 402 1308 468 1309
rect 802 1309 809 1320
rect 861 1350 868 1361
rect 1202 1361 1268 1362
rect 1202 1350 1209 1361
rect 861 1320 1209 1350
rect 861 1309 868 1320
rect 802 1308 868 1309
rect 1202 1309 1209 1320
rect 1261 1350 1268 1361
rect 1602 1361 1668 1362
rect 1602 1350 1609 1361
rect 1261 1320 1609 1350
rect 1261 1309 1268 1320
rect 1202 1308 1268 1309
rect 1602 1309 1609 1320
rect 1661 1350 1668 1361
rect 2002 1361 2068 1362
rect 2002 1350 2009 1361
rect 1661 1320 2009 1350
rect 1661 1309 1668 1320
rect 1602 1308 1668 1309
rect 2002 1309 2009 1320
rect 2061 1350 2068 1361
rect 2402 1361 2468 1362
rect 2402 1350 2409 1361
rect 2061 1320 2409 1350
rect 2061 1309 2068 1320
rect 2002 1308 2068 1309
rect 2402 1309 2409 1320
rect 2461 1350 2468 1361
rect 2802 1361 2868 1362
rect 2802 1350 2809 1361
rect 2461 1320 2809 1350
rect 2461 1309 2468 1320
rect 2402 1308 2468 1309
rect 2802 1309 2809 1320
rect 2861 1350 2868 1361
rect 3202 1361 3268 1362
rect 3202 1350 3209 1361
rect 2861 1320 3209 1350
rect 2861 1309 2868 1320
rect 2802 1308 2868 1309
rect 3202 1309 3209 1320
rect 3261 1350 3268 1361
rect 3602 1361 3668 1362
rect 3602 1350 3609 1361
rect 3261 1320 3609 1350
rect 3261 1309 3268 1320
rect 3202 1308 3268 1309
rect 3602 1309 3609 1320
rect 3661 1350 3668 1361
rect 4002 1361 4068 1362
rect 4002 1350 4009 1361
rect 3661 1320 4009 1350
rect 3661 1309 3668 1320
rect 3602 1308 3668 1309
rect 4002 1309 4009 1320
rect 4061 1350 4068 1361
rect 4402 1361 4468 1362
rect 4402 1350 4409 1361
rect 4061 1320 4409 1350
rect 4061 1309 4068 1320
rect 4002 1308 4068 1309
rect 4402 1309 4409 1320
rect 4461 1350 4468 1361
rect 4802 1361 4868 1362
rect 4802 1350 4809 1361
rect 4461 1320 4809 1350
rect 4461 1309 4468 1320
rect 4402 1308 4468 1309
rect 4802 1309 4809 1320
rect 4861 1350 4868 1361
rect 5202 1361 5268 1362
rect 5202 1350 5209 1361
rect 4861 1320 5209 1350
rect 4861 1309 4868 1320
rect 4802 1308 4868 1309
rect 5202 1309 5209 1320
rect 5261 1350 5268 1361
rect 5602 1361 5668 1362
rect 5602 1350 5609 1361
rect 5261 1320 5609 1350
rect 5261 1309 5268 1320
rect 5202 1308 5268 1309
rect 5602 1309 5609 1320
rect 5661 1350 5668 1361
rect 6002 1361 6068 1362
rect 6002 1350 6009 1361
rect 5661 1320 6009 1350
rect 5661 1309 5668 1320
rect 5602 1308 5668 1309
rect 6002 1309 6009 1320
rect 6061 1350 6068 1361
rect 6402 1361 6468 1362
rect 6402 1350 6409 1361
rect 6061 1320 6409 1350
rect 6061 1309 6068 1320
rect 6002 1308 6068 1309
rect 6402 1309 6409 1320
rect 6461 1350 6468 1361
rect 6500 1361 6566 1362
rect 6500 1350 6507 1361
rect 6461 1320 6507 1350
rect 6461 1309 6468 1320
rect 6402 1308 6468 1309
rect 6500 1309 6507 1320
rect 6559 1309 6566 1361
rect 6500 1308 6566 1309
rect 196 1291 274 1292
rect -4 1275 74 1276
rect -4 1219 7 1275
rect 63 1219 74 1275
rect 196 1235 207 1291
rect 263 1235 274 1291
rect 596 1291 674 1292
rect 196 1234 274 1235
rect 396 1275 474 1276
rect -4 1218 74 1219
rect 396 1219 407 1275
rect 463 1219 474 1275
rect 596 1235 607 1291
rect 663 1235 674 1291
rect 996 1291 1074 1292
rect 596 1234 674 1235
rect 796 1275 874 1276
rect 396 1218 474 1219
rect 796 1219 807 1275
rect 863 1219 874 1275
rect 996 1235 1007 1291
rect 1063 1235 1074 1291
rect 1396 1291 1474 1292
rect 996 1234 1074 1235
rect 1196 1275 1274 1276
rect 796 1218 874 1219
rect 1196 1219 1207 1275
rect 1263 1219 1274 1275
rect 1396 1235 1407 1291
rect 1463 1235 1474 1291
rect 1796 1291 1874 1292
rect 1396 1234 1474 1235
rect 1596 1275 1674 1276
rect 1196 1218 1274 1219
rect 1596 1219 1607 1275
rect 1663 1219 1674 1275
rect 1796 1235 1807 1291
rect 1863 1235 1874 1291
rect 2196 1291 2274 1292
rect 1796 1234 1874 1235
rect 1996 1275 2074 1276
rect 1596 1218 1674 1219
rect 1996 1219 2007 1275
rect 2063 1219 2074 1275
rect 2196 1235 2207 1291
rect 2263 1235 2274 1291
rect 2596 1291 2674 1292
rect 2196 1234 2274 1235
rect 2396 1275 2474 1276
rect 1996 1218 2074 1219
rect 2396 1219 2407 1275
rect 2463 1219 2474 1275
rect 2596 1235 2607 1291
rect 2663 1235 2674 1291
rect 2996 1291 3074 1292
rect 2596 1234 2674 1235
rect 2796 1275 2874 1276
rect 2396 1218 2474 1219
rect 2796 1219 2807 1275
rect 2863 1219 2874 1275
rect 2996 1235 3007 1291
rect 3063 1235 3074 1291
rect 3396 1291 3474 1292
rect 2996 1234 3074 1235
rect 3196 1275 3274 1276
rect 2796 1218 2874 1219
rect 3196 1219 3207 1275
rect 3263 1219 3274 1275
rect 3396 1235 3407 1291
rect 3463 1235 3474 1291
rect 3796 1291 3874 1292
rect 3396 1234 3474 1235
rect 3596 1275 3674 1276
rect 3196 1218 3274 1219
rect 3596 1219 3607 1275
rect 3663 1219 3674 1275
rect 3796 1235 3807 1291
rect 3863 1235 3874 1291
rect 4196 1291 4274 1292
rect 3796 1234 3874 1235
rect 3996 1275 4074 1276
rect 3596 1218 3674 1219
rect 3996 1219 4007 1275
rect 4063 1219 4074 1275
rect 4196 1235 4207 1291
rect 4263 1235 4274 1291
rect 4596 1291 4674 1292
rect 4196 1234 4274 1235
rect 4396 1275 4474 1276
rect 3996 1218 4074 1219
rect 4396 1219 4407 1275
rect 4463 1219 4474 1275
rect 4596 1235 4607 1291
rect 4663 1235 4674 1291
rect 4996 1291 5074 1292
rect 4596 1234 4674 1235
rect 4796 1275 4874 1276
rect 4396 1218 4474 1219
rect 4796 1219 4807 1275
rect 4863 1219 4874 1275
rect 4996 1235 5007 1291
rect 5063 1235 5074 1291
rect 5396 1291 5474 1292
rect 4996 1234 5074 1235
rect 5196 1275 5274 1276
rect 4796 1218 4874 1219
rect 5196 1219 5207 1275
rect 5263 1219 5274 1275
rect 5396 1235 5407 1291
rect 5463 1235 5474 1291
rect 5796 1291 5874 1292
rect 5396 1234 5474 1235
rect 5596 1275 5674 1276
rect 5196 1218 5274 1219
rect 5596 1219 5607 1275
rect 5663 1219 5674 1275
rect 5796 1235 5807 1291
rect 5863 1235 5874 1291
rect 6196 1291 6274 1292
rect 5796 1234 5874 1235
rect 5996 1275 6074 1276
rect 5596 1218 5674 1219
rect 5996 1219 6007 1275
rect 6063 1219 6074 1275
rect 6196 1235 6207 1291
rect 6263 1235 6274 1291
rect 6196 1234 6274 1235
rect 5996 1218 6074 1219
rect 202 1201 268 1202
rect 202 1190 209 1201
rect 0 1160 209 1190
rect 202 1149 209 1160
rect 261 1190 268 1201
rect 602 1201 668 1202
rect 602 1190 609 1201
rect 261 1160 609 1190
rect 261 1149 268 1160
rect 202 1148 268 1149
rect 602 1149 609 1160
rect 661 1190 668 1201
rect 1002 1201 1068 1202
rect 1002 1190 1009 1201
rect 661 1160 1009 1190
rect 661 1149 668 1160
rect 602 1148 668 1149
rect 1002 1149 1009 1160
rect 1061 1190 1068 1201
rect 1402 1201 1468 1202
rect 1402 1190 1409 1201
rect 1061 1160 1409 1190
rect 1061 1149 1068 1160
rect 1002 1148 1068 1149
rect 1402 1149 1409 1160
rect 1461 1190 1468 1201
rect 1802 1201 1868 1202
rect 1802 1190 1809 1201
rect 1461 1160 1809 1190
rect 1461 1149 1468 1160
rect 1402 1148 1468 1149
rect 1802 1149 1809 1160
rect 1861 1190 1868 1201
rect 2202 1201 2268 1202
rect 2202 1190 2209 1201
rect 1861 1160 2209 1190
rect 1861 1149 1868 1160
rect 1802 1148 1868 1149
rect 2202 1149 2209 1160
rect 2261 1190 2268 1201
rect 2602 1201 2668 1202
rect 2602 1190 2609 1201
rect 2261 1160 2609 1190
rect 2261 1149 2268 1160
rect 2202 1148 2268 1149
rect 2602 1149 2609 1160
rect 2661 1190 2668 1201
rect 3002 1201 3068 1202
rect 3002 1190 3009 1201
rect 2661 1160 3009 1190
rect 2661 1149 2668 1160
rect 2602 1148 2668 1149
rect 3002 1149 3009 1160
rect 3061 1190 3068 1201
rect 3402 1201 3468 1202
rect 3402 1190 3409 1201
rect 3061 1160 3409 1190
rect 3061 1149 3068 1160
rect 3002 1148 3068 1149
rect 3402 1149 3409 1160
rect 3461 1190 3468 1201
rect 3802 1201 3868 1202
rect 3802 1190 3809 1201
rect 3461 1160 3809 1190
rect 3461 1149 3468 1160
rect 3402 1148 3468 1149
rect 3802 1149 3809 1160
rect 3861 1190 3868 1201
rect 4202 1201 4268 1202
rect 4202 1190 4209 1201
rect 3861 1160 4209 1190
rect 3861 1149 3868 1160
rect 3802 1148 3868 1149
rect 4202 1149 4209 1160
rect 4261 1190 4268 1201
rect 4602 1201 4668 1202
rect 4602 1190 4609 1201
rect 4261 1160 4609 1190
rect 4261 1149 4268 1160
rect 4202 1148 4268 1149
rect 4602 1149 4609 1160
rect 4661 1190 4668 1201
rect 5002 1201 5068 1202
rect 5002 1190 5009 1201
rect 4661 1160 5009 1190
rect 4661 1149 4668 1160
rect 4602 1148 4668 1149
rect 5002 1149 5009 1160
rect 5061 1190 5068 1201
rect 5402 1201 5468 1202
rect 5402 1190 5409 1201
rect 5061 1160 5409 1190
rect 5061 1149 5068 1160
rect 5002 1148 5068 1149
rect 5402 1149 5409 1160
rect 5461 1190 5468 1201
rect 5802 1201 5868 1202
rect 5802 1190 5809 1201
rect 5461 1160 5809 1190
rect 5461 1149 5468 1160
rect 5402 1148 5468 1149
rect 5802 1149 5809 1160
rect 5861 1190 5868 1201
rect 6202 1201 6268 1202
rect 6202 1190 6209 1201
rect 5861 1160 6209 1190
rect 5861 1149 5868 1160
rect 5802 1148 5868 1149
rect 6202 1149 6209 1160
rect 6261 1190 6268 1201
rect 6704 1201 6770 1202
rect 6704 1190 6711 1201
rect 6261 1160 6711 1190
rect 6261 1149 6268 1160
rect 6202 1148 6268 1149
rect 6704 1149 6711 1160
rect 6763 1149 6770 1201
rect 6704 1148 6770 1149
rect 2 1131 68 1132
rect 2 1120 9 1131
rect 0 1090 9 1120
rect 2 1079 9 1090
rect 61 1120 68 1131
rect 402 1131 468 1132
rect 402 1120 409 1131
rect 61 1090 409 1120
rect 61 1079 68 1090
rect 2 1078 68 1079
rect 402 1079 409 1090
rect 461 1120 468 1131
rect 802 1131 868 1132
rect 802 1120 809 1131
rect 461 1090 809 1120
rect 461 1079 468 1090
rect 402 1078 468 1079
rect 802 1079 809 1090
rect 861 1120 868 1131
rect 1202 1131 1268 1132
rect 1202 1120 1209 1131
rect 861 1090 1209 1120
rect 861 1079 868 1090
rect 802 1078 868 1079
rect 1202 1079 1209 1090
rect 1261 1120 1268 1131
rect 1602 1131 1668 1132
rect 1602 1120 1609 1131
rect 1261 1090 1609 1120
rect 1261 1079 1268 1090
rect 1202 1078 1268 1079
rect 1602 1079 1609 1090
rect 1661 1120 1668 1131
rect 2002 1131 2068 1132
rect 2002 1120 2009 1131
rect 1661 1090 2009 1120
rect 1661 1079 1668 1090
rect 1602 1078 1668 1079
rect 2002 1079 2009 1090
rect 2061 1120 2068 1131
rect 2402 1131 2468 1132
rect 2402 1120 2409 1131
rect 2061 1090 2409 1120
rect 2061 1079 2068 1090
rect 2002 1078 2068 1079
rect 2402 1079 2409 1090
rect 2461 1120 2468 1131
rect 2802 1131 2868 1132
rect 2802 1120 2809 1131
rect 2461 1090 2809 1120
rect 2461 1079 2468 1090
rect 2402 1078 2468 1079
rect 2802 1079 2809 1090
rect 2861 1120 2868 1131
rect 3202 1131 3268 1132
rect 3202 1120 3209 1131
rect 2861 1090 3209 1120
rect 2861 1079 2868 1090
rect 2802 1078 2868 1079
rect 3202 1079 3209 1090
rect 3261 1120 3268 1131
rect 3602 1131 3668 1132
rect 3602 1120 3609 1131
rect 3261 1090 3609 1120
rect 3261 1079 3268 1090
rect 3202 1078 3268 1079
rect 3602 1079 3609 1090
rect 3661 1120 3668 1131
rect 4002 1131 4068 1132
rect 4002 1120 4009 1131
rect 3661 1090 4009 1120
rect 3661 1079 3668 1090
rect 3602 1078 3668 1079
rect 4002 1079 4009 1090
rect 4061 1120 4068 1131
rect 4402 1131 4468 1132
rect 4402 1120 4409 1131
rect 4061 1090 4409 1120
rect 4061 1079 4068 1090
rect 4002 1078 4068 1079
rect 4402 1079 4409 1090
rect 4461 1120 4468 1131
rect 4802 1131 4868 1132
rect 4802 1120 4809 1131
rect 4461 1090 4809 1120
rect 4461 1079 4468 1090
rect 4402 1078 4468 1079
rect 4802 1079 4809 1090
rect 4861 1120 4868 1131
rect 5202 1131 5268 1132
rect 5202 1120 5209 1131
rect 4861 1090 5209 1120
rect 4861 1079 4868 1090
rect 4802 1078 4868 1079
rect 5202 1079 5209 1090
rect 5261 1120 5268 1131
rect 5602 1131 5668 1132
rect 5602 1120 5609 1131
rect 5261 1090 5609 1120
rect 5261 1079 5268 1090
rect 5202 1078 5268 1079
rect 5602 1079 5609 1090
rect 5661 1120 5668 1131
rect 6002 1131 6068 1132
rect 6002 1120 6009 1131
rect 5661 1090 6009 1120
rect 5661 1079 5668 1090
rect 5602 1078 5668 1079
rect 6002 1079 6009 1090
rect 6061 1120 6068 1131
rect 6402 1131 6468 1132
rect 6402 1120 6409 1131
rect 6061 1090 6409 1120
rect 6061 1079 6068 1090
rect 6002 1078 6068 1079
rect 6402 1079 6409 1090
rect 6461 1120 6468 1131
rect 6500 1131 6566 1132
rect 6500 1120 6507 1131
rect 6461 1090 6507 1120
rect 6461 1079 6468 1090
rect 6402 1078 6468 1079
rect 6500 1079 6507 1090
rect 6559 1079 6566 1131
rect 6500 1078 6566 1079
rect 202 1061 268 1062
rect 202 1050 209 1061
rect 0 1020 209 1050
rect 202 1009 209 1020
rect 261 1050 268 1061
rect 602 1061 668 1062
rect 602 1050 609 1061
rect 261 1020 609 1050
rect 261 1009 268 1020
rect 202 1008 268 1009
rect 602 1009 609 1020
rect 661 1050 668 1061
rect 1002 1061 1068 1062
rect 1002 1050 1009 1061
rect 661 1020 1009 1050
rect 661 1009 668 1020
rect 602 1008 668 1009
rect 1002 1009 1009 1020
rect 1061 1050 1068 1061
rect 1402 1061 1468 1062
rect 1402 1050 1409 1061
rect 1061 1020 1409 1050
rect 1061 1009 1068 1020
rect 1002 1008 1068 1009
rect 1402 1009 1409 1020
rect 1461 1050 1468 1061
rect 1802 1061 1868 1062
rect 1802 1050 1809 1061
rect 1461 1020 1809 1050
rect 1461 1009 1468 1020
rect 1402 1008 1468 1009
rect 1802 1009 1809 1020
rect 1861 1050 1868 1061
rect 2202 1061 2268 1062
rect 2202 1050 2209 1061
rect 1861 1020 2209 1050
rect 1861 1009 1868 1020
rect 1802 1008 1868 1009
rect 2202 1009 2209 1020
rect 2261 1050 2268 1061
rect 2602 1061 2668 1062
rect 2602 1050 2609 1061
rect 2261 1020 2609 1050
rect 2261 1009 2268 1020
rect 2202 1008 2268 1009
rect 2602 1009 2609 1020
rect 2661 1050 2668 1061
rect 3002 1061 3068 1062
rect 3002 1050 3009 1061
rect 2661 1020 3009 1050
rect 2661 1009 2668 1020
rect 2602 1008 2668 1009
rect 3002 1009 3009 1020
rect 3061 1050 3068 1061
rect 3402 1061 3468 1062
rect 3402 1050 3409 1061
rect 3061 1020 3409 1050
rect 3061 1009 3068 1020
rect 3002 1008 3068 1009
rect 3402 1009 3409 1020
rect 3461 1050 3468 1061
rect 3802 1061 3868 1062
rect 3802 1050 3809 1061
rect 3461 1020 3809 1050
rect 3461 1009 3468 1020
rect 3402 1008 3468 1009
rect 3802 1009 3809 1020
rect 3861 1050 3868 1061
rect 4202 1061 4268 1062
rect 4202 1050 4209 1061
rect 3861 1020 4209 1050
rect 3861 1009 3868 1020
rect 3802 1008 3868 1009
rect 4202 1009 4209 1020
rect 4261 1050 4268 1061
rect 4602 1061 4668 1062
rect 4602 1050 4609 1061
rect 4261 1020 4609 1050
rect 4261 1009 4268 1020
rect 4202 1008 4268 1009
rect 4602 1009 4609 1020
rect 4661 1050 4668 1061
rect 5002 1061 5068 1062
rect 5002 1050 5009 1061
rect 4661 1020 5009 1050
rect 4661 1009 4668 1020
rect 4602 1008 4668 1009
rect 5002 1009 5009 1020
rect 5061 1050 5068 1061
rect 5402 1061 5468 1062
rect 5402 1050 5409 1061
rect 5061 1020 5409 1050
rect 5061 1009 5068 1020
rect 5002 1008 5068 1009
rect 5402 1009 5409 1020
rect 5461 1050 5468 1061
rect 5802 1061 5868 1062
rect 5802 1050 5809 1061
rect 5461 1020 5809 1050
rect 5461 1009 5468 1020
rect 5402 1008 5468 1009
rect 5802 1009 5809 1020
rect 5861 1050 5868 1061
rect 6202 1061 6268 1062
rect 6202 1050 6209 1061
rect 5861 1020 6209 1050
rect 5861 1009 5868 1020
rect 5802 1008 5868 1009
rect 6202 1009 6209 1020
rect 6261 1050 6268 1061
rect 6704 1061 6770 1062
rect 6704 1050 6711 1061
rect 6261 1020 6711 1050
rect 6261 1009 6268 1020
rect 6202 1008 6268 1009
rect 6704 1009 6711 1020
rect 6763 1009 6770 1061
rect 6704 1008 6770 1009
rect 2 991 68 992
rect 2 980 9 991
rect 0 950 9 980
rect 2 939 9 950
rect 61 980 68 991
rect 402 991 468 992
rect 402 980 409 991
rect 61 950 409 980
rect 61 939 68 950
rect 2 938 68 939
rect 402 939 409 950
rect 461 980 468 991
rect 802 991 868 992
rect 802 980 809 991
rect 461 950 809 980
rect 461 939 468 950
rect 402 938 468 939
rect 802 939 809 950
rect 861 980 868 991
rect 1202 991 1268 992
rect 1202 980 1209 991
rect 861 950 1209 980
rect 861 939 868 950
rect 802 938 868 939
rect 1202 939 1209 950
rect 1261 980 1268 991
rect 1602 991 1668 992
rect 1602 980 1609 991
rect 1261 950 1609 980
rect 1261 939 1268 950
rect 1202 938 1268 939
rect 1602 939 1609 950
rect 1661 980 1668 991
rect 2002 991 2068 992
rect 2002 980 2009 991
rect 1661 950 2009 980
rect 1661 939 1668 950
rect 1602 938 1668 939
rect 2002 939 2009 950
rect 2061 980 2068 991
rect 2402 991 2468 992
rect 2402 980 2409 991
rect 2061 950 2409 980
rect 2061 939 2068 950
rect 2002 938 2068 939
rect 2402 939 2409 950
rect 2461 980 2468 991
rect 2802 991 2868 992
rect 2802 980 2809 991
rect 2461 950 2809 980
rect 2461 939 2468 950
rect 2402 938 2468 939
rect 2802 939 2809 950
rect 2861 980 2868 991
rect 3202 991 3268 992
rect 3202 980 3209 991
rect 2861 950 3209 980
rect 2861 939 2868 950
rect 2802 938 2868 939
rect 3202 939 3209 950
rect 3261 980 3268 991
rect 3602 991 3668 992
rect 3602 980 3609 991
rect 3261 950 3609 980
rect 3261 939 3268 950
rect 3202 938 3268 939
rect 3602 939 3609 950
rect 3661 980 3668 991
rect 4002 991 4068 992
rect 4002 980 4009 991
rect 3661 950 4009 980
rect 3661 939 3668 950
rect 3602 938 3668 939
rect 4002 939 4009 950
rect 4061 980 4068 991
rect 4402 991 4468 992
rect 4402 980 4409 991
rect 4061 950 4409 980
rect 4061 939 4068 950
rect 4002 938 4068 939
rect 4402 939 4409 950
rect 4461 980 4468 991
rect 4802 991 4868 992
rect 4802 980 4809 991
rect 4461 950 4809 980
rect 4461 939 4468 950
rect 4402 938 4468 939
rect 4802 939 4809 950
rect 4861 980 4868 991
rect 5202 991 5268 992
rect 5202 980 5209 991
rect 4861 950 5209 980
rect 4861 939 4868 950
rect 4802 938 4868 939
rect 5202 939 5209 950
rect 5261 980 5268 991
rect 5602 991 5668 992
rect 5602 980 5609 991
rect 5261 950 5609 980
rect 5261 939 5268 950
rect 5202 938 5268 939
rect 5602 939 5609 950
rect 5661 980 5668 991
rect 6002 991 6068 992
rect 6002 980 6009 991
rect 5661 950 6009 980
rect 5661 939 5668 950
rect 5602 938 5668 939
rect 6002 939 6009 950
rect 6061 980 6068 991
rect 6402 991 6468 992
rect 6402 980 6409 991
rect 6061 950 6409 980
rect 6061 939 6068 950
rect 6002 938 6068 939
rect 6402 939 6409 950
rect 6461 980 6468 991
rect 6500 991 6566 992
rect 6500 980 6507 991
rect 6461 950 6507 980
rect 6461 939 6468 950
rect 6402 938 6468 939
rect 6500 939 6507 950
rect 6559 939 6566 991
rect 6500 938 6566 939
rect 202 921 268 922
rect 202 910 209 921
rect 0 880 209 910
rect 202 869 209 880
rect 261 910 268 921
rect 602 921 668 922
rect 602 910 609 921
rect 261 880 609 910
rect 261 869 268 880
rect 202 868 268 869
rect 602 869 609 880
rect 661 910 668 921
rect 1002 921 1068 922
rect 1002 910 1009 921
rect 661 880 1009 910
rect 661 869 668 880
rect 602 868 668 869
rect 1002 869 1009 880
rect 1061 910 1068 921
rect 1402 921 1468 922
rect 1402 910 1409 921
rect 1061 880 1409 910
rect 1061 869 1068 880
rect 1002 868 1068 869
rect 1402 869 1409 880
rect 1461 910 1468 921
rect 1802 921 1868 922
rect 1802 910 1809 921
rect 1461 880 1809 910
rect 1461 869 1468 880
rect 1402 868 1468 869
rect 1802 869 1809 880
rect 1861 910 1868 921
rect 2202 921 2268 922
rect 2202 910 2209 921
rect 1861 880 2209 910
rect 1861 869 1868 880
rect 1802 868 1868 869
rect 2202 869 2209 880
rect 2261 910 2268 921
rect 2602 921 2668 922
rect 2602 910 2609 921
rect 2261 880 2609 910
rect 2261 869 2268 880
rect 2202 868 2268 869
rect 2602 869 2609 880
rect 2661 910 2668 921
rect 3002 921 3068 922
rect 3002 910 3009 921
rect 2661 880 3009 910
rect 2661 869 2668 880
rect 2602 868 2668 869
rect 3002 869 3009 880
rect 3061 910 3068 921
rect 3402 921 3468 922
rect 3402 910 3409 921
rect 3061 880 3409 910
rect 3061 869 3068 880
rect 3002 868 3068 869
rect 3402 869 3409 880
rect 3461 910 3468 921
rect 3802 921 3868 922
rect 3802 910 3809 921
rect 3461 880 3809 910
rect 3461 869 3468 880
rect 3402 868 3468 869
rect 3802 869 3809 880
rect 3861 910 3868 921
rect 4202 921 4268 922
rect 4202 910 4209 921
rect 3861 880 4209 910
rect 3861 869 3868 880
rect 3802 868 3868 869
rect 4202 869 4209 880
rect 4261 910 4268 921
rect 4602 921 4668 922
rect 4602 910 4609 921
rect 4261 880 4609 910
rect 4261 869 4268 880
rect 4202 868 4268 869
rect 4602 869 4609 880
rect 4661 910 4668 921
rect 5002 921 5068 922
rect 5002 910 5009 921
rect 4661 880 5009 910
rect 4661 869 4668 880
rect 4602 868 4668 869
rect 5002 869 5009 880
rect 5061 910 5068 921
rect 5402 921 5468 922
rect 5402 910 5409 921
rect 5061 880 5409 910
rect 5061 869 5068 880
rect 5002 868 5068 869
rect 5402 869 5409 880
rect 5461 910 5468 921
rect 5802 921 5868 922
rect 5802 910 5809 921
rect 5461 880 5809 910
rect 5461 869 5468 880
rect 5402 868 5468 869
rect 5802 869 5809 880
rect 5861 910 5868 921
rect 6202 921 6268 922
rect 6202 910 6209 921
rect 5861 880 6209 910
rect 5861 869 5868 880
rect 5802 868 5868 869
rect 6202 869 6209 880
rect 6261 910 6268 921
rect 6704 921 6770 922
rect 6704 910 6711 921
rect 6261 880 6711 910
rect 6261 869 6268 880
rect 6202 868 6268 869
rect 6704 869 6711 880
rect 6763 869 6770 921
rect 6704 868 6770 869
rect 2 851 68 852
rect 2 840 9 851
rect 0 810 9 840
rect 2 799 9 810
rect 61 840 68 851
rect 402 851 468 852
rect 402 840 409 851
rect 61 810 409 840
rect 61 799 68 810
rect 2 798 68 799
rect 402 799 409 810
rect 461 840 468 851
rect 802 851 868 852
rect 802 840 809 851
rect 461 810 809 840
rect 461 799 468 810
rect 402 798 468 799
rect 802 799 809 810
rect 861 840 868 851
rect 1202 851 1268 852
rect 1202 840 1209 851
rect 861 810 1209 840
rect 861 799 868 810
rect 802 798 868 799
rect 1202 799 1209 810
rect 1261 840 1268 851
rect 1602 851 1668 852
rect 1602 840 1609 851
rect 1261 810 1609 840
rect 1261 799 1268 810
rect 1202 798 1268 799
rect 1602 799 1609 810
rect 1661 840 1668 851
rect 2002 851 2068 852
rect 2002 840 2009 851
rect 1661 810 2009 840
rect 1661 799 1668 810
rect 1602 798 1668 799
rect 2002 799 2009 810
rect 2061 840 2068 851
rect 2402 851 2468 852
rect 2402 840 2409 851
rect 2061 810 2409 840
rect 2061 799 2068 810
rect 2002 798 2068 799
rect 2402 799 2409 810
rect 2461 840 2468 851
rect 2802 851 2868 852
rect 2802 840 2809 851
rect 2461 810 2809 840
rect 2461 799 2468 810
rect 2402 798 2468 799
rect 2802 799 2809 810
rect 2861 840 2868 851
rect 3202 851 3268 852
rect 3202 840 3209 851
rect 2861 810 3209 840
rect 2861 799 2868 810
rect 2802 798 2868 799
rect 3202 799 3209 810
rect 3261 840 3268 851
rect 3602 851 3668 852
rect 3602 840 3609 851
rect 3261 810 3609 840
rect 3261 799 3268 810
rect 3202 798 3268 799
rect 3602 799 3609 810
rect 3661 840 3668 851
rect 4002 851 4068 852
rect 4002 840 4009 851
rect 3661 810 4009 840
rect 3661 799 3668 810
rect 3602 798 3668 799
rect 4002 799 4009 810
rect 4061 840 4068 851
rect 4402 851 4468 852
rect 4402 840 4409 851
rect 4061 810 4409 840
rect 4061 799 4068 810
rect 4002 798 4068 799
rect 4402 799 4409 810
rect 4461 840 4468 851
rect 4802 851 4868 852
rect 4802 840 4809 851
rect 4461 810 4809 840
rect 4461 799 4468 810
rect 4402 798 4468 799
rect 4802 799 4809 810
rect 4861 840 4868 851
rect 5202 851 5268 852
rect 5202 840 5209 851
rect 4861 810 5209 840
rect 4861 799 4868 810
rect 4802 798 4868 799
rect 5202 799 5209 810
rect 5261 840 5268 851
rect 5602 851 5668 852
rect 5602 840 5609 851
rect 5261 810 5609 840
rect 5261 799 5268 810
rect 5202 798 5268 799
rect 5602 799 5609 810
rect 5661 840 5668 851
rect 6002 851 6068 852
rect 6002 840 6009 851
rect 5661 810 6009 840
rect 5661 799 5668 810
rect 5602 798 5668 799
rect 6002 799 6009 810
rect 6061 840 6068 851
rect 6402 851 6468 852
rect 6402 840 6409 851
rect 6061 810 6409 840
rect 6061 799 6068 810
rect 6002 798 6068 799
rect 6402 799 6409 810
rect 6461 840 6468 851
rect 6500 851 6566 852
rect 6500 840 6507 851
rect 6461 810 6507 840
rect 6461 799 6468 810
rect 6402 798 6468 799
rect 6500 799 6507 810
rect 6559 799 6566 851
rect 6500 798 6566 799
rect 202 781 268 782
rect 202 770 209 781
rect 0 740 209 770
rect 202 729 209 740
rect 261 770 268 781
rect 602 781 668 782
rect 602 770 609 781
rect 261 740 609 770
rect 261 729 268 740
rect 202 728 268 729
rect 602 729 609 740
rect 661 770 668 781
rect 1002 781 1068 782
rect 1002 770 1009 781
rect 661 740 1009 770
rect 661 729 668 740
rect 602 728 668 729
rect 1002 729 1009 740
rect 1061 770 1068 781
rect 1402 781 1468 782
rect 1402 770 1409 781
rect 1061 740 1409 770
rect 1061 729 1068 740
rect 1002 728 1068 729
rect 1402 729 1409 740
rect 1461 770 1468 781
rect 1802 781 1868 782
rect 1802 770 1809 781
rect 1461 740 1809 770
rect 1461 729 1468 740
rect 1402 728 1468 729
rect 1802 729 1809 740
rect 1861 770 1868 781
rect 2202 781 2268 782
rect 2202 770 2209 781
rect 1861 740 2209 770
rect 1861 729 1868 740
rect 1802 728 1868 729
rect 2202 729 2209 740
rect 2261 770 2268 781
rect 2602 781 2668 782
rect 2602 770 2609 781
rect 2261 740 2609 770
rect 2261 729 2268 740
rect 2202 728 2268 729
rect 2602 729 2609 740
rect 2661 770 2668 781
rect 3002 781 3068 782
rect 3002 770 3009 781
rect 2661 740 3009 770
rect 2661 729 2668 740
rect 2602 728 2668 729
rect 3002 729 3009 740
rect 3061 770 3068 781
rect 3402 781 3468 782
rect 3402 770 3409 781
rect 3061 740 3409 770
rect 3061 729 3068 740
rect 3002 728 3068 729
rect 3402 729 3409 740
rect 3461 770 3468 781
rect 3802 781 3868 782
rect 3802 770 3809 781
rect 3461 740 3809 770
rect 3461 729 3468 740
rect 3402 728 3468 729
rect 3802 729 3809 740
rect 3861 770 3868 781
rect 4202 781 4268 782
rect 4202 770 4209 781
rect 3861 740 4209 770
rect 3861 729 3868 740
rect 3802 728 3868 729
rect 4202 729 4209 740
rect 4261 770 4268 781
rect 4602 781 4668 782
rect 4602 770 4609 781
rect 4261 740 4609 770
rect 4261 729 4268 740
rect 4202 728 4268 729
rect 4602 729 4609 740
rect 4661 770 4668 781
rect 5002 781 5068 782
rect 5002 770 5009 781
rect 4661 740 5009 770
rect 4661 729 4668 740
rect 4602 728 4668 729
rect 5002 729 5009 740
rect 5061 770 5068 781
rect 5402 781 5468 782
rect 5402 770 5409 781
rect 5061 740 5409 770
rect 5061 729 5068 740
rect 5002 728 5068 729
rect 5402 729 5409 740
rect 5461 770 5468 781
rect 5802 781 5868 782
rect 5802 770 5809 781
rect 5461 740 5809 770
rect 5461 729 5468 740
rect 5402 728 5468 729
rect 5802 729 5809 740
rect 5861 770 5868 781
rect 6202 781 6268 782
rect 6202 770 6209 781
rect 5861 740 6209 770
rect 5861 729 5868 740
rect 5802 728 5868 729
rect 6202 729 6209 740
rect 6261 770 6268 781
rect 6704 781 6770 782
rect 6704 770 6711 781
rect 6261 740 6711 770
rect 6261 729 6268 740
rect 6202 728 6268 729
rect 6704 729 6711 740
rect 6763 729 6770 781
rect 6704 728 6770 729
rect 2 711 68 712
rect 2 700 9 711
rect 0 670 9 700
rect 2 659 9 670
rect 61 700 68 711
rect 402 711 468 712
rect 402 700 409 711
rect 61 670 409 700
rect 61 659 68 670
rect 2 658 68 659
rect 402 659 409 670
rect 461 700 468 711
rect 802 711 868 712
rect 802 700 809 711
rect 461 670 809 700
rect 461 659 468 670
rect 402 658 468 659
rect 802 659 809 670
rect 861 700 868 711
rect 1202 711 1268 712
rect 1202 700 1209 711
rect 861 670 1209 700
rect 861 659 868 670
rect 802 658 868 659
rect 1202 659 1209 670
rect 1261 700 1268 711
rect 1602 711 1668 712
rect 1602 700 1609 711
rect 1261 670 1609 700
rect 1261 659 1268 670
rect 1202 658 1268 659
rect 1602 659 1609 670
rect 1661 700 1668 711
rect 2002 711 2068 712
rect 2002 700 2009 711
rect 1661 670 2009 700
rect 1661 659 1668 670
rect 1602 658 1668 659
rect 2002 659 2009 670
rect 2061 700 2068 711
rect 2402 711 2468 712
rect 2402 700 2409 711
rect 2061 670 2409 700
rect 2061 659 2068 670
rect 2002 658 2068 659
rect 2402 659 2409 670
rect 2461 700 2468 711
rect 2802 711 2868 712
rect 2802 700 2809 711
rect 2461 670 2809 700
rect 2461 659 2468 670
rect 2402 658 2468 659
rect 2802 659 2809 670
rect 2861 700 2868 711
rect 3202 711 3268 712
rect 3202 700 3209 711
rect 2861 670 3209 700
rect 2861 659 2868 670
rect 2802 658 2868 659
rect 3202 659 3209 670
rect 3261 700 3268 711
rect 3602 711 3668 712
rect 3602 700 3609 711
rect 3261 670 3609 700
rect 3261 659 3268 670
rect 3202 658 3268 659
rect 3602 659 3609 670
rect 3661 700 3668 711
rect 4002 711 4068 712
rect 4002 700 4009 711
rect 3661 670 4009 700
rect 3661 659 3668 670
rect 3602 658 3668 659
rect 4002 659 4009 670
rect 4061 700 4068 711
rect 4402 711 4468 712
rect 4402 700 4409 711
rect 4061 670 4409 700
rect 4061 659 4068 670
rect 4002 658 4068 659
rect 4402 659 4409 670
rect 4461 700 4468 711
rect 4802 711 4868 712
rect 4802 700 4809 711
rect 4461 670 4809 700
rect 4461 659 4468 670
rect 4402 658 4468 659
rect 4802 659 4809 670
rect 4861 700 4868 711
rect 5202 711 5268 712
rect 5202 700 5209 711
rect 4861 670 5209 700
rect 4861 659 4868 670
rect 4802 658 4868 659
rect 5202 659 5209 670
rect 5261 700 5268 711
rect 5602 711 5668 712
rect 5602 700 5609 711
rect 5261 670 5609 700
rect 5261 659 5268 670
rect 5202 658 5268 659
rect 5602 659 5609 670
rect 5661 700 5668 711
rect 6002 711 6068 712
rect 6002 700 6009 711
rect 5661 670 6009 700
rect 5661 659 5668 670
rect 5602 658 5668 659
rect 6002 659 6009 670
rect 6061 700 6068 711
rect 6402 711 6468 712
rect 6402 700 6409 711
rect 6061 670 6409 700
rect 6061 659 6068 670
rect 6002 658 6068 659
rect 6402 659 6409 670
rect 6461 700 6468 711
rect 6500 711 6566 712
rect 6500 700 6507 711
rect 6461 670 6507 700
rect 6461 659 6468 670
rect 6402 658 6468 659
rect 6500 659 6507 670
rect 6559 659 6566 711
rect 6500 658 6566 659
rect 202 641 268 642
rect 202 630 209 641
rect 0 600 209 630
rect 202 589 209 600
rect 261 630 268 641
rect 602 641 668 642
rect 602 630 609 641
rect 261 600 609 630
rect 261 589 268 600
rect 202 588 268 589
rect 602 589 609 600
rect 661 630 668 641
rect 1002 641 1068 642
rect 1002 630 1009 641
rect 661 600 1009 630
rect 661 589 668 600
rect 602 588 668 589
rect 1002 589 1009 600
rect 1061 630 1068 641
rect 1402 641 1468 642
rect 1402 630 1409 641
rect 1061 600 1409 630
rect 1061 589 1068 600
rect 1002 588 1068 589
rect 1402 589 1409 600
rect 1461 630 1468 641
rect 1802 641 1868 642
rect 1802 630 1809 641
rect 1461 600 1809 630
rect 1461 589 1468 600
rect 1402 588 1468 589
rect 1802 589 1809 600
rect 1861 630 1868 641
rect 2202 641 2268 642
rect 2202 630 2209 641
rect 1861 600 2209 630
rect 1861 589 1868 600
rect 1802 588 1868 589
rect 2202 589 2209 600
rect 2261 630 2268 641
rect 2602 641 2668 642
rect 2602 630 2609 641
rect 2261 600 2609 630
rect 2261 589 2268 600
rect 2202 588 2268 589
rect 2602 589 2609 600
rect 2661 630 2668 641
rect 3002 641 3068 642
rect 3002 630 3009 641
rect 2661 600 3009 630
rect 2661 589 2668 600
rect 2602 588 2668 589
rect 3002 589 3009 600
rect 3061 630 3068 641
rect 3402 641 3468 642
rect 3402 630 3409 641
rect 3061 600 3409 630
rect 3061 589 3068 600
rect 3002 588 3068 589
rect 3402 589 3409 600
rect 3461 630 3468 641
rect 3802 641 3868 642
rect 3802 630 3809 641
rect 3461 600 3809 630
rect 3461 589 3468 600
rect 3402 588 3468 589
rect 3802 589 3809 600
rect 3861 630 3868 641
rect 4202 641 4268 642
rect 4202 630 4209 641
rect 3861 600 4209 630
rect 3861 589 3868 600
rect 3802 588 3868 589
rect 4202 589 4209 600
rect 4261 630 4268 641
rect 4602 641 4668 642
rect 4602 630 4609 641
rect 4261 600 4609 630
rect 4261 589 4268 600
rect 4202 588 4268 589
rect 4602 589 4609 600
rect 4661 630 4668 641
rect 5002 641 5068 642
rect 5002 630 5009 641
rect 4661 600 5009 630
rect 4661 589 4668 600
rect 4602 588 4668 589
rect 5002 589 5009 600
rect 5061 630 5068 641
rect 5402 641 5468 642
rect 5402 630 5409 641
rect 5061 600 5409 630
rect 5061 589 5068 600
rect 5002 588 5068 589
rect 5402 589 5409 600
rect 5461 630 5468 641
rect 5802 641 5868 642
rect 5802 630 5809 641
rect 5461 600 5809 630
rect 5461 589 5468 600
rect 5402 588 5468 589
rect 5802 589 5809 600
rect 5861 630 5868 641
rect 6202 641 6268 642
rect 6202 630 6209 641
rect 5861 600 6209 630
rect 5861 589 5868 600
rect 5802 588 5868 589
rect 6202 589 6209 600
rect 6261 630 6268 641
rect 6704 641 6770 642
rect 6704 630 6711 641
rect 6261 600 6711 630
rect 6261 589 6268 600
rect 6202 588 6268 589
rect 6704 589 6711 600
rect 6763 589 6770 641
rect 6704 588 6770 589
rect 2 571 68 572
rect 2 560 9 571
rect 0 530 9 560
rect 2 519 9 530
rect 61 560 68 571
rect 402 571 468 572
rect 402 560 409 571
rect 61 530 409 560
rect 61 519 68 530
rect 2 518 68 519
rect 402 519 409 530
rect 461 560 468 571
rect 802 571 868 572
rect 802 560 809 571
rect 461 530 809 560
rect 461 519 468 530
rect 402 518 468 519
rect 802 519 809 530
rect 861 560 868 571
rect 1202 571 1268 572
rect 1202 560 1209 571
rect 861 530 1209 560
rect 861 519 868 530
rect 802 518 868 519
rect 1202 519 1209 530
rect 1261 560 1268 571
rect 1602 571 1668 572
rect 1602 560 1609 571
rect 1261 530 1609 560
rect 1261 519 1268 530
rect 1202 518 1268 519
rect 1602 519 1609 530
rect 1661 560 1668 571
rect 2002 571 2068 572
rect 2002 560 2009 571
rect 1661 530 2009 560
rect 1661 519 1668 530
rect 1602 518 1668 519
rect 2002 519 2009 530
rect 2061 560 2068 571
rect 2402 571 2468 572
rect 2402 560 2409 571
rect 2061 530 2409 560
rect 2061 519 2068 530
rect 2002 518 2068 519
rect 2402 519 2409 530
rect 2461 560 2468 571
rect 2802 571 2868 572
rect 2802 560 2809 571
rect 2461 530 2809 560
rect 2461 519 2468 530
rect 2402 518 2468 519
rect 2802 519 2809 530
rect 2861 560 2868 571
rect 3202 571 3268 572
rect 3202 560 3209 571
rect 2861 530 3209 560
rect 2861 519 2868 530
rect 2802 518 2868 519
rect 3202 519 3209 530
rect 3261 560 3268 571
rect 3602 571 3668 572
rect 3602 560 3609 571
rect 3261 530 3609 560
rect 3261 519 3268 530
rect 3202 518 3268 519
rect 3602 519 3609 530
rect 3661 560 3668 571
rect 4002 571 4068 572
rect 4002 560 4009 571
rect 3661 530 4009 560
rect 3661 519 3668 530
rect 3602 518 3668 519
rect 4002 519 4009 530
rect 4061 560 4068 571
rect 4402 571 4468 572
rect 4402 560 4409 571
rect 4061 530 4409 560
rect 4061 519 4068 530
rect 4002 518 4068 519
rect 4402 519 4409 530
rect 4461 560 4468 571
rect 4802 571 4868 572
rect 4802 560 4809 571
rect 4461 530 4809 560
rect 4461 519 4468 530
rect 4402 518 4468 519
rect 4802 519 4809 530
rect 4861 560 4868 571
rect 5202 571 5268 572
rect 5202 560 5209 571
rect 4861 530 5209 560
rect 4861 519 4868 530
rect 4802 518 4868 519
rect 5202 519 5209 530
rect 5261 560 5268 571
rect 5602 571 5668 572
rect 5602 560 5609 571
rect 5261 530 5609 560
rect 5261 519 5268 530
rect 5202 518 5268 519
rect 5602 519 5609 530
rect 5661 560 5668 571
rect 6002 571 6068 572
rect 6002 560 6009 571
rect 5661 530 6009 560
rect 5661 519 5668 530
rect 5602 518 5668 519
rect 6002 519 6009 530
rect 6061 560 6068 571
rect 6402 571 6468 572
rect 6402 560 6409 571
rect 6061 530 6409 560
rect 6061 519 6068 530
rect 6002 518 6068 519
rect 6402 519 6409 530
rect 6461 560 6468 571
rect 6500 571 6566 572
rect 6500 560 6507 571
rect 6461 530 6507 560
rect 6461 519 6468 530
rect 6402 518 6468 519
rect 6500 519 6507 530
rect 6559 519 6566 571
rect 6500 518 6566 519
rect 202 501 268 502
rect 202 490 209 501
rect 0 460 209 490
rect 202 449 209 460
rect 261 490 268 501
rect 602 501 668 502
rect 602 490 609 501
rect 261 460 609 490
rect 261 449 268 460
rect 202 448 268 449
rect 602 449 609 460
rect 661 490 668 501
rect 1002 501 1068 502
rect 1002 490 1009 501
rect 661 460 1009 490
rect 661 449 668 460
rect 602 448 668 449
rect 1002 449 1009 460
rect 1061 490 1068 501
rect 1402 501 1468 502
rect 1402 490 1409 501
rect 1061 460 1409 490
rect 1061 449 1068 460
rect 1002 448 1068 449
rect 1402 449 1409 460
rect 1461 490 1468 501
rect 1802 501 1868 502
rect 1802 490 1809 501
rect 1461 460 1809 490
rect 1461 449 1468 460
rect 1402 448 1468 449
rect 1802 449 1809 460
rect 1861 490 1868 501
rect 2202 501 2268 502
rect 2202 490 2209 501
rect 1861 460 2209 490
rect 1861 449 1868 460
rect 1802 448 1868 449
rect 2202 449 2209 460
rect 2261 490 2268 501
rect 2602 501 2668 502
rect 2602 490 2609 501
rect 2261 460 2609 490
rect 2261 449 2268 460
rect 2202 448 2268 449
rect 2602 449 2609 460
rect 2661 490 2668 501
rect 3002 501 3068 502
rect 3002 490 3009 501
rect 2661 460 3009 490
rect 2661 449 2668 460
rect 2602 448 2668 449
rect 3002 449 3009 460
rect 3061 490 3068 501
rect 3402 501 3468 502
rect 3402 490 3409 501
rect 3061 460 3409 490
rect 3061 449 3068 460
rect 3002 448 3068 449
rect 3402 449 3409 460
rect 3461 490 3468 501
rect 3802 501 3868 502
rect 3802 490 3809 501
rect 3461 460 3809 490
rect 3461 449 3468 460
rect 3402 448 3468 449
rect 3802 449 3809 460
rect 3861 490 3868 501
rect 4202 501 4268 502
rect 4202 490 4209 501
rect 3861 460 4209 490
rect 3861 449 3868 460
rect 3802 448 3868 449
rect 4202 449 4209 460
rect 4261 490 4268 501
rect 4602 501 4668 502
rect 4602 490 4609 501
rect 4261 460 4609 490
rect 4261 449 4268 460
rect 4202 448 4268 449
rect 4602 449 4609 460
rect 4661 490 4668 501
rect 5002 501 5068 502
rect 5002 490 5009 501
rect 4661 460 5009 490
rect 4661 449 4668 460
rect 4602 448 4668 449
rect 5002 449 5009 460
rect 5061 490 5068 501
rect 5402 501 5468 502
rect 5402 490 5409 501
rect 5061 460 5409 490
rect 5061 449 5068 460
rect 5002 448 5068 449
rect 5402 449 5409 460
rect 5461 490 5468 501
rect 5802 501 5868 502
rect 5802 490 5809 501
rect 5461 460 5809 490
rect 5461 449 5468 460
rect 5402 448 5468 449
rect 5802 449 5809 460
rect 5861 490 5868 501
rect 6202 501 6268 502
rect 6202 490 6209 501
rect 5861 460 6209 490
rect 5861 449 5868 460
rect 5802 448 5868 449
rect 6202 449 6209 460
rect 6261 490 6268 501
rect 6704 501 6770 502
rect 6704 490 6711 501
rect 6261 460 6711 490
rect 6261 449 6268 460
rect 6202 448 6268 449
rect 6704 449 6711 460
rect 6763 449 6770 501
rect 6704 448 6770 449
rect 2 431 68 432
rect 2 420 9 431
rect 0 390 9 420
rect 2 379 9 390
rect 61 420 68 431
rect 402 431 468 432
rect 402 420 409 431
rect 61 390 409 420
rect 61 379 68 390
rect 2 378 68 379
rect 402 379 409 390
rect 461 420 468 431
rect 802 431 868 432
rect 802 420 809 431
rect 461 390 809 420
rect 461 379 468 390
rect 402 378 468 379
rect 802 379 809 390
rect 861 420 868 431
rect 1202 431 1268 432
rect 1202 420 1209 431
rect 861 390 1209 420
rect 861 379 868 390
rect 802 378 868 379
rect 1202 379 1209 390
rect 1261 420 1268 431
rect 1602 431 1668 432
rect 1602 420 1609 431
rect 1261 390 1609 420
rect 1261 379 1268 390
rect 1202 378 1268 379
rect 1602 379 1609 390
rect 1661 420 1668 431
rect 2002 431 2068 432
rect 2002 420 2009 431
rect 1661 390 2009 420
rect 1661 379 1668 390
rect 1602 378 1668 379
rect 2002 379 2009 390
rect 2061 420 2068 431
rect 2402 431 2468 432
rect 2402 420 2409 431
rect 2061 390 2409 420
rect 2061 379 2068 390
rect 2002 378 2068 379
rect 2402 379 2409 390
rect 2461 420 2468 431
rect 2802 431 2868 432
rect 2802 420 2809 431
rect 2461 390 2809 420
rect 2461 379 2468 390
rect 2402 378 2468 379
rect 2802 379 2809 390
rect 2861 420 2868 431
rect 3202 431 3268 432
rect 3202 420 3209 431
rect 2861 390 3209 420
rect 2861 379 2868 390
rect 2802 378 2868 379
rect 3202 379 3209 390
rect 3261 420 3268 431
rect 3602 431 3668 432
rect 3602 420 3609 431
rect 3261 390 3609 420
rect 3261 379 3268 390
rect 3202 378 3268 379
rect 3602 379 3609 390
rect 3661 420 3668 431
rect 4002 431 4068 432
rect 4002 420 4009 431
rect 3661 390 4009 420
rect 3661 379 3668 390
rect 3602 378 3668 379
rect 4002 379 4009 390
rect 4061 420 4068 431
rect 4402 431 4468 432
rect 4402 420 4409 431
rect 4061 390 4409 420
rect 4061 379 4068 390
rect 4002 378 4068 379
rect 4402 379 4409 390
rect 4461 420 4468 431
rect 4802 431 4868 432
rect 4802 420 4809 431
rect 4461 390 4809 420
rect 4461 379 4468 390
rect 4402 378 4468 379
rect 4802 379 4809 390
rect 4861 420 4868 431
rect 5202 431 5268 432
rect 5202 420 5209 431
rect 4861 390 5209 420
rect 4861 379 4868 390
rect 4802 378 4868 379
rect 5202 379 5209 390
rect 5261 420 5268 431
rect 5602 431 5668 432
rect 5602 420 5609 431
rect 5261 390 5609 420
rect 5261 379 5268 390
rect 5202 378 5268 379
rect 5602 379 5609 390
rect 5661 420 5668 431
rect 6002 431 6068 432
rect 6002 420 6009 431
rect 5661 390 6009 420
rect 5661 379 5668 390
rect 5602 378 5668 379
rect 6002 379 6009 390
rect 6061 420 6068 431
rect 6402 431 6468 432
rect 6402 420 6409 431
rect 6061 390 6409 420
rect 6061 379 6068 390
rect 6002 378 6068 379
rect 6402 379 6409 390
rect 6461 420 6468 431
rect 6500 431 6566 432
rect 6500 420 6507 431
rect 6461 390 6507 420
rect 6461 379 6468 390
rect 6402 378 6468 379
rect 6500 379 6507 390
rect 6559 379 6566 431
rect 6500 378 6566 379
rect 202 361 268 362
rect 202 350 209 361
rect 0 320 209 350
rect 202 309 209 320
rect 261 350 268 361
rect 602 361 668 362
rect 602 350 609 361
rect 261 320 609 350
rect 261 309 268 320
rect 202 308 268 309
rect 602 309 609 320
rect 661 350 668 361
rect 1002 361 1068 362
rect 1002 350 1009 361
rect 661 320 1009 350
rect 661 309 668 320
rect 602 308 668 309
rect 1002 309 1009 320
rect 1061 350 1068 361
rect 1402 361 1468 362
rect 1402 350 1409 361
rect 1061 320 1409 350
rect 1061 309 1068 320
rect 1002 308 1068 309
rect 1402 309 1409 320
rect 1461 350 1468 361
rect 1802 361 1868 362
rect 1802 350 1809 361
rect 1461 320 1809 350
rect 1461 309 1468 320
rect 1402 308 1468 309
rect 1802 309 1809 320
rect 1861 350 1868 361
rect 2202 361 2268 362
rect 2202 350 2209 361
rect 1861 320 2209 350
rect 1861 309 1868 320
rect 1802 308 1868 309
rect 2202 309 2209 320
rect 2261 350 2268 361
rect 2602 361 2668 362
rect 2602 350 2609 361
rect 2261 320 2609 350
rect 2261 309 2268 320
rect 2202 308 2268 309
rect 2602 309 2609 320
rect 2661 350 2668 361
rect 3002 361 3068 362
rect 3002 350 3009 361
rect 2661 320 3009 350
rect 2661 309 2668 320
rect 2602 308 2668 309
rect 3002 309 3009 320
rect 3061 350 3068 361
rect 3402 361 3468 362
rect 3402 350 3409 361
rect 3061 320 3409 350
rect 3061 309 3068 320
rect 3002 308 3068 309
rect 3402 309 3409 320
rect 3461 350 3468 361
rect 3802 361 3868 362
rect 3802 350 3809 361
rect 3461 320 3809 350
rect 3461 309 3468 320
rect 3402 308 3468 309
rect 3802 309 3809 320
rect 3861 350 3868 361
rect 4202 361 4268 362
rect 4202 350 4209 361
rect 3861 320 4209 350
rect 3861 309 3868 320
rect 3802 308 3868 309
rect 4202 309 4209 320
rect 4261 350 4268 361
rect 4602 361 4668 362
rect 4602 350 4609 361
rect 4261 320 4609 350
rect 4261 309 4268 320
rect 4202 308 4268 309
rect 4602 309 4609 320
rect 4661 350 4668 361
rect 5002 361 5068 362
rect 5002 350 5009 361
rect 4661 320 5009 350
rect 4661 309 4668 320
rect 4602 308 4668 309
rect 5002 309 5009 320
rect 5061 350 5068 361
rect 5402 361 5468 362
rect 5402 350 5409 361
rect 5061 320 5409 350
rect 5061 309 5068 320
rect 5002 308 5068 309
rect 5402 309 5409 320
rect 5461 350 5468 361
rect 5802 361 5868 362
rect 5802 350 5809 361
rect 5461 320 5809 350
rect 5461 309 5468 320
rect 5402 308 5468 309
rect 5802 309 5809 320
rect 5861 350 5868 361
rect 6202 361 6268 362
rect 6202 350 6209 361
rect 5861 320 6209 350
rect 5861 309 5868 320
rect 5802 308 5868 309
rect 6202 309 6209 320
rect 6261 350 6268 361
rect 6704 361 6770 362
rect 6704 350 6711 361
rect 6261 320 6711 350
rect 6261 309 6268 320
rect 6202 308 6268 309
rect 6704 309 6711 320
rect 6763 309 6770 361
rect 6704 308 6770 309
rect 2 291 68 292
rect 2 280 9 291
rect 0 250 9 280
rect 2 239 9 250
rect 61 280 68 291
rect 402 291 468 292
rect 402 280 409 291
rect 61 250 409 280
rect 61 239 68 250
rect 2 238 68 239
rect 402 239 409 250
rect 461 280 468 291
rect 802 291 868 292
rect 802 280 809 291
rect 461 250 809 280
rect 461 239 468 250
rect 402 238 468 239
rect 802 239 809 250
rect 861 280 868 291
rect 1202 291 1268 292
rect 1202 280 1209 291
rect 861 250 1209 280
rect 861 239 868 250
rect 802 238 868 239
rect 1202 239 1209 250
rect 1261 280 1268 291
rect 1602 291 1668 292
rect 1602 280 1609 291
rect 1261 250 1609 280
rect 1261 239 1268 250
rect 1202 238 1268 239
rect 1602 239 1609 250
rect 1661 280 1668 291
rect 2002 291 2068 292
rect 2002 280 2009 291
rect 1661 250 2009 280
rect 1661 239 1668 250
rect 1602 238 1668 239
rect 2002 239 2009 250
rect 2061 280 2068 291
rect 2402 291 2468 292
rect 2402 280 2409 291
rect 2061 250 2409 280
rect 2061 239 2068 250
rect 2002 238 2068 239
rect 2402 239 2409 250
rect 2461 280 2468 291
rect 2802 291 2868 292
rect 2802 280 2809 291
rect 2461 250 2809 280
rect 2461 239 2468 250
rect 2402 238 2468 239
rect 2802 239 2809 250
rect 2861 280 2868 291
rect 3202 291 3268 292
rect 3202 280 3209 291
rect 2861 250 3209 280
rect 2861 239 2868 250
rect 2802 238 2868 239
rect 3202 239 3209 250
rect 3261 280 3268 291
rect 3602 291 3668 292
rect 3602 280 3609 291
rect 3261 250 3609 280
rect 3261 239 3268 250
rect 3202 238 3268 239
rect 3602 239 3609 250
rect 3661 280 3668 291
rect 4002 291 4068 292
rect 4002 280 4009 291
rect 3661 250 4009 280
rect 3661 239 3668 250
rect 3602 238 3668 239
rect 4002 239 4009 250
rect 4061 280 4068 291
rect 4402 291 4468 292
rect 4402 280 4409 291
rect 4061 250 4409 280
rect 4061 239 4068 250
rect 4002 238 4068 239
rect 4402 239 4409 250
rect 4461 280 4468 291
rect 4802 291 4868 292
rect 4802 280 4809 291
rect 4461 250 4809 280
rect 4461 239 4468 250
rect 4402 238 4468 239
rect 4802 239 4809 250
rect 4861 280 4868 291
rect 5202 291 5268 292
rect 5202 280 5209 291
rect 4861 250 5209 280
rect 4861 239 4868 250
rect 4802 238 4868 239
rect 5202 239 5209 250
rect 5261 280 5268 291
rect 5602 291 5668 292
rect 5602 280 5609 291
rect 5261 250 5609 280
rect 5261 239 5268 250
rect 5202 238 5268 239
rect 5602 239 5609 250
rect 5661 280 5668 291
rect 6002 291 6068 292
rect 6002 280 6009 291
rect 5661 250 6009 280
rect 5661 239 5668 250
rect 5602 238 5668 239
rect 6002 239 6009 250
rect 6061 280 6068 291
rect 6402 291 6468 292
rect 6402 280 6409 291
rect 6061 250 6409 280
rect 6061 239 6068 250
rect 6002 238 6068 239
rect 6402 239 6409 250
rect 6461 280 6468 291
rect 6500 291 6566 292
rect 6500 280 6507 291
rect 6461 250 6507 280
rect 6461 239 6468 250
rect 6402 238 6468 239
rect 6500 239 6507 250
rect 6559 239 6566 291
rect 6500 238 6566 239
rect 202 221 268 222
rect 202 210 209 221
rect 0 180 209 210
rect 202 169 209 180
rect 261 210 268 221
rect 602 221 668 222
rect 602 210 609 221
rect 261 180 609 210
rect 261 169 268 180
rect 202 168 268 169
rect 602 169 609 180
rect 661 210 668 221
rect 1002 221 1068 222
rect 1002 210 1009 221
rect 661 180 1009 210
rect 661 169 668 180
rect 602 168 668 169
rect 1002 169 1009 180
rect 1061 210 1068 221
rect 1402 221 1468 222
rect 1402 210 1409 221
rect 1061 180 1409 210
rect 1061 169 1068 180
rect 1002 168 1068 169
rect 1402 169 1409 180
rect 1461 210 1468 221
rect 1802 221 1868 222
rect 1802 210 1809 221
rect 1461 180 1809 210
rect 1461 169 1468 180
rect 1402 168 1468 169
rect 1802 169 1809 180
rect 1861 210 1868 221
rect 2202 221 2268 222
rect 2202 210 2209 221
rect 1861 180 2209 210
rect 1861 169 1868 180
rect 1802 168 1868 169
rect 2202 169 2209 180
rect 2261 210 2268 221
rect 2602 221 2668 222
rect 2602 210 2609 221
rect 2261 180 2609 210
rect 2261 169 2268 180
rect 2202 168 2268 169
rect 2602 169 2609 180
rect 2661 210 2668 221
rect 3002 221 3068 222
rect 3002 210 3009 221
rect 2661 180 3009 210
rect 2661 169 2668 180
rect 2602 168 2668 169
rect 3002 169 3009 180
rect 3061 210 3068 221
rect 3402 221 3468 222
rect 3402 210 3409 221
rect 3061 180 3409 210
rect 3061 169 3068 180
rect 3002 168 3068 169
rect 3402 169 3409 180
rect 3461 210 3468 221
rect 3802 221 3868 222
rect 3802 210 3809 221
rect 3461 180 3809 210
rect 3461 169 3468 180
rect 3402 168 3468 169
rect 3802 169 3809 180
rect 3861 210 3868 221
rect 4202 221 4268 222
rect 4202 210 4209 221
rect 3861 180 4209 210
rect 3861 169 3868 180
rect 3802 168 3868 169
rect 4202 169 4209 180
rect 4261 210 4268 221
rect 4602 221 4668 222
rect 4602 210 4609 221
rect 4261 180 4609 210
rect 4261 169 4268 180
rect 4202 168 4268 169
rect 4602 169 4609 180
rect 4661 210 4668 221
rect 5002 221 5068 222
rect 5002 210 5009 221
rect 4661 180 5009 210
rect 4661 169 4668 180
rect 4602 168 4668 169
rect 5002 169 5009 180
rect 5061 210 5068 221
rect 5402 221 5468 222
rect 5402 210 5409 221
rect 5061 180 5409 210
rect 5061 169 5068 180
rect 5002 168 5068 169
rect 5402 169 5409 180
rect 5461 210 5468 221
rect 5802 221 5868 222
rect 5802 210 5809 221
rect 5461 180 5809 210
rect 5461 169 5468 180
rect 5402 168 5468 169
rect 5802 169 5809 180
rect 5861 210 5868 221
rect 6202 221 6268 222
rect 6202 210 6209 221
rect 5861 180 6209 210
rect 5861 169 5868 180
rect 5802 168 5868 169
rect 6202 169 6209 180
rect 6261 210 6268 221
rect 6704 221 6770 222
rect 6704 210 6711 221
rect 6261 180 6711 210
rect 6261 169 6268 180
rect 6202 168 6268 169
rect 6704 169 6711 180
rect 6763 169 6770 221
rect 6704 168 6770 169
rect 2 151 68 152
rect 2 140 9 151
rect 0 110 9 140
rect 2 99 9 110
rect 61 140 68 151
rect 402 151 468 152
rect 402 140 409 151
rect 61 110 409 140
rect 61 99 68 110
rect 2 98 68 99
rect 402 99 409 110
rect 461 140 468 151
rect 802 151 868 152
rect 802 140 809 151
rect 461 110 809 140
rect 461 99 468 110
rect 402 98 468 99
rect 802 99 809 110
rect 861 140 868 151
rect 1202 151 1268 152
rect 1202 140 1209 151
rect 861 110 1209 140
rect 861 99 868 110
rect 802 98 868 99
rect 1202 99 1209 110
rect 1261 140 1268 151
rect 1602 151 1668 152
rect 1602 140 1609 151
rect 1261 110 1609 140
rect 1261 99 1268 110
rect 1202 98 1268 99
rect 1602 99 1609 110
rect 1661 140 1668 151
rect 2002 151 2068 152
rect 2002 140 2009 151
rect 1661 110 2009 140
rect 1661 99 1668 110
rect 1602 98 1668 99
rect 2002 99 2009 110
rect 2061 140 2068 151
rect 2402 151 2468 152
rect 2402 140 2409 151
rect 2061 110 2409 140
rect 2061 99 2068 110
rect 2002 98 2068 99
rect 2402 99 2409 110
rect 2461 140 2468 151
rect 2802 151 2868 152
rect 2802 140 2809 151
rect 2461 110 2809 140
rect 2461 99 2468 110
rect 2402 98 2468 99
rect 2802 99 2809 110
rect 2861 140 2868 151
rect 3202 151 3268 152
rect 3202 140 3209 151
rect 2861 110 3209 140
rect 2861 99 2868 110
rect 2802 98 2868 99
rect 3202 99 3209 110
rect 3261 140 3268 151
rect 3602 151 3668 152
rect 3602 140 3609 151
rect 3261 110 3609 140
rect 3261 99 3268 110
rect 3202 98 3268 99
rect 3602 99 3609 110
rect 3661 140 3668 151
rect 4002 151 4068 152
rect 4002 140 4009 151
rect 3661 110 4009 140
rect 3661 99 3668 110
rect 3602 98 3668 99
rect 4002 99 4009 110
rect 4061 140 4068 151
rect 4402 151 4468 152
rect 4402 140 4409 151
rect 4061 110 4409 140
rect 4061 99 4068 110
rect 4002 98 4068 99
rect 4402 99 4409 110
rect 4461 140 4468 151
rect 4802 151 4868 152
rect 4802 140 4809 151
rect 4461 110 4809 140
rect 4461 99 4468 110
rect 4402 98 4468 99
rect 4802 99 4809 110
rect 4861 140 4868 151
rect 5202 151 5268 152
rect 5202 140 5209 151
rect 4861 110 5209 140
rect 4861 99 4868 110
rect 4802 98 4868 99
rect 5202 99 5209 110
rect 5261 140 5268 151
rect 5602 151 5668 152
rect 5602 140 5609 151
rect 5261 110 5609 140
rect 5261 99 5268 110
rect 5202 98 5268 99
rect 5602 99 5609 110
rect 5661 140 5668 151
rect 6002 151 6068 152
rect 6002 140 6009 151
rect 5661 110 6009 140
rect 5661 99 5668 110
rect 5602 98 5668 99
rect 6002 99 6009 110
rect 6061 140 6068 151
rect 6402 151 6468 152
rect 6402 140 6409 151
rect 6061 110 6409 140
rect 6061 99 6068 110
rect 6002 98 6068 99
rect 6402 99 6409 110
rect 6461 140 6468 151
rect 6500 151 6566 152
rect 6500 140 6507 151
rect 6461 110 6507 140
rect 6461 99 6468 110
rect 6402 98 6468 99
rect 6500 99 6507 110
rect 6559 99 6566 151
rect 6500 98 6566 99
rect 196 81 274 82
rect -4 65 74 66
rect -4 9 7 65
rect 63 9 74 65
rect 196 25 207 81
rect 263 25 274 81
rect 596 81 674 82
rect 196 24 274 25
rect 396 65 474 66
rect -4 8 74 9
rect -93 -15 -37 0
rect -93 -67 -91 -15
rect -39 -67 -37 -15
rect -93 -79 -37 -67
rect -93 -110 -91 -79
rect -138 -131 -91 -110
rect -39 -110 -37 -79
rect 7 -16 63 8
rect 7 -74 9 -72
rect 61 -74 63 -72
rect 7 -81 63 -74
rect 107 -15 163 0
rect 107 -67 109 -15
rect 161 -67 163 -15
rect 107 -79 163 -67
rect 107 -110 109 -79
rect -39 -131 109 -110
rect 161 -110 163 -79
rect 207 -16 263 24
rect 396 9 407 65
rect 463 9 474 65
rect 596 25 607 81
rect 663 25 674 81
rect 996 81 1074 82
rect 596 24 674 25
rect 796 65 874 66
rect 396 8 474 9
rect 207 -74 209 -72
rect 261 -74 263 -72
rect 207 -81 263 -74
rect 307 -15 363 0
rect 307 -67 309 -15
rect 361 -67 363 -15
rect 307 -79 363 -67
rect 307 -110 309 -79
rect 161 -131 309 -110
rect 361 -110 363 -79
rect 407 -16 463 8
rect 407 -74 409 -72
rect 461 -74 463 -72
rect 407 -81 463 -74
rect 507 -15 563 0
rect 507 -67 509 -15
rect 561 -67 563 -15
rect 507 -79 563 -67
rect 507 -110 509 -79
rect 361 -131 509 -110
rect 561 -110 563 -79
rect 607 -16 663 24
rect 796 9 807 65
rect 863 9 874 65
rect 996 25 1007 81
rect 1063 25 1074 81
rect 1396 81 1474 82
rect 996 24 1074 25
rect 1196 65 1274 66
rect 796 8 874 9
rect 607 -74 609 -72
rect 661 -74 663 -72
rect 607 -81 663 -74
rect 707 -15 763 0
rect 707 -67 709 -15
rect 761 -67 763 -15
rect 707 -79 763 -67
rect 707 -110 709 -79
rect 561 -131 709 -110
rect 761 -110 763 -79
rect 807 -16 863 8
rect 807 -74 809 -72
rect 861 -74 863 -72
rect 807 -81 863 -74
rect 907 -15 963 0
rect 907 -67 909 -15
rect 961 -67 963 -15
rect 907 -79 963 -67
rect 907 -110 909 -79
rect 761 -131 909 -110
rect 961 -110 963 -79
rect 1007 -16 1063 24
rect 1196 9 1207 65
rect 1263 9 1274 65
rect 1396 25 1407 81
rect 1463 25 1474 81
rect 1796 81 1874 82
rect 1396 24 1474 25
rect 1596 65 1674 66
rect 1196 8 1274 9
rect 1007 -74 1009 -72
rect 1061 -74 1063 -72
rect 1007 -81 1063 -74
rect 1107 -15 1163 0
rect 1107 -67 1109 -15
rect 1161 -67 1163 -15
rect 1107 -79 1163 -67
rect 1107 -110 1109 -79
rect 961 -131 1109 -110
rect 1161 -110 1163 -79
rect 1207 -16 1263 8
rect 1207 -74 1209 -72
rect 1261 -74 1263 -72
rect 1207 -81 1263 -74
rect 1307 -15 1363 0
rect 1307 -67 1309 -15
rect 1361 -67 1363 -15
rect 1307 -79 1363 -67
rect 1307 -110 1309 -79
rect 1161 -131 1309 -110
rect 1361 -110 1363 -79
rect 1407 -16 1463 24
rect 1596 9 1607 65
rect 1663 9 1674 65
rect 1796 25 1807 81
rect 1863 25 1874 81
rect 2196 81 2274 82
rect 1796 24 1874 25
rect 1996 65 2074 66
rect 1596 8 1674 9
rect 1407 -74 1409 -72
rect 1461 -74 1463 -72
rect 1407 -81 1463 -74
rect 1507 -15 1563 0
rect 1507 -67 1509 -15
rect 1561 -67 1563 -15
rect 1507 -79 1563 -67
rect 1507 -110 1509 -79
rect 1361 -131 1509 -110
rect 1561 -110 1563 -79
rect 1607 -16 1663 8
rect 1607 -74 1609 -72
rect 1661 -74 1663 -72
rect 1607 -81 1663 -74
rect 1707 -15 1763 0
rect 1707 -67 1709 -15
rect 1761 -67 1763 -15
rect 1707 -79 1763 -67
rect 1707 -110 1709 -79
rect 1561 -131 1709 -110
rect 1761 -110 1763 -79
rect 1807 -16 1863 24
rect 1996 9 2007 65
rect 2063 9 2074 65
rect 2196 25 2207 81
rect 2263 25 2274 81
rect 2596 81 2674 82
rect 2196 24 2274 25
rect 2396 65 2474 66
rect 1996 8 2074 9
rect 1807 -74 1809 -72
rect 1861 -74 1863 -72
rect 1807 -81 1863 -74
rect 1907 -15 1963 0
rect 1907 -67 1909 -15
rect 1961 -67 1963 -15
rect 1907 -79 1963 -67
rect 1907 -110 1909 -79
rect 1761 -131 1909 -110
rect 1961 -110 1963 -79
rect 2007 -16 2063 8
rect 2007 -74 2009 -72
rect 2061 -74 2063 -72
rect 2007 -81 2063 -74
rect 2107 -15 2163 0
rect 2107 -67 2109 -15
rect 2161 -67 2163 -15
rect 2107 -79 2163 -67
rect 2107 -110 2109 -79
rect 1961 -131 2109 -110
rect 2161 -110 2163 -79
rect 2207 -16 2263 24
rect 2396 9 2407 65
rect 2463 9 2474 65
rect 2596 25 2607 81
rect 2663 25 2674 81
rect 2996 81 3074 82
rect 2596 24 2674 25
rect 2796 65 2874 66
rect 2396 8 2474 9
rect 2207 -74 2209 -72
rect 2261 -74 2263 -72
rect 2207 -81 2263 -74
rect 2307 -15 2363 0
rect 2307 -67 2309 -15
rect 2361 -67 2363 -15
rect 2307 -79 2363 -67
rect 2307 -110 2309 -79
rect 2161 -131 2309 -110
rect 2361 -110 2363 -79
rect 2407 -16 2463 8
rect 2407 -74 2409 -72
rect 2461 -74 2463 -72
rect 2407 -81 2463 -74
rect 2507 -15 2563 0
rect 2507 -67 2509 -15
rect 2561 -67 2563 -15
rect 2507 -79 2563 -67
rect 2507 -110 2509 -79
rect 2361 -131 2509 -110
rect 2561 -110 2563 -79
rect 2607 -16 2663 24
rect 2796 9 2807 65
rect 2863 9 2874 65
rect 2996 25 3007 81
rect 3063 25 3074 81
rect 3396 81 3474 82
rect 2996 24 3074 25
rect 3196 65 3274 66
rect 2796 8 2874 9
rect 2607 -74 2609 -72
rect 2661 -74 2663 -72
rect 2607 -81 2663 -74
rect 2707 -15 2763 0
rect 2707 -67 2709 -15
rect 2761 -67 2763 -15
rect 2707 -79 2763 -67
rect 2707 -110 2709 -79
rect 2561 -131 2709 -110
rect 2761 -110 2763 -79
rect 2807 -16 2863 8
rect 2807 -74 2809 -72
rect 2861 -74 2863 -72
rect 2807 -81 2863 -74
rect 2907 -15 2963 0
rect 2907 -67 2909 -15
rect 2961 -67 2963 -15
rect 2907 -79 2963 -67
rect 2907 -110 2909 -79
rect 2761 -131 2909 -110
rect 2961 -110 2963 -79
rect 3007 -16 3063 24
rect 3196 9 3207 65
rect 3263 9 3274 65
rect 3396 25 3407 81
rect 3463 25 3474 81
rect 3796 81 3874 82
rect 3396 24 3474 25
rect 3596 65 3674 66
rect 3196 8 3274 9
rect 3007 -74 3009 -72
rect 3061 -74 3063 -72
rect 3007 -81 3063 -74
rect 3107 -15 3163 0
rect 3107 -67 3109 -15
rect 3161 -67 3163 -15
rect 3107 -79 3163 -67
rect 3107 -110 3109 -79
rect 2961 -131 3109 -110
rect 3161 -110 3163 -79
rect 3207 -16 3263 8
rect 3207 -74 3209 -72
rect 3261 -74 3263 -72
rect 3207 -81 3263 -74
rect 3307 -15 3363 0
rect 3307 -67 3309 -15
rect 3361 -67 3363 -15
rect 3307 -79 3363 -67
rect 3307 -110 3309 -79
rect 3161 -131 3309 -110
rect 3361 -110 3363 -79
rect 3407 -16 3463 24
rect 3596 9 3607 65
rect 3663 9 3674 65
rect 3796 25 3807 81
rect 3863 25 3874 81
rect 4196 81 4274 82
rect 3796 24 3874 25
rect 3996 65 4074 66
rect 3596 8 3674 9
rect 3407 -74 3409 -72
rect 3461 -74 3463 -72
rect 3407 -81 3463 -74
rect 3507 -15 3563 0
rect 3507 -67 3509 -15
rect 3561 -67 3563 -15
rect 3507 -79 3563 -67
rect 3507 -110 3509 -79
rect 3361 -131 3509 -110
rect 3561 -110 3563 -79
rect 3607 -16 3663 8
rect 3607 -74 3609 -72
rect 3661 -74 3663 -72
rect 3607 -81 3663 -74
rect 3707 -15 3763 0
rect 3707 -67 3709 -15
rect 3761 -67 3763 -15
rect 3707 -79 3763 -67
rect 3707 -110 3709 -79
rect 3561 -131 3709 -110
rect 3761 -110 3763 -79
rect 3807 -16 3863 24
rect 3996 9 4007 65
rect 4063 9 4074 65
rect 4196 25 4207 81
rect 4263 25 4274 81
rect 4596 81 4674 82
rect 4196 24 4274 25
rect 4396 65 4474 66
rect 3996 8 4074 9
rect 3807 -74 3809 -72
rect 3861 -74 3863 -72
rect 3807 -81 3863 -74
rect 3907 -15 3963 0
rect 3907 -67 3909 -15
rect 3961 -67 3963 -15
rect 3907 -79 3963 -67
rect 3907 -110 3909 -79
rect 3761 -131 3909 -110
rect 3961 -110 3963 -79
rect 4007 -16 4063 8
rect 4007 -74 4009 -72
rect 4061 -74 4063 -72
rect 4007 -81 4063 -74
rect 4107 -15 4163 0
rect 4107 -67 4109 -15
rect 4161 -67 4163 -15
rect 4107 -79 4163 -67
rect 4107 -110 4109 -79
rect 3961 -131 4109 -110
rect 4161 -110 4163 -79
rect 4207 -16 4263 24
rect 4396 9 4407 65
rect 4463 9 4474 65
rect 4596 25 4607 81
rect 4663 25 4674 81
rect 4996 81 5074 82
rect 4596 24 4674 25
rect 4796 65 4874 66
rect 4396 8 4474 9
rect 4207 -74 4209 -72
rect 4261 -74 4263 -72
rect 4207 -81 4263 -74
rect 4307 -15 4363 0
rect 4307 -67 4309 -15
rect 4361 -67 4363 -15
rect 4307 -79 4363 -67
rect 4307 -110 4309 -79
rect 4161 -131 4309 -110
rect 4361 -110 4363 -79
rect 4407 -16 4463 8
rect 4407 -74 4409 -72
rect 4461 -74 4463 -72
rect 4407 -81 4463 -74
rect 4507 -15 4563 0
rect 4507 -67 4509 -15
rect 4561 -67 4563 -15
rect 4507 -79 4563 -67
rect 4507 -110 4509 -79
rect 4361 -131 4509 -110
rect 4561 -110 4563 -79
rect 4607 -16 4663 24
rect 4796 9 4807 65
rect 4863 9 4874 65
rect 4996 25 5007 81
rect 5063 25 5074 81
rect 5396 81 5474 82
rect 4996 24 5074 25
rect 5196 65 5274 66
rect 4796 8 4874 9
rect 4607 -74 4609 -72
rect 4661 -74 4663 -72
rect 4607 -81 4663 -74
rect 4707 -15 4763 0
rect 4707 -67 4709 -15
rect 4761 -67 4763 -15
rect 4707 -79 4763 -67
rect 4707 -110 4709 -79
rect 4561 -131 4709 -110
rect 4761 -110 4763 -79
rect 4807 -16 4863 8
rect 4807 -74 4809 -72
rect 4861 -74 4863 -72
rect 4807 -81 4863 -74
rect 4907 -15 4963 0
rect 4907 -67 4909 -15
rect 4961 -67 4963 -15
rect 4907 -79 4963 -67
rect 4907 -110 4909 -79
rect 4761 -131 4909 -110
rect 4961 -110 4963 -79
rect 5007 -16 5063 24
rect 5196 9 5207 65
rect 5263 9 5274 65
rect 5396 25 5407 81
rect 5463 25 5474 81
rect 5796 81 5874 82
rect 5396 24 5474 25
rect 5596 65 5674 66
rect 5196 8 5274 9
rect 5007 -74 5009 -72
rect 5061 -74 5063 -72
rect 5007 -81 5063 -74
rect 5107 -15 5163 0
rect 5107 -67 5109 -15
rect 5161 -67 5163 -15
rect 5107 -79 5163 -67
rect 5107 -110 5109 -79
rect 4961 -131 5109 -110
rect 5161 -110 5163 -79
rect 5207 -16 5263 8
rect 5207 -74 5209 -72
rect 5261 -74 5263 -72
rect 5207 -81 5263 -74
rect 5307 -15 5363 0
rect 5307 -67 5309 -15
rect 5361 -67 5363 -15
rect 5307 -79 5363 -67
rect 5307 -110 5309 -79
rect 5161 -131 5309 -110
rect 5361 -110 5363 -79
rect 5407 -16 5463 24
rect 5596 9 5607 65
rect 5663 9 5674 65
rect 5796 25 5807 81
rect 5863 25 5874 81
rect 6196 81 6274 82
rect 5796 24 5874 25
rect 5996 65 6074 66
rect 5596 8 5674 9
rect 5407 -74 5409 -72
rect 5461 -74 5463 -72
rect 5407 -81 5463 -74
rect 5507 -15 5563 0
rect 5507 -67 5509 -15
rect 5561 -67 5563 -15
rect 5507 -79 5563 -67
rect 5507 -110 5509 -79
rect 5361 -131 5509 -110
rect 5561 -110 5563 -79
rect 5607 -16 5663 8
rect 5607 -74 5609 -72
rect 5661 -74 5663 -72
rect 5607 -81 5663 -74
rect 5707 -15 5763 0
rect 5707 -67 5709 -15
rect 5761 -67 5763 -15
rect 5707 -79 5763 -67
rect 5707 -110 5709 -79
rect 5561 -131 5709 -110
rect 5761 -110 5763 -79
rect 5807 -16 5863 24
rect 5996 9 6007 65
rect 6063 9 6074 65
rect 6196 25 6207 81
rect 6263 25 6274 81
rect 6196 24 6274 25
rect 5996 8 6074 9
rect 5807 -74 5809 -72
rect 5861 -74 5863 -72
rect 5807 -81 5863 -74
rect 5907 -15 5963 0
rect 5907 -67 5909 -15
rect 5961 -67 5963 -15
rect 5907 -79 5963 -67
rect 5907 -110 5909 -79
rect 5761 -131 5909 -110
rect 5961 -110 5963 -79
rect 6007 -16 6063 8
rect 6007 -74 6009 -72
rect 6061 -74 6063 -72
rect 6007 -81 6063 -74
rect 6107 -15 6163 0
rect 6107 -67 6109 -15
rect 6161 -67 6163 -15
rect 6107 -79 6163 -67
rect 6107 -110 6109 -79
rect 5961 -131 6109 -110
rect 6161 -110 6163 -79
rect 6207 -16 6263 24
rect 8126 3 8297 12
rect 6207 -74 6209 -72
rect 6261 -74 6263 -72
rect 6207 -81 6263 -74
rect 6307 -15 6363 0
rect 6307 -67 6309 -15
rect 6361 -67 6363 -15
rect 8126 -53 8143 3
rect 8199 1 8223 3
rect 8205 -51 8217 1
rect 8199 -53 8223 -51
rect 8279 -53 8297 3
rect 8126 -62 8297 -53
rect 8405 3 8736 12
rect 8405 1 8422 3
rect 8478 1 8502 3
rect 8558 1 8582 3
rect 8638 1 8662 3
rect 8718 1 8736 3
rect 8405 -51 8416 1
rect 8478 -51 8480 1
rect 8660 -51 8662 1
rect 8724 -51 8736 1
rect 8405 -53 8422 -51
rect 8478 -53 8502 -51
rect 8558 -53 8582 -51
rect 8638 -53 8662 -51
rect 8718 -53 8736 -51
rect 8405 -62 8736 -53
rect 8806 3 9137 12
rect 8806 1 8823 3
rect 8879 1 8903 3
rect 8959 1 8983 3
rect 9039 1 9063 3
rect 9119 1 9137 3
rect 8806 -51 8817 1
rect 8879 -51 8881 1
rect 9061 -51 9063 1
rect 9125 -51 9137 1
rect 8806 -53 8823 -51
rect 8879 -53 8903 -51
rect 8959 -53 8983 -51
rect 9039 -53 9063 -51
rect 9119 -53 9137 -51
rect 8806 -62 9137 -53
rect 9245 3 9416 12
rect 9245 -53 9262 3
rect 9318 1 9342 3
rect 9324 -51 9336 1
rect 9318 -53 9342 -51
rect 9398 -53 9416 3
rect 9245 -62 9416 -53
rect 6307 -79 6363 -67
rect 6307 -110 6309 -79
rect 6161 -131 6309 -110
rect 6361 -110 6363 -79
rect 6361 -131 6408 -110
rect -138 -143 6408 -131
rect -138 -145 -91 -143
rect -39 -145 109 -143
rect 161 -145 309 -143
rect 361 -145 509 -143
rect 561 -145 709 -143
rect 761 -145 909 -143
rect 961 -145 1109 -143
rect 1161 -145 1309 -143
rect 1361 -145 1509 -143
rect 1561 -145 1709 -143
rect 1761 -145 1909 -143
rect 1961 -145 2109 -143
rect 2161 -145 2309 -143
rect 2361 -145 2509 -143
rect 2561 -145 2709 -143
rect 2761 -145 2909 -143
rect 2961 -145 3109 -143
rect 3161 -145 3309 -143
rect 3361 -145 3509 -143
rect 3561 -145 3709 -143
rect 3761 -145 3909 -143
rect 3961 -145 4109 -143
rect 4161 -145 4309 -143
rect 4361 -145 4509 -143
rect 4561 -145 4709 -143
rect 4761 -145 4909 -143
rect 4961 -145 5109 -143
rect 5161 -145 5309 -143
rect 5361 -145 5509 -143
rect 5561 -145 5709 -143
rect 5761 -145 5909 -143
rect 5961 -145 6109 -143
rect 6161 -145 6309 -143
rect 6361 -145 6408 -143
rect -138 -201 -133 -145
rect -77 -201 -53 -195
rect 3 -201 67 -145
rect 123 -201 147 -195
rect 203 -201 267 -145
rect 323 -201 347 -195
rect 403 -201 467 -145
rect 523 -201 547 -195
rect 603 -201 667 -145
rect 723 -201 747 -195
rect 803 -201 867 -145
rect 923 -201 947 -195
rect 1003 -201 1067 -145
rect 1123 -201 1147 -195
rect 1203 -201 1267 -145
rect 1323 -201 1347 -195
rect 1403 -201 1467 -145
rect 1523 -201 1547 -195
rect 1603 -201 1667 -145
rect 1723 -201 1747 -195
rect 1803 -201 1867 -145
rect 1923 -201 1947 -195
rect 2003 -201 2067 -145
rect 2123 -201 2147 -195
rect 2203 -201 2267 -145
rect 2323 -201 2347 -195
rect 2403 -201 2467 -145
rect 2523 -201 2547 -195
rect 2603 -201 2667 -145
rect 2723 -201 2747 -195
rect 2803 -201 2867 -145
rect 2923 -201 2947 -195
rect 3003 -201 3067 -145
rect 3123 -201 3147 -195
rect 3203 -201 3267 -145
rect 3323 -201 3347 -195
rect 3403 -201 3467 -145
rect 3523 -201 3547 -195
rect 3603 -201 3667 -145
rect 3723 -201 3747 -195
rect 3803 -201 3867 -145
rect 3923 -201 3947 -195
rect 4003 -201 4067 -145
rect 4123 -201 4147 -195
rect 4203 -201 4267 -145
rect 4323 -201 4347 -195
rect 4403 -201 4467 -145
rect 4523 -201 4547 -195
rect 4603 -201 4667 -145
rect 4723 -201 4747 -195
rect 4803 -201 4867 -145
rect 4923 -201 4947 -195
rect 5003 -201 5067 -145
rect 5123 -201 5147 -195
rect 5203 -201 5267 -145
rect 5323 -201 5347 -195
rect 5403 -201 5467 -145
rect 5523 -201 5547 -195
rect 5603 -201 5667 -145
rect 5723 -201 5747 -195
rect 5803 -201 5867 -145
rect 5923 -201 5947 -195
rect 6003 -201 6067 -145
rect 6123 -201 6147 -195
rect 6203 -201 6267 -145
rect 6323 -201 6347 -195
rect 6403 -201 6408 -145
rect -138 -210 6408 -201
rect 8040 -151 8812 -99
rect 8864 -151 8870 -99
rect 9165 -151 9440 -99
rect 8040 -199 8092 -151
rect -81 -291 -75 -239
rect -23 -291 61 -239
rect 119 -291 125 -239
rect 177 -291 261 -239
rect 319 -291 325 -239
rect 377 -291 461 -239
rect 519 -291 525 -239
rect 577 -291 661 -239
rect 719 -291 725 -239
rect 777 -291 861 -239
rect 919 -291 925 -239
rect 977 -291 1061 -239
rect 1119 -291 1125 -239
rect 1177 -291 1261 -239
rect 1319 -291 1325 -239
rect 1377 -291 1461 -239
rect 1519 -291 1525 -239
rect 1577 -291 1661 -239
rect 1719 -291 1725 -239
rect 1777 -291 1861 -239
rect 1919 -291 1925 -239
rect 1977 -291 2061 -239
rect 2119 -291 2125 -239
rect 2177 -291 2261 -239
rect 2319 -291 2325 -239
rect 2377 -291 2461 -239
rect 2519 -291 2525 -239
rect 2577 -291 2661 -239
rect 2719 -291 2725 -239
rect 2777 -291 2861 -239
rect 2919 -291 2925 -239
rect 2977 -291 3061 -239
rect 3119 -291 3125 -239
rect 3177 -291 3261 -239
rect 3319 -291 3325 -239
rect 3377 -291 3461 -239
rect 3519 -291 3525 -239
rect 3577 -291 3661 -239
rect 3719 -291 3725 -239
rect 3777 -291 3861 -239
rect 3919 -291 3925 -239
rect 3977 -291 4061 -239
rect 4119 -291 4125 -239
rect 4177 -291 4261 -239
rect 4319 -291 4325 -239
rect 4377 -291 4461 -239
rect 4519 -291 4525 -239
rect 4577 -291 4661 -239
rect 4719 -291 4725 -239
rect 4777 -291 4861 -239
rect 4919 -291 4925 -239
rect 4977 -291 5061 -239
rect 5119 -291 5125 -239
rect 5177 -291 5261 -239
rect 5319 -291 5325 -239
rect 5377 -291 5461 -239
rect 5519 -291 5525 -239
rect 5577 -291 5661 -239
rect 5719 -291 5725 -239
rect 5777 -291 5861 -239
rect 5919 -291 5925 -239
rect 5977 -291 6061 -239
rect 6119 -291 6125 -239
rect 6177 -291 6261 -239
rect 8040 -257 8092 -251
rect 8126 -197 8297 -188
rect 8126 -253 8143 -197
rect 8199 -199 8223 -197
rect 8205 -251 8217 -199
rect 8199 -253 8223 -251
rect 8279 -253 8297 -197
rect 8126 -262 8297 -253
rect 8325 -199 8377 -151
rect 8325 -257 8377 -251
rect 8405 -197 8736 -188
rect 8405 -199 8422 -197
rect 8478 -199 8502 -197
rect 8558 -199 8582 -197
rect 8638 -199 8662 -197
rect 8718 -199 8736 -197
rect 8405 -251 8416 -199
rect 8478 -251 8480 -199
rect 8660 -251 8662 -199
rect 8724 -251 8736 -199
rect 8405 -253 8422 -251
rect 8478 -253 8502 -251
rect 8558 -253 8582 -251
rect 8638 -253 8662 -251
rect 8718 -253 8736 -251
rect 8405 -262 8736 -253
rect 8806 -197 9137 -188
rect 8806 -199 8823 -197
rect 8879 -199 8903 -197
rect 8959 -199 8983 -197
rect 9039 -199 9063 -197
rect 9119 -199 9137 -197
rect 8806 -251 8817 -199
rect 8879 -251 8881 -199
rect 9061 -251 9063 -199
rect 9125 -251 9137 -199
rect 8806 -253 8823 -251
rect 8879 -253 8903 -251
rect 8959 -253 8983 -251
rect 9039 -253 9063 -251
rect 9119 -253 9137 -251
rect 8806 -262 9137 -253
rect 9165 -199 9217 -151
rect 9165 -257 9217 -251
rect 9245 -197 9416 -188
rect 9245 -253 9262 -197
rect 9318 -199 9342 -197
rect 9324 -251 9336 -199
rect 9318 -253 9342 -251
rect 9398 -253 9416 -197
rect 9245 -262 9416 -253
rect -93 -326 -37 -320
rect -93 -348 -91 -326
rect -39 -348 -37 -326
rect -93 -428 -91 -404
rect -39 -428 -37 -404
rect -93 -506 -91 -484
rect -39 -506 -37 -484
rect -93 -512 -37 -506
rect 9 -828 61 -291
rect 107 -326 163 -320
rect 107 -348 109 -326
rect 161 -348 163 -326
rect 107 -428 109 -404
rect 161 -428 163 -404
rect 107 -506 109 -484
rect 161 -506 163 -484
rect 107 -512 163 -506
rect 209 -828 261 -291
rect 307 -326 363 -320
rect 307 -348 309 -326
rect 361 -348 363 -326
rect 307 -428 309 -404
rect 361 -428 363 -404
rect 307 -506 309 -484
rect 361 -506 363 -484
rect 307 -512 363 -506
rect 409 -828 461 -291
rect 507 -326 563 -320
rect 507 -348 509 -326
rect 561 -348 563 -326
rect 507 -428 509 -404
rect 561 -428 563 -404
rect 507 -506 509 -484
rect 561 -506 563 -484
rect 507 -512 563 -506
rect 609 -828 661 -291
rect 707 -326 763 -320
rect 707 -348 709 -326
rect 761 -348 763 -326
rect 707 -428 709 -404
rect 761 -428 763 -404
rect 707 -506 709 -484
rect 761 -506 763 -484
rect 707 -512 763 -506
rect 809 -828 861 -291
rect 907 -326 963 -320
rect 907 -348 909 -326
rect 961 -348 963 -326
rect 907 -428 909 -404
rect 961 -428 963 -404
rect 907 -506 909 -484
rect 961 -506 963 -484
rect 907 -512 963 -506
rect 1009 -828 1061 -291
rect 1107 -326 1163 -320
rect 1107 -348 1109 -326
rect 1161 -348 1163 -326
rect 1107 -428 1109 -404
rect 1161 -428 1163 -404
rect 1107 -506 1109 -484
rect 1161 -506 1163 -484
rect 1107 -512 1163 -506
rect 1209 -828 1261 -291
rect 1307 -326 1363 -320
rect 1307 -348 1309 -326
rect 1361 -348 1363 -326
rect 1307 -428 1309 -404
rect 1361 -428 1363 -404
rect 1307 -506 1309 -484
rect 1361 -506 1363 -484
rect 1307 -512 1363 -506
rect 1409 -828 1461 -291
rect 1507 -326 1563 -320
rect 1507 -348 1509 -326
rect 1561 -348 1563 -326
rect 1507 -428 1509 -404
rect 1561 -428 1563 -404
rect 1507 -506 1509 -484
rect 1561 -506 1563 -484
rect 1507 -512 1563 -506
rect 1609 -828 1661 -291
rect 1707 -326 1763 -320
rect 1707 -348 1709 -326
rect 1761 -348 1763 -326
rect 1707 -428 1709 -404
rect 1761 -428 1763 -404
rect 1707 -506 1709 -484
rect 1761 -506 1763 -484
rect 1707 -512 1763 -506
rect 1809 -828 1861 -291
rect 1907 -326 1963 -320
rect 1907 -348 1909 -326
rect 1961 -348 1963 -326
rect 1907 -428 1909 -404
rect 1961 -428 1963 -404
rect 1907 -506 1909 -484
rect 1961 -506 1963 -484
rect 1907 -512 1963 -506
rect 2009 -828 2061 -291
rect 2107 -326 2163 -320
rect 2107 -348 2109 -326
rect 2161 -348 2163 -326
rect 2107 -428 2109 -404
rect 2161 -428 2163 -404
rect 2107 -506 2109 -484
rect 2161 -506 2163 -484
rect 2107 -512 2163 -506
rect 2209 -828 2261 -291
rect 2307 -326 2363 -320
rect 2307 -348 2309 -326
rect 2361 -348 2363 -326
rect 2307 -428 2309 -404
rect 2361 -428 2363 -404
rect 2307 -506 2309 -484
rect 2361 -506 2363 -484
rect 2307 -512 2363 -506
rect 2409 -828 2461 -291
rect 2507 -326 2563 -320
rect 2507 -348 2509 -326
rect 2561 -348 2563 -326
rect 2507 -428 2509 -404
rect 2561 -428 2563 -404
rect 2507 -506 2509 -484
rect 2561 -506 2563 -484
rect 2507 -512 2563 -506
rect 2609 -828 2661 -291
rect 2707 -326 2763 -320
rect 2707 -348 2709 -326
rect 2761 -348 2763 -326
rect 2707 -428 2709 -404
rect 2761 -428 2763 -404
rect 2707 -506 2709 -484
rect 2761 -506 2763 -484
rect 2707 -512 2763 -506
rect 2809 -828 2861 -291
rect 2907 -326 2963 -320
rect 2907 -348 2909 -326
rect 2961 -348 2963 -326
rect 2907 -428 2909 -404
rect 2961 -428 2963 -404
rect 2907 -506 2909 -484
rect 2961 -506 2963 -484
rect 2907 -512 2963 -506
rect 3009 -828 3061 -291
rect 3107 -326 3163 -320
rect 3107 -348 3109 -326
rect 3161 -348 3163 -326
rect 3107 -428 3109 -404
rect 3161 -428 3163 -404
rect 3107 -506 3109 -484
rect 3161 -506 3163 -484
rect 3107 -512 3163 -506
rect 3209 -828 3261 -291
rect 3307 -326 3363 -320
rect 3307 -348 3309 -326
rect 3361 -348 3363 -326
rect 3307 -428 3309 -404
rect 3361 -428 3363 -404
rect 3307 -506 3309 -484
rect 3361 -506 3363 -484
rect 3307 -512 3363 -506
rect 3409 -828 3461 -291
rect 3507 -326 3563 -320
rect 3507 -348 3509 -326
rect 3561 -348 3563 -326
rect 3507 -428 3509 -404
rect 3561 -428 3563 -404
rect 3507 -506 3509 -484
rect 3561 -506 3563 -484
rect 3507 -512 3563 -506
rect 3609 -828 3661 -291
rect 3707 -326 3763 -320
rect 3707 -348 3709 -326
rect 3761 -348 3763 -326
rect 3707 -428 3709 -404
rect 3761 -428 3763 -404
rect 3707 -506 3709 -484
rect 3761 -506 3763 -484
rect 3707 -512 3763 -506
rect 3809 -828 3861 -291
rect 3907 -326 3963 -320
rect 3907 -348 3909 -326
rect 3961 -348 3963 -326
rect 3907 -428 3909 -404
rect 3961 -428 3963 -404
rect 3907 -506 3909 -484
rect 3961 -506 3963 -484
rect 3907 -512 3963 -506
rect 4009 -828 4061 -291
rect 4107 -326 4163 -320
rect 4107 -348 4109 -326
rect 4161 -348 4163 -326
rect 4107 -428 4109 -404
rect 4161 -428 4163 -404
rect 4107 -506 4109 -484
rect 4161 -506 4163 -484
rect 4107 -512 4163 -506
rect 4209 -828 4261 -291
rect 4307 -326 4363 -320
rect 4307 -348 4309 -326
rect 4361 -348 4363 -326
rect 4307 -428 4309 -404
rect 4361 -428 4363 -404
rect 4307 -506 4309 -484
rect 4361 -506 4363 -484
rect 4307 -512 4363 -506
rect 4409 -828 4461 -291
rect 4507 -326 4563 -320
rect 4507 -348 4509 -326
rect 4561 -348 4563 -326
rect 4507 -428 4509 -404
rect 4561 -428 4563 -404
rect 4507 -506 4509 -484
rect 4561 -506 4563 -484
rect 4507 -512 4563 -506
rect 4609 -828 4661 -291
rect 4707 -326 4763 -320
rect 4707 -348 4709 -326
rect 4761 -348 4763 -326
rect 4707 -428 4709 -404
rect 4761 -428 4763 -404
rect 4707 -506 4709 -484
rect 4761 -506 4763 -484
rect 4707 -512 4763 -506
rect 4809 -828 4861 -291
rect 4907 -326 4963 -320
rect 4907 -348 4909 -326
rect 4961 -348 4963 -326
rect 4907 -428 4909 -404
rect 4961 -428 4963 -404
rect 4907 -506 4909 -484
rect 4961 -506 4963 -484
rect 4907 -512 4963 -506
rect 5009 -828 5061 -291
rect 5107 -326 5163 -320
rect 5107 -348 5109 -326
rect 5161 -348 5163 -326
rect 5107 -428 5109 -404
rect 5161 -428 5163 -404
rect 5107 -506 5109 -484
rect 5161 -506 5163 -484
rect 5107 -512 5163 -506
rect 5209 -828 5261 -291
rect 5307 -326 5363 -320
rect 5307 -348 5309 -326
rect 5361 -348 5363 -326
rect 5307 -428 5309 -404
rect 5361 -428 5363 -404
rect 5307 -506 5309 -484
rect 5361 -506 5363 -484
rect 5307 -512 5363 -506
rect 5409 -828 5461 -291
rect 5507 -326 5563 -320
rect 5507 -348 5509 -326
rect 5561 -348 5563 -326
rect 5507 -428 5509 -404
rect 5561 -428 5563 -404
rect 5507 -506 5509 -484
rect 5561 -506 5563 -484
rect 5507 -512 5563 -506
rect 5609 -828 5661 -291
rect 5707 -326 5763 -320
rect 5707 -348 5709 -326
rect 5761 -348 5763 -326
rect 5707 -428 5709 -404
rect 5761 -428 5763 -404
rect 5707 -506 5709 -484
rect 5761 -506 5763 -484
rect 5707 -512 5763 -506
rect 5809 -828 5861 -291
rect 5907 -326 5963 -320
rect 5907 -348 5909 -326
rect 5961 -348 5963 -326
rect 5907 -428 5909 -404
rect 5961 -428 5963 -404
rect 5907 -506 5909 -484
rect 5961 -506 5963 -484
rect 5907 -512 5963 -506
rect 6009 -828 6061 -291
rect 6107 -326 6163 -320
rect 6107 -348 6109 -326
rect 6161 -348 6163 -326
rect 6107 -428 6109 -404
rect 6161 -428 6163 -404
rect 6107 -506 6109 -484
rect 6161 -506 6163 -484
rect 6107 -512 6163 -506
rect 6209 -828 6261 -291
rect 6307 -326 6363 -320
rect 6307 -348 6309 -326
rect 6361 -348 6363 -326
rect 6307 -428 6309 -404
rect 6361 -428 6363 -404
rect 8040 -351 8812 -299
rect 8864 -351 8870 -299
rect 9165 -351 9440 -299
rect 8040 -399 8092 -351
rect 8040 -457 8092 -451
rect 8126 -397 8297 -388
rect 8126 -453 8143 -397
rect 8199 -399 8223 -397
rect 8205 -451 8217 -399
rect 8199 -453 8223 -451
rect 8279 -453 8297 -397
rect 8126 -462 8297 -453
rect 8325 -399 8377 -351
rect 8325 -457 8377 -451
rect 8405 -397 8736 -388
rect 8405 -399 8422 -397
rect 8478 -399 8502 -397
rect 8558 -399 8582 -397
rect 8638 -399 8662 -397
rect 8718 -399 8736 -397
rect 8405 -451 8416 -399
rect 8478 -451 8480 -399
rect 8660 -451 8662 -399
rect 8724 -451 8736 -399
rect 8405 -453 8422 -451
rect 8478 -453 8502 -451
rect 8558 -453 8582 -451
rect 8638 -453 8662 -451
rect 8718 -453 8736 -451
rect 8405 -462 8736 -453
rect 8806 -397 9137 -388
rect 8806 -399 8823 -397
rect 8879 -399 8903 -397
rect 8959 -399 8983 -397
rect 9039 -399 9063 -397
rect 9119 -399 9137 -397
rect 8806 -451 8817 -399
rect 8879 -451 8881 -399
rect 9061 -451 9063 -399
rect 9125 -451 9137 -399
rect 8806 -453 8823 -451
rect 8879 -453 8903 -451
rect 8959 -453 8983 -451
rect 9039 -453 9063 -451
rect 9119 -453 9137 -451
rect 8806 -462 9137 -453
rect 9165 -399 9217 -351
rect 9165 -457 9217 -451
rect 9245 -397 9416 -388
rect 9245 -453 9262 -397
rect 9318 -399 9342 -397
rect 9324 -451 9336 -399
rect 9318 -453 9342 -451
rect 9398 -453 9416 -397
rect 9245 -462 9416 -453
rect 6307 -506 6309 -484
rect 6361 -506 6363 -484
rect 6307 -512 6363 -506
rect 8040 -551 8812 -499
rect 8864 -551 8870 -499
rect 9165 -551 9440 -499
rect 8040 -599 8092 -551
rect 8040 -657 8092 -651
rect 8126 -597 8297 -588
rect 8126 -653 8143 -597
rect 8199 -599 8223 -597
rect 8205 -651 8217 -599
rect 8199 -653 8223 -651
rect 8279 -653 8297 -597
rect 8126 -662 8297 -653
rect 8325 -599 8377 -551
rect 8325 -657 8377 -651
rect 8405 -597 8736 -588
rect 8405 -599 8422 -597
rect 8478 -599 8502 -597
rect 8558 -599 8582 -597
rect 8638 -599 8662 -597
rect 8718 -599 8736 -597
rect 8405 -651 8416 -599
rect 8478 -651 8480 -599
rect 8660 -651 8662 -599
rect 8724 -651 8736 -599
rect 8405 -653 8422 -651
rect 8478 -653 8502 -651
rect 8558 -653 8582 -651
rect 8638 -653 8662 -651
rect 8718 -653 8736 -651
rect 8405 -662 8736 -653
rect 8806 -597 9137 -588
rect 8806 -599 8823 -597
rect 8879 -599 8903 -597
rect 8959 -599 8983 -597
rect 9039 -599 9063 -597
rect 9119 -599 9137 -597
rect 8806 -651 8817 -599
rect 8879 -651 8881 -599
rect 9061 -651 9063 -599
rect 9125 -651 9137 -599
rect 8806 -653 8823 -651
rect 8879 -653 8903 -651
rect 8959 -653 8983 -651
rect 9039 -653 9063 -651
rect 9119 -653 9137 -651
rect 8806 -662 9137 -653
rect 9165 -599 9217 -551
rect 9165 -657 9217 -651
rect 9245 -597 9416 -588
rect 9245 -653 9262 -597
rect 9318 -599 9342 -597
rect 9324 -651 9336 -599
rect 9318 -653 9342 -651
rect 9398 -653 9416 -597
rect 9245 -662 9416 -653
rect 8040 -751 8812 -699
rect 8864 -751 8870 -699
rect 9165 -751 9440 -699
rect 8040 -799 8092 -751
rect -18 -880 -9 -828
rect 43 -880 55 -828
rect 107 -880 116 -828
rect 154 -880 163 -828
rect 215 -880 227 -828
rect 279 -880 288 -828
rect 382 -880 391 -828
rect 443 -880 455 -828
rect 507 -880 516 -828
rect 554 -880 563 -828
rect 615 -880 627 -828
rect 679 -880 688 -828
rect 782 -880 791 -828
rect 843 -880 855 -828
rect 907 -880 916 -828
rect 954 -880 963 -828
rect 1015 -880 1027 -828
rect 1079 -880 1088 -828
rect 1182 -880 1191 -828
rect 1243 -880 1255 -828
rect 1307 -880 1316 -828
rect 1354 -880 1363 -828
rect 1415 -880 1427 -828
rect 1479 -880 1488 -828
rect 1582 -880 1591 -828
rect 1643 -880 1655 -828
rect 1707 -880 1716 -828
rect 1754 -880 1763 -828
rect 1815 -880 1827 -828
rect 1879 -880 1888 -828
rect 1982 -880 1991 -828
rect 2043 -880 2055 -828
rect 2107 -880 2116 -828
rect 2154 -880 2163 -828
rect 2215 -880 2227 -828
rect 2279 -880 2288 -828
rect 2382 -880 2391 -828
rect 2443 -880 2455 -828
rect 2507 -880 2516 -828
rect 2554 -880 2563 -828
rect 2615 -880 2627 -828
rect 2679 -880 2688 -828
rect 2782 -880 2791 -828
rect 2843 -880 2855 -828
rect 2907 -880 2916 -828
rect 2954 -880 2963 -828
rect 3015 -880 3027 -828
rect 3079 -880 3088 -828
rect 3182 -880 3191 -828
rect 3243 -880 3255 -828
rect 3307 -880 3316 -828
rect 3354 -880 3363 -828
rect 3415 -880 3427 -828
rect 3479 -880 3488 -828
rect 3582 -880 3591 -828
rect 3643 -880 3655 -828
rect 3707 -880 3716 -828
rect 3754 -880 3763 -828
rect 3815 -880 3827 -828
rect 3879 -880 3888 -828
rect 3982 -880 3991 -828
rect 4043 -880 4055 -828
rect 4107 -880 4116 -828
rect 4154 -880 4163 -828
rect 4215 -880 4227 -828
rect 4279 -880 4288 -828
rect 4382 -880 4391 -828
rect 4443 -880 4455 -828
rect 4507 -880 4516 -828
rect 4554 -880 4563 -828
rect 4615 -880 4627 -828
rect 4679 -880 4688 -828
rect 4782 -880 4791 -828
rect 4843 -880 4855 -828
rect 4907 -880 4916 -828
rect 4954 -880 4963 -828
rect 5015 -880 5027 -828
rect 5079 -880 5088 -828
rect 5182 -880 5191 -828
rect 5243 -880 5255 -828
rect 5307 -880 5316 -828
rect 5354 -880 5363 -828
rect 5415 -880 5427 -828
rect 5479 -880 5488 -828
rect 5582 -880 5591 -828
rect 5643 -880 5655 -828
rect 5707 -880 5716 -828
rect 5754 -880 5763 -828
rect 5815 -880 5827 -828
rect 5879 -880 5888 -828
rect 5982 -880 5991 -828
rect 6043 -880 6055 -828
rect 6107 -880 6116 -828
rect 6154 -880 6163 -828
rect 6215 -880 6227 -828
rect 6279 -880 6288 -828
rect 8040 -857 8092 -851
rect 8126 -797 8297 -788
rect 8126 -853 8143 -797
rect 8199 -799 8223 -797
rect 8205 -851 8217 -799
rect 8199 -853 8223 -851
rect 8279 -853 8297 -797
rect 8126 -862 8297 -853
rect 8325 -799 8377 -751
rect 8325 -857 8377 -851
rect 8405 -797 8736 -788
rect 8405 -799 8422 -797
rect 8478 -799 8502 -797
rect 8558 -799 8582 -797
rect 8638 -799 8662 -797
rect 8718 -799 8736 -797
rect 8405 -851 8416 -799
rect 8478 -851 8480 -799
rect 8660 -851 8662 -799
rect 8724 -851 8736 -799
rect 8405 -853 8422 -851
rect 8478 -853 8502 -851
rect 8558 -853 8582 -851
rect 8638 -853 8662 -851
rect 8718 -853 8736 -851
rect 8405 -862 8736 -853
rect 8806 -797 9137 -788
rect 8806 -799 8823 -797
rect 8879 -799 8903 -797
rect 8959 -799 8983 -797
rect 9039 -799 9063 -797
rect 9119 -799 9137 -797
rect 8806 -851 8817 -799
rect 8879 -851 8881 -799
rect 9061 -851 9063 -799
rect 9125 -851 9137 -799
rect 8806 -853 8823 -851
rect 8879 -853 8903 -851
rect 8959 -853 8983 -851
rect 9039 -853 9063 -851
rect 9119 -853 9137 -851
rect 8806 -862 9137 -853
rect 9165 -799 9217 -751
rect 9165 -857 9217 -851
rect 9245 -797 9416 -788
rect 9245 -853 9262 -797
rect 9318 -799 9342 -797
rect 9324 -851 9336 -799
rect 9318 -853 9342 -851
rect 9398 -853 9416 -797
rect 9245 -862 9416 -853
rect 8040 -951 8812 -899
rect 8864 -951 8870 -899
rect 9165 -951 9440 -899
rect 8040 -999 8092 -951
rect 8040 -1057 8092 -1051
rect 8126 -997 8297 -988
rect 8126 -1053 8143 -997
rect 8199 -999 8223 -997
rect 8205 -1051 8217 -999
rect 8199 -1053 8223 -1051
rect 8279 -1053 8297 -997
rect 8126 -1062 8297 -1053
rect 8325 -999 8377 -951
rect 8325 -1057 8377 -1051
rect 8405 -997 8736 -988
rect 8405 -999 8422 -997
rect 8478 -999 8502 -997
rect 8558 -999 8582 -997
rect 8638 -999 8662 -997
rect 8718 -999 8736 -997
rect 8405 -1051 8416 -999
rect 8478 -1051 8480 -999
rect 8660 -1051 8662 -999
rect 8724 -1051 8736 -999
rect 8405 -1053 8422 -1051
rect 8478 -1053 8502 -1051
rect 8558 -1053 8582 -1051
rect 8638 -1053 8662 -1051
rect 8718 -1053 8736 -1051
rect 8405 -1062 8736 -1053
rect 8806 -997 9137 -988
rect 8806 -999 8823 -997
rect 8879 -999 8903 -997
rect 8959 -999 8983 -997
rect 9039 -999 9063 -997
rect 9119 -999 9137 -997
rect 8806 -1051 8817 -999
rect 8879 -1051 8881 -999
rect 9061 -1051 9063 -999
rect 9125 -1051 9137 -999
rect 8806 -1053 8823 -1051
rect 8879 -1053 8903 -1051
rect 8959 -1053 8983 -1051
rect 9039 -1053 9063 -1051
rect 9119 -1053 9137 -1051
rect 8806 -1062 9137 -1053
rect 9165 -999 9217 -951
rect 9165 -1057 9217 -1051
rect 9245 -997 9416 -988
rect 9245 -1053 9262 -997
rect 9318 -999 9342 -997
rect 9324 -1051 9336 -999
rect 9318 -1053 9342 -1051
rect 9398 -1053 9416 -997
rect 9245 -1062 9416 -1053
rect 8040 -1151 8812 -1099
rect 8864 -1151 8870 -1099
rect 9165 -1151 9440 -1099
rect 8040 -1199 8092 -1151
rect 8040 -1257 8092 -1251
rect 8126 -1197 8297 -1188
rect 8126 -1253 8143 -1197
rect 8199 -1199 8223 -1197
rect 8205 -1251 8217 -1199
rect 8199 -1253 8223 -1251
rect 8279 -1253 8297 -1197
rect 8126 -1262 8297 -1253
rect 8325 -1199 8377 -1151
rect 8325 -1257 8377 -1251
rect 8405 -1197 8736 -1188
rect 8405 -1199 8422 -1197
rect 8478 -1199 8502 -1197
rect 8558 -1199 8582 -1197
rect 8638 -1199 8662 -1197
rect 8718 -1199 8736 -1197
rect 8405 -1251 8416 -1199
rect 8478 -1251 8480 -1199
rect 8660 -1251 8662 -1199
rect 8724 -1251 8736 -1199
rect 8405 -1253 8422 -1251
rect 8478 -1253 8502 -1251
rect 8558 -1253 8582 -1251
rect 8638 -1253 8662 -1251
rect 8718 -1253 8736 -1251
rect 8405 -1262 8736 -1253
rect 8806 -1197 9137 -1188
rect 8806 -1199 8823 -1197
rect 8879 -1199 8903 -1197
rect 8959 -1199 8983 -1197
rect 9039 -1199 9063 -1197
rect 9119 -1199 9137 -1197
rect 8806 -1251 8817 -1199
rect 8879 -1251 8881 -1199
rect 9061 -1251 9063 -1199
rect 9125 -1251 9137 -1199
rect 8806 -1253 8823 -1251
rect 8879 -1253 8903 -1251
rect 8959 -1253 8983 -1251
rect 9039 -1253 9063 -1251
rect 9119 -1253 9137 -1251
rect 8806 -1262 9137 -1253
rect 9165 -1199 9217 -1151
rect 9165 -1257 9217 -1251
rect 9245 -1197 9416 -1188
rect 9245 -1253 9262 -1197
rect 9318 -1199 9342 -1197
rect 9324 -1251 9336 -1199
rect 9318 -1253 9342 -1251
rect 9398 -1253 9416 -1197
rect 9245 -1262 9416 -1253
rect 8040 -1351 8812 -1299
rect 8864 -1351 8870 -1299
rect 9165 -1351 9440 -1299
rect 8040 -1399 8092 -1351
rect 8040 -1457 8092 -1451
rect 8126 -1397 8297 -1388
rect 8126 -1453 8143 -1397
rect 8199 -1399 8223 -1397
rect 8205 -1451 8217 -1399
rect 8199 -1453 8223 -1451
rect 8279 -1453 8297 -1397
rect 8126 -1462 8297 -1453
rect 8325 -1399 8377 -1351
rect 8325 -1457 8377 -1451
rect 8405 -1397 8736 -1388
rect 8405 -1399 8422 -1397
rect 8478 -1399 8502 -1397
rect 8558 -1399 8582 -1397
rect 8638 -1399 8662 -1397
rect 8718 -1399 8736 -1397
rect 8405 -1451 8416 -1399
rect 8478 -1451 8480 -1399
rect 8660 -1451 8662 -1399
rect 8724 -1451 8736 -1399
rect 8405 -1453 8422 -1451
rect 8478 -1453 8502 -1451
rect 8558 -1453 8582 -1451
rect 8638 -1453 8662 -1451
rect 8718 -1453 8736 -1451
rect 8405 -1462 8736 -1453
rect 8806 -1397 9137 -1388
rect 8806 -1399 8823 -1397
rect 8879 -1399 8903 -1397
rect 8959 -1399 8983 -1397
rect 9039 -1399 9063 -1397
rect 9119 -1399 9137 -1397
rect 8806 -1451 8817 -1399
rect 8879 -1451 8881 -1399
rect 9061 -1451 9063 -1399
rect 9125 -1451 9137 -1399
rect 8806 -1453 8823 -1451
rect 8879 -1453 8903 -1451
rect 8959 -1453 8983 -1451
rect 9039 -1453 9063 -1451
rect 9119 -1453 9137 -1451
rect 8806 -1462 9137 -1453
rect 9165 -1399 9217 -1351
rect 9165 -1457 9217 -1451
rect 9245 -1397 9416 -1388
rect 9245 -1453 9262 -1397
rect 9318 -1399 9342 -1397
rect 9324 -1451 9336 -1399
rect 9318 -1453 9342 -1451
rect 9398 -1453 9416 -1397
rect 9245 -1462 9416 -1453
rect 8040 -1551 8812 -1499
rect 8864 -1551 8870 -1499
rect 9165 -1551 9440 -1499
rect 8040 -1599 8092 -1551
rect 8040 -1657 8092 -1651
rect 8126 -1597 8297 -1588
rect 8126 -1653 8143 -1597
rect 8199 -1599 8223 -1597
rect 8205 -1651 8217 -1599
rect 8199 -1653 8223 -1651
rect 8279 -1653 8297 -1597
rect 8126 -1662 8297 -1653
rect 8325 -1599 8377 -1551
rect 8325 -1657 8377 -1651
rect 8405 -1597 8736 -1588
rect 8405 -1599 8422 -1597
rect 8478 -1599 8502 -1597
rect 8558 -1599 8582 -1597
rect 8638 -1599 8662 -1597
rect 8718 -1599 8736 -1597
rect 8405 -1651 8416 -1599
rect 8478 -1651 8480 -1599
rect 8660 -1651 8662 -1599
rect 8724 -1651 8736 -1599
rect 8405 -1653 8422 -1651
rect 8478 -1653 8502 -1651
rect 8558 -1653 8582 -1651
rect 8638 -1653 8662 -1651
rect 8718 -1653 8736 -1651
rect 8405 -1662 8736 -1653
rect 8806 -1597 9137 -1588
rect 8806 -1599 8823 -1597
rect 8879 -1599 8903 -1597
rect 8959 -1599 8983 -1597
rect 9039 -1599 9063 -1597
rect 9119 -1599 9137 -1597
rect 8806 -1651 8817 -1599
rect 8879 -1651 8881 -1599
rect 9061 -1651 9063 -1599
rect 9125 -1651 9137 -1599
rect 8806 -1653 8823 -1651
rect 8879 -1653 8903 -1651
rect 8959 -1653 8983 -1651
rect 9039 -1653 9063 -1651
rect 9119 -1653 9137 -1651
rect 8806 -1662 9137 -1653
rect 9165 -1599 9217 -1551
rect 9165 -1657 9217 -1651
rect 9245 -1597 9416 -1588
rect 9245 -1653 9262 -1597
rect 9318 -1599 9342 -1597
rect 9324 -1651 9336 -1599
rect 9318 -1653 9342 -1651
rect 9398 -1653 9416 -1597
rect 9245 -1662 9416 -1653
rect 8040 -1751 8812 -1699
rect 8864 -1751 8870 -1699
rect 9165 -1751 9440 -1699
rect 8040 -1799 8092 -1751
rect 8040 -1857 8092 -1851
rect 8126 -1797 8297 -1788
rect 8126 -1853 8143 -1797
rect 8199 -1799 8223 -1797
rect 8205 -1851 8217 -1799
rect 8199 -1853 8223 -1851
rect 8279 -1853 8297 -1797
rect 8126 -1862 8297 -1853
rect 8325 -1799 8377 -1751
rect 8325 -1857 8377 -1851
rect 8405 -1797 8736 -1788
rect 8405 -1799 8422 -1797
rect 8478 -1799 8502 -1797
rect 8558 -1799 8582 -1797
rect 8638 -1799 8662 -1797
rect 8718 -1799 8736 -1797
rect 8405 -1851 8416 -1799
rect 8478 -1851 8480 -1799
rect 8660 -1851 8662 -1799
rect 8724 -1851 8736 -1799
rect 8405 -1853 8422 -1851
rect 8478 -1853 8502 -1851
rect 8558 -1853 8582 -1851
rect 8638 -1853 8662 -1851
rect 8718 -1853 8736 -1851
rect 8405 -1862 8736 -1853
rect 8806 -1797 9137 -1788
rect 8806 -1799 8823 -1797
rect 8879 -1799 8903 -1797
rect 8959 -1799 8983 -1797
rect 9039 -1799 9063 -1797
rect 9119 -1799 9137 -1797
rect 8806 -1851 8817 -1799
rect 8879 -1851 8881 -1799
rect 9061 -1851 9063 -1799
rect 9125 -1851 9137 -1799
rect 8806 -1853 8823 -1851
rect 8879 -1853 8903 -1851
rect 8959 -1853 8983 -1851
rect 9039 -1853 9063 -1851
rect 9119 -1853 9137 -1851
rect 8806 -1862 9137 -1853
rect 9165 -1799 9217 -1751
rect 9165 -1857 9217 -1851
rect 9245 -1797 9416 -1788
rect 9245 -1853 9262 -1797
rect 9318 -1799 9342 -1797
rect 9324 -1851 9336 -1799
rect 9318 -1853 9342 -1851
rect 9398 -1853 9416 -1797
rect 9245 -1862 9416 -1853
<< via2 >>
rect 7 9883 63 9885
rect 7 9831 9 9883
rect 9 9831 61 9883
rect 61 9831 63 9883
rect 7 9829 63 9831
rect 207 9899 263 9901
rect 207 9847 209 9899
rect 209 9847 261 9899
rect 261 9847 263 9899
rect 207 9845 263 9847
rect 407 9883 463 9885
rect 407 9831 409 9883
rect 409 9831 461 9883
rect 461 9831 463 9883
rect 407 9829 463 9831
rect 607 9899 663 9901
rect 607 9847 609 9899
rect 609 9847 661 9899
rect 661 9847 663 9899
rect 607 9845 663 9847
rect 807 9883 863 9885
rect 807 9831 809 9883
rect 809 9831 861 9883
rect 861 9831 863 9883
rect 807 9829 863 9831
rect 1007 9899 1063 9901
rect 1007 9847 1009 9899
rect 1009 9847 1061 9899
rect 1061 9847 1063 9899
rect 1007 9845 1063 9847
rect 1207 9883 1263 9885
rect 1207 9831 1209 9883
rect 1209 9831 1261 9883
rect 1261 9831 1263 9883
rect 1207 9829 1263 9831
rect 1407 9899 1463 9901
rect 1407 9847 1409 9899
rect 1409 9847 1461 9899
rect 1461 9847 1463 9899
rect 1407 9845 1463 9847
rect 1607 9883 1663 9885
rect 1607 9831 1609 9883
rect 1609 9831 1661 9883
rect 1661 9831 1663 9883
rect 1607 9829 1663 9831
rect 1807 9899 1863 9901
rect 1807 9847 1809 9899
rect 1809 9847 1861 9899
rect 1861 9847 1863 9899
rect 1807 9845 1863 9847
rect 2007 9883 2063 9885
rect 2007 9831 2009 9883
rect 2009 9831 2061 9883
rect 2061 9831 2063 9883
rect 2007 9829 2063 9831
rect 2207 9899 2263 9901
rect 2207 9847 2209 9899
rect 2209 9847 2261 9899
rect 2261 9847 2263 9899
rect 2207 9845 2263 9847
rect 2407 9883 2463 9885
rect 2407 9831 2409 9883
rect 2409 9831 2461 9883
rect 2461 9831 2463 9883
rect 2407 9829 2463 9831
rect 2607 9899 2663 9901
rect 2607 9847 2609 9899
rect 2609 9847 2661 9899
rect 2661 9847 2663 9899
rect 2607 9845 2663 9847
rect 2807 9883 2863 9885
rect 2807 9831 2809 9883
rect 2809 9831 2861 9883
rect 2861 9831 2863 9883
rect 2807 9829 2863 9831
rect 3007 9899 3063 9901
rect 3007 9847 3009 9899
rect 3009 9847 3061 9899
rect 3061 9847 3063 9899
rect 3007 9845 3063 9847
rect 3207 9883 3263 9885
rect 3207 9831 3209 9883
rect 3209 9831 3261 9883
rect 3261 9831 3263 9883
rect 3207 9829 3263 9831
rect 3407 9899 3463 9901
rect 3407 9847 3409 9899
rect 3409 9847 3461 9899
rect 3461 9847 3463 9899
rect 3407 9845 3463 9847
rect 3607 9883 3663 9885
rect 3607 9831 3609 9883
rect 3609 9831 3661 9883
rect 3661 9831 3663 9883
rect 3607 9829 3663 9831
rect 3807 9899 3863 9901
rect 3807 9847 3809 9899
rect 3809 9847 3861 9899
rect 3861 9847 3863 9899
rect 3807 9845 3863 9847
rect 4007 9883 4063 9885
rect 4007 9831 4009 9883
rect 4009 9831 4061 9883
rect 4061 9831 4063 9883
rect 4007 9829 4063 9831
rect 4207 9899 4263 9901
rect 4207 9847 4209 9899
rect 4209 9847 4261 9899
rect 4261 9847 4263 9899
rect 4207 9845 4263 9847
rect 4407 9883 4463 9885
rect 4407 9831 4409 9883
rect 4409 9831 4461 9883
rect 4461 9831 4463 9883
rect 4407 9829 4463 9831
rect 4607 9899 4663 9901
rect 4607 9847 4609 9899
rect 4609 9847 4661 9899
rect 4661 9847 4663 9899
rect 4607 9845 4663 9847
rect 4807 9883 4863 9885
rect 4807 9831 4809 9883
rect 4809 9831 4861 9883
rect 4861 9831 4863 9883
rect 4807 9829 4863 9831
rect 5007 9899 5063 9901
rect 5007 9847 5009 9899
rect 5009 9847 5061 9899
rect 5061 9847 5063 9899
rect 5007 9845 5063 9847
rect 5207 9883 5263 9885
rect 5207 9831 5209 9883
rect 5209 9831 5261 9883
rect 5261 9831 5263 9883
rect 5207 9829 5263 9831
rect 5407 9899 5463 9901
rect 5407 9847 5409 9899
rect 5409 9847 5461 9899
rect 5461 9847 5463 9899
rect 5407 9845 5463 9847
rect 5607 9883 5663 9885
rect 5607 9831 5609 9883
rect 5609 9831 5661 9883
rect 5661 9831 5663 9883
rect 5607 9829 5663 9831
rect 5807 9899 5863 9901
rect 5807 9847 5809 9899
rect 5809 9847 5861 9899
rect 5861 9847 5863 9899
rect 5807 9845 5863 9847
rect 6007 9883 6063 9885
rect 6007 9831 6009 9883
rect 6009 9831 6061 9883
rect 6061 9831 6063 9883
rect 6007 9829 6063 9831
rect 6207 9899 6263 9901
rect 6207 9847 6209 9899
rect 6209 9847 6261 9899
rect 6261 9847 6263 9899
rect 6207 9845 6263 9847
rect 7 8673 63 8675
rect 7 8621 9 8673
rect 9 8621 61 8673
rect 61 8621 63 8673
rect 7 8619 63 8621
rect 207 8689 263 8691
rect 207 8637 209 8689
rect 209 8637 261 8689
rect 261 8637 263 8689
rect 207 8635 263 8637
rect 407 8673 463 8675
rect 407 8621 409 8673
rect 409 8621 461 8673
rect 461 8621 463 8673
rect 407 8619 463 8621
rect 607 8689 663 8691
rect 607 8637 609 8689
rect 609 8637 661 8689
rect 661 8637 663 8689
rect 607 8635 663 8637
rect 807 8673 863 8675
rect 807 8621 809 8673
rect 809 8621 861 8673
rect 861 8621 863 8673
rect 807 8619 863 8621
rect 1007 8689 1063 8691
rect 1007 8637 1009 8689
rect 1009 8637 1061 8689
rect 1061 8637 1063 8689
rect 1007 8635 1063 8637
rect 1207 8673 1263 8675
rect 1207 8621 1209 8673
rect 1209 8621 1261 8673
rect 1261 8621 1263 8673
rect 1207 8619 1263 8621
rect 1407 8689 1463 8691
rect 1407 8637 1409 8689
rect 1409 8637 1461 8689
rect 1461 8637 1463 8689
rect 1407 8635 1463 8637
rect 1607 8673 1663 8675
rect 1607 8621 1609 8673
rect 1609 8621 1661 8673
rect 1661 8621 1663 8673
rect 1607 8619 1663 8621
rect 1807 8689 1863 8691
rect 1807 8637 1809 8689
rect 1809 8637 1861 8689
rect 1861 8637 1863 8689
rect 1807 8635 1863 8637
rect 2007 8673 2063 8675
rect 2007 8621 2009 8673
rect 2009 8621 2061 8673
rect 2061 8621 2063 8673
rect 2007 8619 2063 8621
rect 2207 8689 2263 8691
rect 2207 8637 2209 8689
rect 2209 8637 2261 8689
rect 2261 8637 2263 8689
rect 2207 8635 2263 8637
rect 2407 8673 2463 8675
rect 2407 8621 2409 8673
rect 2409 8621 2461 8673
rect 2461 8621 2463 8673
rect 2407 8619 2463 8621
rect 2607 8689 2663 8691
rect 2607 8637 2609 8689
rect 2609 8637 2661 8689
rect 2661 8637 2663 8689
rect 2607 8635 2663 8637
rect 2807 8673 2863 8675
rect 2807 8621 2809 8673
rect 2809 8621 2861 8673
rect 2861 8621 2863 8673
rect 2807 8619 2863 8621
rect 3007 8689 3063 8691
rect 3007 8637 3009 8689
rect 3009 8637 3061 8689
rect 3061 8637 3063 8689
rect 3007 8635 3063 8637
rect 3207 8673 3263 8675
rect 3207 8621 3209 8673
rect 3209 8621 3261 8673
rect 3261 8621 3263 8673
rect 3207 8619 3263 8621
rect 3407 8689 3463 8691
rect 3407 8637 3409 8689
rect 3409 8637 3461 8689
rect 3461 8637 3463 8689
rect 3407 8635 3463 8637
rect 3607 8673 3663 8675
rect 3607 8621 3609 8673
rect 3609 8621 3661 8673
rect 3661 8621 3663 8673
rect 3607 8619 3663 8621
rect 3807 8689 3863 8691
rect 3807 8637 3809 8689
rect 3809 8637 3861 8689
rect 3861 8637 3863 8689
rect 3807 8635 3863 8637
rect 4007 8673 4063 8675
rect 4007 8621 4009 8673
rect 4009 8621 4061 8673
rect 4061 8621 4063 8673
rect 4007 8619 4063 8621
rect 4207 8689 4263 8691
rect 4207 8637 4209 8689
rect 4209 8637 4261 8689
rect 4261 8637 4263 8689
rect 4207 8635 4263 8637
rect 4407 8673 4463 8675
rect 4407 8621 4409 8673
rect 4409 8621 4461 8673
rect 4461 8621 4463 8673
rect 4407 8619 4463 8621
rect 4607 8689 4663 8691
rect 4607 8637 4609 8689
rect 4609 8637 4661 8689
rect 4661 8637 4663 8689
rect 4607 8635 4663 8637
rect 4807 8673 4863 8675
rect 4807 8621 4809 8673
rect 4809 8621 4861 8673
rect 4861 8621 4863 8673
rect 4807 8619 4863 8621
rect 5007 8689 5063 8691
rect 5007 8637 5009 8689
rect 5009 8637 5061 8689
rect 5061 8637 5063 8689
rect 5007 8635 5063 8637
rect 5207 8673 5263 8675
rect 5207 8621 5209 8673
rect 5209 8621 5261 8673
rect 5261 8621 5263 8673
rect 5207 8619 5263 8621
rect 5407 8689 5463 8691
rect 5407 8637 5409 8689
rect 5409 8637 5461 8689
rect 5461 8637 5463 8689
rect 5407 8635 5463 8637
rect 5607 8673 5663 8675
rect 5607 8621 5609 8673
rect 5609 8621 5661 8673
rect 5661 8621 5663 8673
rect 5607 8619 5663 8621
rect 5807 8689 5863 8691
rect 5807 8637 5809 8689
rect 5809 8637 5861 8689
rect 5861 8637 5863 8689
rect 5807 8635 5863 8637
rect 6007 8673 6063 8675
rect 6007 8621 6009 8673
rect 6009 8621 6061 8673
rect 6061 8621 6063 8673
rect 6007 8619 6063 8621
rect 6207 8689 6263 8691
rect 6207 8637 6209 8689
rect 6209 8637 6261 8689
rect 6261 8637 6263 8689
rect 6207 8635 6263 8637
rect 7 7463 63 7465
rect 7 7411 9 7463
rect 9 7411 61 7463
rect 61 7411 63 7463
rect 7 7409 63 7411
rect 207 7479 263 7481
rect 207 7427 209 7479
rect 209 7427 261 7479
rect 261 7427 263 7479
rect 207 7425 263 7427
rect 407 7463 463 7465
rect 407 7411 409 7463
rect 409 7411 461 7463
rect 461 7411 463 7463
rect 407 7409 463 7411
rect 607 7479 663 7481
rect 607 7427 609 7479
rect 609 7427 661 7479
rect 661 7427 663 7479
rect 607 7425 663 7427
rect 807 7463 863 7465
rect 807 7411 809 7463
rect 809 7411 861 7463
rect 861 7411 863 7463
rect 807 7409 863 7411
rect 1007 7479 1063 7481
rect 1007 7427 1009 7479
rect 1009 7427 1061 7479
rect 1061 7427 1063 7479
rect 1007 7425 1063 7427
rect 1207 7463 1263 7465
rect 1207 7411 1209 7463
rect 1209 7411 1261 7463
rect 1261 7411 1263 7463
rect 1207 7409 1263 7411
rect 1407 7479 1463 7481
rect 1407 7427 1409 7479
rect 1409 7427 1461 7479
rect 1461 7427 1463 7479
rect 1407 7425 1463 7427
rect 1607 7463 1663 7465
rect 1607 7411 1609 7463
rect 1609 7411 1661 7463
rect 1661 7411 1663 7463
rect 1607 7409 1663 7411
rect 1807 7479 1863 7481
rect 1807 7427 1809 7479
rect 1809 7427 1861 7479
rect 1861 7427 1863 7479
rect 1807 7425 1863 7427
rect 2007 7463 2063 7465
rect 2007 7411 2009 7463
rect 2009 7411 2061 7463
rect 2061 7411 2063 7463
rect 2007 7409 2063 7411
rect 2207 7479 2263 7481
rect 2207 7427 2209 7479
rect 2209 7427 2261 7479
rect 2261 7427 2263 7479
rect 2207 7425 2263 7427
rect 2407 7463 2463 7465
rect 2407 7411 2409 7463
rect 2409 7411 2461 7463
rect 2461 7411 2463 7463
rect 2407 7409 2463 7411
rect 2607 7479 2663 7481
rect 2607 7427 2609 7479
rect 2609 7427 2661 7479
rect 2661 7427 2663 7479
rect 2607 7425 2663 7427
rect 2807 7463 2863 7465
rect 2807 7411 2809 7463
rect 2809 7411 2861 7463
rect 2861 7411 2863 7463
rect 2807 7409 2863 7411
rect 3007 7479 3063 7481
rect 3007 7427 3009 7479
rect 3009 7427 3061 7479
rect 3061 7427 3063 7479
rect 3007 7425 3063 7427
rect 3207 7463 3263 7465
rect 3207 7411 3209 7463
rect 3209 7411 3261 7463
rect 3261 7411 3263 7463
rect 3207 7409 3263 7411
rect 3407 7479 3463 7481
rect 3407 7427 3409 7479
rect 3409 7427 3461 7479
rect 3461 7427 3463 7479
rect 3407 7425 3463 7427
rect 3607 7463 3663 7465
rect 3607 7411 3609 7463
rect 3609 7411 3661 7463
rect 3661 7411 3663 7463
rect 3607 7409 3663 7411
rect 3807 7479 3863 7481
rect 3807 7427 3809 7479
rect 3809 7427 3861 7479
rect 3861 7427 3863 7479
rect 3807 7425 3863 7427
rect 4007 7463 4063 7465
rect 4007 7411 4009 7463
rect 4009 7411 4061 7463
rect 4061 7411 4063 7463
rect 4007 7409 4063 7411
rect 4207 7479 4263 7481
rect 4207 7427 4209 7479
rect 4209 7427 4261 7479
rect 4261 7427 4263 7479
rect 4207 7425 4263 7427
rect 4407 7463 4463 7465
rect 4407 7411 4409 7463
rect 4409 7411 4461 7463
rect 4461 7411 4463 7463
rect 4407 7409 4463 7411
rect 4607 7479 4663 7481
rect 4607 7427 4609 7479
rect 4609 7427 4661 7479
rect 4661 7427 4663 7479
rect 4607 7425 4663 7427
rect 4807 7463 4863 7465
rect 4807 7411 4809 7463
rect 4809 7411 4861 7463
rect 4861 7411 4863 7463
rect 4807 7409 4863 7411
rect 5007 7479 5063 7481
rect 5007 7427 5009 7479
rect 5009 7427 5061 7479
rect 5061 7427 5063 7479
rect 5007 7425 5063 7427
rect 5207 7463 5263 7465
rect 5207 7411 5209 7463
rect 5209 7411 5261 7463
rect 5261 7411 5263 7463
rect 5207 7409 5263 7411
rect 5407 7479 5463 7481
rect 5407 7427 5409 7479
rect 5409 7427 5461 7479
rect 5461 7427 5463 7479
rect 5407 7425 5463 7427
rect 5607 7463 5663 7465
rect 5607 7411 5609 7463
rect 5609 7411 5661 7463
rect 5661 7411 5663 7463
rect 5607 7409 5663 7411
rect 5807 7479 5863 7481
rect 5807 7427 5809 7479
rect 5809 7427 5861 7479
rect 5861 7427 5863 7479
rect 5807 7425 5863 7427
rect 6007 7463 6063 7465
rect 6007 7411 6009 7463
rect 6009 7411 6061 7463
rect 6061 7411 6063 7463
rect 6007 7409 6063 7411
rect 6207 7479 6263 7481
rect 6207 7427 6209 7479
rect 6209 7427 6261 7479
rect 6261 7427 6263 7479
rect 6207 7425 6263 7427
rect 7 6253 63 6255
rect 7 6201 9 6253
rect 9 6201 61 6253
rect 61 6201 63 6253
rect 7 6199 63 6201
rect 207 6269 263 6271
rect 207 6217 209 6269
rect 209 6217 261 6269
rect 261 6217 263 6269
rect 207 6215 263 6217
rect 407 6253 463 6255
rect 407 6201 409 6253
rect 409 6201 461 6253
rect 461 6201 463 6253
rect 407 6199 463 6201
rect 607 6269 663 6271
rect 607 6217 609 6269
rect 609 6217 661 6269
rect 661 6217 663 6269
rect 607 6215 663 6217
rect 807 6253 863 6255
rect 807 6201 809 6253
rect 809 6201 861 6253
rect 861 6201 863 6253
rect 807 6199 863 6201
rect 1007 6269 1063 6271
rect 1007 6217 1009 6269
rect 1009 6217 1061 6269
rect 1061 6217 1063 6269
rect 1007 6215 1063 6217
rect 1207 6253 1263 6255
rect 1207 6201 1209 6253
rect 1209 6201 1261 6253
rect 1261 6201 1263 6253
rect 1207 6199 1263 6201
rect 1407 6269 1463 6271
rect 1407 6217 1409 6269
rect 1409 6217 1461 6269
rect 1461 6217 1463 6269
rect 1407 6215 1463 6217
rect 1607 6253 1663 6255
rect 1607 6201 1609 6253
rect 1609 6201 1661 6253
rect 1661 6201 1663 6253
rect 1607 6199 1663 6201
rect 1807 6269 1863 6271
rect 1807 6217 1809 6269
rect 1809 6217 1861 6269
rect 1861 6217 1863 6269
rect 1807 6215 1863 6217
rect 2007 6253 2063 6255
rect 2007 6201 2009 6253
rect 2009 6201 2061 6253
rect 2061 6201 2063 6253
rect 2007 6199 2063 6201
rect 2207 6269 2263 6271
rect 2207 6217 2209 6269
rect 2209 6217 2261 6269
rect 2261 6217 2263 6269
rect 2207 6215 2263 6217
rect 2407 6253 2463 6255
rect 2407 6201 2409 6253
rect 2409 6201 2461 6253
rect 2461 6201 2463 6253
rect 2407 6199 2463 6201
rect 2607 6269 2663 6271
rect 2607 6217 2609 6269
rect 2609 6217 2661 6269
rect 2661 6217 2663 6269
rect 2607 6215 2663 6217
rect 2807 6253 2863 6255
rect 2807 6201 2809 6253
rect 2809 6201 2861 6253
rect 2861 6201 2863 6253
rect 2807 6199 2863 6201
rect 3007 6269 3063 6271
rect 3007 6217 3009 6269
rect 3009 6217 3061 6269
rect 3061 6217 3063 6269
rect 3007 6215 3063 6217
rect 3207 6253 3263 6255
rect 3207 6201 3209 6253
rect 3209 6201 3261 6253
rect 3261 6201 3263 6253
rect 3207 6199 3263 6201
rect 3407 6269 3463 6271
rect 3407 6217 3409 6269
rect 3409 6217 3461 6269
rect 3461 6217 3463 6269
rect 3407 6215 3463 6217
rect 3607 6253 3663 6255
rect 3607 6201 3609 6253
rect 3609 6201 3661 6253
rect 3661 6201 3663 6253
rect 3607 6199 3663 6201
rect 3807 6269 3863 6271
rect 3807 6217 3809 6269
rect 3809 6217 3861 6269
rect 3861 6217 3863 6269
rect 3807 6215 3863 6217
rect 4007 6253 4063 6255
rect 4007 6201 4009 6253
rect 4009 6201 4061 6253
rect 4061 6201 4063 6253
rect 4007 6199 4063 6201
rect 4207 6269 4263 6271
rect 4207 6217 4209 6269
rect 4209 6217 4261 6269
rect 4261 6217 4263 6269
rect 4207 6215 4263 6217
rect 4407 6253 4463 6255
rect 4407 6201 4409 6253
rect 4409 6201 4461 6253
rect 4461 6201 4463 6253
rect 4407 6199 4463 6201
rect 4607 6269 4663 6271
rect 4607 6217 4609 6269
rect 4609 6217 4661 6269
rect 4661 6217 4663 6269
rect 4607 6215 4663 6217
rect 4807 6253 4863 6255
rect 4807 6201 4809 6253
rect 4809 6201 4861 6253
rect 4861 6201 4863 6253
rect 4807 6199 4863 6201
rect 5007 6269 5063 6271
rect 5007 6217 5009 6269
rect 5009 6217 5061 6269
rect 5061 6217 5063 6269
rect 5007 6215 5063 6217
rect 5207 6253 5263 6255
rect 5207 6201 5209 6253
rect 5209 6201 5261 6253
rect 5261 6201 5263 6253
rect 5207 6199 5263 6201
rect 5407 6269 5463 6271
rect 5407 6217 5409 6269
rect 5409 6217 5461 6269
rect 5461 6217 5463 6269
rect 5407 6215 5463 6217
rect 5607 6253 5663 6255
rect 5607 6201 5609 6253
rect 5609 6201 5661 6253
rect 5661 6201 5663 6253
rect 5607 6199 5663 6201
rect 5807 6269 5863 6271
rect 5807 6217 5809 6269
rect 5809 6217 5861 6269
rect 5861 6217 5863 6269
rect 5807 6215 5863 6217
rect 6007 6253 6063 6255
rect 6007 6201 6009 6253
rect 6009 6201 6061 6253
rect 6061 6201 6063 6253
rect 6007 6199 6063 6201
rect 6207 6269 6263 6271
rect 6207 6217 6209 6269
rect 6209 6217 6261 6269
rect 6261 6217 6263 6269
rect 6207 6215 6263 6217
rect 7 4903 63 4905
rect 7 4851 9 4903
rect 9 4851 61 4903
rect 61 4851 63 4903
rect 7 4849 63 4851
rect 207 4919 263 4921
rect 207 4867 209 4919
rect 209 4867 261 4919
rect 261 4867 263 4919
rect 207 4865 263 4867
rect 407 4903 463 4905
rect 407 4851 409 4903
rect 409 4851 461 4903
rect 461 4851 463 4903
rect 407 4849 463 4851
rect 607 4919 663 4921
rect 607 4867 609 4919
rect 609 4867 661 4919
rect 661 4867 663 4919
rect 607 4865 663 4867
rect 807 4903 863 4905
rect 807 4851 809 4903
rect 809 4851 861 4903
rect 861 4851 863 4903
rect 807 4849 863 4851
rect 1007 4919 1063 4921
rect 1007 4867 1009 4919
rect 1009 4867 1061 4919
rect 1061 4867 1063 4919
rect 1007 4865 1063 4867
rect 1207 4903 1263 4905
rect 1207 4851 1209 4903
rect 1209 4851 1261 4903
rect 1261 4851 1263 4903
rect 1207 4849 1263 4851
rect 1407 4919 1463 4921
rect 1407 4867 1409 4919
rect 1409 4867 1461 4919
rect 1461 4867 1463 4919
rect 1407 4865 1463 4867
rect 1607 4903 1663 4905
rect 1607 4851 1609 4903
rect 1609 4851 1661 4903
rect 1661 4851 1663 4903
rect 1607 4849 1663 4851
rect 1807 4919 1863 4921
rect 1807 4867 1809 4919
rect 1809 4867 1861 4919
rect 1861 4867 1863 4919
rect 1807 4865 1863 4867
rect 2007 4903 2063 4905
rect 2007 4851 2009 4903
rect 2009 4851 2061 4903
rect 2061 4851 2063 4903
rect 2007 4849 2063 4851
rect 2207 4919 2263 4921
rect 2207 4867 2209 4919
rect 2209 4867 2261 4919
rect 2261 4867 2263 4919
rect 2207 4865 2263 4867
rect 2407 4903 2463 4905
rect 2407 4851 2409 4903
rect 2409 4851 2461 4903
rect 2461 4851 2463 4903
rect 2407 4849 2463 4851
rect 2607 4919 2663 4921
rect 2607 4867 2609 4919
rect 2609 4867 2661 4919
rect 2661 4867 2663 4919
rect 2607 4865 2663 4867
rect 2807 4903 2863 4905
rect 2807 4851 2809 4903
rect 2809 4851 2861 4903
rect 2861 4851 2863 4903
rect 2807 4849 2863 4851
rect 3007 4919 3063 4921
rect 3007 4867 3009 4919
rect 3009 4867 3061 4919
rect 3061 4867 3063 4919
rect 3007 4865 3063 4867
rect 3207 4903 3263 4905
rect 3207 4851 3209 4903
rect 3209 4851 3261 4903
rect 3261 4851 3263 4903
rect 3207 4849 3263 4851
rect 3407 4919 3463 4921
rect 3407 4867 3409 4919
rect 3409 4867 3461 4919
rect 3461 4867 3463 4919
rect 3407 4865 3463 4867
rect 3607 4903 3663 4905
rect 3607 4851 3609 4903
rect 3609 4851 3661 4903
rect 3661 4851 3663 4903
rect 3607 4849 3663 4851
rect 3807 4919 3863 4921
rect 3807 4867 3809 4919
rect 3809 4867 3861 4919
rect 3861 4867 3863 4919
rect 3807 4865 3863 4867
rect 4007 4903 4063 4905
rect 4007 4851 4009 4903
rect 4009 4851 4061 4903
rect 4061 4851 4063 4903
rect 4007 4849 4063 4851
rect 4207 4919 4263 4921
rect 4207 4867 4209 4919
rect 4209 4867 4261 4919
rect 4261 4867 4263 4919
rect 4207 4865 4263 4867
rect 4407 4903 4463 4905
rect 4407 4851 4409 4903
rect 4409 4851 4461 4903
rect 4461 4851 4463 4903
rect 4407 4849 4463 4851
rect 4607 4919 4663 4921
rect 4607 4867 4609 4919
rect 4609 4867 4661 4919
rect 4661 4867 4663 4919
rect 4607 4865 4663 4867
rect 4807 4903 4863 4905
rect 4807 4851 4809 4903
rect 4809 4851 4861 4903
rect 4861 4851 4863 4903
rect 4807 4849 4863 4851
rect 5007 4919 5063 4921
rect 5007 4867 5009 4919
rect 5009 4867 5061 4919
rect 5061 4867 5063 4919
rect 5007 4865 5063 4867
rect 5207 4903 5263 4905
rect 5207 4851 5209 4903
rect 5209 4851 5261 4903
rect 5261 4851 5263 4903
rect 5207 4849 5263 4851
rect 5407 4919 5463 4921
rect 5407 4867 5409 4919
rect 5409 4867 5461 4919
rect 5461 4867 5463 4919
rect 5407 4865 5463 4867
rect 5607 4903 5663 4905
rect 5607 4851 5609 4903
rect 5609 4851 5661 4903
rect 5661 4851 5663 4903
rect 5607 4849 5663 4851
rect 5807 4919 5863 4921
rect 5807 4867 5809 4919
rect 5809 4867 5861 4919
rect 5861 4867 5863 4919
rect 5807 4865 5863 4867
rect 6007 4903 6063 4905
rect 6007 4851 6009 4903
rect 6009 4851 6061 4903
rect 6061 4851 6063 4903
rect 6007 4849 6063 4851
rect 6207 4919 6263 4921
rect 6207 4867 6209 4919
rect 6209 4867 6261 4919
rect 6261 4867 6263 4919
rect 6207 4865 6263 4867
rect 7 3693 63 3695
rect 7 3641 9 3693
rect 9 3641 61 3693
rect 61 3641 63 3693
rect 7 3639 63 3641
rect 207 3709 263 3711
rect 207 3657 209 3709
rect 209 3657 261 3709
rect 261 3657 263 3709
rect 207 3655 263 3657
rect 407 3693 463 3695
rect 407 3641 409 3693
rect 409 3641 461 3693
rect 461 3641 463 3693
rect 407 3639 463 3641
rect 607 3709 663 3711
rect 607 3657 609 3709
rect 609 3657 661 3709
rect 661 3657 663 3709
rect 607 3655 663 3657
rect 807 3693 863 3695
rect 807 3641 809 3693
rect 809 3641 861 3693
rect 861 3641 863 3693
rect 807 3639 863 3641
rect 1007 3709 1063 3711
rect 1007 3657 1009 3709
rect 1009 3657 1061 3709
rect 1061 3657 1063 3709
rect 1007 3655 1063 3657
rect 1207 3693 1263 3695
rect 1207 3641 1209 3693
rect 1209 3641 1261 3693
rect 1261 3641 1263 3693
rect 1207 3639 1263 3641
rect 1407 3709 1463 3711
rect 1407 3657 1409 3709
rect 1409 3657 1461 3709
rect 1461 3657 1463 3709
rect 1407 3655 1463 3657
rect 1607 3693 1663 3695
rect 1607 3641 1609 3693
rect 1609 3641 1661 3693
rect 1661 3641 1663 3693
rect 1607 3639 1663 3641
rect 1807 3709 1863 3711
rect 1807 3657 1809 3709
rect 1809 3657 1861 3709
rect 1861 3657 1863 3709
rect 1807 3655 1863 3657
rect 2007 3693 2063 3695
rect 2007 3641 2009 3693
rect 2009 3641 2061 3693
rect 2061 3641 2063 3693
rect 2007 3639 2063 3641
rect 2207 3709 2263 3711
rect 2207 3657 2209 3709
rect 2209 3657 2261 3709
rect 2261 3657 2263 3709
rect 2207 3655 2263 3657
rect 2407 3693 2463 3695
rect 2407 3641 2409 3693
rect 2409 3641 2461 3693
rect 2461 3641 2463 3693
rect 2407 3639 2463 3641
rect 2607 3709 2663 3711
rect 2607 3657 2609 3709
rect 2609 3657 2661 3709
rect 2661 3657 2663 3709
rect 2607 3655 2663 3657
rect 2807 3693 2863 3695
rect 2807 3641 2809 3693
rect 2809 3641 2861 3693
rect 2861 3641 2863 3693
rect 2807 3639 2863 3641
rect 3007 3709 3063 3711
rect 3007 3657 3009 3709
rect 3009 3657 3061 3709
rect 3061 3657 3063 3709
rect 3007 3655 3063 3657
rect 3207 3693 3263 3695
rect 3207 3641 3209 3693
rect 3209 3641 3261 3693
rect 3261 3641 3263 3693
rect 3207 3639 3263 3641
rect 3407 3709 3463 3711
rect 3407 3657 3409 3709
rect 3409 3657 3461 3709
rect 3461 3657 3463 3709
rect 3407 3655 3463 3657
rect 3607 3693 3663 3695
rect 3607 3641 3609 3693
rect 3609 3641 3661 3693
rect 3661 3641 3663 3693
rect 3607 3639 3663 3641
rect 3807 3709 3863 3711
rect 3807 3657 3809 3709
rect 3809 3657 3861 3709
rect 3861 3657 3863 3709
rect 3807 3655 3863 3657
rect 4007 3693 4063 3695
rect 4007 3641 4009 3693
rect 4009 3641 4061 3693
rect 4061 3641 4063 3693
rect 4007 3639 4063 3641
rect 4207 3709 4263 3711
rect 4207 3657 4209 3709
rect 4209 3657 4261 3709
rect 4261 3657 4263 3709
rect 4207 3655 4263 3657
rect 4407 3693 4463 3695
rect 4407 3641 4409 3693
rect 4409 3641 4461 3693
rect 4461 3641 4463 3693
rect 4407 3639 4463 3641
rect 4607 3709 4663 3711
rect 4607 3657 4609 3709
rect 4609 3657 4661 3709
rect 4661 3657 4663 3709
rect 4607 3655 4663 3657
rect 4807 3693 4863 3695
rect 4807 3641 4809 3693
rect 4809 3641 4861 3693
rect 4861 3641 4863 3693
rect 4807 3639 4863 3641
rect 5007 3709 5063 3711
rect 5007 3657 5009 3709
rect 5009 3657 5061 3709
rect 5061 3657 5063 3709
rect 5007 3655 5063 3657
rect 5207 3693 5263 3695
rect 5207 3641 5209 3693
rect 5209 3641 5261 3693
rect 5261 3641 5263 3693
rect 5207 3639 5263 3641
rect 5407 3709 5463 3711
rect 5407 3657 5409 3709
rect 5409 3657 5461 3709
rect 5461 3657 5463 3709
rect 5407 3655 5463 3657
rect 5607 3693 5663 3695
rect 5607 3641 5609 3693
rect 5609 3641 5661 3693
rect 5661 3641 5663 3693
rect 5607 3639 5663 3641
rect 5807 3709 5863 3711
rect 5807 3657 5809 3709
rect 5809 3657 5861 3709
rect 5861 3657 5863 3709
rect 5807 3655 5863 3657
rect 6007 3693 6063 3695
rect 6007 3641 6009 3693
rect 6009 3641 6061 3693
rect 6061 3641 6063 3693
rect 6007 3639 6063 3641
rect 6207 3709 6263 3711
rect 6207 3657 6209 3709
rect 6209 3657 6261 3709
rect 6261 3657 6263 3709
rect 6207 3655 6263 3657
rect 7 2483 63 2485
rect 7 2431 9 2483
rect 9 2431 61 2483
rect 61 2431 63 2483
rect 7 2429 63 2431
rect 207 2499 263 2501
rect 207 2447 209 2499
rect 209 2447 261 2499
rect 261 2447 263 2499
rect 207 2445 263 2447
rect 407 2483 463 2485
rect 407 2431 409 2483
rect 409 2431 461 2483
rect 461 2431 463 2483
rect 407 2429 463 2431
rect 607 2499 663 2501
rect 607 2447 609 2499
rect 609 2447 661 2499
rect 661 2447 663 2499
rect 607 2445 663 2447
rect 807 2483 863 2485
rect 807 2431 809 2483
rect 809 2431 861 2483
rect 861 2431 863 2483
rect 807 2429 863 2431
rect 1007 2499 1063 2501
rect 1007 2447 1009 2499
rect 1009 2447 1061 2499
rect 1061 2447 1063 2499
rect 1007 2445 1063 2447
rect 1207 2483 1263 2485
rect 1207 2431 1209 2483
rect 1209 2431 1261 2483
rect 1261 2431 1263 2483
rect 1207 2429 1263 2431
rect 1407 2499 1463 2501
rect 1407 2447 1409 2499
rect 1409 2447 1461 2499
rect 1461 2447 1463 2499
rect 1407 2445 1463 2447
rect 1607 2483 1663 2485
rect 1607 2431 1609 2483
rect 1609 2431 1661 2483
rect 1661 2431 1663 2483
rect 1607 2429 1663 2431
rect 1807 2499 1863 2501
rect 1807 2447 1809 2499
rect 1809 2447 1861 2499
rect 1861 2447 1863 2499
rect 1807 2445 1863 2447
rect 2007 2483 2063 2485
rect 2007 2431 2009 2483
rect 2009 2431 2061 2483
rect 2061 2431 2063 2483
rect 2007 2429 2063 2431
rect 2207 2499 2263 2501
rect 2207 2447 2209 2499
rect 2209 2447 2261 2499
rect 2261 2447 2263 2499
rect 2207 2445 2263 2447
rect 2407 2483 2463 2485
rect 2407 2431 2409 2483
rect 2409 2431 2461 2483
rect 2461 2431 2463 2483
rect 2407 2429 2463 2431
rect 2607 2499 2663 2501
rect 2607 2447 2609 2499
rect 2609 2447 2661 2499
rect 2661 2447 2663 2499
rect 2607 2445 2663 2447
rect 2807 2483 2863 2485
rect 2807 2431 2809 2483
rect 2809 2431 2861 2483
rect 2861 2431 2863 2483
rect 2807 2429 2863 2431
rect 3007 2499 3063 2501
rect 3007 2447 3009 2499
rect 3009 2447 3061 2499
rect 3061 2447 3063 2499
rect 3007 2445 3063 2447
rect 3207 2483 3263 2485
rect 3207 2431 3209 2483
rect 3209 2431 3261 2483
rect 3261 2431 3263 2483
rect 3207 2429 3263 2431
rect 3407 2499 3463 2501
rect 3407 2447 3409 2499
rect 3409 2447 3461 2499
rect 3461 2447 3463 2499
rect 3407 2445 3463 2447
rect 3607 2483 3663 2485
rect 3607 2431 3609 2483
rect 3609 2431 3661 2483
rect 3661 2431 3663 2483
rect 3607 2429 3663 2431
rect 3807 2499 3863 2501
rect 3807 2447 3809 2499
rect 3809 2447 3861 2499
rect 3861 2447 3863 2499
rect 3807 2445 3863 2447
rect 4007 2483 4063 2485
rect 4007 2431 4009 2483
rect 4009 2431 4061 2483
rect 4061 2431 4063 2483
rect 4007 2429 4063 2431
rect 4207 2499 4263 2501
rect 4207 2447 4209 2499
rect 4209 2447 4261 2499
rect 4261 2447 4263 2499
rect 4207 2445 4263 2447
rect 4407 2483 4463 2485
rect 4407 2431 4409 2483
rect 4409 2431 4461 2483
rect 4461 2431 4463 2483
rect 4407 2429 4463 2431
rect 4607 2499 4663 2501
rect 4607 2447 4609 2499
rect 4609 2447 4661 2499
rect 4661 2447 4663 2499
rect 4607 2445 4663 2447
rect 4807 2483 4863 2485
rect 4807 2431 4809 2483
rect 4809 2431 4861 2483
rect 4861 2431 4863 2483
rect 4807 2429 4863 2431
rect 5007 2499 5063 2501
rect 5007 2447 5009 2499
rect 5009 2447 5061 2499
rect 5061 2447 5063 2499
rect 5007 2445 5063 2447
rect 5207 2483 5263 2485
rect 5207 2431 5209 2483
rect 5209 2431 5261 2483
rect 5261 2431 5263 2483
rect 5207 2429 5263 2431
rect 5407 2499 5463 2501
rect 5407 2447 5409 2499
rect 5409 2447 5461 2499
rect 5461 2447 5463 2499
rect 5407 2445 5463 2447
rect 5607 2483 5663 2485
rect 5607 2431 5609 2483
rect 5609 2431 5661 2483
rect 5661 2431 5663 2483
rect 5607 2429 5663 2431
rect 5807 2499 5863 2501
rect 5807 2447 5809 2499
rect 5809 2447 5861 2499
rect 5861 2447 5863 2499
rect 5807 2445 5863 2447
rect 6007 2483 6063 2485
rect 6007 2431 6009 2483
rect 6009 2431 6061 2483
rect 6061 2431 6063 2483
rect 6007 2429 6063 2431
rect 6207 2499 6263 2501
rect 6207 2447 6209 2499
rect 6209 2447 6261 2499
rect 6261 2447 6263 2499
rect 6207 2445 6263 2447
rect 7 1273 63 1275
rect 7 1221 9 1273
rect 9 1221 61 1273
rect 61 1221 63 1273
rect 7 1219 63 1221
rect 207 1289 263 1291
rect 207 1237 209 1289
rect 209 1237 261 1289
rect 261 1237 263 1289
rect 207 1235 263 1237
rect 407 1273 463 1275
rect 407 1221 409 1273
rect 409 1221 461 1273
rect 461 1221 463 1273
rect 407 1219 463 1221
rect 607 1289 663 1291
rect 607 1237 609 1289
rect 609 1237 661 1289
rect 661 1237 663 1289
rect 607 1235 663 1237
rect 807 1273 863 1275
rect 807 1221 809 1273
rect 809 1221 861 1273
rect 861 1221 863 1273
rect 807 1219 863 1221
rect 1007 1289 1063 1291
rect 1007 1237 1009 1289
rect 1009 1237 1061 1289
rect 1061 1237 1063 1289
rect 1007 1235 1063 1237
rect 1207 1273 1263 1275
rect 1207 1221 1209 1273
rect 1209 1221 1261 1273
rect 1261 1221 1263 1273
rect 1207 1219 1263 1221
rect 1407 1289 1463 1291
rect 1407 1237 1409 1289
rect 1409 1237 1461 1289
rect 1461 1237 1463 1289
rect 1407 1235 1463 1237
rect 1607 1273 1663 1275
rect 1607 1221 1609 1273
rect 1609 1221 1661 1273
rect 1661 1221 1663 1273
rect 1607 1219 1663 1221
rect 1807 1289 1863 1291
rect 1807 1237 1809 1289
rect 1809 1237 1861 1289
rect 1861 1237 1863 1289
rect 1807 1235 1863 1237
rect 2007 1273 2063 1275
rect 2007 1221 2009 1273
rect 2009 1221 2061 1273
rect 2061 1221 2063 1273
rect 2007 1219 2063 1221
rect 2207 1289 2263 1291
rect 2207 1237 2209 1289
rect 2209 1237 2261 1289
rect 2261 1237 2263 1289
rect 2207 1235 2263 1237
rect 2407 1273 2463 1275
rect 2407 1221 2409 1273
rect 2409 1221 2461 1273
rect 2461 1221 2463 1273
rect 2407 1219 2463 1221
rect 2607 1289 2663 1291
rect 2607 1237 2609 1289
rect 2609 1237 2661 1289
rect 2661 1237 2663 1289
rect 2607 1235 2663 1237
rect 2807 1273 2863 1275
rect 2807 1221 2809 1273
rect 2809 1221 2861 1273
rect 2861 1221 2863 1273
rect 2807 1219 2863 1221
rect 3007 1289 3063 1291
rect 3007 1237 3009 1289
rect 3009 1237 3061 1289
rect 3061 1237 3063 1289
rect 3007 1235 3063 1237
rect 3207 1273 3263 1275
rect 3207 1221 3209 1273
rect 3209 1221 3261 1273
rect 3261 1221 3263 1273
rect 3207 1219 3263 1221
rect 3407 1289 3463 1291
rect 3407 1237 3409 1289
rect 3409 1237 3461 1289
rect 3461 1237 3463 1289
rect 3407 1235 3463 1237
rect 3607 1273 3663 1275
rect 3607 1221 3609 1273
rect 3609 1221 3661 1273
rect 3661 1221 3663 1273
rect 3607 1219 3663 1221
rect 3807 1289 3863 1291
rect 3807 1237 3809 1289
rect 3809 1237 3861 1289
rect 3861 1237 3863 1289
rect 3807 1235 3863 1237
rect 4007 1273 4063 1275
rect 4007 1221 4009 1273
rect 4009 1221 4061 1273
rect 4061 1221 4063 1273
rect 4007 1219 4063 1221
rect 4207 1289 4263 1291
rect 4207 1237 4209 1289
rect 4209 1237 4261 1289
rect 4261 1237 4263 1289
rect 4207 1235 4263 1237
rect 4407 1273 4463 1275
rect 4407 1221 4409 1273
rect 4409 1221 4461 1273
rect 4461 1221 4463 1273
rect 4407 1219 4463 1221
rect 4607 1289 4663 1291
rect 4607 1237 4609 1289
rect 4609 1237 4661 1289
rect 4661 1237 4663 1289
rect 4607 1235 4663 1237
rect 4807 1273 4863 1275
rect 4807 1221 4809 1273
rect 4809 1221 4861 1273
rect 4861 1221 4863 1273
rect 4807 1219 4863 1221
rect 5007 1289 5063 1291
rect 5007 1237 5009 1289
rect 5009 1237 5061 1289
rect 5061 1237 5063 1289
rect 5007 1235 5063 1237
rect 5207 1273 5263 1275
rect 5207 1221 5209 1273
rect 5209 1221 5261 1273
rect 5261 1221 5263 1273
rect 5207 1219 5263 1221
rect 5407 1289 5463 1291
rect 5407 1237 5409 1289
rect 5409 1237 5461 1289
rect 5461 1237 5463 1289
rect 5407 1235 5463 1237
rect 5607 1273 5663 1275
rect 5607 1221 5609 1273
rect 5609 1221 5661 1273
rect 5661 1221 5663 1273
rect 5607 1219 5663 1221
rect 5807 1289 5863 1291
rect 5807 1237 5809 1289
rect 5809 1237 5861 1289
rect 5861 1237 5863 1289
rect 5807 1235 5863 1237
rect 6007 1273 6063 1275
rect 6007 1221 6009 1273
rect 6009 1221 6061 1273
rect 6061 1221 6063 1273
rect 6007 1219 6063 1221
rect 6207 1289 6263 1291
rect 6207 1237 6209 1289
rect 6209 1237 6261 1289
rect 6261 1237 6263 1289
rect 6207 1235 6263 1237
rect 7 63 63 65
rect 7 11 9 63
rect 9 11 61 63
rect 61 11 63 63
rect 7 9 63 11
rect 207 79 263 81
rect 207 27 209 79
rect 209 27 261 79
rect 261 27 263 79
rect 207 25 263 27
rect 7 -22 63 -16
rect 7 -72 9 -22
rect 9 -72 61 -22
rect 61 -72 63 -22
rect 407 63 463 65
rect 407 11 409 63
rect 409 11 461 63
rect 461 11 463 63
rect 407 9 463 11
rect 607 79 663 81
rect 607 27 609 79
rect 609 27 661 79
rect 661 27 663 79
rect 607 25 663 27
rect 207 -22 263 -16
rect 207 -72 209 -22
rect 209 -72 261 -22
rect 261 -72 263 -22
rect 407 -22 463 -16
rect 407 -72 409 -22
rect 409 -72 461 -22
rect 461 -72 463 -22
rect 807 63 863 65
rect 807 11 809 63
rect 809 11 861 63
rect 861 11 863 63
rect 807 9 863 11
rect 1007 79 1063 81
rect 1007 27 1009 79
rect 1009 27 1061 79
rect 1061 27 1063 79
rect 1007 25 1063 27
rect 607 -22 663 -16
rect 607 -72 609 -22
rect 609 -72 661 -22
rect 661 -72 663 -22
rect 807 -22 863 -16
rect 807 -72 809 -22
rect 809 -72 861 -22
rect 861 -72 863 -22
rect 1207 63 1263 65
rect 1207 11 1209 63
rect 1209 11 1261 63
rect 1261 11 1263 63
rect 1207 9 1263 11
rect 1407 79 1463 81
rect 1407 27 1409 79
rect 1409 27 1461 79
rect 1461 27 1463 79
rect 1407 25 1463 27
rect 1007 -22 1063 -16
rect 1007 -72 1009 -22
rect 1009 -72 1061 -22
rect 1061 -72 1063 -22
rect 1207 -22 1263 -16
rect 1207 -72 1209 -22
rect 1209 -72 1261 -22
rect 1261 -72 1263 -22
rect 1607 63 1663 65
rect 1607 11 1609 63
rect 1609 11 1661 63
rect 1661 11 1663 63
rect 1607 9 1663 11
rect 1807 79 1863 81
rect 1807 27 1809 79
rect 1809 27 1861 79
rect 1861 27 1863 79
rect 1807 25 1863 27
rect 1407 -22 1463 -16
rect 1407 -72 1409 -22
rect 1409 -72 1461 -22
rect 1461 -72 1463 -22
rect 1607 -22 1663 -16
rect 1607 -72 1609 -22
rect 1609 -72 1661 -22
rect 1661 -72 1663 -22
rect 2007 63 2063 65
rect 2007 11 2009 63
rect 2009 11 2061 63
rect 2061 11 2063 63
rect 2007 9 2063 11
rect 2207 79 2263 81
rect 2207 27 2209 79
rect 2209 27 2261 79
rect 2261 27 2263 79
rect 2207 25 2263 27
rect 1807 -22 1863 -16
rect 1807 -72 1809 -22
rect 1809 -72 1861 -22
rect 1861 -72 1863 -22
rect 2007 -22 2063 -16
rect 2007 -72 2009 -22
rect 2009 -72 2061 -22
rect 2061 -72 2063 -22
rect 2407 63 2463 65
rect 2407 11 2409 63
rect 2409 11 2461 63
rect 2461 11 2463 63
rect 2407 9 2463 11
rect 2607 79 2663 81
rect 2607 27 2609 79
rect 2609 27 2661 79
rect 2661 27 2663 79
rect 2607 25 2663 27
rect 2207 -22 2263 -16
rect 2207 -72 2209 -22
rect 2209 -72 2261 -22
rect 2261 -72 2263 -22
rect 2407 -22 2463 -16
rect 2407 -72 2409 -22
rect 2409 -72 2461 -22
rect 2461 -72 2463 -22
rect 2807 63 2863 65
rect 2807 11 2809 63
rect 2809 11 2861 63
rect 2861 11 2863 63
rect 2807 9 2863 11
rect 3007 79 3063 81
rect 3007 27 3009 79
rect 3009 27 3061 79
rect 3061 27 3063 79
rect 3007 25 3063 27
rect 2607 -22 2663 -16
rect 2607 -72 2609 -22
rect 2609 -72 2661 -22
rect 2661 -72 2663 -22
rect 2807 -22 2863 -16
rect 2807 -72 2809 -22
rect 2809 -72 2861 -22
rect 2861 -72 2863 -22
rect 3207 63 3263 65
rect 3207 11 3209 63
rect 3209 11 3261 63
rect 3261 11 3263 63
rect 3207 9 3263 11
rect 3407 79 3463 81
rect 3407 27 3409 79
rect 3409 27 3461 79
rect 3461 27 3463 79
rect 3407 25 3463 27
rect 3007 -22 3063 -16
rect 3007 -72 3009 -22
rect 3009 -72 3061 -22
rect 3061 -72 3063 -22
rect 3207 -22 3263 -16
rect 3207 -72 3209 -22
rect 3209 -72 3261 -22
rect 3261 -72 3263 -22
rect 3607 63 3663 65
rect 3607 11 3609 63
rect 3609 11 3661 63
rect 3661 11 3663 63
rect 3607 9 3663 11
rect 3807 79 3863 81
rect 3807 27 3809 79
rect 3809 27 3861 79
rect 3861 27 3863 79
rect 3807 25 3863 27
rect 3407 -22 3463 -16
rect 3407 -72 3409 -22
rect 3409 -72 3461 -22
rect 3461 -72 3463 -22
rect 3607 -22 3663 -16
rect 3607 -72 3609 -22
rect 3609 -72 3661 -22
rect 3661 -72 3663 -22
rect 4007 63 4063 65
rect 4007 11 4009 63
rect 4009 11 4061 63
rect 4061 11 4063 63
rect 4007 9 4063 11
rect 4207 79 4263 81
rect 4207 27 4209 79
rect 4209 27 4261 79
rect 4261 27 4263 79
rect 4207 25 4263 27
rect 3807 -22 3863 -16
rect 3807 -72 3809 -22
rect 3809 -72 3861 -22
rect 3861 -72 3863 -22
rect 4007 -22 4063 -16
rect 4007 -72 4009 -22
rect 4009 -72 4061 -22
rect 4061 -72 4063 -22
rect 4407 63 4463 65
rect 4407 11 4409 63
rect 4409 11 4461 63
rect 4461 11 4463 63
rect 4407 9 4463 11
rect 4607 79 4663 81
rect 4607 27 4609 79
rect 4609 27 4661 79
rect 4661 27 4663 79
rect 4607 25 4663 27
rect 4207 -22 4263 -16
rect 4207 -72 4209 -22
rect 4209 -72 4261 -22
rect 4261 -72 4263 -22
rect 4407 -22 4463 -16
rect 4407 -72 4409 -22
rect 4409 -72 4461 -22
rect 4461 -72 4463 -22
rect 4807 63 4863 65
rect 4807 11 4809 63
rect 4809 11 4861 63
rect 4861 11 4863 63
rect 4807 9 4863 11
rect 5007 79 5063 81
rect 5007 27 5009 79
rect 5009 27 5061 79
rect 5061 27 5063 79
rect 5007 25 5063 27
rect 4607 -22 4663 -16
rect 4607 -72 4609 -22
rect 4609 -72 4661 -22
rect 4661 -72 4663 -22
rect 4807 -22 4863 -16
rect 4807 -72 4809 -22
rect 4809 -72 4861 -22
rect 4861 -72 4863 -22
rect 5207 63 5263 65
rect 5207 11 5209 63
rect 5209 11 5261 63
rect 5261 11 5263 63
rect 5207 9 5263 11
rect 5407 79 5463 81
rect 5407 27 5409 79
rect 5409 27 5461 79
rect 5461 27 5463 79
rect 5407 25 5463 27
rect 5007 -22 5063 -16
rect 5007 -72 5009 -22
rect 5009 -72 5061 -22
rect 5061 -72 5063 -22
rect 5207 -22 5263 -16
rect 5207 -72 5209 -22
rect 5209 -72 5261 -22
rect 5261 -72 5263 -22
rect 5607 63 5663 65
rect 5607 11 5609 63
rect 5609 11 5661 63
rect 5661 11 5663 63
rect 5607 9 5663 11
rect 5807 79 5863 81
rect 5807 27 5809 79
rect 5809 27 5861 79
rect 5861 27 5863 79
rect 5807 25 5863 27
rect 5407 -22 5463 -16
rect 5407 -72 5409 -22
rect 5409 -72 5461 -22
rect 5461 -72 5463 -22
rect 5607 -22 5663 -16
rect 5607 -72 5609 -22
rect 5609 -72 5661 -22
rect 5661 -72 5663 -22
rect 6007 63 6063 65
rect 6007 11 6009 63
rect 6009 11 6061 63
rect 6061 11 6063 63
rect 6007 9 6063 11
rect 6207 79 6263 81
rect 6207 27 6209 79
rect 6209 27 6261 79
rect 6261 27 6263 79
rect 6207 25 6263 27
rect 5807 -22 5863 -16
rect 5807 -72 5809 -22
rect 5809 -72 5861 -22
rect 5861 -72 5863 -22
rect 6007 -22 6063 -16
rect 6007 -72 6009 -22
rect 6009 -72 6061 -22
rect 6061 -72 6063 -22
rect 6207 -22 6263 -16
rect 6207 -72 6209 -22
rect 6209 -72 6261 -22
rect 6261 -72 6263 -22
rect 8143 1 8199 3
rect 8223 1 8279 3
rect 8143 -51 8153 1
rect 8153 -51 8199 1
rect 8223 -51 8269 1
rect 8269 -51 8279 1
rect 8143 -53 8199 -51
rect 8223 -53 8279 -51
rect 8422 1 8478 3
rect 8502 1 8558 3
rect 8582 1 8638 3
rect 8662 1 8718 3
rect 8422 -51 8468 1
rect 8468 -51 8478 1
rect 8502 -51 8532 1
rect 8532 -51 8544 1
rect 8544 -51 8558 1
rect 8582 -51 8596 1
rect 8596 -51 8608 1
rect 8608 -51 8638 1
rect 8662 -51 8672 1
rect 8672 -51 8718 1
rect 8422 -53 8478 -51
rect 8502 -53 8558 -51
rect 8582 -53 8638 -51
rect 8662 -53 8718 -51
rect 8823 1 8879 3
rect 8903 1 8959 3
rect 8983 1 9039 3
rect 9063 1 9119 3
rect 8823 -51 8869 1
rect 8869 -51 8879 1
rect 8903 -51 8933 1
rect 8933 -51 8945 1
rect 8945 -51 8959 1
rect 8983 -51 8997 1
rect 8997 -51 9009 1
rect 9009 -51 9039 1
rect 9063 -51 9073 1
rect 9073 -51 9119 1
rect 8823 -53 8879 -51
rect 8903 -53 8959 -51
rect 8983 -53 9039 -51
rect 9063 -53 9119 -51
rect 9262 1 9318 3
rect 9342 1 9398 3
rect 9262 -51 9272 1
rect 9272 -51 9318 1
rect 9342 -51 9388 1
rect 9388 -51 9398 1
rect 9262 -53 9318 -51
rect 9342 -53 9398 -51
rect -133 -195 -91 -145
rect -91 -195 -77 -145
rect -53 -195 -39 -145
rect -39 -195 3 -145
rect -133 -201 -77 -195
rect -53 -201 3 -195
rect 67 -195 109 -145
rect 109 -195 123 -145
rect 147 -195 161 -145
rect 161 -195 203 -145
rect 67 -201 123 -195
rect 147 -201 203 -195
rect 267 -195 309 -145
rect 309 -195 323 -145
rect 347 -195 361 -145
rect 361 -195 403 -145
rect 267 -201 323 -195
rect 347 -201 403 -195
rect 467 -195 509 -145
rect 509 -195 523 -145
rect 547 -195 561 -145
rect 561 -195 603 -145
rect 467 -201 523 -195
rect 547 -201 603 -195
rect 667 -195 709 -145
rect 709 -195 723 -145
rect 747 -195 761 -145
rect 761 -195 803 -145
rect 667 -201 723 -195
rect 747 -201 803 -195
rect 867 -195 909 -145
rect 909 -195 923 -145
rect 947 -195 961 -145
rect 961 -195 1003 -145
rect 867 -201 923 -195
rect 947 -201 1003 -195
rect 1067 -195 1109 -145
rect 1109 -195 1123 -145
rect 1147 -195 1161 -145
rect 1161 -195 1203 -145
rect 1067 -201 1123 -195
rect 1147 -201 1203 -195
rect 1267 -195 1309 -145
rect 1309 -195 1323 -145
rect 1347 -195 1361 -145
rect 1361 -195 1403 -145
rect 1267 -201 1323 -195
rect 1347 -201 1403 -195
rect 1467 -195 1509 -145
rect 1509 -195 1523 -145
rect 1547 -195 1561 -145
rect 1561 -195 1603 -145
rect 1467 -201 1523 -195
rect 1547 -201 1603 -195
rect 1667 -195 1709 -145
rect 1709 -195 1723 -145
rect 1747 -195 1761 -145
rect 1761 -195 1803 -145
rect 1667 -201 1723 -195
rect 1747 -201 1803 -195
rect 1867 -195 1909 -145
rect 1909 -195 1923 -145
rect 1947 -195 1961 -145
rect 1961 -195 2003 -145
rect 1867 -201 1923 -195
rect 1947 -201 2003 -195
rect 2067 -195 2109 -145
rect 2109 -195 2123 -145
rect 2147 -195 2161 -145
rect 2161 -195 2203 -145
rect 2067 -201 2123 -195
rect 2147 -201 2203 -195
rect 2267 -195 2309 -145
rect 2309 -195 2323 -145
rect 2347 -195 2361 -145
rect 2361 -195 2403 -145
rect 2267 -201 2323 -195
rect 2347 -201 2403 -195
rect 2467 -195 2509 -145
rect 2509 -195 2523 -145
rect 2547 -195 2561 -145
rect 2561 -195 2603 -145
rect 2467 -201 2523 -195
rect 2547 -201 2603 -195
rect 2667 -195 2709 -145
rect 2709 -195 2723 -145
rect 2747 -195 2761 -145
rect 2761 -195 2803 -145
rect 2667 -201 2723 -195
rect 2747 -201 2803 -195
rect 2867 -195 2909 -145
rect 2909 -195 2923 -145
rect 2947 -195 2961 -145
rect 2961 -195 3003 -145
rect 2867 -201 2923 -195
rect 2947 -201 3003 -195
rect 3067 -195 3109 -145
rect 3109 -195 3123 -145
rect 3147 -195 3161 -145
rect 3161 -195 3203 -145
rect 3067 -201 3123 -195
rect 3147 -201 3203 -195
rect 3267 -195 3309 -145
rect 3309 -195 3323 -145
rect 3347 -195 3361 -145
rect 3361 -195 3403 -145
rect 3267 -201 3323 -195
rect 3347 -201 3403 -195
rect 3467 -195 3509 -145
rect 3509 -195 3523 -145
rect 3547 -195 3561 -145
rect 3561 -195 3603 -145
rect 3467 -201 3523 -195
rect 3547 -201 3603 -195
rect 3667 -195 3709 -145
rect 3709 -195 3723 -145
rect 3747 -195 3761 -145
rect 3761 -195 3803 -145
rect 3667 -201 3723 -195
rect 3747 -201 3803 -195
rect 3867 -195 3909 -145
rect 3909 -195 3923 -145
rect 3947 -195 3961 -145
rect 3961 -195 4003 -145
rect 3867 -201 3923 -195
rect 3947 -201 4003 -195
rect 4067 -195 4109 -145
rect 4109 -195 4123 -145
rect 4147 -195 4161 -145
rect 4161 -195 4203 -145
rect 4067 -201 4123 -195
rect 4147 -201 4203 -195
rect 4267 -195 4309 -145
rect 4309 -195 4323 -145
rect 4347 -195 4361 -145
rect 4361 -195 4403 -145
rect 4267 -201 4323 -195
rect 4347 -201 4403 -195
rect 4467 -195 4509 -145
rect 4509 -195 4523 -145
rect 4547 -195 4561 -145
rect 4561 -195 4603 -145
rect 4467 -201 4523 -195
rect 4547 -201 4603 -195
rect 4667 -195 4709 -145
rect 4709 -195 4723 -145
rect 4747 -195 4761 -145
rect 4761 -195 4803 -145
rect 4667 -201 4723 -195
rect 4747 -201 4803 -195
rect 4867 -195 4909 -145
rect 4909 -195 4923 -145
rect 4947 -195 4961 -145
rect 4961 -195 5003 -145
rect 4867 -201 4923 -195
rect 4947 -201 5003 -195
rect 5067 -195 5109 -145
rect 5109 -195 5123 -145
rect 5147 -195 5161 -145
rect 5161 -195 5203 -145
rect 5067 -201 5123 -195
rect 5147 -201 5203 -195
rect 5267 -195 5309 -145
rect 5309 -195 5323 -145
rect 5347 -195 5361 -145
rect 5361 -195 5403 -145
rect 5267 -201 5323 -195
rect 5347 -201 5403 -195
rect 5467 -195 5509 -145
rect 5509 -195 5523 -145
rect 5547 -195 5561 -145
rect 5561 -195 5603 -145
rect 5467 -201 5523 -195
rect 5547 -201 5603 -195
rect 5667 -195 5709 -145
rect 5709 -195 5723 -145
rect 5747 -195 5761 -145
rect 5761 -195 5803 -145
rect 5667 -201 5723 -195
rect 5747 -201 5803 -195
rect 5867 -195 5909 -145
rect 5909 -195 5923 -145
rect 5947 -195 5961 -145
rect 5961 -195 6003 -145
rect 5867 -201 5923 -195
rect 5947 -201 6003 -195
rect 6067 -195 6109 -145
rect 6109 -195 6123 -145
rect 6147 -195 6161 -145
rect 6161 -195 6203 -145
rect 6067 -201 6123 -195
rect 6147 -201 6203 -195
rect 6267 -195 6309 -145
rect 6309 -195 6323 -145
rect 6347 -195 6361 -145
rect 6361 -195 6403 -145
rect 6267 -201 6323 -195
rect 6347 -201 6403 -195
rect 8143 -199 8199 -197
rect 8223 -199 8279 -197
rect 8143 -251 8153 -199
rect 8153 -251 8199 -199
rect 8223 -251 8269 -199
rect 8269 -251 8279 -199
rect 8143 -253 8199 -251
rect 8223 -253 8279 -251
rect 8422 -199 8478 -197
rect 8502 -199 8558 -197
rect 8582 -199 8638 -197
rect 8662 -199 8718 -197
rect 8422 -251 8468 -199
rect 8468 -251 8478 -199
rect 8502 -251 8532 -199
rect 8532 -251 8544 -199
rect 8544 -251 8558 -199
rect 8582 -251 8596 -199
rect 8596 -251 8608 -199
rect 8608 -251 8638 -199
rect 8662 -251 8672 -199
rect 8672 -251 8718 -199
rect 8422 -253 8478 -251
rect 8502 -253 8558 -251
rect 8582 -253 8638 -251
rect 8662 -253 8718 -251
rect 8823 -199 8879 -197
rect 8903 -199 8959 -197
rect 8983 -199 9039 -197
rect 9063 -199 9119 -197
rect 8823 -251 8869 -199
rect 8869 -251 8879 -199
rect 8903 -251 8933 -199
rect 8933 -251 8945 -199
rect 8945 -251 8959 -199
rect 8983 -251 8997 -199
rect 8997 -251 9009 -199
rect 9009 -251 9039 -199
rect 9063 -251 9073 -199
rect 9073 -251 9119 -199
rect 8823 -253 8879 -251
rect 8903 -253 8959 -251
rect 8983 -253 9039 -251
rect 9063 -253 9119 -251
rect 9262 -199 9318 -197
rect 9342 -199 9398 -197
rect 9262 -251 9272 -199
rect 9272 -251 9318 -199
rect 9342 -251 9388 -199
rect 9388 -251 9398 -199
rect 9262 -253 9318 -251
rect 9342 -253 9398 -251
rect -93 -378 -91 -348
rect -91 -378 -39 -348
rect -39 -378 -37 -348
rect -93 -390 -37 -378
rect -93 -404 -91 -390
rect -91 -404 -39 -390
rect -39 -404 -37 -390
rect -93 -442 -91 -428
rect -91 -442 -39 -428
rect -39 -442 -37 -428
rect -93 -454 -37 -442
rect -93 -484 -91 -454
rect -91 -484 -39 -454
rect -39 -484 -37 -454
rect 107 -378 109 -348
rect 109 -378 161 -348
rect 161 -378 163 -348
rect 107 -390 163 -378
rect 107 -404 109 -390
rect 109 -404 161 -390
rect 161 -404 163 -390
rect 107 -442 109 -428
rect 109 -442 161 -428
rect 161 -442 163 -428
rect 107 -454 163 -442
rect 107 -484 109 -454
rect 109 -484 161 -454
rect 161 -484 163 -454
rect 307 -378 309 -348
rect 309 -378 361 -348
rect 361 -378 363 -348
rect 307 -390 363 -378
rect 307 -404 309 -390
rect 309 -404 361 -390
rect 361 -404 363 -390
rect 307 -442 309 -428
rect 309 -442 361 -428
rect 361 -442 363 -428
rect 307 -454 363 -442
rect 307 -484 309 -454
rect 309 -484 361 -454
rect 361 -484 363 -454
rect 507 -378 509 -348
rect 509 -378 561 -348
rect 561 -378 563 -348
rect 507 -390 563 -378
rect 507 -404 509 -390
rect 509 -404 561 -390
rect 561 -404 563 -390
rect 507 -442 509 -428
rect 509 -442 561 -428
rect 561 -442 563 -428
rect 507 -454 563 -442
rect 507 -484 509 -454
rect 509 -484 561 -454
rect 561 -484 563 -454
rect 707 -378 709 -348
rect 709 -378 761 -348
rect 761 -378 763 -348
rect 707 -390 763 -378
rect 707 -404 709 -390
rect 709 -404 761 -390
rect 761 -404 763 -390
rect 707 -442 709 -428
rect 709 -442 761 -428
rect 761 -442 763 -428
rect 707 -454 763 -442
rect 707 -484 709 -454
rect 709 -484 761 -454
rect 761 -484 763 -454
rect 907 -378 909 -348
rect 909 -378 961 -348
rect 961 -378 963 -348
rect 907 -390 963 -378
rect 907 -404 909 -390
rect 909 -404 961 -390
rect 961 -404 963 -390
rect 907 -442 909 -428
rect 909 -442 961 -428
rect 961 -442 963 -428
rect 907 -454 963 -442
rect 907 -484 909 -454
rect 909 -484 961 -454
rect 961 -484 963 -454
rect 1107 -378 1109 -348
rect 1109 -378 1161 -348
rect 1161 -378 1163 -348
rect 1107 -390 1163 -378
rect 1107 -404 1109 -390
rect 1109 -404 1161 -390
rect 1161 -404 1163 -390
rect 1107 -442 1109 -428
rect 1109 -442 1161 -428
rect 1161 -442 1163 -428
rect 1107 -454 1163 -442
rect 1107 -484 1109 -454
rect 1109 -484 1161 -454
rect 1161 -484 1163 -454
rect 1307 -378 1309 -348
rect 1309 -378 1361 -348
rect 1361 -378 1363 -348
rect 1307 -390 1363 -378
rect 1307 -404 1309 -390
rect 1309 -404 1361 -390
rect 1361 -404 1363 -390
rect 1307 -442 1309 -428
rect 1309 -442 1361 -428
rect 1361 -442 1363 -428
rect 1307 -454 1363 -442
rect 1307 -484 1309 -454
rect 1309 -484 1361 -454
rect 1361 -484 1363 -454
rect 1507 -378 1509 -348
rect 1509 -378 1561 -348
rect 1561 -378 1563 -348
rect 1507 -390 1563 -378
rect 1507 -404 1509 -390
rect 1509 -404 1561 -390
rect 1561 -404 1563 -390
rect 1507 -442 1509 -428
rect 1509 -442 1561 -428
rect 1561 -442 1563 -428
rect 1507 -454 1563 -442
rect 1507 -484 1509 -454
rect 1509 -484 1561 -454
rect 1561 -484 1563 -454
rect 1707 -378 1709 -348
rect 1709 -378 1761 -348
rect 1761 -378 1763 -348
rect 1707 -390 1763 -378
rect 1707 -404 1709 -390
rect 1709 -404 1761 -390
rect 1761 -404 1763 -390
rect 1707 -442 1709 -428
rect 1709 -442 1761 -428
rect 1761 -442 1763 -428
rect 1707 -454 1763 -442
rect 1707 -484 1709 -454
rect 1709 -484 1761 -454
rect 1761 -484 1763 -454
rect 1907 -378 1909 -348
rect 1909 -378 1961 -348
rect 1961 -378 1963 -348
rect 1907 -390 1963 -378
rect 1907 -404 1909 -390
rect 1909 -404 1961 -390
rect 1961 -404 1963 -390
rect 1907 -442 1909 -428
rect 1909 -442 1961 -428
rect 1961 -442 1963 -428
rect 1907 -454 1963 -442
rect 1907 -484 1909 -454
rect 1909 -484 1961 -454
rect 1961 -484 1963 -454
rect 2107 -378 2109 -348
rect 2109 -378 2161 -348
rect 2161 -378 2163 -348
rect 2107 -390 2163 -378
rect 2107 -404 2109 -390
rect 2109 -404 2161 -390
rect 2161 -404 2163 -390
rect 2107 -442 2109 -428
rect 2109 -442 2161 -428
rect 2161 -442 2163 -428
rect 2107 -454 2163 -442
rect 2107 -484 2109 -454
rect 2109 -484 2161 -454
rect 2161 -484 2163 -454
rect 2307 -378 2309 -348
rect 2309 -378 2361 -348
rect 2361 -378 2363 -348
rect 2307 -390 2363 -378
rect 2307 -404 2309 -390
rect 2309 -404 2361 -390
rect 2361 -404 2363 -390
rect 2307 -442 2309 -428
rect 2309 -442 2361 -428
rect 2361 -442 2363 -428
rect 2307 -454 2363 -442
rect 2307 -484 2309 -454
rect 2309 -484 2361 -454
rect 2361 -484 2363 -454
rect 2507 -378 2509 -348
rect 2509 -378 2561 -348
rect 2561 -378 2563 -348
rect 2507 -390 2563 -378
rect 2507 -404 2509 -390
rect 2509 -404 2561 -390
rect 2561 -404 2563 -390
rect 2507 -442 2509 -428
rect 2509 -442 2561 -428
rect 2561 -442 2563 -428
rect 2507 -454 2563 -442
rect 2507 -484 2509 -454
rect 2509 -484 2561 -454
rect 2561 -484 2563 -454
rect 2707 -378 2709 -348
rect 2709 -378 2761 -348
rect 2761 -378 2763 -348
rect 2707 -390 2763 -378
rect 2707 -404 2709 -390
rect 2709 -404 2761 -390
rect 2761 -404 2763 -390
rect 2707 -442 2709 -428
rect 2709 -442 2761 -428
rect 2761 -442 2763 -428
rect 2707 -454 2763 -442
rect 2707 -484 2709 -454
rect 2709 -484 2761 -454
rect 2761 -484 2763 -454
rect 2907 -378 2909 -348
rect 2909 -378 2961 -348
rect 2961 -378 2963 -348
rect 2907 -390 2963 -378
rect 2907 -404 2909 -390
rect 2909 -404 2961 -390
rect 2961 -404 2963 -390
rect 2907 -442 2909 -428
rect 2909 -442 2961 -428
rect 2961 -442 2963 -428
rect 2907 -454 2963 -442
rect 2907 -484 2909 -454
rect 2909 -484 2961 -454
rect 2961 -484 2963 -454
rect 3107 -378 3109 -348
rect 3109 -378 3161 -348
rect 3161 -378 3163 -348
rect 3107 -390 3163 -378
rect 3107 -404 3109 -390
rect 3109 -404 3161 -390
rect 3161 -404 3163 -390
rect 3107 -442 3109 -428
rect 3109 -442 3161 -428
rect 3161 -442 3163 -428
rect 3107 -454 3163 -442
rect 3107 -484 3109 -454
rect 3109 -484 3161 -454
rect 3161 -484 3163 -454
rect 3307 -378 3309 -348
rect 3309 -378 3361 -348
rect 3361 -378 3363 -348
rect 3307 -390 3363 -378
rect 3307 -404 3309 -390
rect 3309 -404 3361 -390
rect 3361 -404 3363 -390
rect 3307 -442 3309 -428
rect 3309 -442 3361 -428
rect 3361 -442 3363 -428
rect 3307 -454 3363 -442
rect 3307 -484 3309 -454
rect 3309 -484 3361 -454
rect 3361 -484 3363 -454
rect 3507 -378 3509 -348
rect 3509 -378 3561 -348
rect 3561 -378 3563 -348
rect 3507 -390 3563 -378
rect 3507 -404 3509 -390
rect 3509 -404 3561 -390
rect 3561 -404 3563 -390
rect 3507 -442 3509 -428
rect 3509 -442 3561 -428
rect 3561 -442 3563 -428
rect 3507 -454 3563 -442
rect 3507 -484 3509 -454
rect 3509 -484 3561 -454
rect 3561 -484 3563 -454
rect 3707 -378 3709 -348
rect 3709 -378 3761 -348
rect 3761 -378 3763 -348
rect 3707 -390 3763 -378
rect 3707 -404 3709 -390
rect 3709 -404 3761 -390
rect 3761 -404 3763 -390
rect 3707 -442 3709 -428
rect 3709 -442 3761 -428
rect 3761 -442 3763 -428
rect 3707 -454 3763 -442
rect 3707 -484 3709 -454
rect 3709 -484 3761 -454
rect 3761 -484 3763 -454
rect 3907 -378 3909 -348
rect 3909 -378 3961 -348
rect 3961 -378 3963 -348
rect 3907 -390 3963 -378
rect 3907 -404 3909 -390
rect 3909 -404 3961 -390
rect 3961 -404 3963 -390
rect 3907 -442 3909 -428
rect 3909 -442 3961 -428
rect 3961 -442 3963 -428
rect 3907 -454 3963 -442
rect 3907 -484 3909 -454
rect 3909 -484 3961 -454
rect 3961 -484 3963 -454
rect 4107 -378 4109 -348
rect 4109 -378 4161 -348
rect 4161 -378 4163 -348
rect 4107 -390 4163 -378
rect 4107 -404 4109 -390
rect 4109 -404 4161 -390
rect 4161 -404 4163 -390
rect 4107 -442 4109 -428
rect 4109 -442 4161 -428
rect 4161 -442 4163 -428
rect 4107 -454 4163 -442
rect 4107 -484 4109 -454
rect 4109 -484 4161 -454
rect 4161 -484 4163 -454
rect 4307 -378 4309 -348
rect 4309 -378 4361 -348
rect 4361 -378 4363 -348
rect 4307 -390 4363 -378
rect 4307 -404 4309 -390
rect 4309 -404 4361 -390
rect 4361 -404 4363 -390
rect 4307 -442 4309 -428
rect 4309 -442 4361 -428
rect 4361 -442 4363 -428
rect 4307 -454 4363 -442
rect 4307 -484 4309 -454
rect 4309 -484 4361 -454
rect 4361 -484 4363 -454
rect 4507 -378 4509 -348
rect 4509 -378 4561 -348
rect 4561 -378 4563 -348
rect 4507 -390 4563 -378
rect 4507 -404 4509 -390
rect 4509 -404 4561 -390
rect 4561 -404 4563 -390
rect 4507 -442 4509 -428
rect 4509 -442 4561 -428
rect 4561 -442 4563 -428
rect 4507 -454 4563 -442
rect 4507 -484 4509 -454
rect 4509 -484 4561 -454
rect 4561 -484 4563 -454
rect 4707 -378 4709 -348
rect 4709 -378 4761 -348
rect 4761 -378 4763 -348
rect 4707 -390 4763 -378
rect 4707 -404 4709 -390
rect 4709 -404 4761 -390
rect 4761 -404 4763 -390
rect 4707 -442 4709 -428
rect 4709 -442 4761 -428
rect 4761 -442 4763 -428
rect 4707 -454 4763 -442
rect 4707 -484 4709 -454
rect 4709 -484 4761 -454
rect 4761 -484 4763 -454
rect 4907 -378 4909 -348
rect 4909 -378 4961 -348
rect 4961 -378 4963 -348
rect 4907 -390 4963 -378
rect 4907 -404 4909 -390
rect 4909 -404 4961 -390
rect 4961 -404 4963 -390
rect 4907 -442 4909 -428
rect 4909 -442 4961 -428
rect 4961 -442 4963 -428
rect 4907 -454 4963 -442
rect 4907 -484 4909 -454
rect 4909 -484 4961 -454
rect 4961 -484 4963 -454
rect 5107 -378 5109 -348
rect 5109 -378 5161 -348
rect 5161 -378 5163 -348
rect 5107 -390 5163 -378
rect 5107 -404 5109 -390
rect 5109 -404 5161 -390
rect 5161 -404 5163 -390
rect 5107 -442 5109 -428
rect 5109 -442 5161 -428
rect 5161 -442 5163 -428
rect 5107 -454 5163 -442
rect 5107 -484 5109 -454
rect 5109 -484 5161 -454
rect 5161 -484 5163 -454
rect 5307 -378 5309 -348
rect 5309 -378 5361 -348
rect 5361 -378 5363 -348
rect 5307 -390 5363 -378
rect 5307 -404 5309 -390
rect 5309 -404 5361 -390
rect 5361 -404 5363 -390
rect 5307 -442 5309 -428
rect 5309 -442 5361 -428
rect 5361 -442 5363 -428
rect 5307 -454 5363 -442
rect 5307 -484 5309 -454
rect 5309 -484 5361 -454
rect 5361 -484 5363 -454
rect 5507 -378 5509 -348
rect 5509 -378 5561 -348
rect 5561 -378 5563 -348
rect 5507 -390 5563 -378
rect 5507 -404 5509 -390
rect 5509 -404 5561 -390
rect 5561 -404 5563 -390
rect 5507 -442 5509 -428
rect 5509 -442 5561 -428
rect 5561 -442 5563 -428
rect 5507 -454 5563 -442
rect 5507 -484 5509 -454
rect 5509 -484 5561 -454
rect 5561 -484 5563 -454
rect 5707 -378 5709 -348
rect 5709 -378 5761 -348
rect 5761 -378 5763 -348
rect 5707 -390 5763 -378
rect 5707 -404 5709 -390
rect 5709 -404 5761 -390
rect 5761 -404 5763 -390
rect 5707 -442 5709 -428
rect 5709 -442 5761 -428
rect 5761 -442 5763 -428
rect 5707 -454 5763 -442
rect 5707 -484 5709 -454
rect 5709 -484 5761 -454
rect 5761 -484 5763 -454
rect 5907 -378 5909 -348
rect 5909 -378 5961 -348
rect 5961 -378 5963 -348
rect 5907 -390 5963 -378
rect 5907 -404 5909 -390
rect 5909 -404 5961 -390
rect 5961 -404 5963 -390
rect 5907 -442 5909 -428
rect 5909 -442 5961 -428
rect 5961 -442 5963 -428
rect 5907 -454 5963 -442
rect 5907 -484 5909 -454
rect 5909 -484 5961 -454
rect 5961 -484 5963 -454
rect 6107 -378 6109 -348
rect 6109 -378 6161 -348
rect 6161 -378 6163 -348
rect 6107 -390 6163 -378
rect 6107 -404 6109 -390
rect 6109 -404 6161 -390
rect 6161 -404 6163 -390
rect 6107 -442 6109 -428
rect 6109 -442 6161 -428
rect 6161 -442 6163 -428
rect 6107 -454 6163 -442
rect 6107 -484 6109 -454
rect 6109 -484 6161 -454
rect 6161 -484 6163 -454
rect 6307 -378 6309 -348
rect 6309 -378 6361 -348
rect 6361 -378 6363 -348
rect 6307 -390 6363 -378
rect 6307 -404 6309 -390
rect 6309 -404 6361 -390
rect 6361 -404 6363 -390
rect 6307 -442 6309 -428
rect 6309 -442 6361 -428
rect 6361 -442 6363 -428
rect 6307 -454 6363 -442
rect 6307 -484 6309 -454
rect 6309 -484 6361 -454
rect 6361 -484 6363 -454
rect 8143 -399 8199 -397
rect 8223 -399 8279 -397
rect 8143 -451 8153 -399
rect 8153 -451 8199 -399
rect 8223 -451 8269 -399
rect 8269 -451 8279 -399
rect 8143 -453 8199 -451
rect 8223 -453 8279 -451
rect 8422 -399 8478 -397
rect 8502 -399 8558 -397
rect 8582 -399 8638 -397
rect 8662 -399 8718 -397
rect 8422 -451 8468 -399
rect 8468 -451 8478 -399
rect 8502 -451 8532 -399
rect 8532 -451 8544 -399
rect 8544 -451 8558 -399
rect 8582 -451 8596 -399
rect 8596 -451 8608 -399
rect 8608 -451 8638 -399
rect 8662 -451 8672 -399
rect 8672 -451 8718 -399
rect 8422 -453 8478 -451
rect 8502 -453 8558 -451
rect 8582 -453 8638 -451
rect 8662 -453 8718 -451
rect 8823 -399 8879 -397
rect 8903 -399 8959 -397
rect 8983 -399 9039 -397
rect 9063 -399 9119 -397
rect 8823 -451 8869 -399
rect 8869 -451 8879 -399
rect 8903 -451 8933 -399
rect 8933 -451 8945 -399
rect 8945 -451 8959 -399
rect 8983 -451 8997 -399
rect 8997 -451 9009 -399
rect 9009 -451 9039 -399
rect 9063 -451 9073 -399
rect 9073 -451 9119 -399
rect 8823 -453 8879 -451
rect 8903 -453 8959 -451
rect 8983 -453 9039 -451
rect 9063 -453 9119 -451
rect 9262 -399 9318 -397
rect 9342 -399 9398 -397
rect 9262 -451 9272 -399
rect 9272 -451 9318 -399
rect 9342 -451 9388 -399
rect 9388 -451 9398 -399
rect 9262 -453 9318 -451
rect 9342 -453 9398 -451
rect 8143 -599 8199 -597
rect 8223 -599 8279 -597
rect 8143 -651 8153 -599
rect 8153 -651 8199 -599
rect 8223 -651 8269 -599
rect 8269 -651 8279 -599
rect 8143 -653 8199 -651
rect 8223 -653 8279 -651
rect 8422 -599 8478 -597
rect 8502 -599 8558 -597
rect 8582 -599 8638 -597
rect 8662 -599 8718 -597
rect 8422 -651 8468 -599
rect 8468 -651 8478 -599
rect 8502 -651 8532 -599
rect 8532 -651 8544 -599
rect 8544 -651 8558 -599
rect 8582 -651 8596 -599
rect 8596 -651 8608 -599
rect 8608 -651 8638 -599
rect 8662 -651 8672 -599
rect 8672 -651 8718 -599
rect 8422 -653 8478 -651
rect 8502 -653 8558 -651
rect 8582 -653 8638 -651
rect 8662 -653 8718 -651
rect 8823 -599 8879 -597
rect 8903 -599 8959 -597
rect 8983 -599 9039 -597
rect 9063 -599 9119 -597
rect 8823 -651 8869 -599
rect 8869 -651 8879 -599
rect 8903 -651 8933 -599
rect 8933 -651 8945 -599
rect 8945 -651 8959 -599
rect 8983 -651 8997 -599
rect 8997 -651 9009 -599
rect 9009 -651 9039 -599
rect 9063 -651 9073 -599
rect 9073 -651 9119 -599
rect 8823 -653 8879 -651
rect 8903 -653 8959 -651
rect 8983 -653 9039 -651
rect 9063 -653 9119 -651
rect 9262 -599 9318 -597
rect 9342 -599 9398 -597
rect 9262 -651 9272 -599
rect 9272 -651 9318 -599
rect 9342 -651 9388 -599
rect 9388 -651 9398 -599
rect 9262 -653 9318 -651
rect 9342 -653 9398 -651
rect 8143 -799 8199 -797
rect 8223 -799 8279 -797
rect 8143 -851 8153 -799
rect 8153 -851 8199 -799
rect 8223 -851 8269 -799
rect 8269 -851 8279 -799
rect 8143 -853 8199 -851
rect 8223 -853 8279 -851
rect 8422 -799 8478 -797
rect 8502 -799 8558 -797
rect 8582 -799 8638 -797
rect 8662 -799 8718 -797
rect 8422 -851 8468 -799
rect 8468 -851 8478 -799
rect 8502 -851 8532 -799
rect 8532 -851 8544 -799
rect 8544 -851 8558 -799
rect 8582 -851 8596 -799
rect 8596 -851 8608 -799
rect 8608 -851 8638 -799
rect 8662 -851 8672 -799
rect 8672 -851 8718 -799
rect 8422 -853 8478 -851
rect 8502 -853 8558 -851
rect 8582 -853 8638 -851
rect 8662 -853 8718 -851
rect 8823 -799 8879 -797
rect 8903 -799 8959 -797
rect 8983 -799 9039 -797
rect 9063 -799 9119 -797
rect 8823 -851 8869 -799
rect 8869 -851 8879 -799
rect 8903 -851 8933 -799
rect 8933 -851 8945 -799
rect 8945 -851 8959 -799
rect 8983 -851 8997 -799
rect 8997 -851 9009 -799
rect 9009 -851 9039 -799
rect 9063 -851 9073 -799
rect 9073 -851 9119 -799
rect 8823 -853 8879 -851
rect 8903 -853 8959 -851
rect 8983 -853 9039 -851
rect 9063 -853 9119 -851
rect 9262 -799 9318 -797
rect 9342 -799 9398 -797
rect 9262 -851 9272 -799
rect 9272 -851 9318 -799
rect 9342 -851 9388 -799
rect 9388 -851 9398 -799
rect 9262 -853 9318 -851
rect 9342 -853 9398 -851
rect 8143 -999 8199 -997
rect 8223 -999 8279 -997
rect 8143 -1051 8153 -999
rect 8153 -1051 8199 -999
rect 8223 -1051 8269 -999
rect 8269 -1051 8279 -999
rect 8143 -1053 8199 -1051
rect 8223 -1053 8279 -1051
rect 8422 -999 8478 -997
rect 8502 -999 8558 -997
rect 8582 -999 8638 -997
rect 8662 -999 8718 -997
rect 8422 -1051 8468 -999
rect 8468 -1051 8478 -999
rect 8502 -1051 8532 -999
rect 8532 -1051 8544 -999
rect 8544 -1051 8558 -999
rect 8582 -1051 8596 -999
rect 8596 -1051 8608 -999
rect 8608 -1051 8638 -999
rect 8662 -1051 8672 -999
rect 8672 -1051 8718 -999
rect 8422 -1053 8478 -1051
rect 8502 -1053 8558 -1051
rect 8582 -1053 8638 -1051
rect 8662 -1053 8718 -1051
rect 8823 -999 8879 -997
rect 8903 -999 8959 -997
rect 8983 -999 9039 -997
rect 9063 -999 9119 -997
rect 8823 -1051 8869 -999
rect 8869 -1051 8879 -999
rect 8903 -1051 8933 -999
rect 8933 -1051 8945 -999
rect 8945 -1051 8959 -999
rect 8983 -1051 8997 -999
rect 8997 -1051 9009 -999
rect 9009 -1051 9039 -999
rect 9063 -1051 9073 -999
rect 9073 -1051 9119 -999
rect 8823 -1053 8879 -1051
rect 8903 -1053 8959 -1051
rect 8983 -1053 9039 -1051
rect 9063 -1053 9119 -1051
rect 9262 -999 9318 -997
rect 9342 -999 9398 -997
rect 9262 -1051 9272 -999
rect 9272 -1051 9318 -999
rect 9342 -1051 9388 -999
rect 9388 -1051 9398 -999
rect 9262 -1053 9318 -1051
rect 9342 -1053 9398 -1051
rect 8143 -1199 8199 -1197
rect 8223 -1199 8279 -1197
rect 8143 -1251 8153 -1199
rect 8153 -1251 8199 -1199
rect 8223 -1251 8269 -1199
rect 8269 -1251 8279 -1199
rect 8143 -1253 8199 -1251
rect 8223 -1253 8279 -1251
rect 8422 -1199 8478 -1197
rect 8502 -1199 8558 -1197
rect 8582 -1199 8638 -1197
rect 8662 -1199 8718 -1197
rect 8422 -1251 8468 -1199
rect 8468 -1251 8478 -1199
rect 8502 -1251 8532 -1199
rect 8532 -1251 8544 -1199
rect 8544 -1251 8558 -1199
rect 8582 -1251 8596 -1199
rect 8596 -1251 8608 -1199
rect 8608 -1251 8638 -1199
rect 8662 -1251 8672 -1199
rect 8672 -1251 8718 -1199
rect 8422 -1253 8478 -1251
rect 8502 -1253 8558 -1251
rect 8582 -1253 8638 -1251
rect 8662 -1253 8718 -1251
rect 8823 -1199 8879 -1197
rect 8903 -1199 8959 -1197
rect 8983 -1199 9039 -1197
rect 9063 -1199 9119 -1197
rect 8823 -1251 8869 -1199
rect 8869 -1251 8879 -1199
rect 8903 -1251 8933 -1199
rect 8933 -1251 8945 -1199
rect 8945 -1251 8959 -1199
rect 8983 -1251 8997 -1199
rect 8997 -1251 9009 -1199
rect 9009 -1251 9039 -1199
rect 9063 -1251 9073 -1199
rect 9073 -1251 9119 -1199
rect 8823 -1253 8879 -1251
rect 8903 -1253 8959 -1251
rect 8983 -1253 9039 -1251
rect 9063 -1253 9119 -1251
rect 9262 -1199 9318 -1197
rect 9342 -1199 9398 -1197
rect 9262 -1251 9272 -1199
rect 9272 -1251 9318 -1199
rect 9342 -1251 9388 -1199
rect 9388 -1251 9398 -1199
rect 9262 -1253 9318 -1251
rect 9342 -1253 9398 -1251
rect 8143 -1399 8199 -1397
rect 8223 -1399 8279 -1397
rect 8143 -1451 8153 -1399
rect 8153 -1451 8199 -1399
rect 8223 -1451 8269 -1399
rect 8269 -1451 8279 -1399
rect 8143 -1453 8199 -1451
rect 8223 -1453 8279 -1451
rect 8422 -1399 8478 -1397
rect 8502 -1399 8558 -1397
rect 8582 -1399 8638 -1397
rect 8662 -1399 8718 -1397
rect 8422 -1451 8468 -1399
rect 8468 -1451 8478 -1399
rect 8502 -1451 8532 -1399
rect 8532 -1451 8544 -1399
rect 8544 -1451 8558 -1399
rect 8582 -1451 8596 -1399
rect 8596 -1451 8608 -1399
rect 8608 -1451 8638 -1399
rect 8662 -1451 8672 -1399
rect 8672 -1451 8718 -1399
rect 8422 -1453 8478 -1451
rect 8502 -1453 8558 -1451
rect 8582 -1453 8638 -1451
rect 8662 -1453 8718 -1451
rect 8823 -1399 8879 -1397
rect 8903 -1399 8959 -1397
rect 8983 -1399 9039 -1397
rect 9063 -1399 9119 -1397
rect 8823 -1451 8869 -1399
rect 8869 -1451 8879 -1399
rect 8903 -1451 8933 -1399
rect 8933 -1451 8945 -1399
rect 8945 -1451 8959 -1399
rect 8983 -1451 8997 -1399
rect 8997 -1451 9009 -1399
rect 9009 -1451 9039 -1399
rect 9063 -1451 9073 -1399
rect 9073 -1451 9119 -1399
rect 8823 -1453 8879 -1451
rect 8903 -1453 8959 -1451
rect 8983 -1453 9039 -1451
rect 9063 -1453 9119 -1451
rect 9262 -1399 9318 -1397
rect 9342 -1399 9398 -1397
rect 9262 -1451 9272 -1399
rect 9272 -1451 9318 -1399
rect 9342 -1451 9388 -1399
rect 9388 -1451 9398 -1399
rect 9262 -1453 9318 -1451
rect 9342 -1453 9398 -1451
rect 8143 -1599 8199 -1597
rect 8223 -1599 8279 -1597
rect 8143 -1651 8153 -1599
rect 8153 -1651 8199 -1599
rect 8223 -1651 8269 -1599
rect 8269 -1651 8279 -1599
rect 8143 -1653 8199 -1651
rect 8223 -1653 8279 -1651
rect 8422 -1599 8478 -1597
rect 8502 -1599 8558 -1597
rect 8582 -1599 8638 -1597
rect 8662 -1599 8718 -1597
rect 8422 -1651 8468 -1599
rect 8468 -1651 8478 -1599
rect 8502 -1651 8532 -1599
rect 8532 -1651 8544 -1599
rect 8544 -1651 8558 -1599
rect 8582 -1651 8596 -1599
rect 8596 -1651 8608 -1599
rect 8608 -1651 8638 -1599
rect 8662 -1651 8672 -1599
rect 8672 -1651 8718 -1599
rect 8422 -1653 8478 -1651
rect 8502 -1653 8558 -1651
rect 8582 -1653 8638 -1651
rect 8662 -1653 8718 -1651
rect 8823 -1599 8879 -1597
rect 8903 -1599 8959 -1597
rect 8983 -1599 9039 -1597
rect 9063 -1599 9119 -1597
rect 8823 -1651 8869 -1599
rect 8869 -1651 8879 -1599
rect 8903 -1651 8933 -1599
rect 8933 -1651 8945 -1599
rect 8945 -1651 8959 -1599
rect 8983 -1651 8997 -1599
rect 8997 -1651 9009 -1599
rect 9009 -1651 9039 -1599
rect 9063 -1651 9073 -1599
rect 9073 -1651 9119 -1599
rect 8823 -1653 8879 -1651
rect 8903 -1653 8959 -1651
rect 8983 -1653 9039 -1651
rect 9063 -1653 9119 -1651
rect 9262 -1599 9318 -1597
rect 9342 -1599 9398 -1597
rect 9262 -1651 9272 -1599
rect 9272 -1651 9318 -1599
rect 9342 -1651 9388 -1599
rect 9388 -1651 9398 -1599
rect 9262 -1653 9318 -1651
rect 9342 -1653 9398 -1651
rect 8143 -1799 8199 -1797
rect 8223 -1799 8279 -1797
rect 8143 -1851 8153 -1799
rect 8153 -1851 8199 -1799
rect 8223 -1851 8269 -1799
rect 8269 -1851 8279 -1799
rect 8143 -1853 8199 -1851
rect 8223 -1853 8279 -1851
rect 8422 -1799 8478 -1797
rect 8502 -1799 8558 -1797
rect 8582 -1799 8638 -1797
rect 8662 -1799 8718 -1797
rect 8422 -1851 8468 -1799
rect 8468 -1851 8478 -1799
rect 8502 -1851 8532 -1799
rect 8532 -1851 8544 -1799
rect 8544 -1851 8558 -1799
rect 8582 -1851 8596 -1799
rect 8596 -1851 8608 -1799
rect 8608 -1851 8638 -1799
rect 8662 -1851 8672 -1799
rect 8672 -1851 8718 -1799
rect 8422 -1853 8478 -1851
rect 8502 -1853 8558 -1851
rect 8582 -1853 8638 -1851
rect 8662 -1853 8718 -1851
rect 8823 -1799 8879 -1797
rect 8903 -1799 8959 -1797
rect 8983 -1799 9039 -1797
rect 9063 -1799 9119 -1797
rect 8823 -1851 8869 -1799
rect 8869 -1851 8879 -1799
rect 8903 -1851 8933 -1799
rect 8933 -1851 8945 -1799
rect 8945 -1851 8959 -1799
rect 8983 -1851 8997 -1799
rect 8997 -1851 9009 -1799
rect 9009 -1851 9039 -1799
rect 9063 -1851 9073 -1799
rect 9073 -1851 9119 -1799
rect 8823 -1853 8879 -1851
rect 8903 -1853 8959 -1851
rect 8983 -1853 9039 -1851
rect 9063 -1853 9119 -1851
rect 9262 -1799 9318 -1797
rect 9342 -1799 9398 -1797
rect 9262 -1851 9272 -1799
rect 9272 -1851 9318 -1799
rect 9342 -1851 9388 -1799
rect 9388 -1851 9398 -1799
rect 9262 -1853 9318 -1851
rect 9342 -1853 9398 -1851
<< metal3 >>
rect 0 9885 70 10050
rect 0 9829 7 9885
rect 63 9829 70 9885
rect 0 8675 70 9829
rect 0 8619 7 8675
rect 63 8619 70 8675
rect 0 7465 70 8619
rect 0 7409 7 7465
rect 63 7409 70 7465
rect 0 6255 70 7409
rect 0 6199 7 6255
rect 63 6199 70 6255
rect 0 4905 70 6199
rect 0 4849 7 4905
rect 63 4849 70 4905
rect 0 3695 70 4849
rect 0 3639 7 3695
rect 63 3639 70 3695
rect 0 2485 70 3639
rect 0 2429 7 2485
rect 63 2429 70 2485
rect 0 1275 70 2429
rect 0 1219 7 1275
rect 63 1219 70 1275
rect 0 65 70 1219
rect 0 9 7 65
rect 63 9 70 65
rect 0 -16 70 9
rect 0 -72 7 -16
rect 63 -72 70 -16
rect 0 -77 70 -72
rect 200 9901 270 10050
rect 200 9845 207 9901
rect 263 9845 270 9901
rect 200 8691 270 9845
rect 200 8635 207 8691
rect 263 8635 270 8691
rect 200 7481 270 8635
rect 200 7425 207 7481
rect 263 7425 270 7481
rect 200 6271 270 7425
rect 200 6215 207 6271
rect 263 6215 270 6271
rect 200 4921 270 6215
rect 200 4865 207 4921
rect 263 4865 270 4921
rect 200 3711 270 4865
rect 200 3655 207 3711
rect 263 3655 270 3711
rect 200 2501 270 3655
rect 200 2445 207 2501
rect 263 2445 270 2501
rect 200 1291 270 2445
rect 200 1235 207 1291
rect 263 1235 270 1291
rect 200 81 270 1235
rect 200 25 207 81
rect 263 25 270 81
rect 200 -16 270 25
rect 200 -72 207 -16
rect 263 -72 270 -16
rect 200 -77 270 -72
rect 400 9885 470 10050
rect 400 9829 407 9885
rect 463 9829 470 9885
rect 400 8675 470 9829
rect 400 8619 407 8675
rect 463 8619 470 8675
rect 400 7465 470 8619
rect 400 7409 407 7465
rect 463 7409 470 7465
rect 400 6255 470 7409
rect 400 6199 407 6255
rect 463 6199 470 6255
rect 400 4905 470 6199
rect 400 4849 407 4905
rect 463 4849 470 4905
rect 400 3695 470 4849
rect 400 3639 407 3695
rect 463 3639 470 3695
rect 400 2485 470 3639
rect 400 2429 407 2485
rect 463 2429 470 2485
rect 400 1275 470 2429
rect 400 1219 407 1275
rect 463 1219 470 1275
rect 400 65 470 1219
rect 400 9 407 65
rect 463 9 470 65
rect 400 -16 470 9
rect 400 -72 407 -16
rect 463 -72 470 -16
rect 400 -77 470 -72
rect 600 9901 670 10050
rect 600 9845 607 9901
rect 663 9845 670 9901
rect 600 8691 670 9845
rect 600 8635 607 8691
rect 663 8635 670 8691
rect 600 7481 670 8635
rect 600 7425 607 7481
rect 663 7425 670 7481
rect 600 6271 670 7425
rect 600 6215 607 6271
rect 663 6215 670 6271
rect 600 4921 670 6215
rect 600 4865 607 4921
rect 663 4865 670 4921
rect 600 3711 670 4865
rect 600 3655 607 3711
rect 663 3655 670 3711
rect 600 2501 670 3655
rect 600 2445 607 2501
rect 663 2445 670 2501
rect 600 1291 670 2445
rect 600 1235 607 1291
rect 663 1235 670 1291
rect 600 81 670 1235
rect 600 25 607 81
rect 663 25 670 81
rect 600 -16 670 25
rect 600 -72 607 -16
rect 663 -72 670 -16
rect 600 -77 670 -72
rect 800 9885 870 10050
rect 800 9829 807 9885
rect 863 9829 870 9885
rect 800 8675 870 9829
rect 800 8619 807 8675
rect 863 8619 870 8675
rect 800 7465 870 8619
rect 800 7409 807 7465
rect 863 7409 870 7465
rect 800 6255 870 7409
rect 800 6199 807 6255
rect 863 6199 870 6255
rect 800 4905 870 6199
rect 800 4849 807 4905
rect 863 4849 870 4905
rect 800 3695 870 4849
rect 800 3639 807 3695
rect 863 3639 870 3695
rect 800 2485 870 3639
rect 800 2429 807 2485
rect 863 2429 870 2485
rect 800 1275 870 2429
rect 800 1219 807 1275
rect 863 1219 870 1275
rect 800 65 870 1219
rect 800 9 807 65
rect 863 9 870 65
rect 800 -16 870 9
rect 800 -72 807 -16
rect 863 -72 870 -16
rect 800 -77 870 -72
rect 1000 9901 1070 10050
rect 1000 9845 1007 9901
rect 1063 9845 1070 9901
rect 1000 8691 1070 9845
rect 1000 8635 1007 8691
rect 1063 8635 1070 8691
rect 1000 7481 1070 8635
rect 1000 7425 1007 7481
rect 1063 7425 1070 7481
rect 1000 6271 1070 7425
rect 1000 6215 1007 6271
rect 1063 6215 1070 6271
rect 1000 4921 1070 6215
rect 1000 4865 1007 4921
rect 1063 4865 1070 4921
rect 1000 3711 1070 4865
rect 1000 3655 1007 3711
rect 1063 3655 1070 3711
rect 1000 2501 1070 3655
rect 1000 2445 1007 2501
rect 1063 2445 1070 2501
rect 1000 1291 1070 2445
rect 1000 1235 1007 1291
rect 1063 1235 1070 1291
rect 1000 81 1070 1235
rect 1000 25 1007 81
rect 1063 25 1070 81
rect 1000 -16 1070 25
rect 1000 -72 1007 -16
rect 1063 -72 1070 -16
rect 1000 -77 1070 -72
rect 1200 9885 1270 10050
rect 1200 9829 1207 9885
rect 1263 9829 1270 9885
rect 1200 8675 1270 9829
rect 1200 8619 1207 8675
rect 1263 8619 1270 8675
rect 1200 7465 1270 8619
rect 1200 7409 1207 7465
rect 1263 7409 1270 7465
rect 1200 6255 1270 7409
rect 1200 6199 1207 6255
rect 1263 6199 1270 6255
rect 1200 4905 1270 6199
rect 1200 4849 1207 4905
rect 1263 4849 1270 4905
rect 1200 3695 1270 4849
rect 1200 3639 1207 3695
rect 1263 3639 1270 3695
rect 1200 2485 1270 3639
rect 1200 2429 1207 2485
rect 1263 2429 1270 2485
rect 1200 1275 1270 2429
rect 1200 1219 1207 1275
rect 1263 1219 1270 1275
rect 1200 65 1270 1219
rect 1200 9 1207 65
rect 1263 9 1270 65
rect 1200 -16 1270 9
rect 1200 -72 1207 -16
rect 1263 -72 1270 -16
rect 1200 -77 1270 -72
rect 1400 9901 1470 10050
rect 1400 9845 1407 9901
rect 1463 9845 1470 9901
rect 1400 8691 1470 9845
rect 1400 8635 1407 8691
rect 1463 8635 1470 8691
rect 1400 7481 1470 8635
rect 1400 7425 1407 7481
rect 1463 7425 1470 7481
rect 1400 6271 1470 7425
rect 1400 6215 1407 6271
rect 1463 6215 1470 6271
rect 1400 4921 1470 6215
rect 1400 4865 1407 4921
rect 1463 4865 1470 4921
rect 1400 3711 1470 4865
rect 1400 3655 1407 3711
rect 1463 3655 1470 3711
rect 1400 2501 1470 3655
rect 1400 2445 1407 2501
rect 1463 2445 1470 2501
rect 1400 1291 1470 2445
rect 1400 1235 1407 1291
rect 1463 1235 1470 1291
rect 1400 81 1470 1235
rect 1400 25 1407 81
rect 1463 25 1470 81
rect 1400 -16 1470 25
rect 1400 -72 1407 -16
rect 1463 -72 1470 -16
rect 1400 -77 1470 -72
rect 1600 9885 1670 10050
rect 1600 9829 1607 9885
rect 1663 9829 1670 9885
rect 1600 8675 1670 9829
rect 1600 8619 1607 8675
rect 1663 8619 1670 8675
rect 1600 7465 1670 8619
rect 1600 7409 1607 7465
rect 1663 7409 1670 7465
rect 1600 6255 1670 7409
rect 1600 6199 1607 6255
rect 1663 6199 1670 6255
rect 1600 4905 1670 6199
rect 1600 4849 1607 4905
rect 1663 4849 1670 4905
rect 1600 3695 1670 4849
rect 1600 3639 1607 3695
rect 1663 3639 1670 3695
rect 1600 2485 1670 3639
rect 1600 2429 1607 2485
rect 1663 2429 1670 2485
rect 1600 1275 1670 2429
rect 1600 1219 1607 1275
rect 1663 1219 1670 1275
rect 1600 65 1670 1219
rect 1600 9 1607 65
rect 1663 9 1670 65
rect 1600 -16 1670 9
rect 1600 -72 1607 -16
rect 1663 -72 1670 -16
rect 1600 -77 1670 -72
rect 1800 9901 1870 10050
rect 1800 9845 1807 9901
rect 1863 9845 1870 9901
rect 1800 8691 1870 9845
rect 1800 8635 1807 8691
rect 1863 8635 1870 8691
rect 1800 7481 1870 8635
rect 1800 7425 1807 7481
rect 1863 7425 1870 7481
rect 1800 6271 1870 7425
rect 1800 6215 1807 6271
rect 1863 6215 1870 6271
rect 1800 4921 1870 6215
rect 1800 4865 1807 4921
rect 1863 4865 1870 4921
rect 1800 3711 1870 4865
rect 1800 3655 1807 3711
rect 1863 3655 1870 3711
rect 1800 2501 1870 3655
rect 1800 2445 1807 2501
rect 1863 2445 1870 2501
rect 1800 1291 1870 2445
rect 1800 1235 1807 1291
rect 1863 1235 1870 1291
rect 1800 81 1870 1235
rect 1800 25 1807 81
rect 1863 25 1870 81
rect 1800 -16 1870 25
rect 1800 -72 1807 -16
rect 1863 -72 1870 -16
rect 1800 -77 1870 -72
rect 2000 9885 2070 10050
rect 2000 9829 2007 9885
rect 2063 9829 2070 9885
rect 2000 8675 2070 9829
rect 2000 8619 2007 8675
rect 2063 8619 2070 8675
rect 2000 7465 2070 8619
rect 2000 7409 2007 7465
rect 2063 7409 2070 7465
rect 2000 6255 2070 7409
rect 2000 6199 2007 6255
rect 2063 6199 2070 6255
rect 2000 4905 2070 6199
rect 2000 4849 2007 4905
rect 2063 4849 2070 4905
rect 2000 3695 2070 4849
rect 2000 3639 2007 3695
rect 2063 3639 2070 3695
rect 2000 2485 2070 3639
rect 2000 2429 2007 2485
rect 2063 2429 2070 2485
rect 2000 1275 2070 2429
rect 2000 1219 2007 1275
rect 2063 1219 2070 1275
rect 2000 65 2070 1219
rect 2000 9 2007 65
rect 2063 9 2070 65
rect 2000 -16 2070 9
rect 2000 -72 2007 -16
rect 2063 -72 2070 -16
rect 2000 -77 2070 -72
rect 2200 9901 2270 10050
rect 2200 9845 2207 9901
rect 2263 9845 2270 9901
rect 2200 8691 2270 9845
rect 2200 8635 2207 8691
rect 2263 8635 2270 8691
rect 2200 7481 2270 8635
rect 2200 7425 2207 7481
rect 2263 7425 2270 7481
rect 2200 6271 2270 7425
rect 2200 6215 2207 6271
rect 2263 6215 2270 6271
rect 2200 4921 2270 6215
rect 2200 4865 2207 4921
rect 2263 4865 2270 4921
rect 2200 3711 2270 4865
rect 2200 3655 2207 3711
rect 2263 3655 2270 3711
rect 2200 2501 2270 3655
rect 2200 2445 2207 2501
rect 2263 2445 2270 2501
rect 2200 1291 2270 2445
rect 2200 1235 2207 1291
rect 2263 1235 2270 1291
rect 2200 81 2270 1235
rect 2200 25 2207 81
rect 2263 25 2270 81
rect 2200 -16 2270 25
rect 2200 -72 2207 -16
rect 2263 -72 2270 -16
rect 2200 -77 2270 -72
rect 2400 9885 2470 10050
rect 2400 9829 2407 9885
rect 2463 9829 2470 9885
rect 2400 8675 2470 9829
rect 2400 8619 2407 8675
rect 2463 8619 2470 8675
rect 2400 7465 2470 8619
rect 2400 7409 2407 7465
rect 2463 7409 2470 7465
rect 2400 6255 2470 7409
rect 2400 6199 2407 6255
rect 2463 6199 2470 6255
rect 2400 4905 2470 6199
rect 2400 4849 2407 4905
rect 2463 4849 2470 4905
rect 2400 3695 2470 4849
rect 2400 3639 2407 3695
rect 2463 3639 2470 3695
rect 2400 2485 2470 3639
rect 2400 2429 2407 2485
rect 2463 2429 2470 2485
rect 2400 1275 2470 2429
rect 2400 1219 2407 1275
rect 2463 1219 2470 1275
rect 2400 65 2470 1219
rect 2400 9 2407 65
rect 2463 9 2470 65
rect 2400 -16 2470 9
rect 2400 -72 2407 -16
rect 2463 -72 2470 -16
rect 2400 -77 2470 -72
rect 2600 9901 2670 10050
rect 2600 9845 2607 9901
rect 2663 9845 2670 9901
rect 2600 8691 2670 9845
rect 2600 8635 2607 8691
rect 2663 8635 2670 8691
rect 2600 7481 2670 8635
rect 2600 7425 2607 7481
rect 2663 7425 2670 7481
rect 2600 6271 2670 7425
rect 2600 6215 2607 6271
rect 2663 6215 2670 6271
rect 2600 4921 2670 6215
rect 2600 4865 2607 4921
rect 2663 4865 2670 4921
rect 2600 3711 2670 4865
rect 2600 3655 2607 3711
rect 2663 3655 2670 3711
rect 2600 2501 2670 3655
rect 2600 2445 2607 2501
rect 2663 2445 2670 2501
rect 2600 1291 2670 2445
rect 2600 1235 2607 1291
rect 2663 1235 2670 1291
rect 2600 81 2670 1235
rect 2600 25 2607 81
rect 2663 25 2670 81
rect 2600 -16 2670 25
rect 2600 -72 2607 -16
rect 2663 -72 2670 -16
rect 2600 -77 2670 -72
rect 2800 9885 2870 10050
rect 2800 9829 2807 9885
rect 2863 9829 2870 9885
rect 2800 8675 2870 9829
rect 2800 8619 2807 8675
rect 2863 8619 2870 8675
rect 2800 7465 2870 8619
rect 2800 7409 2807 7465
rect 2863 7409 2870 7465
rect 2800 6255 2870 7409
rect 2800 6199 2807 6255
rect 2863 6199 2870 6255
rect 2800 4905 2870 6199
rect 2800 4849 2807 4905
rect 2863 4849 2870 4905
rect 2800 3695 2870 4849
rect 2800 3639 2807 3695
rect 2863 3639 2870 3695
rect 2800 2485 2870 3639
rect 2800 2429 2807 2485
rect 2863 2429 2870 2485
rect 2800 1275 2870 2429
rect 2800 1219 2807 1275
rect 2863 1219 2870 1275
rect 2800 65 2870 1219
rect 2800 9 2807 65
rect 2863 9 2870 65
rect 2800 -16 2870 9
rect 2800 -72 2807 -16
rect 2863 -72 2870 -16
rect 2800 -77 2870 -72
rect 3000 9901 3070 10050
rect 3000 9845 3007 9901
rect 3063 9845 3070 9901
rect 3000 8691 3070 9845
rect 3000 8635 3007 8691
rect 3063 8635 3070 8691
rect 3000 7481 3070 8635
rect 3000 7425 3007 7481
rect 3063 7425 3070 7481
rect 3000 6271 3070 7425
rect 3000 6215 3007 6271
rect 3063 6215 3070 6271
rect 3000 4921 3070 6215
rect 3000 4865 3007 4921
rect 3063 4865 3070 4921
rect 3000 3711 3070 4865
rect 3000 3655 3007 3711
rect 3063 3655 3070 3711
rect 3000 2501 3070 3655
rect 3000 2445 3007 2501
rect 3063 2445 3070 2501
rect 3000 1291 3070 2445
rect 3000 1235 3007 1291
rect 3063 1235 3070 1291
rect 3000 81 3070 1235
rect 3000 25 3007 81
rect 3063 25 3070 81
rect 3000 -16 3070 25
rect 3000 -72 3007 -16
rect 3063 -72 3070 -16
rect 3000 -77 3070 -72
rect 3200 9885 3270 10050
rect 3200 9829 3207 9885
rect 3263 9829 3270 9885
rect 3200 8675 3270 9829
rect 3200 8619 3207 8675
rect 3263 8619 3270 8675
rect 3200 7465 3270 8619
rect 3200 7409 3207 7465
rect 3263 7409 3270 7465
rect 3200 6255 3270 7409
rect 3200 6199 3207 6255
rect 3263 6199 3270 6255
rect 3200 4905 3270 6199
rect 3200 4849 3207 4905
rect 3263 4849 3270 4905
rect 3200 3695 3270 4849
rect 3200 3639 3207 3695
rect 3263 3639 3270 3695
rect 3200 2485 3270 3639
rect 3200 2429 3207 2485
rect 3263 2429 3270 2485
rect 3200 1275 3270 2429
rect 3200 1219 3207 1275
rect 3263 1219 3270 1275
rect 3200 65 3270 1219
rect 3200 9 3207 65
rect 3263 9 3270 65
rect 3200 -16 3270 9
rect 3200 -72 3207 -16
rect 3263 -72 3270 -16
rect 3200 -77 3270 -72
rect 3400 9901 3470 10050
rect 3400 9845 3407 9901
rect 3463 9845 3470 9901
rect 3400 8691 3470 9845
rect 3400 8635 3407 8691
rect 3463 8635 3470 8691
rect 3400 7481 3470 8635
rect 3400 7425 3407 7481
rect 3463 7425 3470 7481
rect 3400 6271 3470 7425
rect 3400 6215 3407 6271
rect 3463 6215 3470 6271
rect 3400 4921 3470 6215
rect 3400 4865 3407 4921
rect 3463 4865 3470 4921
rect 3400 3711 3470 4865
rect 3400 3655 3407 3711
rect 3463 3655 3470 3711
rect 3400 2501 3470 3655
rect 3400 2445 3407 2501
rect 3463 2445 3470 2501
rect 3400 1291 3470 2445
rect 3400 1235 3407 1291
rect 3463 1235 3470 1291
rect 3400 81 3470 1235
rect 3400 25 3407 81
rect 3463 25 3470 81
rect 3400 -16 3470 25
rect 3400 -72 3407 -16
rect 3463 -72 3470 -16
rect 3400 -77 3470 -72
rect 3600 9885 3670 10050
rect 3600 9829 3607 9885
rect 3663 9829 3670 9885
rect 3600 8675 3670 9829
rect 3600 8619 3607 8675
rect 3663 8619 3670 8675
rect 3600 7465 3670 8619
rect 3600 7409 3607 7465
rect 3663 7409 3670 7465
rect 3600 6255 3670 7409
rect 3600 6199 3607 6255
rect 3663 6199 3670 6255
rect 3600 4905 3670 6199
rect 3600 4849 3607 4905
rect 3663 4849 3670 4905
rect 3600 3695 3670 4849
rect 3600 3639 3607 3695
rect 3663 3639 3670 3695
rect 3600 2485 3670 3639
rect 3600 2429 3607 2485
rect 3663 2429 3670 2485
rect 3600 1275 3670 2429
rect 3600 1219 3607 1275
rect 3663 1219 3670 1275
rect 3600 65 3670 1219
rect 3600 9 3607 65
rect 3663 9 3670 65
rect 3600 -16 3670 9
rect 3600 -72 3607 -16
rect 3663 -72 3670 -16
rect 3600 -77 3670 -72
rect 3800 9901 3870 10050
rect 3800 9845 3807 9901
rect 3863 9845 3870 9901
rect 3800 8691 3870 9845
rect 3800 8635 3807 8691
rect 3863 8635 3870 8691
rect 3800 7481 3870 8635
rect 3800 7425 3807 7481
rect 3863 7425 3870 7481
rect 3800 6271 3870 7425
rect 3800 6215 3807 6271
rect 3863 6215 3870 6271
rect 3800 4921 3870 6215
rect 3800 4865 3807 4921
rect 3863 4865 3870 4921
rect 3800 3711 3870 4865
rect 3800 3655 3807 3711
rect 3863 3655 3870 3711
rect 3800 2501 3870 3655
rect 3800 2445 3807 2501
rect 3863 2445 3870 2501
rect 3800 1291 3870 2445
rect 3800 1235 3807 1291
rect 3863 1235 3870 1291
rect 3800 81 3870 1235
rect 3800 25 3807 81
rect 3863 25 3870 81
rect 3800 -16 3870 25
rect 3800 -72 3807 -16
rect 3863 -72 3870 -16
rect 3800 -77 3870 -72
rect 4000 9885 4070 10050
rect 4000 9829 4007 9885
rect 4063 9829 4070 9885
rect 4000 8675 4070 9829
rect 4000 8619 4007 8675
rect 4063 8619 4070 8675
rect 4000 7465 4070 8619
rect 4000 7409 4007 7465
rect 4063 7409 4070 7465
rect 4000 6255 4070 7409
rect 4000 6199 4007 6255
rect 4063 6199 4070 6255
rect 4000 4905 4070 6199
rect 4000 4849 4007 4905
rect 4063 4849 4070 4905
rect 4000 3695 4070 4849
rect 4000 3639 4007 3695
rect 4063 3639 4070 3695
rect 4000 2485 4070 3639
rect 4000 2429 4007 2485
rect 4063 2429 4070 2485
rect 4000 1275 4070 2429
rect 4000 1219 4007 1275
rect 4063 1219 4070 1275
rect 4000 65 4070 1219
rect 4000 9 4007 65
rect 4063 9 4070 65
rect 4000 -16 4070 9
rect 4000 -72 4007 -16
rect 4063 -72 4070 -16
rect 4000 -77 4070 -72
rect 4200 9901 4270 10050
rect 4200 9845 4207 9901
rect 4263 9845 4270 9901
rect 4200 8691 4270 9845
rect 4200 8635 4207 8691
rect 4263 8635 4270 8691
rect 4200 7481 4270 8635
rect 4200 7425 4207 7481
rect 4263 7425 4270 7481
rect 4200 6271 4270 7425
rect 4200 6215 4207 6271
rect 4263 6215 4270 6271
rect 4200 4921 4270 6215
rect 4200 4865 4207 4921
rect 4263 4865 4270 4921
rect 4200 3711 4270 4865
rect 4200 3655 4207 3711
rect 4263 3655 4270 3711
rect 4200 2501 4270 3655
rect 4200 2445 4207 2501
rect 4263 2445 4270 2501
rect 4200 1291 4270 2445
rect 4200 1235 4207 1291
rect 4263 1235 4270 1291
rect 4200 81 4270 1235
rect 4200 25 4207 81
rect 4263 25 4270 81
rect 4200 -16 4270 25
rect 4200 -72 4207 -16
rect 4263 -72 4270 -16
rect 4200 -77 4270 -72
rect 4400 9885 4470 10050
rect 4400 9829 4407 9885
rect 4463 9829 4470 9885
rect 4400 8675 4470 9829
rect 4400 8619 4407 8675
rect 4463 8619 4470 8675
rect 4400 7465 4470 8619
rect 4400 7409 4407 7465
rect 4463 7409 4470 7465
rect 4400 6255 4470 7409
rect 4400 6199 4407 6255
rect 4463 6199 4470 6255
rect 4400 4905 4470 6199
rect 4400 4849 4407 4905
rect 4463 4849 4470 4905
rect 4400 3695 4470 4849
rect 4400 3639 4407 3695
rect 4463 3639 4470 3695
rect 4400 2485 4470 3639
rect 4400 2429 4407 2485
rect 4463 2429 4470 2485
rect 4400 1275 4470 2429
rect 4400 1219 4407 1275
rect 4463 1219 4470 1275
rect 4400 65 4470 1219
rect 4400 9 4407 65
rect 4463 9 4470 65
rect 4400 -16 4470 9
rect 4400 -72 4407 -16
rect 4463 -72 4470 -16
rect 4400 -77 4470 -72
rect 4600 9901 4670 10050
rect 4600 9845 4607 9901
rect 4663 9845 4670 9901
rect 4600 8691 4670 9845
rect 4600 8635 4607 8691
rect 4663 8635 4670 8691
rect 4600 7481 4670 8635
rect 4600 7425 4607 7481
rect 4663 7425 4670 7481
rect 4600 6271 4670 7425
rect 4600 6215 4607 6271
rect 4663 6215 4670 6271
rect 4600 4921 4670 6215
rect 4600 4865 4607 4921
rect 4663 4865 4670 4921
rect 4600 3711 4670 4865
rect 4600 3655 4607 3711
rect 4663 3655 4670 3711
rect 4600 2501 4670 3655
rect 4600 2445 4607 2501
rect 4663 2445 4670 2501
rect 4600 1291 4670 2445
rect 4600 1235 4607 1291
rect 4663 1235 4670 1291
rect 4600 81 4670 1235
rect 4600 25 4607 81
rect 4663 25 4670 81
rect 4600 -16 4670 25
rect 4600 -72 4607 -16
rect 4663 -72 4670 -16
rect 4600 -77 4670 -72
rect 4800 9885 4870 10050
rect 4800 9829 4807 9885
rect 4863 9829 4870 9885
rect 4800 8675 4870 9829
rect 4800 8619 4807 8675
rect 4863 8619 4870 8675
rect 4800 7465 4870 8619
rect 4800 7409 4807 7465
rect 4863 7409 4870 7465
rect 4800 6255 4870 7409
rect 4800 6199 4807 6255
rect 4863 6199 4870 6255
rect 4800 4905 4870 6199
rect 4800 4849 4807 4905
rect 4863 4849 4870 4905
rect 4800 3695 4870 4849
rect 4800 3639 4807 3695
rect 4863 3639 4870 3695
rect 4800 2485 4870 3639
rect 4800 2429 4807 2485
rect 4863 2429 4870 2485
rect 4800 1275 4870 2429
rect 4800 1219 4807 1275
rect 4863 1219 4870 1275
rect 4800 65 4870 1219
rect 4800 9 4807 65
rect 4863 9 4870 65
rect 4800 -16 4870 9
rect 4800 -72 4807 -16
rect 4863 -72 4870 -16
rect 4800 -77 4870 -72
rect 5000 9901 5070 10050
rect 5000 9845 5007 9901
rect 5063 9845 5070 9901
rect 5000 8691 5070 9845
rect 5000 8635 5007 8691
rect 5063 8635 5070 8691
rect 5000 7481 5070 8635
rect 5000 7425 5007 7481
rect 5063 7425 5070 7481
rect 5000 6271 5070 7425
rect 5000 6215 5007 6271
rect 5063 6215 5070 6271
rect 5000 4921 5070 6215
rect 5000 4865 5007 4921
rect 5063 4865 5070 4921
rect 5000 3711 5070 4865
rect 5000 3655 5007 3711
rect 5063 3655 5070 3711
rect 5000 2501 5070 3655
rect 5000 2445 5007 2501
rect 5063 2445 5070 2501
rect 5000 1291 5070 2445
rect 5000 1235 5007 1291
rect 5063 1235 5070 1291
rect 5000 81 5070 1235
rect 5000 25 5007 81
rect 5063 25 5070 81
rect 5000 -16 5070 25
rect 5000 -72 5007 -16
rect 5063 -72 5070 -16
rect 5000 -77 5070 -72
rect 5200 9885 5270 10050
rect 5200 9829 5207 9885
rect 5263 9829 5270 9885
rect 5200 8675 5270 9829
rect 5200 8619 5207 8675
rect 5263 8619 5270 8675
rect 5200 7465 5270 8619
rect 5200 7409 5207 7465
rect 5263 7409 5270 7465
rect 5200 6255 5270 7409
rect 5200 6199 5207 6255
rect 5263 6199 5270 6255
rect 5200 4905 5270 6199
rect 5200 4849 5207 4905
rect 5263 4849 5270 4905
rect 5200 3695 5270 4849
rect 5200 3639 5207 3695
rect 5263 3639 5270 3695
rect 5200 2485 5270 3639
rect 5200 2429 5207 2485
rect 5263 2429 5270 2485
rect 5200 1275 5270 2429
rect 5200 1219 5207 1275
rect 5263 1219 5270 1275
rect 5200 65 5270 1219
rect 5200 9 5207 65
rect 5263 9 5270 65
rect 5200 -16 5270 9
rect 5200 -72 5207 -16
rect 5263 -72 5270 -16
rect 5200 -77 5270 -72
rect 5400 9901 5470 10050
rect 5400 9845 5407 9901
rect 5463 9845 5470 9901
rect 5400 8691 5470 9845
rect 5400 8635 5407 8691
rect 5463 8635 5470 8691
rect 5400 7481 5470 8635
rect 5400 7425 5407 7481
rect 5463 7425 5470 7481
rect 5400 6271 5470 7425
rect 5400 6215 5407 6271
rect 5463 6215 5470 6271
rect 5400 4921 5470 6215
rect 5400 4865 5407 4921
rect 5463 4865 5470 4921
rect 5400 3711 5470 4865
rect 5400 3655 5407 3711
rect 5463 3655 5470 3711
rect 5400 2501 5470 3655
rect 5400 2445 5407 2501
rect 5463 2445 5470 2501
rect 5400 1291 5470 2445
rect 5400 1235 5407 1291
rect 5463 1235 5470 1291
rect 5400 81 5470 1235
rect 5400 25 5407 81
rect 5463 25 5470 81
rect 5400 -16 5470 25
rect 5400 -72 5407 -16
rect 5463 -72 5470 -16
rect 5400 -77 5470 -72
rect 5600 9885 5670 10050
rect 5600 9829 5607 9885
rect 5663 9829 5670 9885
rect 5600 8675 5670 9829
rect 5600 8619 5607 8675
rect 5663 8619 5670 8675
rect 5600 7465 5670 8619
rect 5600 7409 5607 7465
rect 5663 7409 5670 7465
rect 5600 6255 5670 7409
rect 5600 6199 5607 6255
rect 5663 6199 5670 6255
rect 5600 4905 5670 6199
rect 5600 4849 5607 4905
rect 5663 4849 5670 4905
rect 5600 3695 5670 4849
rect 5600 3639 5607 3695
rect 5663 3639 5670 3695
rect 5600 2485 5670 3639
rect 5600 2429 5607 2485
rect 5663 2429 5670 2485
rect 5600 1275 5670 2429
rect 5600 1219 5607 1275
rect 5663 1219 5670 1275
rect 5600 65 5670 1219
rect 5600 9 5607 65
rect 5663 9 5670 65
rect 5600 -16 5670 9
rect 5600 -72 5607 -16
rect 5663 -72 5670 -16
rect 5600 -77 5670 -72
rect 5800 9901 5870 10050
rect 5800 9845 5807 9901
rect 5863 9845 5870 9901
rect 5800 8691 5870 9845
rect 5800 8635 5807 8691
rect 5863 8635 5870 8691
rect 5800 7481 5870 8635
rect 5800 7425 5807 7481
rect 5863 7425 5870 7481
rect 5800 6271 5870 7425
rect 5800 6215 5807 6271
rect 5863 6215 5870 6271
rect 5800 4921 5870 6215
rect 5800 4865 5807 4921
rect 5863 4865 5870 4921
rect 5800 3711 5870 4865
rect 5800 3655 5807 3711
rect 5863 3655 5870 3711
rect 5800 2501 5870 3655
rect 5800 2445 5807 2501
rect 5863 2445 5870 2501
rect 5800 1291 5870 2445
rect 5800 1235 5807 1291
rect 5863 1235 5870 1291
rect 5800 81 5870 1235
rect 5800 25 5807 81
rect 5863 25 5870 81
rect 5800 -16 5870 25
rect 5800 -72 5807 -16
rect 5863 -72 5870 -16
rect 5800 -77 5870 -72
rect 6000 9885 6070 10050
rect 6000 9829 6007 9885
rect 6063 9829 6070 9885
rect 6000 8675 6070 9829
rect 6000 8619 6007 8675
rect 6063 8619 6070 8675
rect 6000 7465 6070 8619
rect 6000 7409 6007 7465
rect 6063 7409 6070 7465
rect 6000 6255 6070 7409
rect 6000 6199 6007 6255
rect 6063 6199 6070 6255
rect 6000 4905 6070 6199
rect 6000 4849 6007 4905
rect 6063 4849 6070 4905
rect 6000 3695 6070 4849
rect 6000 3639 6007 3695
rect 6063 3639 6070 3695
rect 6000 2485 6070 3639
rect 6000 2429 6007 2485
rect 6063 2429 6070 2485
rect 6000 1275 6070 2429
rect 6000 1219 6007 1275
rect 6063 1219 6070 1275
rect 6000 65 6070 1219
rect 6000 9 6007 65
rect 6063 9 6070 65
rect 6000 -16 6070 9
rect 6000 -72 6007 -16
rect 6063 -72 6070 -16
rect 6000 -77 6070 -72
rect 6200 9901 6270 10050
rect 6200 9845 6207 9901
rect 6263 9845 6270 9901
rect 6200 8691 6270 9845
rect 6200 8635 6207 8691
rect 6263 8635 6270 8691
rect 6200 7481 6270 8635
rect 6200 7425 6207 7481
rect 6263 7425 6270 7481
rect 6200 6271 6270 7425
rect 6200 6215 6207 6271
rect 6263 6215 6270 6271
rect 6200 4921 6270 6215
rect 6200 4865 6207 4921
rect 6263 4865 6270 4921
rect 6200 3711 6270 4865
rect 6200 3655 6207 3711
rect 6263 3655 6270 3711
rect 6200 2501 6270 3655
rect 6200 2445 6207 2501
rect 6263 2445 6270 2501
rect 6200 1291 6270 2445
rect 6200 1235 6207 1291
rect 6263 1235 6270 1291
rect 6200 81 6270 1235
rect 6200 25 6207 81
rect 6263 25 6270 81
rect 6200 -16 6270 25
rect 6200 -72 6207 -16
rect 6263 -72 6270 -16
rect 6200 -77 6270 -72
rect 8121 3 8302 40
rect 8121 -53 8143 3
rect 8199 -53 8223 3
rect 8279 -53 8302 3
rect -138 -145 6408 -140
rect -138 -201 -133 -145
rect -77 -201 -53 -145
rect 3 -201 67 -145
rect 123 -201 147 -145
rect 203 -201 267 -145
rect 323 -201 347 -145
rect 403 -201 467 -145
rect 523 -201 547 -145
rect 603 -201 667 -145
rect 723 -201 747 -145
rect 803 -201 867 -145
rect 923 -201 947 -145
rect 1003 -201 1067 -145
rect 1123 -201 1147 -145
rect 1203 -201 1267 -145
rect 1323 -201 1347 -145
rect 1403 -201 1467 -145
rect 1523 -201 1547 -145
rect 1603 -201 1667 -145
rect 1723 -201 1747 -145
rect 1803 -201 1867 -145
rect 1923 -201 1947 -145
rect 2003 -201 2067 -145
rect 2123 -201 2147 -145
rect 2203 -201 2267 -145
rect 2323 -201 2347 -145
rect 2403 -201 2467 -145
rect 2523 -201 2547 -145
rect 2603 -201 2667 -145
rect 2723 -201 2747 -145
rect 2803 -201 2867 -145
rect 2923 -201 2947 -145
rect 3003 -201 3067 -145
rect 3123 -201 3147 -145
rect 3203 -201 3267 -145
rect 3323 -201 3347 -145
rect 3403 -201 3467 -145
rect 3523 -201 3547 -145
rect 3603 -201 3667 -145
rect 3723 -201 3747 -145
rect 3803 -201 3867 -145
rect 3923 -201 3947 -145
rect 4003 -201 4067 -145
rect 4123 -201 4147 -145
rect 4203 -201 4267 -145
rect 4323 -201 4347 -145
rect 4403 -201 4467 -145
rect 4523 -201 4547 -145
rect 4603 -201 4667 -145
rect 4723 -201 4747 -145
rect 4803 -201 4867 -145
rect 4923 -201 4947 -145
rect 5003 -201 5067 -145
rect 5123 -201 5147 -145
rect 5203 -201 5267 -145
rect 5323 -201 5347 -145
rect 5403 -201 5467 -145
rect 5523 -201 5547 -145
rect 5603 -201 5667 -145
rect 5723 -201 5747 -145
rect 5803 -201 5867 -145
rect 5923 -201 5947 -145
rect 6003 -201 6067 -145
rect 6123 -201 6147 -145
rect 6203 -201 6267 -145
rect 6323 -201 6347 -145
rect 6403 -201 6408 -145
rect -138 -240 6408 -201
rect 8121 -197 8302 -53
rect 8121 -253 8143 -197
rect 8199 -253 8223 -197
rect 8279 -253 8302 -197
rect -98 -348 6368 -324
rect -98 -404 -93 -348
rect -37 -404 107 -348
rect 163 -404 307 -348
rect 363 -404 507 -348
rect 563 -404 707 -348
rect 763 -404 907 -348
rect 963 -404 1107 -348
rect 1163 -404 1307 -348
rect 1363 -404 1507 -348
rect 1563 -404 1707 -348
rect 1763 -404 1907 -348
rect 1963 -404 2107 -348
rect 2163 -404 2307 -348
rect 2363 -404 2507 -348
rect 2563 -404 2707 -348
rect 2763 -404 2907 -348
rect 2963 -404 3107 -348
rect 3163 -404 3307 -348
rect 3363 -404 3507 -348
rect 3563 -404 3707 -348
rect 3763 -404 3907 -348
rect 3963 -404 4107 -348
rect 4163 -404 4307 -348
rect 4363 -404 4507 -348
rect 4563 -404 4707 -348
rect 4763 -404 4907 -348
rect 4963 -404 5107 -348
rect 5163 -404 5307 -348
rect 5363 -404 5507 -348
rect 5563 -404 5707 -348
rect 5763 -404 5907 -348
rect 5963 -404 6107 -348
rect 6163 -404 6307 -348
rect 6363 -404 6368 -348
rect -98 -428 6368 -404
rect -98 -484 -93 -428
rect -37 -484 107 -428
rect 163 -484 307 -428
rect 363 -484 507 -428
rect 563 -484 707 -428
rect 763 -484 907 -428
rect 963 -484 1107 -428
rect 1163 -484 1307 -428
rect 1363 -484 1507 -428
rect 1563 -484 1707 -428
rect 1763 -484 1907 -428
rect 1963 -484 2107 -428
rect 2163 -484 2307 -428
rect 2363 -484 2507 -428
rect 2563 -484 2707 -428
rect 2763 -484 2907 -428
rect 2963 -484 3107 -428
rect 3163 -484 3307 -428
rect 3363 -484 3507 -428
rect 3563 -484 3707 -428
rect 3763 -484 3907 -428
rect 3963 -484 4107 -428
rect 4163 -484 4307 -428
rect 4363 -484 4507 -428
rect 4563 -484 4707 -428
rect 4763 -484 4907 -428
rect 4963 -484 5107 -428
rect 5163 -484 5307 -428
rect 5363 -484 5507 -428
rect 5563 -484 5707 -428
rect 5763 -484 5907 -428
rect 5963 -484 6107 -428
rect 6163 -484 6307 -428
rect 6363 -484 6368 -428
rect -98 -508 6368 -484
rect 8121 -397 8302 -253
rect 8121 -453 8143 -397
rect 8199 -453 8223 -397
rect 8279 -453 8302 -397
rect 8121 -597 8302 -453
rect 8121 -653 8143 -597
rect 8199 -653 8223 -597
rect 8279 -653 8302 -597
rect 8121 -797 8302 -653
rect 8121 -853 8143 -797
rect 8199 -853 8223 -797
rect 8279 -853 8302 -797
rect 8121 -997 8302 -853
rect 8121 -1053 8143 -997
rect 8199 -1053 8223 -997
rect 8279 -1053 8302 -997
rect 8121 -1197 8302 -1053
rect 8121 -1253 8143 -1197
rect 8199 -1253 8223 -1197
rect 8279 -1253 8302 -1197
rect 8121 -1397 8302 -1253
rect 8121 -1453 8143 -1397
rect 8199 -1453 8223 -1397
rect 8279 -1453 8302 -1397
rect 8121 -1597 8302 -1453
rect 8121 -1653 8143 -1597
rect 8199 -1653 8223 -1597
rect 8279 -1653 8302 -1597
rect 8121 -1797 8302 -1653
rect 8121 -1853 8143 -1797
rect 8199 -1853 8223 -1797
rect 8279 -1853 8302 -1797
rect 8121 -1890 8302 -1853
rect 8400 3 8741 40
rect 8400 -53 8422 3
rect 8478 -53 8502 3
rect 8558 -53 8582 3
rect 8638 -53 8662 3
rect 8718 -53 8741 3
rect 8400 -197 8741 -53
rect 8400 -253 8422 -197
rect 8478 -253 8502 -197
rect 8558 -253 8582 -197
rect 8638 -253 8662 -197
rect 8718 -253 8741 -197
rect 8400 -397 8741 -253
rect 8400 -453 8422 -397
rect 8478 -453 8502 -397
rect 8558 -453 8582 -397
rect 8638 -453 8662 -397
rect 8718 -453 8741 -397
rect 8400 -597 8741 -453
rect 8400 -653 8422 -597
rect 8478 -653 8502 -597
rect 8558 -653 8582 -597
rect 8638 -653 8662 -597
rect 8718 -653 8741 -597
rect 8400 -797 8741 -653
rect 8400 -853 8422 -797
rect 8478 -853 8502 -797
rect 8558 -853 8582 -797
rect 8638 -853 8662 -797
rect 8718 -853 8741 -797
rect 8400 -997 8741 -853
rect 8400 -1053 8422 -997
rect 8478 -1053 8502 -997
rect 8558 -1053 8582 -997
rect 8638 -1053 8662 -997
rect 8718 -1053 8741 -997
rect 8400 -1197 8741 -1053
rect 8400 -1253 8422 -1197
rect 8478 -1253 8502 -1197
rect 8558 -1253 8582 -1197
rect 8638 -1253 8662 -1197
rect 8718 -1253 8741 -1197
rect 8400 -1397 8741 -1253
rect 8400 -1453 8422 -1397
rect 8478 -1453 8502 -1397
rect 8558 -1453 8582 -1397
rect 8638 -1453 8662 -1397
rect 8718 -1453 8741 -1397
rect 8400 -1597 8741 -1453
rect 8400 -1653 8422 -1597
rect 8478 -1653 8502 -1597
rect 8558 -1653 8582 -1597
rect 8638 -1653 8662 -1597
rect 8718 -1653 8741 -1597
rect 8400 -1797 8741 -1653
rect 8400 -1853 8422 -1797
rect 8478 -1853 8502 -1797
rect 8558 -1853 8582 -1797
rect 8638 -1853 8662 -1797
rect 8718 -1853 8741 -1797
rect 8400 -1890 8741 -1853
rect 8801 3 9142 40
rect 8801 -53 8823 3
rect 8879 -53 8903 3
rect 8959 -53 8983 3
rect 9039 -53 9063 3
rect 9119 -53 9142 3
rect 8801 -197 9142 -53
rect 8801 -253 8823 -197
rect 8879 -253 8903 -197
rect 8959 -253 8983 -197
rect 9039 -253 9063 -197
rect 9119 -253 9142 -197
rect 8801 -397 9142 -253
rect 8801 -453 8823 -397
rect 8879 -453 8903 -397
rect 8959 -453 8983 -397
rect 9039 -453 9063 -397
rect 9119 -453 9142 -397
rect 8801 -597 9142 -453
rect 8801 -653 8823 -597
rect 8879 -653 8903 -597
rect 8959 -653 8983 -597
rect 9039 -653 9063 -597
rect 9119 -653 9142 -597
rect 8801 -797 9142 -653
rect 8801 -853 8823 -797
rect 8879 -853 8903 -797
rect 8959 -853 8983 -797
rect 9039 -853 9063 -797
rect 9119 -853 9142 -797
rect 8801 -997 9142 -853
rect 8801 -1053 8823 -997
rect 8879 -1053 8903 -997
rect 8959 -1053 8983 -997
rect 9039 -1053 9063 -997
rect 9119 -1053 9142 -997
rect 8801 -1197 9142 -1053
rect 8801 -1253 8823 -1197
rect 8879 -1253 8903 -1197
rect 8959 -1253 8983 -1197
rect 9039 -1253 9063 -1197
rect 9119 -1253 9142 -1197
rect 8801 -1397 9142 -1253
rect 8801 -1453 8823 -1397
rect 8879 -1453 8903 -1397
rect 8959 -1453 8983 -1397
rect 9039 -1453 9063 -1397
rect 9119 -1453 9142 -1397
rect 8801 -1597 9142 -1453
rect 8801 -1653 8823 -1597
rect 8879 -1653 8903 -1597
rect 8959 -1653 8983 -1597
rect 9039 -1653 9063 -1597
rect 9119 -1653 9142 -1597
rect 8801 -1797 9142 -1653
rect 8801 -1853 8823 -1797
rect 8879 -1853 8903 -1797
rect 8959 -1853 8983 -1797
rect 9039 -1853 9063 -1797
rect 9119 -1853 9142 -1797
rect 8801 -1890 9142 -1853
rect 9240 3 9421 40
rect 9240 -53 9262 3
rect 9318 -53 9342 3
rect 9398 -53 9421 3
rect 9240 -197 9421 -53
rect 9240 -253 9262 -197
rect 9318 -253 9342 -197
rect 9398 -253 9421 -197
rect 9240 -397 9421 -253
rect 9240 -453 9262 -397
rect 9318 -453 9342 -397
rect 9398 -453 9421 -397
rect 9240 -597 9421 -453
rect 9240 -653 9262 -597
rect 9318 -653 9342 -597
rect 9398 -653 9421 -597
rect 9240 -797 9421 -653
rect 9240 -853 9262 -797
rect 9318 -853 9342 -797
rect 9398 -853 9421 -797
rect 9240 -997 9421 -853
rect 9240 -1053 9262 -997
rect 9318 -1053 9342 -997
rect 9398 -1053 9421 -997
rect 9240 -1197 9421 -1053
rect 9240 -1253 9262 -1197
rect 9318 -1253 9342 -1197
rect 9398 -1253 9421 -1197
rect 9240 -1397 9421 -1253
rect 9240 -1453 9262 -1397
rect 9318 -1453 9342 -1397
rect 9398 -1453 9421 -1397
rect 9240 -1597 9421 -1453
rect 9240 -1653 9262 -1597
rect 9318 -1653 9342 -1597
rect 9398 -1653 9421 -1597
rect 9240 -1797 9421 -1653
rect 9240 -1853 9262 -1797
rect 9318 -1853 9342 -1797
rect 9398 -1853 9421 -1797
rect 9240 -1890 9421 -1853
<< properties >>
string GDS_END 4783668
string GDS_FILE ../gds/rom_4k_0_core.gds
string GDS_START 112
<< end >>
