magic
tech sky130A
magscale 1 2
timestamp 1730748763
<< nwell >>
rect 14465 2550 14973 7080
<< locali >>
rect 13911 7000 13945 7016
rect 13911 6950 13945 6966
rect 13911 6860 13945 6876
rect 13911 6810 13945 6826
rect 13911 6720 13945 6736
rect 13911 6670 13945 6686
rect 13911 6580 13945 6596
rect 13911 6530 13945 6546
rect 13911 6440 13945 6456
rect 13911 6390 13945 6406
rect 13911 6300 13945 6316
rect 13911 6250 13945 6266
rect 13911 6160 13945 6176
rect 13911 6110 13945 6126
rect 13911 6020 13945 6036
rect 13911 5970 13945 5986
rect 13911 5790 13945 5806
rect 13911 5740 13945 5756
rect 13911 5650 13945 5666
rect 13911 5600 13945 5616
rect 13911 5510 13945 5526
rect 13911 5460 13945 5476
rect 13911 5370 13945 5386
rect 13911 5320 13945 5336
rect 13911 5230 13945 5246
rect 13911 5180 13945 5196
rect 13911 5090 13945 5106
rect 13911 5040 13945 5056
rect 13911 4950 13945 4966
rect 13911 4900 13945 4916
rect 13911 4810 13945 4826
rect 13911 4760 13945 4776
rect 13911 4580 13945 4596
rect 13911 4530 13945 4546
rect 13911 4440 13945 4456
rect 13911 4390 13945 4406
rect 13911 4300 13945 4316
rect 13911 4250 13945 4266
rect 13911 4160 13945 4176
rect 13911 4110 13945 4126
rect 13911 4020 13945 4036
rect 13911 3970 13945 3986
rect 13911 3880 13945 3896
rect 13911 3830 13945 3846
rect 13911 3740 13945 3756
rect 13911 3690 13945 3706
rect 13911 3600 13945 3616
rect 13911 3550 13945 3566
rect 13911 3370 13945 3386
rect 13911 3320 13945 3336
rect 13911 3230 13945 3246
rect 13911 3180 13945 3196
rect 13911 3090 13945 3106
rect 13911 3040 13945 3056
rect 13911 2950 13945 2966
rect 13911 2900 13945 2916
rect 13911 2810 13945 2826
rect 13911 2760 13945 2776
rect 13911 2670 13945 2686
rect 13911 2620 13945 2636
rect 13911 2530 13945 2546
rect 13911 2480 13945 2496
rect 13911 2390 13945 2406
rect 13911 2340 13945 2356
<< viali >>
rect 13911 6966 13945 7000
rect 13911 6826 13945 6860
rect 13911 6686 13945 6720
rect 13911 6546 13945 6580
rect 13911 6406 13945 6440
rect 13911 6266 13945 6300
rect 13911 6126 13945 6160
rect 13911 5986 13945 6020
rect 13911 5756 13945 5790
rect 13911 5616 13945 5650
rect 13911 5476 13945 5510
rect 13911 5336 13945 5370
rect 13911 5196 13945 5230
rect 13911 5056 13945 5090
rect 13911 4916 13945 4950
rect 13911 4776 13945 4810
rect 13911 4546 13945 4580
rect 13911 4406 13945 4440
rect 13911 4266 13945 4300
rect 13911 4126 13945 4160
rect 13911 3986 13945 4020
rect 13911 3846 13945 3880
rect 13911 3706 13945 3740
rect 13911 3566 13945 3600
rect 13911 3336 13945 3370
rect 13911 3196 13945 3230
rect 13911 3056 13945 3090
rect 13911 2916 13945 2950
rect 13911 2776 13945 2810
rect 13911 2636 13945 2670
rect 13911 2496 13945 2530
rect 13911 2356 13945 2390
<< metal1 >>
rect 13911 7015 13945 7023
rect 13902 7009 13954 7015
rect 13902 6951 13954 6957
rect 13911 6872 13945 6951
rect 13905 6860 13951 6872
rect 13905 6826 13911 6860
rect 13945 6826 13951 6860
rect 13905 6814 13951 6826
rect 13911 6732 13945 6814
rect 13905 6720 13951 6732
rect 13905 6686 13911 6720
rect 13945 6686 13951 6720
rect 13905 6674 13951 6686
rect 13911 6592 13945 6674
rect 13905 6580 13951 6592
rect 13905 6546 13911 6580
rect 13945 6546 13951 6580
rect 13905 6534 13951 6546
rect 13911 6524 13945 6534
rect 13911 6455 13945 6463
rect 13902 6449 13954 6455
rect 13902 6391 13954 6397
rect 13911 6312 13945 6391
rect 13905 6300 13951 6312
rect 13905 6266 13911 6300
rect 13945 6266 13951 6300
rect 13905 6254 13951 6266
rect 13911 6172 13945 6254
rect 13905 6160 13951 6172
rect 13905 6126 13911 6160
rect 13945 6126 13951 6160
rect 13905 6114 13951 6126
rect 13911 6032 13945 6114
rect 13905 6020 13951 6032
rect 13905 5986 13911 6020
rect 13945 5986 13951 6020
rect 13905 5974 13951 5986
rect 13911 5964 13945 5974
rect 13911 5805 13945 5813
rect 13902 5799 13954 5805
rect 13902 5741 13954 5747
rect 13911 5662 13945 5741
rect 13905 5650 13951 5662
rect 13905 5616 13911 5650
rect 13945 5616 13951 5650
rect 13905 5604 13951 5616
rect 13911 5522 13945 5604
rect 13905 5510 13951 5522
rect 13905 5476 13911 5510
rect 13945 5476 13951 5510
rect 13905 5464 13951 5476
rect 13911 5382 13945 5464
rect 13905 5370 13951 5382
rect 13905 5336 13911 5370
rect 13945 5336 13951 5370
rect 13905 5324 13951 5336
rect 13911 5314 13945 5324
rect 13911 5245 13945 5253
rect 13902 5239 13954 5245
rect 13902 5181 13954 5187
rect 13911 5102 13945 5181
rect 13905 5090 13951 5102
rect 13905 5056 13911 5090
rect 13945 5056 13951 5090
rect 13905 5044 13951 5056
rect 13911 4962 13945 5044
rect 13905 4950 13951 4962
rect 13905 4916 13911 4950
rect 13945 4916 13951 4950
rect 13905 4904 13951 4916
rect 13911 4822 13945 4904
rect 13905 4810 13951 4822
rect 13905 4776 13911 4810
rect 13945 4776 13951 4810
rect 13905 4764 13951 4776
rect 13911 4754 13945 4764
rect 13911 4595 13945 4603
rect 13902 4589 13954 4595
rect 13902 4531 13954 4537
rect 13911 4452 13945 4531
rect 13905 4440 13951 4452
rect 13905 4406 13911 4440
rect 13945 4406 13951 4440
rect 13905 4394 13951 4406
rect 13911 4312 13945 4394
rect 13905 4300 13951 4312
rect 13905 4266 13911 4300
rect 13945 4266 13951 4300
rect 13905 4254 13951 4266
rect 13911 4172 13945 4254
rect 13905 4160 13951 4172
rect 13905 4126 13911 4160
rect 13945 4126 13951 4160
rect 13905 4114 13951 4126
rect 13911 4104 13945 4114
rect 13911 4035 13945 4043
rect 13902 4029 13954 4035
rect 13902 3971 13954 3977
rect 13911 3892 13945 3971
rect 13905 3880 13951 3892
rect 13905 3846 13911 3880
rect 13945 3846 13951 3880
rect 13905 3834 13951 3846
rect 13911 3752 13945 3834
rect 13905 3740 13951 3752
rect 13905 3706 13911 3740
rect 13945 3706 13951 3740
rect 13905 3694 13951 3706
rect 13911 3612 13945 3694
rect 13905 3600 13951 3612
rect 13905 3566 13911 3600
rect 13945 3566 13951 3600
rect 13905 3554 13951 3566
rect 13911 3544 13945 3554
rect 13911 3385 13945 3393
rect 13902 3379 13954 3385
rect 13902 3321 13954 3327
rect 13911 3242 13945 3321
rect 13905 3230 13951 3242
rect 13905 3196 13911 3230
rect 13945 3196 13951 3230
rect 13905 3184 13951 3196
rect 13911 3102 13945 3184
rect 13905 3090 13951 3102
rect 13905 3056 13911 3090
rect 13945 3056 13951 3090
rect 13905 3044 13951 3056
rect 13911 2962 13945 3044
rect 13905 2950 13951 2962
rect 13905 2916 13911 2950
rect 13945 2916 13951 2950
rect 13905 2904 13951 2916
rect 13911 2894 13945 2904
rect 13911 2825 13945 2833
rect 13902 2819 13954 2825
rect 13902 2761 13954 2767
rect 13911 2682 13945 2761
rect 13905 2670 13951 2682
rect 13905 2636 13911 2670
rect 13945 2636 13951 2670
rect 13905 2624 13951 2636
rect 13911 2542 13945 2624
rect 14420 2583 14454 7053
rect 15200 6887 15206 6939
rect 15274 6887 15280 6939
rect 15200 6327 15206 6379
rect 15274 6327 15280 6379
rect 15200 5677 15206 5729
rect 15274 5677 15280 5729
rect 15200 5117 15206 5169
rect 15274 5117 15280 5169
rect 15200 4467 15206 4519
rect 15274 4467 15280 4519
rect 15200 3907 15206 3959
rect 15274 3907 15280 3959
rect 15200 3257 15206 3309
rect 15274 3257 15280 3309
rect 15200 2697 15206 2749
rect 15274 2697 15280 2749
rect 13905 2530 13951 2542
rect 13905 2496 13911 2530
rect 13945 2496 13951 2530
rect 13905 2484 13951 2496
rect 13911 2402 13945 2484
rect 13905 2390 13951 2402
rect 13905 2356 13911 2390
rect 13945 2356 13951 2390
rect 13905 2344 13951 2356
rect 13911 2334 13945 2344
rect 41 2003 157 2033
rect 13011 2003 13127 2033
rect 41 1581 71 2003
rect 13097 1581 13127 2003
rect 41 1551 101 1581
rect 13067 1551 13127 1581
rect 13239 1403 13269 2213
rect 13299 1503 13329 2213
rect 13529 1603 13559 2213
rect 13629 1703 13659 2213
rect 13729 1803 13759 2213
rect 13829 1903 13859 2213
rect 13829 1873 14649 1903
rect 13729 1773 14649 1803
rect 13629 1673 14649 1703
rect 13529 1573 14649 1603
rect 13299 1473 14649 1503
rect 13239 1373 14649 1403
rect 13025 1273 14649 1303
rect 13025 1173 14649 1203
rect 13025 1073 14649 1103
rect 13025 973 14649 1003
rect 13025 873 14649 903
rect 13025 773 14649 803
rect 13025 673 14649 703
rect 13025 573 14649 603
rect 13025 473 14649 503
rect 13025 373 14649 403
rect 13025 273 14649 303
rect 13025 173 14649 203
rect 11 90 211 96
rect 11 32 17 90
rect 205 32 211 90
rect 11 26 211 32
rect 12957 90 13157 96
rect 12957 32 12963 90
rect 13151 32 13157 90
rect 12957 26 13157 32
<< via1 >>
rect 13902 7000 13954 7009
rect 13902 6966 13911 7000
rect 13911 6966 13945 7000
rect 13945 6966 13954 7000
rect 13902 6957 13954 6966
rect 13902 6440 13954 6449
rect 13902 6406 13911 6440
rect 13911 6406 13945 6440
rect 13945 6406 13954 6440
rect 13902 6397 13954 6406
rect 13902 5790 13954 5799
rect 13902 5756 13911 5790
rect 13911 5756 13945 5790
rect 13945 5756 13954 5790
rect 13902 5747 13954 5756
rect 13902 5230 13954 5239
rect 13902 5196 13911 5230
rect 13911 5196 13945 5230
rect 13945 5196 13954 5230
rect 13902 5187 13954 5196
rect 13902 4580 13954 4589
rect 13902 4546 13911 4580
rect 13911 4546 13945 4580
rect 13945 4546 13954 4580
rect 13902 4537 13954 4546
rect 13902 4020 13954 4029
rect 13902 3986 13911 4020
rect 13911 3986 13945 4020
rect 13945 3986 13954 4020
rect 13902 3977 13954 3986
rect 13902 3370 13954 3379
rect 13902 3336 13911 3370
rect 13911 3336 13945 3370
rect 13945 3336 13954 3370
rect 13902 3327 13954 3336
rect 13902 2810 13954 2819
rect 13902 2776 13911 2810
rect 13911 2776 13945 2810
rect 13945 2776 13954 2810
rect 13902 2767 13954 2776
rect 15206 6887 15274 6939
rect 15206 6327 15274 6379
rect 15206 5677 15274 5729
rect 15206 5117 15274 5169
rect 15206 4467 15274 4519
rect 15206 3907 15274 3959
rect 15206 3257 15274 3309
rect 15206 2697 15274 2749
rect 17 32 205 90
rect 12963 32 13151 90
<< metal2 >>
rect 13902 7009 13954 7015
rect 13902 6936 13954 6957
rect 13902 6890 14400 6936
rect 15200 6887 15206 6939
rect 15274 6887 16180 6939
rect 13902 6449 13954 6455
rect 13902 6376 13954 6397
rect 13902 6330 14400 6376
rect 15200 6327 15206 6379
rect 15274 6327 16180 6379
rect 13902 5799 13954 5805
rect 13902 5726 13954 5747
rect 13902 5680 14400 5726
rect 15200 5677 15206 5729
rect 15274 5677 16180 5729
rect 13902 5239 13954 5245
rect 13902 5166 13954 5187
rect 13902 5120 14400 5166
rect 15200 5117 15206 5169
rect 15274 5117 16180 5169
rect 13902 4589 13954 4595
rect 13902 4516 13954 4537
rect 13902 4470 14400 4516
rect 15200 4467 15206 4519
rect 15274 4467 16180 4519
rect 13902 4029 13954 4035
rect 13902 3956 13954 3977
rect 13902 3910 14400 3956
rect 15200 3907 15206 3959
rect 15274 3907 16180 3959
rect 13902 3379 13954 3385
rect 13902 3306 13954 3327
rect 13902 3260 14400 3306
rect 15200 3257 15206 3309
rect 15274 3257 16180 3309
rect 13902 2819 13954 2825
rect 13902 2746 13954 2767
rect 13902 2700 14400 2746
rect 15200 2697 15206 2749
rect 15274 2697 16180 2749
rect 14417 2103 14426 2253
rect 14665 2248 15795 2253
rect 14665 2108 15054 2248
rect 15786 2108 15795 2248
rect 14665 2103 15795 2108
rect 11 1534 111 2103
rect 11 1294 16 1534
rect 106 1294 111 1534
rect 11 96 111 1294
rect 13057 2068 13257 2103
rect 13057 1978 13076 2068
rect 13252 1978 13257 2068
rect 13057 1534 13257 1978
rect 16089 1862 16180 1914
rect 16089 1662 16180 1714
rect 13057 1294 13062 1534
rect 13252 1294 13257 1534
rect 16089 1462 16180 1514
rect 13057 1285 13257 1294
rect 13057 96 13157 1285
rect 16089 1262 16180 1314
rect 16089 1062 16180 1114
rect 16089 862 16180 914
rect 16089 662 16180 714
rect 16089 462 16180 514
rect 16089 262 16180 314
rect 11 90 211 96
rect 11 32 17 90
rect 205 32 211 90
rect 11 26 211 32
rect 12957 90 13157 96
rect 12957 32 12963 90
rect 13151 32 13157 90
rect 12957 26 13157 32
<< via2 >>
rect 14426 2103 14665 2253
rect 15054 2108 15786 2248
rect 16 1294 106 1534
rect 13076 1978 13252 2068
rect 13062 1294 13252 1534
<< metal3 >>
rect 14675 2902 14943 7053
rect 14421 2653 14943 2902
rect 14421 2583 14675 2653
rect 14421 2253 14670 2583
rect 15059 2553 15169 7053
rect 15059 2523 16070 2553
rect 14421 2103 14426 2253
rect 14665 2103 14670 2253
rect 111 2068 13257 2073
rect 111 1978 13076 2068
rect 13252 1978 13257 2068
rect 111 1973 13257 1978
rect 14421 1889 14670 2103
rect 14770 2353 16070 2523
rect 14770 2053 14951 2353
rect 15049 2248 15791 2253
rect 15049 2108 15054 2248
rect 15786 2108 15791 2248
rect 15049 2053 15791 2108
rect 15889 2053 16070 2353
rect 151 1639 14670 1889
rect 11 1534 14770 1539
rect 11 1294 16 1534
rect 106 1294 13062 1534
rect 13252 1294 14770 1534
rect 11 1289 14770 1294
use out_drive  out_drive_0
timestamp 1728730538
transform 1 0 9700 0 1 6633
box 4700 -55 5500 474
use out_drive  out_drive_1
timestamp 1728730538
transform 1 0 9700 0 1 2443
box 4700 -55 5500 474
use out_drive  out_drive_2
timestamp 1728730538
transform 1 0 9700 0 1 3003
box 4700 -55 5500 474
use out_drive  out_drive_3
timestamp 1728730538
transform 1 0 9700 0 1 3653
box 4700 -55 5500 474
use out_drive  out_drive_4
timestamp 1728730538
transform 1 0 9700 0 1 4213
box 4700 -55 5500 474
use out_drive  out_drive_5
timestamp 1728730538
transform 1 0 9700 0 1 4863
box 4700 -55 5500 474
use out_drive  out_drive_6
timestamp 1728730538
transform 1 0 9700 0 1 5423
box 4700 -55 5500 474
use out_drive  out_drive_7
timestamp 1728730538
transform 1 0 9700 0 1 6073
box 4700 -55 5500 474
use rom_4k_1_core  rom_4k_1_core_0
timestamp 1730660070
transform 1 0 249 0 1 2213
box -169 -2213 15840 5070
<< labels >>
flabel metal3 s 151 1639 14670 1889 0 FreeSans 400 0 0 0 VPWR
port 21 nsew power bidirectional
flabel metal3 s 111 1973 13257 2073 0 FreeSans 400 0 0 0 VGND
port 20 nsew ground bidirectional
flabel metal3 s 11 1289 14951 1539 0 FreeSans 400 0 0 0 VGND
port 20 nsew ground bidirectional
flabel metal2 s 16120 262 16180 314 0 FreeSans 160 0 0 0 addr[8]
port 10 nsew signal input
flabel metal2 s 16120 462 16180 514 0 FreeSans 160 0 0 0 addr[7]
port 9 nsew signal input
flabel metal2 s 16120 662 16180 714 0 FreeSans 160 0 0 0 addr[6]
port 8 nsew signal input
flabel metal2 s 16120 862 16180 914 0 FreeSans 160 0 0 0 addr[5]
port 7 nsew signal input
flabel metal2 s 16120 1062 16180 1114 0 FreeSans 160 0 0 0 addr[4]
port 6 nsew signal input
flabel metal2 s 16120 1262 16180 1314 0 FreeSans 160 0 0 0 addr[3]
port 5 nsew signal input
flabel metal2 s 16120 1862 16180 1914 0 FreeSans 160 0 0 0 addr[2]
port 2 nsew signal input
flabel metal2 s 16120 1662 16180 1714 0 FreeSans 160 0 0 0 addr[1]
port 1 nsew signal input
flabel metal2 s 16120 1462 16180 1514 0 FreeSans 160 0 0 0 addr[0]
port 0 nsew signal input
flabel metal2 s 16120 2697 16180 2749 0 FreeSans 160 0 0 0 q[0]
port 12 nsew signal output
flabel metal2 s 16120 3257 16180 3309 0 FreeSans 160 0 0 0 q[1]
port 13 nsew signal output
flabel metal2 s 16120 3907 16180 3959 0 FreeSans 160 0 0 0 q[2]
port 14 nsew signal output
flabel metal2 s 16120 4467 16180 4519 0 FreeSans 160 0 0 0 q[3]
port 15 nsew signal output
flabel metal2 s 16120 5117 16180 5169 0 FreeSans 160 0 0 0 q[4]
port 16 nsew signal output
flabel metal2 s 16120 5677 16180 5729 0 FreeSans 160 0 0 0 q[5]
port 17 nsew signal output
flabel metal2 s 16120 6327 16180 6379 0 FreeSans 160 0 0 0 q[6]
port 18 nsew signal output
flabel metal2 s 16120 6887 16180 6939 0 FreeSans 160 0 0 0 q[7]
port 19 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 16180 7283
<< end >>
