magic
tech sky130A
magscale 1 2
timestamp 1728730538
<< nwell >>
rect 4765 -55 5273 460
<< nmos >>
rect 5357 308 5457 338
rect 5357 222 5457 252
<< pmos >>
rect 4801 234 4885 326
rect 4987 308 5237 338
rect 4987 222 5237 252
<< ndiff >>
rect 5357 383 5457 391
rect 5357 349 5369 383
rect 5445 349 5457 383
rect 5357 338 5457 349
rect 5357 297 5457 308
rect 5357 263 5368 297
rect 5449 263 5457 297
rect 5357 252 5457 263
rect 5357 211 5457 222
rect 5357 177 5369 211
rect 5445 177 5457 211
rect 5357 169 5457 177
<< pdiff >>
rect 4801 383 4885 391
rect 4801 349 4826 383
rect 4860 349 4885 383
rect 4801 326 4885 349
rect 4987 383 5237 391
rect 4987 349 4999 383
rect 5225 349 5237 383
rect 4987 338 5237 349
rect 4987 297 5237 308
rect 4987 263 4995 297
rect 5229 263 5237 297
rect 4987 252 5237 263
rect 4801 211 4885 234
rect 4801 177 4826 211
rect 4860 177 4885 211
rect 4801 169 4885 177
rect 4987 211 5237 222
rect 4987 177 4999 211
rect 5225 177 5237 211
rect 4987 169 5237 177
<< ndiffc >>
rect 5369 349 5445 383
rect 5368 263 5449 297
rect 5369 177 5445 211
<< pdiffc >>
rect 4826 349 4860 383
rect 4999 349 5225 383
rect 4995 263 5229 297
rect 4826 177 4860 211
rect 4999 177 5225 211
<< psubdiff >>
rect 5299 -19 5323 15
rect 5433 -19 5457 15
<< nsubdiff >>
rect 4801 -19 4825 15
rect 5213 -19 5237 15
<< psubdiffcont >>
rect 5323 -19 5433 15
<< nsubdiffcont >>
rect 4825 -19 5213 15
<< poly >>
rect 4710 297 4801 326
rect 4710 263 4720 297
rect 4754 263 4801 297
rect 4710 234 4801 263
rect 4885 234 4911 326
rect 4953 308 4987 338
rect 5237 322 5357 338
rect 5237 308 5284 322
rect 5274 252 5284 308
rect 4953 222 4987 252
rect 5237 238 5284 252
rect 5318 308 5357 322
rect 5457 308 5483 338
rect 5318 252 5328 308
rect 5318 238 5357 252
rect 5237 222 5357 238
rect 5457 222 5483 252
<< polycont >>
rect 4720 263 4754 297
rect 5284 238 5318 322
<< locali >>
rect 4810 349 4826 383
rect 4860 349 4876 383
rect 5235 349 5241 383
rect 5353 349 5367 383
rect 5284 322 5318 338
rect 4720 297 4754 313
rect 4720 247 4754 263
rect 5284 211 5318 238
rect 4809 177 4826 211
rect 4860 177 4983 211
rect 5235 177 5241 211
rect 4809 15 5241 177
rect 5284 165 5318 177
rect 5353 177 5367 211
rect 5353 15 5461 177
rect 4809 -19 4825 15
rect 5213 -19 5241 15
rect 5307 -19 5323 15
rect 5433 -19 5461 15
<< viali >>
rect 4826 349 4860 383
rect 4983 349 4999 383
rect 4999 349 5225 383
rect 5225 349 5235 383
rect 5367 349 5369 383
rect 5369 349 5445 383
rect 5445 349 5461 383
rect 4720 263 4754 297
rect 4979 263 4995 297
rect 4995 263 5229 297
rect 5229 263 5245 297
rect 5352 263 5368 297
rect 5368 263 5449 297
rect 5449 263 5465 297
rect 4983 177 4999 211
rect 4999 177 5225 211
rect 5225 177 5235 211
rect 5284 177 5318 211
rect 5367 177 5369 211
rect 5369 177 5445 211
rect 5445 177 5461 211
<< metal1 >>
rect 4720 440 5389 474
rect 4720 309 4754 440
rect 5355 395 5389 440
rect 4820 383 4866 395
rect 4820 349 4826 383
rect 4860 349 4866 383
rect 4820 312 4866 349
rect 4971 343 4977 395
rect 5241 343 5247 395
rect 5355 343 5361 395
rect 5467 343 5473 395
rect 4714 297 4760 309
rect 4714 263 4720 297
rect 4754 263 4760 297
rect 4714 251 4760 263
rect 4817 306 4869 312
rect 4967 297 5500 303
rect 4967 263 4979 297
rect 5245 263 5352 297
rect 5465 263 5500 297
rect 4967 257 5500 263
rect 4720 140 4754 251
rect 4817 248 4869 254
rect 5275 217 5327 223
rect 4971 165 4977 217
rect 5241 165 5247 217
rect 5355 165 5361 217
rect 5467 165 5473 217
rect 5275 159 5327 165
<< via1 >>
rect 4977 383 5241 395
rect 4977 349 4983 383
rect 4983 349 5235 383
rect 5235 349 5241 383
rect 4977 343 5241 349
rect 5361 383 5467 395
rect 5361 349 5367 383
rect 5367 349 5461 383
rect 5461 349 5467 383
rect 5361 343 5467 349
rect 4817 254 4869 306
rect 4977 211 5241 217
rect 4977 177 4983 211
rect 4983 177 5235 211
rect 5235 177 5241 211
rect 4977 165 5241 177
rect 5275 211 5327 217
rect 5275 177 5284 211
rect 5284 177 5318 211
rect 5318 177 5327 211
rect 5275 165 5327 177
rect 5361 211 5467 217
rect 5361 177 5367 211
rect 5367 177 5461 211
rect 5461 177 5467 211
rect 5361 165 5467 177
<< metal2 >>
rect 4971 395 4980 399
rect 5238 395 5247 399
rect 4971 343 4977 395
rect 5241 343 5247 395
rect 5355 395 5364 399
rect 5464 395 5473 399
rect 5355 343 5361 395
rect 5467 343 5473 395
rect 4811 303 4817 306
rect 4700 257 4817 303
rect 4811 254 4817 257
rect 4869 303 4875 306
rect 4869 257 5327 303
rect 4869 254 4875 257
rect 5275 217 5327 257
rect 4971 165 4977 217
rect 5241 165 5247 217
rect 4971 161 4980 165
rect 5238 161 5247 165
rect 5275 159 5327 165
rect 5355 165 5361 217
rect 5467 165 5473 217
rect 5355 161 5364 165
rect 5464 161 5473 165
<< via2 >>
rect 4980 395 5238 399
rect 4980 343 5238 395
rect 5364 395 5464 399
rect 5364 343 5464 395
rect 4980 165 5238 217
rect 4980 161 5238 165
rect 5364 165 5464 217
rect 5364 161 5464 165
<< metal3 >>
rect 4975 399 5243 420
rect 4975 343 4980 399
rect 5238 343 5243 399
rect 4975 217 5243 343
rect 4975 161 4980 217
rect 5238 161 5243 217
rect 4975 140 5243 161
rect 5359 399 5469 420
rect 5359 343 5364 399
rect 5464 343 5469 399
rect 5359 217 5469 343
rect 5359 161 5364 217
rect 5464 161 5469 217
rect 5359 140 5469 161
<< end >>
