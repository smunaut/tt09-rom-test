magic
tech sky130A
magscale 1 2
timestamp 1730749399
<< nwell >>
rect 8065 2910 8573 11860
<< locali >>
rect 7711 11780 7745 11796
rect 7711 11730 7745 11746
rect 7711 11640 7745 11656
rect 7711 11590 7745 11606
rect 7711 11500 7745 11516
rect 7711 11450 7745 11466
rect 7711 11360 7745 11376
rect 7711 11310 7745 11326
rect 7711 11220 7745 11236
rect 7711 11170 7745 11186
rect 7711 11080 7745 11096
rect 7711 11030 7745 11046
rect 7711 10940 7745 10956
rect 7711 10890 7745 10906
rect 7711 10800 7745 10816
rect 7711 10750 7745 10766
rect 7711 10570 7745 10586
rect 7711 10520 7745 10536
rect 7711 10430 7745 10446
rect 7711 10380 7745 10396
rect 7711 10290 7745 10306
rect 7711 10240 7745 10256
rect 7711 10150 7745 10166
rect 7711 10100 7745 10116
rect 7711 10010 7745 10026
rect 7711 9960 7745 9976
rect 7711 9870 7745 9886
rect 7711 9820 7745 9836
rect 7711 9730 7745 9746
rect 7711 9680 7745 9696
rect 7711 9590 7745 9606
rect 7711 9540 7745 9556
rect 7711 9360 7745 9376
rect 7711 9310 7745 9326
rect 7711 9220 7745 9236
rect 7711 9170 7745 9186
rect 7711 9080 7745 9096
rect 7711 9030 7745 9046
rect 7711 8940 7745 8956
rect 7711 8890 7745 8906
rect 7711 8800 7745 8816
rect 7711 8750 7745 8766
rect 7711 8660 7745 8676
rect 7711 8610 7745 8626
rect 7711 8520 7745 8536
rect 7711 8470 7745 8486
rect 7711 8380 7745 8396
rect 7711 8330 7745 8346
rect 7711 8150 7745 8166
rect 7711 8100 7745 8116
rect 7711 8010 7745 8026
rect 7711 7960 7745 7976
rect 7711 7870 7745 7886
rect 7711 7820 7745 7836
rect 7711 7730 7745 7746
rect 7711 7680 7745 7696
rect 7711 7590 7745 7606
rect 7711 7540 7745 7556
rect 7711 7450 7745 7466
rect 7711 7400 7745 7416
rect 7711 7310 7745 7326
rect 7711 7260 7745 7276
rect 7711 7170 7745 7186
rect 7711 7120 7745 7136
rect 7711 6800 7745 6816
rect 7711 6750 7745 6766
rect 7711 6660 7745 6676
rect 7711 6610 7745 6626
rect 7711 6520 7745 6536
rect 7711 6470 7745 6486
rect 7711 6380 7745 6396
rect 7711 6330 7745 6346
rect 7711 6240 7745 6256
rect 7711 6190 7745 6206
rect 7711 6100 7745 6116
rect 7711 6050 7745 6066
rect 7711 5960 7745 5976
rect 7711 5910 7745 5926
rect 7711 5820 7745 5836
rect 7711 5770 7745 5786
rect 7711 5590 7745 5606
rect 7711 5540 7745 5556
rect 7711 5450 7745 5466
rect 7711 5400 7745 5416
rect 7711 5310 7745 5326
rect 7711 5260 7745 5276
rect 7711 5170 7745 5186
rect 7711 5120 7745 5136
rect 7711 5030 7745 5046
rect 7711 4980 7745 4996
rect 7711 4890 7745 4906
rect 7711 4840 7745 4856
rect 7711 4750 7745 4766
rect 7711 4700 7745 4716
rect 7711 4610 7745 4626
rect 7711 4560 7745 4576
rect 7711 4380 7745 4396
rect 7711 4330 7745 4346
rect 7711 4240 7745 4256
rect 7711 4190 7745 4206
rect 7711 4100 7745 4116
rect 7711 4050 7745 4066
rect 7711 3960 7745 3976
rect 7711 3910 7745 3926
rect 7711 3820 7745 3836
rect 7711 3770 7745 3786
rect 7711 3680 7745 3696
rect 7711 3630 7745 3646
rect 7711 3540 7745 3556
rect 7711 3490 7745 3506
rect 7711 3400 7745 3416
rect 7711 3350 7745 3366
rect 7711 3170 7745 3186
rect 7711 3120 7745 3136
rect 7711 3030 7745 3046
rect 7711 2980 7745 2996
rect 7711 2890 7745 2906
rect 7711 2840 7745 2856
rect 7711 2750 7745 2766
rect 7711 2700 7745 2716
rect 7711 2610 7745 2626
rect 7711 2560 7745 2576
rect 7711 2470 7745 2486
rect 7711 2420 7745 2436
rect 7711 2330 7745 2346
rect 7711 2280 7745 2296
rect 7711 2190 7745 2206
rect 7711 2140 7745 2156
<< viali >>
rect 7711 11746 7745 11780
rect 7711 11606 7745 11640
rect 7711 11466 7745 11500
rect 7711 11326 7745 11360
rect 7711 11186 7745 11220
rect 7711 11046 7745 11080
rect 7711 10906 7745 10940
rect 7711 10766 7745 10800
rect 7711 10536 7745 10570
rect 7711 10396 7745 10430
rect 7711 10256 7745 10290
rect 7711 10116 7745 10150
rect 7711 9976 7745 10010
rect 7711 9836 7745 9870
rect 7711 9696 7745 9730
rect 7711 9556 7745 9590
rect 7711 9326 7745 9360
rect 7711 9186 7745 9220
rect 7711 9046 7745 9080
rect 7711 8906 7745 8940
rect 7711 8766 7745 8800
rect 7711 8626 7745 8660
rect 7711 8486 7745 8520
rect 7711 8346 7745 8380
rect 7711 8116 7745 8150
rect 7711 7976 7745 8010
rect 7711 7836 7745 7870
rect 7711 7696 7745 7730
rect 7711 7556 7745 7590
rect 7711 7416 7745 7450
rect 7711 7276 7745 7310
rect 7711 7136 7745 7170
rect 7711 6766 7745 6800
rect 7711 6626 7745 6660
rect 7711 6486 7745 6520
rect 7711 6346 7745 6380
rect 7711 6206 7745 6240
rect 7711 6066 7745 6100
rect 7711 5926 7745 5960
rect 7711 5786 7745 5820
rect 7711 5556 7745 5590
rect 7711 5416 7745 5450
rect 7711 5276 7745 5310
rect 7711 5136 7745 5170
rect 7711 4996 7745 5030
rect 7711 4856 7745 4890
rect 7711 4716 7745 4750
rect 7711 4576 7745 4610
rect 7711 4346 7745 4380
rect 7711 4206 7745 4240
rect 7711 4066 7745 4100
rect 7711 3926 7745 3960
rect 7711 3786 7745 3820
rect 7711 3646 7745 3680
rect 7711 3506 7745 3540
rect 7711 3366 7745 3400
rect 7711 3136 7745 3170
rect 7711 2996 7745 3030
rect 7711 2856 7745 2890
rect 7711 2716 7745 2750
rect 7711 2576 7745 2610
rect 7711 2436 7745 2470
rect 7711 2296 7745 2330
rect 7711 2156 7745 2190
<< metal1 >>
rect 7711 11795 7745 11803
rect 7702 11789 7754 11795
rect 7702 11731 7754 11737
rect 7711 11652 7745 11731
rect 7705 11640 7751 11652
rect 7705 11606 7711 11640
rect 7745 11606 7751 11640
rect 7705 11594 7751 11606
rect 7711 11512 7745 11594
rect 7705 11500 7751 11512
rect 7705 11466 7711 11500
rect 7745 11466 7751 11500
rect 7705 11454 7751 11466
rect 7711 11372 7745 11454
rect 7705 11360 7751 11372
rect 7705 11326 7711 11360
rect 7745 11326 7751 11360
rect 7705 11314 7751 11326
rect 7711 11232 7745 11314
rect 7705 11220 7751 11232
rect 7705 11186 7711 11220
rect 7745 11186 7751 11220
rect 7705 11174 7751 11186
rect 7711 11092 7745 11174
rect 7705 11080 7751 11092
rect 7705 11046 7711 11080
rect 7745 11046 7751 11080
rect 7705 11034 7751 11046
rect 7711 10952 7745 11034
rect 7705 10940 7751 10952
rect 7705 10906 7711 10940
rect 7745 10906 7751 10940
rect 7705 10894 7751 10906
rect 7711 10812 7745 10894
rect 7705 10800 7751 10812
rect 7705 10766 7711 10800
rect 7745 10766 7751 10800
rect 7705 10754 7751 10766
rect 7711 10744 7745 10754
rect 7711 10585 7745 10593
rect 7702 10579 7754 10585
rect 7702 10521 7754 10527
rect 7711 10442 7745 10521
rect 7705 10430 7751 10442
rect 7705 10396 7711 10430
rect 7745 10396 7751 10430
rect 7705 10384 7751 10396
rect 7711 10302 7745 10384
rect 7705 10290 7751 10302
rect 7705 10256 7711 10290
rect 7745 10256 7751 10290
rect 7705 10244 7751 10256
rect 7711 10162 7745 10244
rect 7705 10150 7751 10162
rect 7705 10116 7711 10150
rect 7745 10116 7751 10150
rect 7705 10104 7751 10116
rect 7711 10022 7745 10104
rect 7705 10010 7751 10022
rect 7705 9976 7711 10010
rect 7745 9976 7751 10010
rect 7705 9964 7751 9976
rect 7711 9882 7745 9964
rect 7705 9870 7751 9882
rect 7705 9836 7711 9870
rect 7745 9836 7751 9870
rect 7705 9824 7751 9836
rect 7711 9742 7745 9824
rect 7705 9730 7751 9742
rect 7705 9696 7711 9730
rect 7745 9696 7751 9730
rect 7705 9684 7751 9696
rect 7711 9602 7745 9684
rect 7705 9590 7751 9602
rect 7705 9556 7711 9590
rect 7745 9556 7751 9590
rect 7705 9544 7751 9556
rect 7711 9534 7745 9544
rect 7711 9375 7745 9383
rect 7702 9369 7754 9375
rect 7702 9311 7754 9317
rect 7711 9232 7745 9311
rect 7705 9220 7751 9232
rect 7705 9186 7711 9220
rect 7745 9186 7751 9220
rect 7705 9174 7751 9186
rect 7711 9092 7745 9174
rect 7705 9080 7751 9092
rect 7705 9046 7711 9080
rect 7745 9046 7751 9080
rect 7705 9034 7751 9046
rect 7711 8952 7745 9034
rect 7705 8940 7751 8952
rect 7705 8906 7711 8940
rect 7745 8906 7751 8940
rect 7705 8894 7751 8906
rect 7711 8812 7745 8894
rect 7705 8800 7751 8812
rect 7705 8766 7711 8800
rect 7745 8766 7751 8800
rect 7705 8754 7751 8766
rect 7711 8672 7745 8754
rect 7705 8660 7751 8672
rect 7705 8626 7711 8660
rect 7745 8626 7751 8660
rect 7705 8614 7751 8626
rect 7711 8532 7745 8614
rect 7705 8520 7751 8532
rect 7705 8486 7711 8520
rect 7745 8486 7751 8520
rect 7705 8474 7751 8486
rect 7711 8392 7745 8474
rect 7705 8380 7751 8392
rect 7705 8346 7711 8380
rect 7745 8346 7751 8380
rect 7705 8334 7751 8346
rect 7711 8324 7745 8334
rect 7711 8165 7745 8173
rect 7702 8159 7754 8165
rect 7702 8101 7754 8107
rect 7711 8022 7745 8101
rect 7705 8010 7751 8022
rect 7705 7976 7711 8010
rect 7745 7976 7751 8010
rect 7705 7964 7751 7976
rect 7711 7882 7745 7964
rect 7705 7870 7751 7882
rect 7705 7836 7711 7870
rect 7745 7836 7751 7870
rect 7705 7824 7751 7836
rect 7711 7742 7745 7824
rect 7705 7730 7751 7742
rect 7705 7696 7711 7730
rect 7745 7696 7751 7730
rect 7705 7684 7751 7696
rect 7711 7602 7745 7684
rect 7705 7590 7751 7602
rect 7705 7556 7711 7590
rect 7745 7556 7751 7590
rect 7705 7544 7751 7556
rect 7711 7462 7745 7544
rect 7705 7450 7751 7462
rect 7705 7416 7711 7450
rect 7745 7416 7751 7450
rect 7705 7404 7751 7416
rect 7711 7322 7745 7404
rect 7705 7310 7751 7322
rect 7705 7276 7711 7310
rect 7745 7276 7751 7310
rect 7705 7264 7751 7276
rect 7711 7182 7745 7264
rect 7705 7170 7751 7182
rect 7705 7136 7711 7170
rect 7745 7136 7751 7170
rect 7705 7124 7751 7136
rect 7711 7114 7745 7124
rect 7711 6815 7745 6823
rect 7702 6809 7754 6815
rect 7702 6751 7754 6757
rect 7711 6672 7745 6751
rect 7705 6660 7751 6672
rect 7705 6626 7711 6660
rect 7745 6626 7751 6660
rect 7705 6614 7751 6626
rect 7711 6532 7745 6614
rect 7705 6520 7751 6532
rect 7705 6486 7711 6520
rect 7745 6486 7751 6520
rect 7705 6474 7751 6486
rect 7711 6392 7745 6474
rect 7705 6380 7751 6392
rect 7705 6346 7711 6380
rect 7745 6346 7751 6380
rect 7705 6334 7751 6346
rect 7711 6252 7745 6334
rect 7705 6240 7751 6252
rect 7705 6206 7711 6240
rect 7745 6206 7751 6240
rect 7705 6194 7751 6206
rect 7711 6112 7745 6194
rect 7705 6100 7751 6112
rect 7705 6066 7711 6100
rect 7745 6066 7751 6100
rect 7705 6054 7751 6066
rect 7711 5972 7745 6054
rect 7705 5960 7751 5972
rect 7705 5926 7711 5960
rect 7745 5926 7751 5960
rect 7705 5914 7751 5926
rect 7711 5832 7745 5914
rect 7705 5820 7751 5832
rect 7705 5786 7711 5820
rect 7745 5786 7751 5820
rect 7705 5774 7751 5786
rect 7711 5764 7745 5774
rect 7711 5605 7745 5613
rect 7702 5599 7754 5605
rect 7702 5541 7754 5547
rect 7711 5462 7745 5541
rect 7705 5450 7751 5462
rect 7705 5416 7711 5450
rect 7745 5416 7751 5450
rect 7705 5404 7751 5416
rect 7711 5322 7745 5404
rect 7705 5310 7751 5322
rect 7705 5276 7711 5310
rect 7745 5276 7751 5310
rect 7705 5264 7751 5276
rect 7711 5182 7745 5264
rect 7705 5170 7751 5182
rect 7705 5136 7711 5170
rect 7745 5136 7751 5170
rect 7705 5124 7751 5136
rect 7711 5042 7745 5124
rect 7705 5030 7751 5042
rect 7705 4996 7711 5030
rect 7745 4996 7751 5030
rect 7705 4984 7751 4996
rect 7711 4902 7745 4984
rect 7705 4890 7751 4902
rect 7705 4856 7711 4890
rect 7745 4856 7751 4890
rect 7705 4844 7751 4856
rect 7711 4762 7745 4844
rect 7705 4750 7751 4762
rect 7705 4716 7711 4750
rect 7745 4716 7751 4750
rect 7705 4704 7751 4716
rect 7711 4622 7745 4704
rect 7705 4610 7751 4622
rect 7705 4576 7711 4610
rect 7745 4576 7751 4610
rect 7705 4564 7751 4576
rect 7711 4554 7745 4564
rect 7711 4395 7745 4403
rect 7702 4389 7754 4395
rect 7702 4331 7754 4337
rect 7711 4252 7745 4331
rect 7705 4240 7751 4252
rect 7705 4206 7711 4240
rect 7745 4206 7751 4240
rect 7705 4194 7751 4206
rect 7711 4112 7745 4194
rect 7705 4100 7751 4112
rect 7705 4066 7711 4100
rect 7745 4066 7751 4100
rect 7705 4054 7751 4066
rect 7711 3972 7745 4054
rect 7705 3960 7751 3972
rect 7705 3926 7711 3960
rect 7745 3926 7751 3960
rect 7705 3914 7751 3926
rect 7711 3832 7745 3914
rect 7705 3820 7751 3832
rect 7705 3786 7711 3820
rect 7745 3786 7751 3820
rect 7705 3774 7751 3786
rect 7711 3692 7745 3774
rect 7705 3680 7751 3692
rect 7705 3646 7711 3680
rect 7745 3646 7751 3680
rect 7705 3634 7751 3646
rect 7711 3552 7745 3634
rect 7705 3540 7751 3552
rect 7705 3506 7711 3540
rect 7745 3506 7751 3540
rect 7705 3494 7751 3506
rect 7711 3412 7745 3494
rect 7705 3400 7751 3412
rect 7705 3366 7711 3400
rect 7745 3366 7751 3400
rect 7705 3354 7751 3366
rect 7711 3344 7745 3354
rect 7711 3185 7745 3193
rect 7702 3179 7754 3185
rect 7702 3121 7754 3127
rect 7711 3042 7745 3121
rect 7705 3030 7751 3042
rect 7705 2996 7711 3030
rect 7745 2996 7751 3030
rect 7705 2984 7751 2996
rect 7711 2902 7745 2984
rect 8020 2943 8054 11833
rect 8800 11667 8806 11719
rect 8874 11667 8880 11719
rect 8800 10457 8806 10509
rect 8874 10457 8880 10509
rect 8800 9247 8806 9299
rect 8874 9247 8880 9299
rect 8800 8037 8806 8089
rect 8874 8037 8880 8089
rect 8800 6687 8806 6739
rect 8874 6687 8880 6739
rect 8800 5477 8806 5529
rect 8874 5477 8880 5529
rect 8800 4267 8806 4319
rect 8874 4267 8880 4319
rect 8800 3057 8806 3109
rect 8874 3057 8880 3109
rect 7705 2890 7751 2902
rect 7705 2856 7711 2890
rect 7745 2856 7751 2890
rect 7705 2844 7751 2856
rect 7711 2762 7745 2844
rect 7705 2750 7751 2762
rect 7705 2716 7711 2750
rect 7745 2716 7751 2750
rect 7705 2704 7751 2716
rect 7711 2622 7745 2704
rect 7705 2610 7751 2622
rect 7705 2576 7711 2610
rect 7745 2576 7751 2610
rect 7705 2564 7751 2576
rect 7711 2482 7745 2564
rect 7705 2470 7751 2482
rect 7705 2436 7711 2470
rect 7745 2436 7751 2470
rect 7705 2424 7751 2436
rect 7711 2342 7745 2424
rect 7705 2330 7751 2342
rect 7705 2296 7711 2330
rect 7745 2296 7751 2330
rect 7705 2284 7751 2296
rect 7711 2202 7745 2284
rect 7705 2190 7751 2202
rect 7705 2156 7711 2190
rect 7745 2156 7751 2190
rect 7705 2144 7751 2156
rect 7711 2134 7745 2144
rect 41 1803 157 1833
rect 6611 1803 6727 1833
rect 41 1381 71 1803
rect 6697 1381 6727 1803
rect 41 1351 101 1381
rect 6667 1351 6727 1381
rect 6839 1203 6869 2013
rect 6899 1303 6929 2013
rect 7129 1403 7159 2013
rect 7229 1503 7259 2013
rect 7329 1603 7359 2013
rect 7429 1703 7459 2013
rect 7529 1803 7559 2013
rect 7629 1887 7659 2013
rect 8190 1887 8249 1903
rect 7629 1873 8249 1887
rect 7629 1857 8220 1873
rect 7529 1773 8249 1803
rect 7429 1673 8249 1703
rect 7329 1573 8249 1603
rect 7229 1473 8249 1503
rect 7129 1373 8249 1403
rect 6899 1273 8249 1303
rect 6839 1173 8249 1203
rect 6625 1073 8249 1103
rect 6625 973 8249 1003
rect 6625 873 8249 903
rect 6625 773 8249 803
rect 6625 673 8249 703
rect 6625 573 8249 603
rect 6625 473 8249 503
rect 6625 373 8249 403
rect 6625 273 8249 303
rect 6625 173 8249 203
rect 11 90 211 96
rect 11 32 17 90
rect 205 32 211 90
rect 11 26 211 32
rect 6557 90 6757 96
rect 6557 32 6563 90
rect 6751 32 6757 90
rect 6557 26 6757 32
<< via1 >>
rect 7702 11780 7754 11789
rect 7702 11746 7711 11780
rect 7711 11746 7745 11780
rect 7745 11746 7754 11780
rect 7702 11737 7754 11746
rect 7702 10570 7754 10579
rect 7702 10536 7711 10570
rect 7711 10536 7745 10570
rect 7745 10536 7754 10570
rect 7702 10527 7754 10536
rect 7702 9360 7754 9369
rect 7702 9326 7711 9360
rect 7711 9326 7745 9360
rect 7745 9326 7754 9360
rect 7702 9317 7754 9326
rect 7702 8150 7754 8159
rect 7702 8116 7711 8150
rect 7711 8116 7745 8150
rect 7745 8116 7754 8150
rect 7702 8107 7754 8116
rect 7702 6800 7754 6809
rect 7702 6766 7711 6800
rect 7711 6766 7745 6800
rect 7745 6766 7754 6800
rect 7702 6757 7754 6766
rect 7702 5590 7754 5599
rect 7702 5556 7711 5590
rect 7711 5556 7745 5590
rect 7745 5556 7754 5590
rect 7702 5547 7754 5556
rect 7702 4380 7754 4389
rect 7702 4346 7711 4380
rect 7711 4346 7745 4380
rect 7745 4346 7754 4380
rect 7702 4337 7754 4346
rect 7702 3170 7754 3179
rect 7702 3136 7711 3170
rect 7711 3136 7745 3170
rect 7745 3136 7754 3170
rect 7702 3127 7754 3136
rect 8806 11667 8874 11719
rect 8806 10457 8874 10509
rect 8806 9247 8874 9299
rect 8806 8037 8874 8089
rect 8806 6687 8874 6739
rect 8806 5477 8874 5529
rect 8806 4267 8874 4319
rect 8806 3057 8874 3109
rect 17 32 205 90
rect 6563 32 6751 90
<< metal2 >>
rect 7702 11789 7754 11795
rect 7702 11716 7754 11737
rect 7702 11670 8000 11716
rect 8800 11667 8806 11719
rect 8874 11667 9780 11719
rect 7702 10579 7754 10585
rect 7702 10506 7754 10527
rect 7702 10460 8000 10506
rect 8800 10457 8806 10509
rect 8874 10457 9780 10509
rect 7702 9369 7754 9375
rect 7702 9296 7754 9317
rect 7702 9250 8000 9296
rect 8800 9247 8806 9299
rect 8874 9247 9780 9299
rect 7702 8159 7754 8165
rect 7702 8086 7754 8107
rect 7702 8040 8000 8086
rect 8800 8037 8806 8089
rect 8874 8037 9780 8089
rect 7702 6809 7754 6815
rect 7702 6736 7754 6757
rect 7702 6690 8000 6736
rect 8800 6687 8806 6739
rect 8874 6687 9780 6739
rect 7702 5599 7754 5605
rect 7702 5526 7754 5547
rect 7702 5480 8000 5526
rect 8800 5477 8806 5529
rect 8874 5477 9780 5529
rect 7702 4389 7754 4395
rect 7702 4316 7754 4337
rect 7702 4270 8000 4316
rect 8800 4267 8806 4319
rect 8874 4267 9780 4319
rect 7702 3179 7754 3185
rect 7702 3106 7754 3127
rect 7702 3060 8000 3106
rect 8800 3057 8806 3109
rect 8874 3057 9780 3109
rect 8017 2103 8026 2253
rect 8265 2248 9395 2253
rect 8265 2108 8654 2248
rect 9386 2108 9395 2248
rect 8265 2103 9395 2108
rect 11 1334 111 1903
rect 11 1094 16 1334
rect 106 1094 111 1334
rect 11 96 111 1094
rect 6657 1868 6857 1903
rect 6657 1778 6676 1868
rect 6852 1778 6857 1868
rect 9689 1862 9780 1914
rect 6657 1334 6857 1778
rect 9689 1662 9780 1714
rect 9689 1462 9780 1514
rect 6657 1094 6662 1334
rect 6852 1094 6857 1334
rect 9689 1262 9780 1314
rect 6657 1085 6857 1094
rect 6657 96 6757 1085
rect 9689 1062 9780 1114
rect 9689 862 9780 914
rect 9689 662 9780 714
rect 9689 462 9780 514
rect 9689 262 9780 314
rect 11 90 211 96
rect 11 32 17 90
rect 205 32 211 90
rect 11 26 211 32
rect 6557 90 6757 96
rect 6557 32 6563 90
rect 6751 32 6757 90
rect 6557 26 6757 32
<< via2 >>
rect 8026 2103 8265 2253
rect 8654 2108 9386 2248
rect 16 1094 106 1334
rect 6676 1778 6852 1868
rect 6662 1094 6852 1334
<< metal3 >>
rect 8275 2902 8543 11833
rect 8021 2653 8543 2902
rect 8021 2253 8270 2653
rect 8659 2553 8769 11833
rect 8021 2103 8026 2253
rect 8265 2103 8270 2253
rect 111 1868 6857 1873
rect 111 1778 6676 1868
rect 6852 1778 6857 1868
rect 111 1773 6857 1778
rect 8021 1689 8270 2103
rect 8370 2353 9670 2553
rect 8370 2053 8551 2353
rect 8649 2248 9391 2253
rect 8649 2108 8654 2248
rect 9386 2108 9391 2248
rect 8649 2053 9391 2108
rect 9489 2053 9670 2353
rect 151 1439 8270 1689
rect 11 1334 8370 1339
rect 11 1094 16 1334
rect 106 1094 6662 1334
rect 6852 1094 8370 1334
rect 11 1089 8370 1094
use out_drive  out_drive_0
timestamp 1728730538
transform 1 0 3300 0 1 11413
box 4700 -55 5500 474
use out_drive  out_drive_1
timestamp 1728730538
transform 1 0 3300 0 1 2803
box 4700 -55 5500 474
use out_drive  out_drive_2
timestamp 1728730538
transform 1 0 3300 0 1 4013
box 4700 -55 5500 474
use out_drive  out_drive_3
timestamp 1728730538
transform 1 0 3300 0 1 5223
box 4700 -55 5500 474
use out_drive  out_drive_4
timestamp 1728730538
transform 1 0 3300 0 1 6433
box 4700 -55 5500 474
use out_drive  out_drive_5
timestamp 1728730538
transform 1 0 3300 0 1 7783
box 4700 -55 5500 474
use out_drive  out_drive_6
timestamp 1728730538
transform 1 0 3300 0 1 8993
box 4700 -55 5500 474
use out_drive  out_drive_7
timestamp 1728730538
transform 1 0 3300 0 1 10203
box 4700 -55 5500 474
use rom_4k_0_core  rom_4k_0_core_0
timestamp 1730660070
transform 1 0 249 0 1 2013
box -169 -2013 9440 10050
<< labels >>
flabel metal3 s 151 1439 8270 1689 0 FreeSans 400 0 0 0 VPWR
port 21 nsew power bidirectional
flabel metal3 s 111 1773 6857 1873 0 FreeSans 400 0 0 0 VGND
port 20 nsew ground bidirectional
flabel metal3 s 11 1089 8551 1339 0 FreeSans 400 0 0 0 VGND
port 20 nsew ground bidirectional
flabel metal2 s 9720 1262 9780 1314 0 FreeSans 160 0 0 0 addr[0]
port 0 nsew signal input
flabel metal2 s 9720 1462 9780 1514 0 FreeSans 160 0 0 0 addr[1]
port 1 nsew signal input
flabel metal2 s 9720 1662 9780 1714 0 FreeSans 160 0 0 0 addr[2]
port 2 nsew signal input
flabel metal2 s 9720 1862 9780 1914 0 FreeSans 160 0 0 0 addr[3]
port 3 nsew signal input
flabel metal2 s 9720 1062 9780 1114 0 FreeSans 160 0 0 0 addr[4]
port 5 nsew signal input
flabel metal2 s 9720 862 9780 914 0 FreeSans 160 0 0 0 addr[5]
port 6 nsew signal input
flabel metal2 s 9720 662 9780 714 0 FreeSans 160 0 0 0 addr[6]
port 7 nsew signal input
flabel metal2 s 9720 462 9780 514 0 FreeSans 160 0 0 0 addr[7]
port 8 nsew signal input
flabel metal2 s 9720 262 9780 314 0 FreeSans 160 0 0 0 addr[8]
port 9 nsew signal input
flabel metal2 s 9720 3057 9780 3109 0 FreeSans 160 0 0 0 q[0]
port 12 nsew signal output
flabel metal2 s 9720 4267 9780 4319 0 FreeSans 160 0 0 0 q[1]
port 13 nsew signal output
flabel metal2 s 9720 5477 9780 5529 0 FreeSans 160 0 0 0 q[2]
port 14 nsew signal output
flabel metal2 s 9720 6687 9780 6739 0 FreeSans 160 0 0 0 q[3]
port 15 nsew signal output
flabel metal2 s 9720 8037 9780 8089 0 FreeSans 160 0 0 0 q[4]
port 16 nsew signal output
flabel metal2 s 9720 9247 9780 9299 0 FreeSans 160 0 0 0 q[5]
port 17 nsew signal output
flabel metal2 s 9720 10457 9780 10509 0 FreeSans 160 0 0 0 q[6]
port 18 nsew signal output
flabel metal2 s 9720 11667 9780 11719 0 FreeSans 160 0 0 0 q[7]
port 19 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 9780 12063
<< end >>
