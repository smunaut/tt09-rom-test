magic
tech sky130A
magscale 1 2
timestamp 1730660070
<< nwell >>
rect -169 -778 12839 -294
rect 14780 -2173 15562 -77
<< pwell >>
rect 90 4839 12780 5067
rect -10 91 13696 4839
rect -10 -1 12836 91
rect -166 -87 12836 -1
rect -120 -236 12790 -87
rect -36 -2213 12706 -820
rect 14514 -2163 14716 -87
rect 15626 -2163 15828 -87
<< nmos >>
rect -30 -210 0 -126
rect 70 -210 100 -126
rect 170 -210 200 -126
rect 270 -210 300 -126
rect 370 -210 400 -126
rect 470 -210 500 -126
rect 570 -210 600 -126
rect 670 -210 700 -126
rect 770 -210 800 -126
rect 870 -210 900 -126
rect 970 -210 1000 -126
rect 1070 -210 1100 -126
rect 1170 -210 1200 -126
rect 1270 -210 1300 -126
rect 1370 -210 1400 -126
rect 1470 -210 1500 -126
rect 1570 -210 1600 -126
rect 1670 -210 1700 -126
rect 1770 -210 1800 -126
rect 1870 -210 1900 -126
rect 1970 -210 2000 -126
rect 2070 -210 2100 -126
rect 2170 -210 2200 -126
rect 2270 -210 2300 -126
rect 2370 -210 2400 -126
rect 2470 -210 2500 -126
rect 2570 -210 2600 -126
rect 2670 -210 2700 -126
rect 2770 -210 2800 -126
rect 2870 -210 2900 -126
rect 2970 -210 3000 -126
rect 3070 -210 3100 -126
rect 3170 -210 3200 -126
rect 3270 -210 3300 -126
rect 3370 -210 3400 -126
rect 3470 -210 3500 -126
rect 3570 -210 3600 -126
rect 3670 -210 3700 -126
rect 3770 -210 3800 -126
rect 3870 -210 3900 -126
rect 3970 -210 4000 -126
rect 4070 -210 4100 -126
rect 4170 -210 4200 -126
rect 4270 -210 4300 -126
rect 4370 -210 4400 -126
rect 4470 -210 4500 -126
rect 4570 -210 4600 -126
rect 4670 -210 4700 -126
rect 4770 -210 4800 -126
rect 4870 -210 4900 -126
rect 4970 -210 5000 -126
rect 5070 -210 5100 -126
rect 5170 -210 5200 -126
rect 5270 -210 5300 -126
rect 5370 -210 5400 -126
rect 5470 -210 5500 -126
rect 5570 -210 5600 -126
rect 5670 -210 5700 -126
rect 5770 -210 5800 -126
rect 5870 -210 5900 -126
rect 5970 -210 6000 -126
rect 6070 -210 6100 -126
rect 6170 -210 6200 -126
rect 6270 -210 6300 -126
rect 6370 -210 6400 -126
rect 6470 -210 6500 -126
rect 6570 -210 6600 -126
rect 6670 -210 6700 -126
rect 6770 -210 6800 -126
rect 6870 -210 6900 -126
rect 6970 -210 7000 -126
rect 7070 -210 7100 -126
rect 7170 -210 7200 -126
rect 7270 -210 7300 -126
rect 7370 -210 7400 -126
rect 7470 -210 7500 -126
rect 7570 -210 7600 -126
rect 7670 -210 7700 -126
rect 7770 -210 7800 -126
rect 7870 -210 7900 -126
rect 7970 -210 8000 -126
rect 8070 -210 8100 -126
rect 8170 -210 8200 -126
rect 8270 -210 8300 -126
rect 8370 -210 8400 -126
rect 8470 -210 8500 -126
rect 8570 -210 8600 -126
rect 8670 -210 8700 -126
rect 8770 -210 8800 -126
rect 8870 -210 8900 -126
rect 8970 -210 9000 -126
rect 9070 -210 9100 -126
rect 9170 -210 9200 -126
rect 9270 -210 9300 -126
rect 9370 -210 9400 -126
rect 9470 -210 9500 -126
rect 9570 -210 9600 -126
rect 9670 -210 9700 -126
rect 9770 -210 9800 -126
rect 9870 -210 9900 -126
rect 9970 -210 10000 -126
rect 10070 -210 10100 -126
rect 10170 -210 10200 -126
rect 10270 -210 10300 -126
rect 10370 -210 10400 -126
rect 10470 -210 10500 -126
rect 10570 -210 10600 -126
rect 10670 -210 10700 -126
rect 10770 -210 10800 -126
rect 10870 -210 10900 -126
rect 10970 -210 11000 -126
rect 11070 -210 11100 -126
rect 11170 -210 11200 -126
rect 11270 -210 11300 -126
rect 11370 -210 11400 -126
rect 11470 -210 11500 -126
rect 11570 -210 11600 -126
rect 11670 -210 11700 -126
rect 11770 -210 11800 -126
rect 11870 -210 11900 -126
rect 11970 -210 12000 -126
rect 12070 -210 12100 -126
rect 12170 -210 12200 -126
rect 12270 -210 12300 -126
rect 12370 -210 12400 -126
rect 12470 -210 12500 -126
rect 12570 -210 12600 -126
rect 12670 -210 12700 -126
rect 14540 -290 14690 -260
rect 15652 -290 15802 -260
rect 14540 -390 14690 -360
rect 15652 -390 15802 -360
rect 14540 -490 14690 -460
rect 15652 -490 15802 -460
rect 14540 -590 14690 -560
rect 15652 -590 15802 -560
rect 14540 -690 14690 -660
rect 15652 -690 15802 -660
rect 14540 -790 14690 -760
rect 15652 -790 15802 -760
rect 14540 -890 14690 -860
rect 15652 -890 15802 -860
rect 14540 -990 14690 -960
rect 15652 -990 15802 -960
rect 14540 -1090 14690 -1060
rect 15652 -1090 15802 -1060
rect 14540 -1190 14690 -1160
rect 15652 -1190 15802 -1160
rect 14540 -1290 14690 -1260
rect 15652 -1290 15802 -1260
rect 14540 -1390 14690 -1360
rect 15652 -1390 15802 -1360
rect 14540 -1490 14690 -1460
rect 15652 -1490 15802 -1460
rect 14540 -1590 14690 -1560
rect 15652 -1590 15802 -1560
rect 14540 -1690 14690 -1660
rect 15652 -1690 15802 -1660
rect 14540 -1790 14690 -1760
rect 15652 -1790 15802 -1760
rect 14540 -1890 14690 -1860
rect 15652 -1890 15802 -1860
rect 14540 -1990 14690 -1960
rect 15652 -1990 15802 -1960
<< pmos >>
rect 14816 -290 15116 -260
rect 15226 -290 15526 -260
rect 14816 -390 15116 -360
rect 15226 -390 15526 -360
rect 14816 -490 15116 -460
rect 15226 -490 15526 -460
rect 14816 -590 15116 -560
rect 15226 -590 15526 -560
rect 15 -742 107 -658
rect 163 -742 255 -658
rect 415 -742 507 -658
rect 563 -742 655 -658
rect 815 -742 907 -658
rect 963 -742 1055 -658
rect 1215 -742 1307 -658
rect 1363 -742 1455 -658
rect 1615 -742 1707 -658
rect 1763 -742 1855 -658
rect 2015 -742 2107 -658
rect 2163 -742 2255 -658
rect 2415 -742 2507 -658
rect 2563 -742 2655 -658
rect 2815 -742 2907 -658
rect 2963 -742 3055 -658
rect 3215 -742 3307 -658
rect 3363 -742 3455 -658
rect 3615 -742 3707 -658
rect 3763 -742 3855 -658
rect 4015 -742 4107 -658
rect 4163 -742 4255 -658
rect 4415 -742 4507 -658
rect 4563 -742 4655 -658
rect 4815 -742 4907 -658
rect 4963 -742 5055 -658
rect 5215 -742 5307 -658
rect 5363 -742 5455 -658
rect 5615 -742 5707 -658
rect 5763 -742 5855 -658
rect 6015 -742 6107 -658
rect 6163 -742 6255 -658
rect 6415 -742 6507 -658
rect 6563 -742 6655 -658
rect 6815 -742 6907 -658
rect 6963 -742 7055 -658
rect 7215 -742 7307 -658
rect 7363 -742 7455 -658
rect 7615 -742 7707 -658
rect 7763 -742 7855 -658
rect 8015 -742 8107 -658
rect 8163 -742 8255 -658
rect 8415 -742 8507 -658
rect 8563 -742 8655 -658
rect 8815 -742 8907 -658
rect 8963 -742 9055 -658
rect 9215 -742 9307 -658
rect 9363 -742 9455 -658
rect 9615 -742 9707 -658
rect 9763 -742 9855 -658
rect 10015 -742 10107 -658
rect 10163 -742 10255 -658
rect 10415 -742 10507 -658
rect 10563 -742 10655 -658
rect 10815 -742 10907 -658
rect 10963 -742 11055 -658
rect 11215 -742 11307 -658
rect 11363 -742 11455 -658
rect 11615 -742 11707 -658
rect 11763 -742 11855 -658
rect 12015 -742 12107 -658
rect 12163 -742 12255 -658
rect 12415 -742 12507 -658
rect 12563 -742 12655 -658
rect 14816 -690 15116 -660
rect 15226 -690 15526 -660
rect 14816 -790 15116 -760
rect 15226 -790 15526 -760
rect 14816 -890 15116 -860
rect 15226 -890 15526 -860
rect 14816 -990 15116 -960
rect 15226 -990 15526 -960
rect 14816 -1090 15116 -1060
rect 15226 -1090 15526 -1060
rect 14816 -1190 15116 -1160
rect 15226 -1190 15526 -1160
rect 14816 -1290 15116 -1260
rect 15226 -1290 15526 -1260
rect 14816 -1390 15116 -1360
rect 15226 -1390 15526 -1360
rect 14816 -1490 15116 -1460
rect 15226 -1490 15526 -1460
rect 14816 -1590 15116 -1560
rect 15226 -1590 15526 -1560
rect 14816 -1690 15116 -1660
rect 15226 -1690 15526 -1660
rect 14816 -1790 15116 -1760
rect 15226 -1790 15526 -1760
rect 14816 -1890 15116 -1860
rect 15226 -1890 15526 -1860
rect 14816 -1990 15116 -1960
rect 15226 -1990 15526 -1960
<< pmoshvt >>
rect -30 -498 0 -330
rect 70 -498 100 -330
rect 170 -498 200 -330
rect 270 -498 300 -330
rect 370 -498 400 -330
rect 470 -498 500 -330
rect 570 -498 600 -330
rect 670 -498 700 -330
rect 770 -498 800 -330
rect 870 -498 900 -330
rect 970 -498 1000 -330
rect 1070 -498 1100 -330
rect 1170 -498 1200 -330
rect 1270 -498 1300 -330
rect 1370 -498 1400 -330
rect 1470 -498 1500 -330
rect 1570 -498 1600 -330
rect 1670 -498 1700 -330
rect 1770 -498 1800 -330
rect 1870 -498 1900 -330
rect 1970 -498 2000 -330
rect 2070 -498 2100 -330
rect 2170 -498 2200 -330
rect 2270 -498 2300 -330
rect 2370 -498 2400 -330
rect 2470 -498 2500 -330
rect 2570 -498 2600 -330
rect 2670 -498 2700 -330
rect 2770 -498 2800 -330
rect 2870 -498 2900 -330
rect 2970 -498 3000 -330
rect 3070 -498 3100 -330
rect 3170 -498 3200 -330
rect 3270 -498 3300 -330
rect 3370 -498 3400 -330
rect 3470 -498 3500 -330
rect 3570 -498 3600 -330
rect 3670 -498 3700 -330
rect 3770 -498 3800 -330
rect 3870 -498 3900 -330
rect 3970 -498 4000 -330
rect 4070 -498 4100 -330
rect 4170 -498 4200 -330
rect 4270 -498 4300 -330
rect 4370 -498 4400 -330
rect 4470 -498 4500 -330
rect 4570 -498 4600 -330
rect 4670 -498 4700 -330
rect 4770 -498 4800 -330
rect 4870 -498 4900 -330
rect 4970 -498 5000 -330
rect 5070 -498 5100 -330
rect 5170 -498 5200 -330
rect 5270 -498 5300 -330
rect 5370 -498 5400 -330
rect 5470 -498 5500 -330
rect 5570 -498 5600 -330
rect 5670 -498 5700 -330
rect 5770 -498 5800 -330
rect 5870 -498 5900 -330
rect 5970 -498 6000 -330
rect 6070 -498 6100 -330
rect 6170 -498 6200 -330
rect 6270 -498 6300 -330
rect 6370 -498 6400 -330
rect 6470 -498 6500 -330
rect 6570 -498 6600 -330
rect 6670 -498 6700 -330
rect 6770 -498 6800 -330
rect 6870 -498 6900 -330
rect 6970 -498 7000 -330
rect 7070 -498 7100 -330
rect 7170 -498 7200 -330
rect 7270 -498 7300 -330
rect 7370 -498 7400 -330
rect 7470 -498 7500 -330
rect 7570 -498 7600 -330
rect 7670 -498 7700 -330
rect 7770 -498 7800 -330
rect 7870 -498 7900 -330
rect 7970 -498 8000 -330
rect 8070 -498 8100 -330
rect 8170 -498 8200 -330
rect 8270 -498 8300 -330
rect 8370 -498 8400 -330
rect 8470 -498 8500 -330
rect 8570 -498 8600 -330
rect 8670 -498 8700 -330
rect 8770 -498 8800 -330
rect 8870 -498 8900 -330
rect 8970 -498 9000 -330
rect 9070 -498 9100 -330
rect 9170 -498 9200 -330
rect 9270 -498 9300 -330
rect 9370 -498 9400 -330
rect 9470 -498 9500 -330
rect 9570 -498 9600 -330
rect 9670 -498 9700 -330
rect 9770 -498 9800 -330
rect 9870 -498 9900 -330
rect 9970 -498 10000 -330
rect 10070 -498 10100 -330
rect 10170 -498 10200 -330
rect 10270 -498 10300 -330
rect 10370 -498 10400 -330
rect 10470 -498 10500 -330
rect 10570 -498 10600 -330
rect 10670 -498 10700 -330
rect 10770 -498 10800 -330
rect 10870 -498 10900 -330
rect 10970 -498 11000 -330
rect 11070 -498 11100 -330
rect 11170 -498 11200 -330
rect 11270 -498 11300 -330
rect 11370 -498 11400 -330
rect 11470 -498 11500 -330
rect 11570 -498 11600 -330
rect 11670 -498 11700 -330
rect 11770 -498 11800 -330
rect 11870 -498 11900 -330
rect 11970 -498 12000 -330
rect 12070 -498 12100 -330
rect 12170 -498 12200 -330
rect 12270 -498 12300 -330
rect 12370 -498 12400 -330
rect 12470 -498 12500 -330
rect 12570 -498 12600 -330
rect 12670 -498 12700 -330
<< nmoslvt >>
rect 70 4727 100 4813
rect 170 4727 200 4813
rect 270 4727 300 4813
rect 470 4727 500 4813
rect 570 4727 600 4813
rect 670 4727 700 4813
rect 770 4727 800 4813
rect 870 4727 900 4813
rect 970 4727 1000 4813
rect 1070 4727 1100 4813
rect 70 4587 100 4673
rect 170 4587 200 4673
rect 270 4587 300 4673
rect 370 4587 400 4673
rect 470 4587 500 4673
rect 570 4587 600 4673
rect 670 4587 700 4673
rect 770 4587 800 4673
rect 870 4587 900 4673
rect 970 4587 1000 4673
rect 1070 4587 1100 4673
rect 70 4447 100 4533
rect 170 4447 200 4533
rect 270 4447 300 4533
rect 1270 4727 1300 4813
rect 1370 4727 1400 4813
rect 1470 4727 1500 4813
rect 1570 4727 1600 4813
rect 1670 4727 1700 4813
rect 1770 4727 1800 4813
rect 1870 4727 1900 4813
rect 1970 4727 2000 4813
rect 2070 4727 2100 4813
rect 2170 4727 2200 4813
rect 2270 4727 2300 4813
rect 2470 4727 2500 4813
rect 2570 4727 2600 4813
rect 2670 4727 2700 4813
rect 2770 4727 2800 4813
rect 2870 4727 2900 4813
rect 2970 4727 3000 4813
rect 3070 4727 3100 4813
rect 1270 4587 1300 4673
rect 1370 4587 1400 4673
rect 1470 4587 1500 4673
rect 1570 4587 1600 4673
rect 1670 4587 1700 4673
rect 1770 4587 1800 4673
rect 1870 4587 1900 4673
rect 1970 4587 2000 4673
rect 2070 4587 2100 4673
rect 2170 4587 2200 4673
rect 2270 4587 2300 4673
rect 2370 4587 2400 4673
rect 2470 4587 2500 4673
rect 2570 4587 2600 4673
rect 2670 4587 2700 4673
rect 2770 4587 2800 4673
rect 2870 4587 2900 4673
rect 470 4447 500 4533
rect 570 4447 600 4533
rect 670 4447 700 4533
rect 770 4447 800 4533
rect 870 4447 900 4533
rect 970 4447 1000 4533
rect 1070 4447 1100 4533
rect 1170 4447 1200 4533
rect 1270 4447 1300 4533
rect 1370 4447 1400 4533
rect 1470 4447 1500 4533
rect 1570 4447 1600 4533
rect 70 4307 100 4393
rect 170 4307 200 4393
rect 270 4307 300 4393
rect 370 4307 400 4393
rect 470 4307 500 4393
rect 570 4307 600 4393
rect 670 4307 700 4393
rect 770 4307 800 4393
rect 870 4307 900 4393
rect 970 4307 1000 4393
rect 1070 4307 1100 4393
rect 1170 4307 1200 4393
rect 70 4167 100 4253
rect 170 4167 200 4253
rect 270 4167 300 4253
rect 370 4167 400 4253
rect 470 4167 500 4253
rect 70 4027 100 4113
rect 170 4027 200 4113
rect 370 4027 400 4113
rect 670 4167 700 4253
rect 770 4167 800 4253
rect 870 4167 900 4253
rect 970 4167 1000 4253
rect 1070 4167 1100 4253
rect 1770 4447 1800 4533
rect 1970 4447 2000 4533
rect 2070 4447 2100 4533
rect 2170 4447 2200 4533
rect 2270 4447 2300 4533
rect 1370 4307 1400 4393
rect 1470 4307 1500 4393
rect 1570 4307 1600 4393
rect 1670 4307 1700 4393
rect 1770 4307 1800 4393
rect 1870 4307 1900 4393
rect 1270 4167 1300 4253
rect 1370 4167 1400 4253
rect 1470 4167 1500 4253
rect 1570 4167 1600 4253
rect 1670 4167 1700 4253
rect 1770 4167 1800 4253
rect 1870 4167 1900 4253
rect 570 4027 600 4113
rect 670 4027 700 4113
rect 770 4027 800 4113
rect 870 4027 900 4113
rect 970 4027 1000 4113
rect 1070 4027 1100 4113
rect 1170 4027 1200 4113
rect 1270 4027 1300 4113
rect 1470 4027 1500 4113
rect 1570 4027 1600 4113
rect 2470 4447 2500 4533
rect 2570 4447 2600 4533
rect 2770 4447 2800 4533
rect 3270 4727 3300 4813
rect 3370 4727 3400 4813
rect 3570 4727 3600 4813
rect 3670 4727 3700 4813
rect 3770 4727 3800 4813
rect 3870 4727 3900 4813
rect 3970 4727 4000 4813
rect 4070 4727 4100 4813
rect 4170 4727 4200 4813
rect 3070 4587 3100 4673
rect 3170 4587 3200 4673
rect 3270 4587 3300 4673
rect 3370 4587 3400 4673
rect 3470 4587 3500 4673
rect 3570 4587 3600 4673
rect 4370 4727 4400 4813
rect 4470 4727 4500 4813
rect 4570 4727 4600 4813
rect 4670 4727 4700 4813
rect 4770 4727 4800 4813
rect 4870 4727 4900 4813
rect 4970 4727 5000 4813
rect 5070 4727 5100 4813
rect 5170 4727 5200 4813
rect 5270 4727 5300 4813
rect 5370 4727 5400 4813
rect 5470 4727 5500 4813
rect 5570 4727 5600 4813
rect 5670 4727 5700 4813
rect 5770 4727 5800 4813
rect 5870 4727 5900 4813
rect 5970 4727 6000 4813
rect 6070 4727 6100 4813
rect 6170 4727 6200 4813
rect 6270 4727 6300 4813
rect 6370 4727 6400 4813
rect 3770 4587 3800 4673
rect 3870 4587 3900 4673
rect 3970 4587 4000 4673
rect 4070 4587 4100 4673
rect 4170 4587 4200 4673
rect 4270 4587 4300 4673
rect 4370 4587 4400 4673
rect 4470 4587 4500 4673
rect 4570 4587 4600 4673
rect 4670 4587 4700 4673
rect 2970 4447 3000 4533
rect 3070 4447 3100 4533
rect 3170 4447 3200 4533
rect 3270 4447 3300 4533
rect 3370 4447 3400 4533
rect 3470 4447 3500 4533
rect 3570 4447 3600 4533
rect 3670 4447 3700 4533
rect 2070 4307 2100 4393
rect 2170 4307 2200 4393
rect 2270 4307 2300 4393
rect 2370 4307 2400 4393
rect 2470 4307 2500 4393
rect 2570 4307 2600 4393
rect 2670 4307 2700 4393
rect 2770 4307 2800 4393
rect 2870 4307 2900 4393
rect 2970 4307 3000 4393
rect 3070 4307 3100 4393
rect 3170 4307 3200 4393
rect 3270 4307 3300 4393
rect 3370 4307 3400 4393
rect 3470 4307 3500 4393
rect 3570 4307 3600 4393
rect 3670 4307 3700 4393
rect 4870 4587 4900 4673
rect 4970 4587 5000 4673
rect 3870 4447 3900 4533
rect 3970 4447 4000 4533
rect 4070 4447 4100 4533
rect 4170 4447 4200 4533
rect 4270 4447 4300 4533
rect 4370 4447 4400 4533
rect 4470 4447 4500 4533
rect 4570 4447 4600 4533
rect 4670 4447 4700 4533
rect 4770 4447 4800 4533
rect 4870 4447 4900 4533
rect 4970 4447 5000 4533
rect 5170 4587 5200 4673
rect 5270 4587 5300 4673
rect 5370 4587 5400 4673
rect 5470 4587 5500 4673
rect 5570 4587 5600 4673
rect 5670 4587 5700 4673
rect 5770 4587 5800 4673
rect 5170 4447 5200 4533
rect 5270 4447 5300 4533
rect 5970 4587 6000 4673
rect 6070 4587 6100 4673
rect 6170 4587 6200 4673
rect 6270 4587 6300 4673
rect 6370 4587 6400 4673
rect 5470 4447 5500 4533
rect 5570 4447 5600 4533
rect 5670 4447 5700 4533
rect 5770 4447 5800 4533
rect 5870 4447 5900 4533
rect 5970 4447 6000 4533
rect 3870 4307 3900 4393
rect 3970 4307 4000 4393
rect 4070 4307 4100 4393
rect 4170 4307 4200 4393
rect 4270 4307 4300 4393
rect 4370 4307 4400 4393
rect 4470 4307 4500 4393
rect 4570 4307 4600 4393
rect 4670 4307 4700 4393
rect 4770 4307 4800 4393
rect 4870 4307 4900 4393
rect 4970 4307 5000 4393
rect 5070 4307 5100 4393
rect 5170 4307 5200 4393
rect 5270 4307 5300 4393
rect 5370 4307 5400 4393
rect 5470 4307 5500 4393
rect 5570 4307 5600 4393
rect 5670 4307 5700 4393
rect 5770 4307 5800 4393
rect 5870 4307 5900 4393
rect 5970 4307 6000 4393
rect 2070 4167 2100 4253
rect 2170 4167 2200 4253
rect 2270 4167 2300 4253
rect 2370 4167 2400 4253
rect 2470 4167 2500 4253
rect 2570 4167 2600 4253
rect 2670 4167 2700 4253
rect 2770 4167 2800 4253
rect 2870 4167 2900 4253
rect 2970 4167 3000 4253
rect 3070 4167 3100 4253
rect 3170 4167 3200 4253
rect 3270 4167 3300 4253
rect 3370 4167 3400 4253
rect 3470 4167 3500 4253
rect 3570 4167 3600 4253
rect 3670 4167 3700 4253
rect 3770 4167 3800 4253
rect 3870 4167 3900 4253
rect 3970 4167 4000 4253
rect 1770 4027 1800 4113
rect 1870 4027 1900 4113
rect 1970 4027 2000 4113
rect 2070 4027 2100 4113
rect 2170 4027 2200 4113
rect 70 3887 100 3973
rect 170 3887 200 3973
rect 270 3887 300 3973
rect 370 3887 400 3973
rect 470 3887 500 3973
rect 570 3887 600 3973
rect 670 3887 700 3973
rect 770 3887 800 3973
rect 870 3887 900 3973
rect 970 3887 1000 3973
rect 1070 3887 1100 3973
rect 1170 3887 1200 3973
rect 1270 3887 1300 3973
rect 1370 3887 1400 3973
rect 1470 3887 1500 3973
rect 1570 3887 1600 3973
rect 1670 3887 1700 3973
rect 1770 3887 1800 3973
rect 1870 3887 1900 3973
rect 2370 4027 2400 4113
rect 2470 4027 2500 4113
rect 2570 4027 2600 4113
rect 2770 4027 2800 4113
rect 2870 4027 2900 4113
rect 3070 4027 3100 4113
rect 3170 4027 3200 4113
rect 4170 4167 4200 4253
rect 3370 4027 3400 4113
rect 3470 4027 3500 4113
rect 3570 4027 3600 4113
rect 3670 4027 3700 4113
rect 3770 4027 3800 4113
rect 3870 4027 3900 4113
rect 3970 4027 4000 4113
rect 4070 4027 4100 4113
rect 2070 3887 2100 3973
rect 2170 3887 2200 3973
rect 2270 3887 2300 3973
rect 2370 3887 2400 3973
rect 2470 3887 2500 3973
rect 2570 3887 2600 3973
rect 2670 3887 2700 3973
rect 2770 3887 2800 3973
rect 2870 3887 2900 3973
rect 2970 3887 3000 3973
rect 3070 3887 3100 3973
rect 3170 3887 3200 3973
rect 3270 3887 3300 3973
rect 3370 3887 3400 3973
rect 3470 3887 3500 3973
rect 3570 3887 3600 3973
rect 3670 3887 3700 3973
rect 3770 3887 3800 3973
rect 3870 3887 3900 3973
rect 70 3747 100 3833
rect 170 3747 200 3833
rect 270 3747 300 3833
rect 370 3747 400 3833
rect 470 3747 500 3833
rect 570 3747 600 3833
rect 670 3747 700 3833
rect 770 3747 800 3833
rect 870 3747 900 3833
rect 970 3747 1000 3833
rect 1070 3747 1100 3833
rect 1170 3747 1200 3833
rect 1270 3747 1300 3833
rect 1370 3747 1400 3833
rect 1470 3747 1500 3833
rect 1570 3747 1600 3833
rect 1670 3747 1700 3833
rect 1770 3747 1800 3833
rect 1870 3747 1900 3833
rect 1970 3747 2000 3833
rect 2070 3747 2100 3833
rect 70 3517 100 3603
rect 170 3517 200 3603
rect 270 3517 300 3603
rect 370 3517 400 3603
rect 470 3517 500 3603
rect 570 3517 600 3603
rect 670 3517 700 3603
rect 770 3517 800 3603
rect 70 3377 100 3463
rect 170 3377 200 3463
rect 270 3377 300 3463
rect 470 3377 500 3463
rect 670 3377 700 3463
rect 70 3237 100 3323
rect 170 3237 200 3323
rect 270 3237 300 3323
rect 370 3237 400 3323
rect 470 3237 500 3323
rect 570 3237 600 3323
rect 670 3237 700 3323
rect 70 3097 100 3183
rect 970 3517 1000 3603
rect 870 3377 900 3463
rect 870 3237 900 3323
rect 2270 3747 2300 3833
rect 2370 3747 2400 3833
rect 2470 3747 2500 3833
rect 2670 3747 2700 3833
rect 1170 3517 1200 3603
rect 1270 3517 1300 3603
rect 1370 3517 1400 3603
rect 1470 3517 1500 3603
rect 1570 3517 1600 3603
rect 1670 3517 1700 3603
rect 1770 3517 1800 3603
rect 1870 3517 1900 3603
rect 1970 3517 2000 3603
rect 2070 3517 2100 3603
rect 2170 3517 2200 3603
rect 2270 3517 2300 3603
rect 2370 3517 2400 3603
rect 2470 3517 2500 3603
rect 2870 3747 2900 3833
rect 2970 3747 3000 3833
rect 3070 3747 3100 3833
rect 4070 3887 4100 3973
rect 4370 4167 4400 4253
rect 4270 4027 4300 4113
rect 4570 4167 4600 4253
rect 4470 4027 4500 4113
rect 4770 4167 4800 4253
rect 4670 4027 4700 4113
rect 4970 4167 5000 4253
rect 5070 4167 5100 4253
rect 5170 4167 5200 4253
rect 5270 4167 5300 4253
rect 5370 4167 5400 4253
rect 5470 4167 5500 4253
rect 4870 4027 4900 4113
rect 5070 4027 5100 4113
rect 5170 4027 5200 4113
rect 4270 3887 4300 3973
rect 4370 3887 4400 3973
rect 4470 3887 4500 3973
rect 4570 3887 4600 3973
rect 4670 3887 4700 3973
rect 4770 3887 4800 3973
rect 4870 3887 4900 3973
rect 4970 3887 5000 3973
rect 3270 3747 3300 3833
rect 3370 3747 3400 3833
rect 3470 3747 3500 3833
rect 3570 3747 3600 3833
rect 3670 3747 3700 3833
rect 3770 3747 3800 3833
rect 3870 3747 3900 3833
rect 3970 3747 4000 3833
rect 4070 3747 4100 3833
rect 4170 3747 4200 3833
rect 4270 3747 4300 3833
rect 4370 3747 4400 3833
rect 4470 3747 4500 3833
rect 2670 3517 2700 3603
rect 2770 3517 2800 3603
rect 2870 3517 2900 3603
rect 2970 3517 3000 3603
rect 3070 3517 3100 3603
rect 5170 3887 5200 3973
rect 5670 4167 5700 4253
rect 5770 4167 5800 4253
rect 5870 4167 5900 4253
rect 5970 4167 6000 4253
rect 5370 4027 5400 4113
rect 5470 4027 5500 4113
rect 5570 4027 5600 4113
rect 5370 3887 5400 3973
rect 5470 3887 5500 3973
rect 4670 3747 4700 3833
rect 4770 3747 4800 3833
rect 4870 3747 4900 3833
rect 4970 3747 5000 3833
rect 5070 3747 5100 3833
rect 5170 3747 5200 3833
rect 5270 3747 5300 3833
rect 5370 3747 5400 3833
rect 3270 3517 3300 3603
rect 3370 3517 3400 3603
rect 3470 3517 3500 3603
rect 3570 3517 3600 3603
rect 3670 3517 3700 3603
rect 3770 3517 3800 3603
rect 3870 3517 3900 3603
rect 3970 3517 4000 3603
rect 4070 3517 4100 3603
rect 4170 3517 4200 3603
rect 4270 3517 4300 3603
rect 4370 3517 4400 3603
rect 1070 3377 1100 3463
rect 1170 3377 1200 3463
rect 1270 3377 1300 3463
rect 1370 3377 1400 3463
rect 1470 3377 1500 3463
rect 1570 3377 1600 3463
rect 1670 3377 1700 3463
rect 1770 3377 1800 3463
rect 1870 3377 1900 3463
rect 1970 3377 2000 3463
rect 2070 3377 2100 3463
rect 2170 3377 2200 3463
rect 2270 3377 2300 3463
rect 2370 3377 2400 3463
rect 2470 3377 2500 3463
rect 2570 3377 2600 3463
rect 2670 3377 2700 3463
rect 2770 3377 2800 3463
rect 2870 3377 2900 3463
rect 2970 3377 3000 3463
rect 3070 3377 3100 3463
rect 3170 3377 3200 3463
rect 3270 3377 3300 3463
rect 3370 3377 3400 3463
rect 3470 3377 3500 3463
rect 3570 3377 3600 3463
rect 3670 3377 3700 3463
rect 3770 3377 3800 3463
rect 1070 3237 1100 3323
rect 1170 3237 1200 3323
rect 1270 3237 1300 3323
rect 1370 3237 1400 3323
rect 1470 3237 1500 3323
rect 1570 3237 1600 3323
rect 1670 3237 1700 3323
rect 1770 3237 1800 3323
rect 1870 3237 1900 3323
rect 1970 3237 2000 3323
rect 2070 3237 2100 3323
rect 2170 3237 2200 3323
rect 2270 3237 2300 3323
rect 2370 3237 2400 3323
rect 2470 3237 2500 3323
rect 2570 3237 2600 3323
rect 2670 3237 2700 3323
rect 270 3097 300 3183
rect 370 3097 400 3183
rect 470 3097 500 3183
rect 570 3097 600 3183
rect 670 3097 700 3183
rect 770 3097 800 3183
rect 870 3097 900 3183
rect 970 3097 1000 3183
rect 1070 3097 1100 3183
rect 1170 3097 1200 3183
rect 1270 3097 1300 3183
rect 70 2957 100 3043
rect 170 2957 200 3043
rect 270 2957 300 3043
rect 370 2957 400 3043
rect 470 2957 500 3043
rect 570 2957 600 3043
rect 1470 3097 1500 3183
rect 1570 3097 1600 3183
rect 1670 3097 1700 3183
rect 1770 3097 1800 3183
rect 1870 3097 1900 3183
rect 1970 3097 2000 3183
rect 2070 3097 2100 3183
rect 2170 3097 2200 3183
rect 2270 3097 2300 3183
rect 2370 3097 2400 3183
rect 2470 3097 2500 3183
rect 770 2957 800 3043
rect 870 2957 900 3043
rect 970 2957 1000 3043
rect 1070 2957 1100 3043
rect 1170 2957 1200 3043
rect 1270 2957 1300 3043
rect 1370 2957 1400 3043
rect 1470 2957 1500 3043
rect 1570 2957 1600 3043
rect 1670 2957 1700 3043
rect 1770 2957 1800 3043
rect 1870 2957 1900 3043
rect 1970 2957 2000 3043
rect 70 2817 100 2903
rect 170 2817 200 2903
rect 270 2817 300 2903
rect 370 2817 400 2903
rect 470 2817 500 2903
rect 570 2817 600 2903
rect 670 2817 700 2903
rect 770 2817 800 2903
rect 2870 3237 2900 3323
rect 2970 3237 3000 3323
rect 3070 3237 3100 3323
rect 3170 3237 3200 3323
rect 2670 3097 2700 3183
rect 2770 3097 2800 3183
rect 2870 3097 2900 3183
rect 2970 3097 3000 3183
rect 3070 3097 3100 3183
rect 3170 3097 3200 3183
rect 2170 2957 2200 3043
rect 2270 2957 2300 3043
rect 2370 2957 2400 3043
rect 2470 2957 2500 3043
rect 2570 2957 2600 3043
rect 2670 2957 2700 3043
rect 2770 2957 2800 3043
rect 2870 2957 2900 3043
rect 2970 2957 3000 3043
rect 970 2817 1000 2903
rect 1070 2817 1100 2903
rect 1170 2817 1200 2903
rect 1270 2817 1300 2903
rect 1370 2817 1400 2903
rect 1470 2817 1500 2903
rect 1570 2817 1600 2903
rect 1670 2817 1700 2903
rect 1770 2817 1800 2903
rect 1870 2817 1900 2903
rect 1970 2817 2000 2903
rect 2070 2817 2100 2903
rect 2170 2817 2200 2903
rect 2270 2817 2300 2903
rect 2370 2817 2400 2903
rect 2470 2817 2500 2903
rect 2570 2817 2600 2903
rect 70 2677 100 2763
rect 170 2677 200 2763
rect 270 2677 300 2763
rect 370 2677 400 2763
rect 470 2677 500 2763
rect 570 2677 600 2763
rect 670 2677 700 2763
rect 770 2677 800 2763
rect 870 2677 900 2763
rect 970 2677 1000 2763
rect 1070 2677 1100 2763
rect 1270 2677 1300 2763
rect 1370 2677 1400 2763
rect 1470 2677 1500 2763
rect 1570 2677 1600 2763
rect 1670 2677 1700 2763
rect 1770 2677 1800 2763
rect 1870 2677 1900 2763
rect 1970 2677 2000 2763
rect 2070 2677 2100 2763
rect 2170 2677 2200 2763
rect 2270 2677 2300 2763
rect 2770 2817 2800 2903
rect 2870 2817 2900 2903
rect 3370 3237 3400 3323
rect 3970 3377 4000 3463
rect 4070 3377 4100 3463
rect 4170 3377 4200 3463
rect 4270 3377 4300 3463
rect 4370 3377 4400 3463
rect 6570 4727 6600 4813
rect 6670 4727 6700 4813
rect 6770 4727 6800 4813
rect 6870 4727 6900 4813
rect 6970 4727 7000 4813
rect 7070 4727 7100 4813
rect 7170 4727 7200 4813
rect 7270 4727 7300 4813
rect 7370 4727 7400 4813
rect 7470 4727 7500 4813
rect 7570 4727 7600 4813
rect 7670 4727 7700 4813
rect 7770 4727 7800 4813
rect 7870 4727 7900 4813
rect 7970 4727 8000 4813
rect 8070 4727 8100 4813
rect 8170 4727 8200 4813
rect 8270 4727 8300 4813
rect 8370 4727 8400 4813
rect 8470 4727 8500 4813
rect 8570 4727 8600 4813
rect 8670 4727 8700 4813
rect 8770 4727 8800 4813
rect 8870 4727 8900 4813
rect 8970 4727 9000 4813
rect 9070 4727 9100 4813
rect 9170 4727 9200 4813
rect 9270 4727 9300 4813
rect 9370 4727 9400 4813
rect 9470 4727 9500 4813
rect 9570 4727 9600 4813
rect 9670 4727 9700 4813
rect 9770 4727 9800 4813
rect 6570 4587 6600 4673
rect 6670 4587 6700 4673
rect 6770 4587 6800 4673
rect 6870 4587 6900 4673
rect 6970 4587 7000 4673
rect 7070 4587 7100 4673
rect 7170 4587 7200 4673
rect 7270 4587 7300 4673
rect 7370 4587 7400 4673
rect 7470 4587 7500 4673
rect 7570 4587 7600 4673
rect 7670 4587 7700 4673
rect 7770 4587 7800 4673
rect 7870 4587 7900 4673
rect 7970 4587 8000 4673
rect 8070 4587 8100 4673
rect 8170 4587 8200 4673
rect 8270 4587 8300 4673
rect 8370 4587 8400 4673
rect 8470 4587 8500 4673
rect 8570 4587 8600 4673
rect 8670 4587 8700 4673
rect 6170 4447 6200 4533
rect 6270 4447 6300 4533
rect 6370 4447 6400 4533
rect 6470 4447 6500 4533
rect 6570 4447 6600 4533
rect 6670 4447 6700 4533
rect 6770 4447 6800 4533
rect 6870 4447 6900 4533
rect 6970 4447 7000 4533
rect 7070 4447 7100 4533
rect 7170 4447 7200 4533
rect 7270 4447 7300 4533
rect 7370 4447 7400 4533
rect 7470 4447 7500 4533
rect 7570 4447 7600 4533
rect 7670 4447 7700 4533
rect 7770 4447 7800 4533
rect 7870 4447 7900 4533
rect 7970 4447 8000 4533
rect 6170 4307 6200 4393
rect 6270 4307 6300 4393
rect 6370 4307 6400 4393
rect 6470 4307 6500 4393
rect 6570 4307 6600 4393
rect 6170 4167 6200 4253
rect 6370 4167 6400 4253
rect 6570 4167 6600 4253
rect 6770 4307 6800 4393
rect 6870 4307 6900 4393
rect 6970 4307 7000 4393
rect 7070 4307 7100 4393
rect 7170 4307 7200 4393
rect 7270 4307 7300 4393
rect 6770 4167 6800 4253
rect 6870 4167 6900 4253
rect 6970 4167 7000 4253
rect 7070 4167 7100 4253
rect 8170 4447 8200 4533
rect 8270 4447 8300 4533
rect 9970 4727 10000 4813
rect 10070 4727 10100 4813
rect 10170 4727 10200 4813
rect 10270 4727 10300 4813
rect 10370 4727 10400 4813
rect 10470 4727 10500 4813
rect 10570 4727 10600 4813
rect 10670 4727 10700 4813
rect 10870 4727 10900 4813
rect 10970 4727 11000 4813
rect 11070 4727 11100 4813
rect 11170 4727 11200 4813
rect 11270 4727 11300 4813
rect 11370 4727 11400 4813
rect 11470 4727 11500 4813
rect 11570 4727 11600 4813
rect 11770 4727 11800 4813
rect 11870 4727 11900 4813
rect 11970 4727 12000 4813
rect 12070 4727 12100 4813
rect 12170 4727 12200 4813
rect 12270 4727 12300 4813
rect 12370 4727 12400 4813
rect 12570 4727 12600 4813
rect 12670 4727 12700 4813
rect 12770 4727 12800 4813
rect 12970 4727 13000 4813
rect 13070 4727 13100 4813
rect 13280 4727 13310 4813
rect 13380 4727 13410 4813
rect 13480 4727 13510 4813
rect 13580 4727 13610 4813
rect 8870 4587 8900 4673
rect 8970 4587 9000 4673
rect 9070 4587 9100 4673
rect 9170 4587 9200 4673
rect 9270 4587 9300 4673
rect 9370 4587 9400 4673
rect 9470 4587 9500 4673
rect 9570 4587 9600 4673
rect 9670 4587 9700 4673
rect 9770 4587 9800 4673
rect 9870 4587 9900 4673
rect 9970 4587 10000 4673
rect 10070 4587 10100 4673
rect 10170 4587 10200 4673
rect 10270 4587 10300 4673
rect 10370 4587 10400 4673
rect 10470 4587 10500 4673
rect 10570 4587 10600 4673
rect 10670 4587 10700 4673
rect 10770 4587 10800 4673
rect 10870 4587 10900 4673
rect 10970 4587 11000 4673
rect 11070 4587 11100 4673
rect 11170 4587 11200 4673
rect 11270 4587 11300 4673
rect 11370 4587 11400 4673
rect 11470 4587 11500 4673
rect 11570 4587 11600 4673
rect 11670 4587 11700 4673
rect 11770 4587 11800 4673
rect 11870 4587 11900 4673
rect 11970 4587 12000 4673
rect 12070 4587 12100 4673
rect 12170 4587 12200 4673
rect 12270 4587 12300 4673
rect 12370 4587 12400 4673
rect 12470 4587 12500 4673
rect 12570 4587 12600 4673
rect 8470 4447 8500 4533
rect 8570 4447 8600 4533
rect 8670 4447 8700 4533
rect 8770 4447 8800 4533
rect 8970 4447 9000 4533
rect 9170 4447 9200 4533
rect 9270 4447 9300 4533
rect 9470 4447 9500 4533
rect 9570 4447 9600 4533
rect 9770 4447 9800 4533
rect 9870 4447 9900 4533
rect 10070 4447 10100 4533
rect 10170 4447 10200 4533
rect 10370 4447 10400 4533
rect 10470 4447 10500 4533
rect 10670 4447 10700 4533
rect 10870 4447 10900 4533
rect 7470 4307 7500 4393
rect 7570 4307 7600 4393
rect 7670 4307 7700 4393
rect 7770 4307 7800 4393
rect 7870 4307 7900 4393
rect 7970 4307 8000 4393
rect 8070 4307 8100 4393
rect 8170 4307 8200 4393
rect 8270 4307 8300 4393
rect 8370 4307 8400 4393
rect 8470 4307 8500 4393
rect 8570 4307 8600 4393
rect 8670 4307 8700 4393
rect 8770 4307 8800 4393
rect 8870 4307 8900 4393
rect 8970 4307 9000 4393
rect 9070 4307 9100 4393
rect 9170 4307 9200 4393
rect 9270 4307 9300 4393
rect 9370 4307 9400 4393
rect 9470 4307 9500 4393
rect 9570 4307 9600 4393
rect 9670 4307 9700 4393
rect 9770 4307 9800 4393
rect 9870 4307 9900 4393
rect 9970 4307 10000 4393
rect 10070 4307 10100 4393
rect 10170 4307 10200 4393
rect 10270 4307 10300 4393
rect 10370 4307 10400 4393
rect 10470 4307 10500 4393
rect 10570 4307 10600 4393
rect 10670 4307 10700 4393
rect 10770 4307 10800 4393
rect 7270 4167 7300 4253
rect 7370 4167 7400 4253
rect 7470 4167 7500 4253
rect 7570 4167 7600 4253
rect 7670 4167 7700 4253
rect 7770 4167 7800 4253
rect 7870 4167 7900 4253
rect 7970 4167 8000 4253
rect 8070 4167 8100 4253
rect 5770 4027 5800 4113
rect 5870 4027 5900 4113
rect 5970 4027 6000 4113
rect 6070 4027 6100 4113
rect 6170 4027 6200 4113
rect 6270 4027 6300 4113
rect 6370 4027 6400 4113
rect 6470 4027 6500 4113
rect 6570 4027 6600 4113
rect 6670 4027 6700 4113
rect 6770 4027 6800 4113
rect 6870 4027 6900 4113
rect 6970 4027 7000 4113
rect 7070 4027 7100 4113
rect 7170 4027 7200 4113
rect 7270 4027 7300 4113
rect 5670 3887 5700 3973
rect 5770 3887 5800 3973
rect 5870 3887 5900 3973
rect 5570 3747 5600 3833
rect 5670 3747 5700 3833
rect 5770 3747 5800 3833
rect 5870 3747 5900 3833
rect 4570 3517 4600 3603
rect 4670 3517 4700 3603
rect 4770 3517 4800 3603
rect 4870 3517 4900 3603
rect 4970 3517 5000 3603
rect 5070 3517 5100 3603
rect 5170 3517 5200 3603
rect 5270 3517 5300 3603
rect 5370 3517 5400 3603
rect 5470 3517 5500 3603
rect 5570 3517 5600 3603
rect 5670 3517 5700 3603
rect 4570 3377 4600 3463
rect 4670 3377 4700 3463
rect 4770 3377 4800 3463
rect 4970 3377 5000 3463
rect 6070 3887 6100 3973
rect 6170 3887 6200 3973
rect 6270 3887 6300 3973
rect 6370 3887 6400 3973
rect 6470 3887 6500 3973
rect 6570 3887 6600 3973
rect 6670 3887 6700 3973
rect 6770 3887 6800 3973
rect 6870 3887 6900 3973
rect 7070 3887 7100 3973
rect 7470 4027 7500 4113
rect 7570 4027 7600 4113
rect 7770 4027 7800 4113
rect 8270 4167 8300 4253
rect 8470 4167 8500 4253
rect 8670 4167 8700 4253
rect 7970 4027 8000 4113
rect 8070 4027 8100 4113
rect 8170 4027 8200 4113
rect 8270 4027 8300 4113
rect 8370 4027 8400 4113
rect 8470 4027 8500 4113
rect 8570 4027 8600 4113
rect 8670 4027 8700 4113
rect 7270 3887 7300 3973
rect 7370 3887 7400 3973
rect 7470 3887 7500 3973
rect 7570 3887 7600 3973
rect 7670 3887 7700 3973
rect 7770 3887 7800 3973
rect 7870 3887 7900 3973
rect 7970 3887 8000 3973
rect 8070 3887 8100 3973
rect 8170 3887 8200 3973
rect 8270 3887 8300 3973
rect 8370 3887 8400 3973
rect 8470 3887 8500 3973
rect 8570 3887 8600 3973
rect 8670 3887 8700 3973
rect 6070 3747 6100 3833
rect 6170 3747 6200 3833
rect 6270 3747 6300 3833
rect 6370 3747 6400 3833
rect 6470 3747 6500 3833
rect 6570 3747 6600 3833
rect 6670 3747 6700 3833
rect 6770 3747 6800 3833
rect 6870 3747 6900 3833
rect 6970 3747 7000 3833
rect 7070 3747 7100 3833
rect 7170 3747 7200 3833
rect 7270 3747 7300 3833
rect 7370 3747 7400 3833
rect 7470 3747 7500 3833
rect 7570 3747 7600 3833
rect 8870 4167 8900 4253
rect 8870 4027 8900 4113
rect 9070 4167 9100 4253
rect 9170 4167 9200 4253
rect 9270 4167 9300 4253
rect 9470 4167 9500 4253
rect 9070 4027 9100 4113
rect 9170 4027 9200 4113
rect 9270 4027 9300 4113
rect 9370 4027 9400 4113
rect 9470 4027 9500 4113
rect 8870 3887 8900 3973
rect 8970 3887 9000 3973
rect 9070 3887 9100 3973
rect 9170 3887 9200 3973
rect 9270 3887 9300 3973
rect 9370 3887 9400 3973
rect 9470 3887 9500 3973
rect 7770 3747 7800 3833
rect 7870 3747 7900 3833
rect 7970 3747 8000 3833
rect 8070 3747 8100 3833
rect 8170 3747 8200 3833
rect 8270 3747 8300 3833
rect 8370 3747 8400 3833
rect 8470 3747 8500 3833
rect 8570 3747 8600 3833
rect 8670 3747 8700 3833
rect 8770 3747 8800 3833
rect 8870 3747 8900 3833
rect 8970 3747 9000 3833
rect 9070 3747 9100 3833
rect 9170 3747 9200 3833
rect 9270 3747 9300 3833
rect 9370 3747 9400 3833
rect 5870 3517 5900 3603
rect 5970 3517 6000 3603
rect 6070 3517 6100 3603
rect 6170 3517 6200 3603
rect 6270 3517 6300 3603
rect 6370 3517 6400 3603
rect 6470 3517 6500 3603
rect 6570 3517 6600 3603
rect 6670 3517 6700 3603
rect 6770 3517 6800 3603
rect 6870 3517 6900 3603
rect 6970 3517 7000 3603
rect 7070 3517 7100 3603
rect 7170 3517 7200 3603
rect 7270 3517 7300 3603
rect 7370 3517 7400 3603
rect 7470 3517 7500 3603
rect 7570 3517 7600 3603
rect 7670 3517 7700 3603
rect 7770 3517 7800 3603
rect 7870 3517 7900 3603
rect 7970 3517 8000 3603
rect 8070 3517 8100 3603
rect 8170 3517 8200 3603
rect 8270 3517 8300 3603
rect 8370 3517 8400 3603
rect 8470 3517 8500 3603
rect 8570 3517 8600 3603
rect 8670 3517 8700 3603
rect 8770 3517 8800 3603
rect 8870 3517 8900 3603
rect 5170 3377 5200 3463
rect 5270 3377 5300 3463
rect 5370 3377 5400 3463
rect 5470 3377 5500 3463
rect 5570 3377 5600 3463
rect 5670 3377 5700 3463
rect 5770 3377 5800 3463
rect 5870 3377 5900 3463
rect 5970 3377 6000 3463
rect 6170 3377 6200 3463
rect 6270 3377 6300 3463
rect 6370 3377 6400 3463
rect 6570 3377 6600 3463
rect 6670 3377 6700 3463
rect 9070 3517 9100 3603
rect 9270 3517 9300 3603
rect 9670 4167 9700 4253
rect 9870 4167 9900 4253
rect 9970 4167 10000 4253
rect 11070 4447 11100 4533
rect 11170 4447 11200 4533
rect 10970 4307 11000 4393
rect 11070 4307 11100 4393
rect 10170 4167 10200 4253
rect 10270 4167 10300 4253
rect 10370 4167 10400 4253
rect 10470 4167 10500 4253
rect 10570 4167 10600 4253
rect 10670 4167 10700 4253
rect 10770 4167 10800 4253
rect 10870 4167 10900 4253
rect 9670 4027 9700 4113
rect 9770 4027 9800 4113
rect 9870 4027 9900 4113
rect 9970 4027 10000 4113
rect 10070 4027 10100 4113
rect 10170 4027 10200 4113
rect 10270 4027 10300 4113
rect 10370 4027 10400 4113
rect 10470 4027 10500 4113
rect 10570 4027 10600 4113
rect 10770 4027 10800 4113
rect 11370 4447 11400 4533
rect 11470 4447 11500 4533
rect 11570 4447 11600 4533
rect 11670 4447 11700 4533
rect 11770 4447 11800 4533
rect 11870 4447 11900 4533
rect 11970 4447 12000 4533
rect 12070 4447 12100 4533
rect 12170 4447 12200 4533
rect 12270 4447 12300 4533
rect 12370 4447 12400 4533
rect 11270 4307 11300 4393
rect 11370 4307 11400 4393
rect 11470 4307 11500 4393
rect 11570 4307 11600 4393
rect 11670 4307 11700 4393
rect 11770 4307 11800 4393
rect 11870 4307 11900 4393
rect 11070 4167 11100 4253
rect 11170 4167 11200 4253
rect 11270 4167 11300 4253
rect 10970 4027 11000 4113
rect 11070 4027 11100 4113
rect 11170 4027 11200 4113
rect 11270 4027 11300 4113
rect 9670 3887 9700 3973
rect 9770 3887 9800 3973
rect 9870 3887 9900 3973
rect 9970 3887 10000 3973
rect 10070 3887 10100 3973
rect 10170 3887 10200 3973
rect 10270 3887 10300 3973
rect 10370 3887 10400 3973
rect 10470 3887 10500 3973
rect 10570 3887 10600 3973
rect 10670 3887 10700 3973
rect 10770 3887 10800 3973
rect 10870 3887 10900 3973
rect 10970 3887 11000 3973
rect 9570 3747 9600 3833
rect 9670 3747 9700 3833
rect 9770 3747 9800 3833
rect 9870 3747 9900 3833
rect 9970 3747 10000 3833
rect 11470 4167 11500 4253
rect 11470 4027 11500 4113
rect 12770 4587 12800 4673
rect 12970 4587 13000 4673
rect 13070 4587 13100 4673
rect 13280 4587 13310 4673
rect 13380 4587 13410 4673
rect 13480 4587 13510 4673
rect 13580 4587 13610 4673
rect 12570 4447 12600 4533
rect 12670 4447 12700 4533
rect 12770 4447 12800 4533
rect 12970 4447 13000 4533
rect 13070 4447 13100 4533
rect 13280 4447 13310 4533
rect 13380 4447 13410 4533
rect 13480 4447 13510 4533
rect 13580 4447 13610 4533
rect 12070 4307 12100 4393
rect 12170 4307 12200 4393
rect 12270 4307 12300 4393
rect 12370 4307 12400 4393
rect 12470 4307 12500 4393
rect 12570 4307 12600 4393
rect 12670 4307 12700 4393
rect 12770 4307 12800 4393
rect 12970 4307 13000 4393
rect 13070 4307 13100 4393
rect 13280 4307 13310 4393
rect 13380 4307 13410 4393
rect 13480 4307 13510 4393
rect 13580 4307 13610 4393
rect 11670 4167 11700 4253
rect 11770 4167 11800 4253
rect 11870 4167 11900 4253
rect 11970 4167 12000 4253
rect 12070 4167 12100 4253
rect 12170 4167 12200 4253
rect 12270 4167 12300 4253
rect 12370 4167 12400 4253
rect 12470 4167 12500 4253
rect 12570 4167 12600 4253
rect 12670 4167 12700 4253
rect 12770 4167 12800 4253
rect 12970 4167 13000 4253
rect 13070 4167 13100 4253
rect 13280 4167 13310 4253
rect 13380 4167 13410 4253
rect 13480 4167 13510 4253
rect 13580 4167 13610 4253
rect 11670 4027 11700 4113
rect 11770 4027 11800 4113
rect 11970 4027 12000 4113
rect 12070 4027 12100 4113
rect 12170 4027 12200 4113
rect 12270 4027 12300 4113
rect 12370 4027 12400 4113
rect 12470 4027 12500 4113
rect 12570 4027 12600 4113
rect 12770 4027 12800 4113
rect 12970 4027 13000 4113
rect 13070 4027 13100 4113
rect 13280 4027 13310 4113
rect 13380 4027 13410 4113
rect 13480 4027 13510 4113
rect 13580 4027 13610 4113
rect 11170 3887 11200 3973
rect 11270 3887 11300 3973
rect 11370 3887 11400 3973
rect 11470 3887 11500 3973
rect 11570 3887 11600 3973
rect 11670 3887 11700 3973
rect 11770 3887 11800 3973
rect 11870 3887 11900 3973
rect 11970 3887 12000 3973
rect 12070 3887 12100 3973
rect 12170 3887 12200 3973
rect 12270 3887 12300 3973
rect 12370 3887 12400 3973
rect 12470 3887 12500 3973
rect 12570 3887 12600 3973
rect 12670 3887 12700 3973
rect 12770 3887 12800 3973
rect 12970 3887 13000 3973
rect 13070 3887 13100 3973
rect 13280 3887 13310 3973
rect 13380 3887 13410 3973
rect 13480 3887 13510 3973
rect 13580 3887 13610 3973
rect 10170 3747 10200 3833
rect 10270 3747 10300 3833
rect 10370 3747 10400 3833
rect 10470 3747 10500 3833
rect 10570 3747 10600 3833
rect 10670 3747 10700 3833
rect 10770 3747 10800 3833
rect 10870 3747 10900 3833
rect 10970 3747 11000 3833
rect 11070 3747 11100 3833
rect 9470 3517 9500 3603
rect 9570 3517 9600 3603
rect 9670 3517 9700 3603
rect 9770 3517 9800 3603
rect 9870 3517 9900 3603
rect 9970 3517 10000 3603
rect 6870 3377 6900 3463
rect 6970 3377 7000 3463
rect 7070 3377 7100 3463
rect 7170 3377 7200 3463
rect 7270 3377 7300 3463
rect 7370 3377 7400 3463
rect 7470 3377 7500 3463
rect 7570 3377 7600 3463
rect 7670 3377 7700 3463
rect 7770 3377 7800 3463
rect 7870 3377 7900 3463
rect 7970 3377 8000 3463
rect 8070 3377 8100 3463
rect 8170 3377 8200 3463
rect 8270 3377 8300 3463
rect 8370 3377 8400 3463
rect 8470 3377 8500 3463
rect 8570 3377 8600 3463
rect 8670 3377 8700 3463
rect 8770 3377 8800 3463
rect 8870 3377 8900 3463
rect 8970 3377 9000 3463
rect 9070 3377 9100 3463
rect 9170 3377 9200 3463
rect 9270 3377 9300 3463
rect 9370 3377 9400 3463
rect 3570 3237 3600 3323
rect 3670 3237 3700 3323
rect 3770 3237 3800 3323
rect 3870 3237 3900 3323
rect 3970 3237 4000 3323
rect 4070 3237 4100 3323
rect 4170 3237 4200 3323
rect 4270 3237 4300 3323
rect 4370 3237 4400 3323
rect 4470 3237 4500 3323
rect 4570 3237 4600 3323
rect 4670 3237 4700 3323
rect 4770 3237 4800 3323
rect 4870 3237 4900 3323
rect 4970 3237 5000 3323
rect 5070 3237 5100 3323
rect 5170 3237 5200 3323
rect 5270 3237 5300 3323
rect 5370 3237 5400 3323
rect 5470 3237 5500 3323
rect 5570 3237 5600 3323
rect 5670 3237 5700 3323
rect 5770 3237 5800 3323
rect 5870 3237 5900 3323
rect 5970 3237 6000 3323
rect 6070 3237 6100 3323
rect 6170 3237 6200 3323
rect 6270 3237 6300 3323
rect 6370 3237 6400 3323
rect 6470 3237 6500 3323
rect 6570 3237 6600 3323
rect 6670 3237 6700 3323
rect 6770 3237 6800 3323
rect 6870 3237 6900 3323
rect 6970 3237 7000 3323
rect 7070 3237 7100 3323
rect 7170 3237 7200 3323
rect 7270 3237 7300 3323
rect 3370 3097 3400 3183
rect 3470 3097 3500 3183
rect 3570 3097 3600 3183
rect 3770 3097 3800 3183
rect 3870 3097 3900 3183
rect 3970 3097 4000 3183
rect 4070 3097 4100 3183
rect 4170 3097 4200 3183
rect 4270 3097 4300 3183
rect 4370 3097 4400 3183
rect 4470 3097 4500 3183
rect 4570 3097 4600 3183
rect 4670 3097 4700 3183
rect 4770 3097 4800 3183
rect 4870 3097 4900 3183
rect 4970 3097 5000 3183
rect 5070 3097 5100 3183
rect 5170 3097 5200 3183
rect 5270 3097 5300 3183
rect 5370 3097 5400 3183
rect 3170 2957 3200 3043
rect 3270 2957 3300 3043
rect 3370 2957 3400 3043
rect 3470 2957 3500 3043
rect 3570 2957 3600 3043
rect 3670 2957 3700 3043
rect 3770 2957 3800 3043
rect 3070 2817 3100 2903
rect 3170 2817 3200 2903
rect 3270 2817 3300 2903
rect 3970 2957 4000 3043
rect 4070 2957 4100 3043
rect 4170 2957 4200 3043
rect 4270 2957 4300 3043
rect 4370 2957 4400 3043
rect 4470 2957 4500 3043
rect 3470 2817 3500 2903
rect 3570 2817 3600 2903
rect 3670 2817 3700 2903
rect 3770 2817 3800 2903
rect 3870 2817 3900 2903
rect 4670 2957 4700 3043
rect 4770 2957 4800 3043
rect 4870 2957 4900 3043
rect 5570 3097 5600 3183
rect 5770 3097 5800 3183
rect 5970 3097 6000 3183
rect 6070 3097 6100 3183
rect 6170 3097 6200 3183
rect 6270 3097 6300 3183
rect 5070 2957 5100 3043
rect 5170 2957 5200 3043
rect 5270 2957 5300 3043
rect 5370 2957 5400 3043
rect 5470 2957 5500 3043
rect 5570 2957 5600 3043
rect 5670 2957 5700 3043
rect 5770 2957 5800 3043
rect 5870 2957 5900 3043
rect 4070 2817 4100 2903
rect 4170 2817 4200 2903
rect 4270 2817 4300 2903
rect 4370 2817 4400 2903
rect 4470 2817 4500 2903
rect 4570 2817 4600 2903
rect 4670 2817 4700 2903
rect 4770 2817 4800 2903
rect 4870 2817 4900 2903
rect 4970 2817 5000 2903
rect 5070 2817 5100 2903
rect 5170 2817 5200 2903
rect 5270 2817 5300 2903
rect 2470 2677 2500 2763
rect 2570 2677 2600 2763
rect 2670 2677 2700 2763
rect 2770 2677 2800 2763
rect 2870 2677 2900 2763
rect 2970 2677 3000 2763
rect 3070 2677 3100 2763
rect 3170 2677 3200 2763
rect 3270 2677 3300 2763
rect 3370 2677 3400 2763
rect 3470 2677 3500 2763
rect 3570 2677 3600 2763
rect 3670 2677 3700 2763
rect 3770 2677 3800 2763
rect 3870 2677 3900 2763
rect 3970 2677 4000 2763
rect 4070 2677 4100 2763
rect 70 2537 100 2623
rect 170 2537 200 2623
rect 270 2537 300 2623
rect 370 2537 400 2623
rect 470 2537 500 2623
rect 570 2537 600 2623
rect 670 2537 700 2623
rect 770 2537 800 2623
rect 870 2537 900 2623
rect 970 2537 1000 2623
rect 1070 2537 1100 2623
rect 1170 2537 1200 2623
rect 1270 2537 1300 2623
rect 1370 2537 1400 2623
rect 1470 2537 1500 2623
rect 1570 2537 1600 2623
rect 1670 2537 1700 2623
rect 1770 2537 1800 2623
rect 1870 2537 1900 2623
rect 1970 2537 2000 2623
rect 2070 2537 2100 2623
rect 2170 2537 2200 2623
rect 2270 2537 2300 2623
rect 2370 2537 2400 2623
rect 2470 2537 2500 2623
rect 70 2307 100 2393
rect 270 2307 300 2393
rect 370 2307 400 2393
rect 570 2307 600 2393
rect 770 2307 800 2393
rect 870 2307 900 2393
rect 970 2307 1000 2393
rect 1070 2307 1100 2393
rect 1170 2307 1200 2393
rect 1270 2307 1300 2393
rect 1370 2307 1400 2393
rect 1470 2307 1500 2393
rect 1570 2307 1600 2393
rect 1670 2307 1700 2393
rect 1770 2307 1800 2393
rect 1870 2307 1900 2393
rect 1970 2307 2000 2393
rect 2070 2307 2100 2393
rect 2170 2307 2200 2393
rect 2270 2307 2300 2393
rect 70 2167 100 2253
rect 170 2167 200 2253
rect 270 2167 300 2253
rect 370 2167 400 2253
rect 470 2167 500 2253
rect 570 2167 600 2253
rect 670 2167 700 2253
rect 770 2167 800 2253
rect 70 2027 100 2113
rect 170 2027 200 2113
rect 270 2027 300 2113
rect 370 2027 400 2113
rect 470 2027 500 2113
rect 570 2027 600 2113
rect 670 2027 700 2113
rect 970 2167 1000 2253
rect 2670 2537 2700 2623
rect 2770 2537 2800 2623
rect 2870 2537 2900 2623
rect 2970 2537 3000 2623
rect 3070 2537 3100 2623
rect 3170 2537 3200 2623
rect 3270 2537 3300 2623
rect 2470 2307 2500 2393
rect 2570 2307 2600 2393
rect 1170 2167 1200 2253
rect 1270 2167 1300 2253
rect 1370 2167 1400 2253
rect 1470 2167 1500 2253
rect 1570 2167 1600 2253
rect 1670 2167 1700 2253
rect 1770 2167 1800 2253
rect 1870 2167 1900 2253
rect 1970 2167 2000 2253
rect 2070 2167 2100 2253
rect 2170 2167 2200 2253
rect 2270 2167 2300 2253
rect 2370 2167 2400 2253
rect 2470 2167 2500 2253
rect 2570 2167 2600 2253
rect 870 2027 900 2113
rect 970 2027 1000 2113
rect 1070 2027 1100 2113
rect 1170 2027 1200 2113
rect 1270 2027 1300 2113
rect 1370 2027 1400 2113
rect 70 1887 100 1973
rect 170 1887 200 1973
rect 270 1887 300 1973
rect 370 1887 400 1973
rect 470 1887 500 1973
rect 570 1887 600 1973
rect 670 1887 700 1973
rect 770 1887 800 1973
rect 870 1887 900 1973
rect 3470 2537 3500 2623
rect 3570 2537 3600 2623
rect 3670 2537 3700 2623
rect 3770 2537 3800 2623
rect 3870 2537 3900 2623
rect 4070 2537 4100 2623
rect 4270 2677 4300 2763
rect 4370 2677 4400 2763
rect 4470 2677 4500 2763
rect 4570 2677 4600 2763
rect 4670 2677 4700 2763
rect 4270 2537 4300 2623
rect 4470 2537 4500 2623
rect 4570 2537 4600 2623
rect 4670 2537 4700 2623
rect 4870 2677 4900 2763
rect 4970 2677 5000 2763
rect 5070 2677 5100 2763
rect 5270 2677 5300 2763
rect 6470 3097 6500 3183
rect 6670 3097 6700 3183
rect 6770 3097 6800 3183
rect 6870 3097 6900 3183
rect 6970 3097 7000 3183
rect 9570 3377 9600 3463
rect 9670 3377 9700 3463
rect 7470 3237 7500 3323
rect 7570 3237 7600 3323
rect 7670 3237 7700 3323
rect 7770 3237 7800 3323
rect 7870 3237 7900 3323
rect 7970 3237 8000 3323
rect 8070 3237 8100 3323
rect 8170 3237 8200 3323
rect 8270 3237 8300 3323
rect 8370 3237 8400 3323
rect 8470 3237 8500 3323
rect 8570 3237 8600 3323
rect 8670 3237 8700 3323
rect 8770 3237 8800 3323
rect 8870 3237 8900 3323
rect 8970 3237 9000 3323
rect 9070 3237 9100 3323
rect 9170 3237 9200 3323
rect 9270 3237 9300 3323
rect 9370 3237 9400 3323
rect 9470 3237 9500 3323
rect 7170 3097 7200 3183
rect 7270 3097 7300 3183
rect 7370 3097 7400 3183
rect 7470 3097 7500 3183
rect 7570 3097 7600 3183
rect 7670 3097 7700 3183
rect 7770 3097 7800 3183
rect 7870 3097 7900 3183
rect 7970 3097 8000 3183
rect 8070 3097 8100 3183
rect 6070 2957 6100 3043
rect 6170 2957 6200 3043
rect 6270 2957 6300 3043
rect 6370 2957 6400 3043
rect 6470 2957 6500 3043
rect 6570 2957 6600 3043
rect 6670 2957 6700 3043
rect 6770 2957 6800 3043
rect 6870 2957 6900 3043
rect 6970 2957 7000 3043
rect 7070 2957 7100 3043
rect 7170 2957 7200 3043
rect 7270 2957 7300 3043
rect 7370 2957 7400 3043
rect 7470 2957 7500 3043
rect 7570 2957 7600 3043
rect 7670 2957 7700 3043
rect 7770 2957 7800 3043
rect 7870 2957 7900 3043
rect 7970 2957 8000 3043
rect 5470 2817 5500 2903
rect 5570 2817 5600 2903
rect 5670 2817 5700 2903
rect 5770 2817 5800 2903
rect 5870 2817 5900 2903
rect 5970 2817 6000 2903
rect 5470 2677 5500 2763
rect 5570 2677 5600 2763
rect 5670 2677 5700 2763
rect 5770 2677 5800 2763
rect 5870 2677 5900 2763
rect 5970 2677 6000 2763
rect 6170 2817 6200 2903
rect 6270 2817 6300 2903
rect 6370 2817 6400 2903
rect 6470 2817 6500 2903
rect 6570 2817 6600 2903
rect 6670 2817 6700 2903
rect 6770 2817 6800 2903
rect 6870 2817 6900 2903
rect 6170 2677 6200 2763
rect 4870 2537 4900 2623
rect 4970 2537 5000 2623
rect 5070 2537 5100 2623
rect 5170 2537 5200 2623
rect 5270 2537 5300 2623
rect 5370 2537 5400 2623
rect 5470 2537 5500 2623
rect 5570 2537 5600 2623
rect 5670 2537 5700 2623
rect 5770 2537 5800 2623
rect 5870 2537 5900 2623
rect 5970 2537 6000 2623
rect 6070 2537 6100 2623
rect 6170 2537 6200 2623
rect 6370 2677 6400 2763
rect 6470 2677 6500 2763
rect 7070 2817 7100 2903
rect 7170 2817 7200 2903
rect 7270 2817 7300 2903
rect 7470 2817 7500 2903
rect 7570 2817 7600 2903
rect 7670 2817 7700 2903
rect 7770 2817 7800 2903
rect 7870 2817 7900 2903
rect 8270 3097 8300 3183
rect 8370 3097 8400 3183
rect 8470 3097 8500 3183
rect 8570 3097 8600 3183
rect 8670 3097 8700 3183
rect 8770 3097 8800 3183
rect 8170 2957 8200 3043
rect 8270 2957 8300 3043
rect 8370 2957 8400 3043
rect 8470 2957 8500 3043
rect 8570 2957 8600 3043
rect 8670 2957 8700 3043
rect 8770 2957 8800 3043
rect 8070 2817 8100 2903
rect 8170 2817 8200 2903
rect 8270 2817 8300 2903
rect 8370 2817 8400 2903
rect 8470 2817 8500 2903
rect 8570 2817 8600 2903
rect 8670 2817 8700 2903
rect 6670 2677 6700 2763
rect 6770 2677 6800 2763
rect 6870 2677 6900 2763
rect 6970 2677 7000 2763
rect 7070 2677 7100 2763
rect 7170 2677 7200 2763
rect 7270 2677 7300 2763
rect 7370 2677 7400 2763
rect 7470 2677 7500 2763
rect 7570 2677 7600 2763
rect 7670 2677 7700 2763
rect 7770 2677 7800 2763
rect 7870 2677 7900 2763
rect 7970 2677 8000 2763
rect 8070 2677 8100 2763
rect 8170 2677 8200 2763
rect 6370 2537 6400 2623
rect 6470 2537 6500 2623
rect 6570 2537 6600 2623
rect 6670 2537 6700 2623
rect 6870 2537 6900 2623
rect 6970 2537 7000 2623
rect 7070 2537 7100 2623
rect 7170 2537 7200 2623
rect 7270 2537 7300 2623
rect 7370 2537 7400 2623
rect 7470 2537 7500 2623
rect 7570 2537 7600 2623
rect 7670 2537 7700 2623
rect 7770 2537 7800 2623
rect 7870 2537 7900 2623
rect 7970 2537 8000 2623
rect 8070 2537 8100 2623
rect 8170 2537 8200 2623
rect 2770 2307 2800 2393
rect 2870 2307 2900 2393
rect 2970 2307 3000 2393
rect 3070 2307 3100 2393
rect 3170 2307 3200 2393
rect 3270 2307 3300 2393
rect 3370 2307 3400 2393
rect 3470 2307 3500 2393
rect 3570 2307 3600 2393
rect 3670 2307 3700 2393
rect 3770 2307 3800 2393
rect 3870 2307 3900 2393
rect 3970 2307 4000 2393
rect 4070 2307 4100 2393
rect 4170 2307 4200 2393
rect 4270 2307 4300 2393
rect 4370 2307 4400 2393
rect 4470 2307 4500 2393
rect 4570 2307 4600 2393
rect 4670 2307 4700 2393
rect 4770 2307 4800 2393
rect 4870 2307 4900 2393
rect 4970 2307 5000 2393
rect 5070 2307 5100 2393
rect 5170 2307 5200 2393
rect 5270 2307 5300 2393
rect 5370 2307 5400 2393
rect 5470 2307 5500 2393
rect 5570 2307 5600 2393
rect 5670 2307 5700 2393
rect 5770 2307 5800 2393
rect 5870 2307 5900 2393
rect 5970 2307 6000 2393
rect 6070 2307 6100 2393
rect 6170 2307 6200 2393
rect 6270 2307 6300 2393
rect 6370 2307 6400 2393
rect 6470 2307 6500 2393
rect 6570 2307 6600 2393
rect 6670 2307 6700 2393
rect 6770 2307 6800 2393
rect 6870 2307 6900 2393
rect 2770 2167 2800 2253
rect 1570 2027 1600 2113
rect 1670 2027 1700 2113
rect 1770 2027 1800 2113
rect 1870 2027 1900 2113
rect 1970 2027 2000 2113
rect 2070 2027 2100 2113
rect 2170 2027 2200 2113
rect 2270 2027 2300 2113
rect 2370 2027 2400 2113
rect 2470 2027 2500 2113
rect 2570 2027 2600 2113
rect 2670 2027 2700 2113
rect 1070 1887 1100 1973
rect 1170 1887 1200 1973
rect 1270 1887 1300 1973
rect 1370 1887 1400 1973
rect 1470 1887 1500 1973
rect 2970 2167 3000 2253
rect 2870 2027 2900 2113
rect 3170 2167 3200 2253
rect 3270 2167 3300 2253
rect 3470 2167 3500 2253
rect 3570 2167 3600 2253
rect 3070 2027 3100 2113
rect 3170 2027 3200 2113
rect 3270 2027 3300 2113
rect 3370 2027 3400 2113
rect 3470 2027 3500 2113
rect 3770 2167 3800 2253
rect 3970 2167 4000 2253
rect 4070 2167 4100 2253
rect 4170 2167 4200 2253
rect 4270 2167 4300 2253
rect 4470 2167 4500 2253
rect 4570 2167 4600 2253
rect 4670 2167 4700 2253
rect 4770 2167 4800 2253
rect 4870 2167 4900 2253
rect 4970 2167 5000 2253
rect 5070 2167 5100 2253
rect 5170 2167 5200 2253
rect 5270 2167 5300 2253
rect 5370 2167 5400 2253
rect 5470 2167 5500 2253
rect 5570 2167 5600 2253
rect 5670 2167 5700 2253
rect 5770 2167 5800 2253
rect 5870 2167 5900 2253
rect 5970 2167 6000 2253
rect 6070 2167 6100 2253
rect 3670 2027 3700 2113
rect 3770 2027 3800 2113
rect 3870 2027 3900 2113
rect 3970 2027 4000 2113
rect 4070 2027 4100 2113
rect 4170 2027 4200 2113
rect 4270 2027 4300 2113
rect 4370 2027 4400 2113
rect 4470 2027 4500 2113
rect 4570 2027 4600 2113
rect 1670 1887 1700 1973
rect 1770 1887 1800 1973
rect 1870 1887 1900 1973
rect 1970 1887 2000 1973
rect 2070 1887 2100 1973
rect 2170 1887 2200 1973
rect 2270 1887 2300 1973
rect 2370 1887 2400 1973
rect 2470 1887 2500 1973
rect 2570 1887 2600 1973
rect 2670 1887 2700 1973
rect 2770 1887 2800 1973
rect 2870 1887 2900 1973
rect 2970 1887 3000 1973
rect 3070 1887 3100 1973
rect 3170 1887 3200 1973
rect 3270 1887 3300 1973
rect 3370 1887 3400 1973
rect 3470 1887 3500 1973
rect 3570 1887 3600 1973
rect 70 1747 100 1833
rect 170 1747 200 1833
rect 270 1747 300 1833
rect 370 1747 400 1833
rect 470 1747 500 1833
rect 570 1747 600 1833
rect 670 1747 700 1833
rect 770 1747 800 1833
rect 870 1747 900 1833
rect 970 1747 1000 1833
rect 1070 1747 1100 1833
rect 1170 1747 1200 1833
rect 1270 1747 1300 1833
rect 1370 1747 1400 1833
rect 1470 1747 1500 1833
rect 1570 1747 1600 1833
rect 1670 1747 1700 1833
rect 1770 1747 1800 1833
rect 1870 1747 1900 1833
rect 1970 1747 2000 1833
rect 2070 1747 2100 1833
rect 2170 1747 2200 1833
rect 2270 1747 2300 1833
rect 2370 1747 2400 1833
rect 2470 1747 2500 1833
rect 2570 1747 2600 1833
rect 2670 1747 2700 1833
rect 2770 1747 2800 1833
rect 2870 1747 2900 1833
rect 2970 1747 3000 1833
rect 3070 1747 3100 1833
rect 70 1607 100 1693
rect 170 1607 200 1693
rect 270 1607 300 1693
rect 370 1607 400 1693
rect 470 1607 500 1693
rect 570 1607 600 1693
rect 70 1467 100 1553
rect 170 1467 200 1553
rect 270 1467 300 1553
rect 370 1467 400 1553
rect 770 1607 800 1693
rect 870 1607 900 1693
rect 970 1607 1000 1693
rect 1170 1607 1200 1693
rect 1370 1607 1400 1693
rect 1470 1607 1500 1693
rect 1670 1607 1700 1693
rect 1770 1607 1800 1693
rect 1870 1607 1900 1693
rect 1970 1607 2000 1693
rect 2070 1607 2100 1693
rect 2170 1607 2200 1693
rect 2270 1607 2300 1693
rect 2370 1607 2400 1693
rect 2470 1607 2500 1693
rect 2570 1607 2600 1693
rect 570 1467 600 1553
rect 670 1467 700 1553
rect 770 1467 800 1553
rect 870 1467 900 1553
rect 970 1467 1000 1553
rect 1070 1467 1100 1553
rect 1170 1467 1200 1553
rect 1270 1467 1300 1553
rect 1370 1467 1400 1553
rect 1470 1467 1500 1553
rect 1570 1467 1600 1553
rect 1670 1467 1700 1553
rect 1770 1467 1800 1553
rect 1870 1467 1900 1553
rect 1970 1467 2000 1553
rect 2070 1467 2100 1553
rect 2170 1467 2200 1553
rect 2270 1467 2300 1553
rect 2370 1467 2400 1553
rect 2470 1467 2500 1553
rect 70 1327 100 1413
rect 170 1327 200 1413
rect 270 1327 300 1413
rect 370 1327 400 1413
rect 470 1327 500 1413
rect 570 1327 600 1413
rect 670 1327 700 1413
rect 770 1327 800 1413
rect 3270 1747 3300 1833
rect 3770 1887 3800 1973
rect 3870 1887 3900 1973
rect 3970 1887 4000 1973
rect 4070 1887 4100 1973
rect 4170 1887 4200 1973
rect 3470 1747 3500 1833
rect 3570 1747 3600 1833
rect 3670 1747 3700 1833
rect 3770 1747 3800 1833
rect 3870 1747 3900 1833
rect 2770 1607 2800 1693
rect 2870 1607 2900 1693
rect 2970 1607 3000 1693
rect 3070 1607 3100 1693
rect 3170 1607 3200 1693
rect 3270 1607 3300 1693
rect 3370 1607 3400 1693
rect 3470 1607 3500 1693
rect 3570 1607 3600 1693
rect 3670 1607 3700 1693
rect 2670 1467 2700 1553
rect 2770 1467 2800 1553
rect 2870 1467 2900 1553
rect 2970 1467 3000 1553
rect 3070 1467 3100 1553
rect 970 1327 1000 1413
rect 1070 1327 1100 1413
rect 1170 1327 1200 1413
rect 1270 1327 1300 1413
rect 1370 1327 1400 1413
rect 1470 1327 1500 1413
rect 1570 1327 1600 1413
rect 1670 1327 1700 1413
rect 1770 1327 1800 1413
rect 1870 1327 1900 1413
rect 1970 1327 2000 1413
rect 2070 1327 2100 1413
rect 2170 1327 2200 1413
rect 2270 1327 2300 1413
rect 2370 1327 2400 1413
rect 2470 1327 2500 1413
rect 2570 1327 2600 1413
rect 2670 1327 2700 1413
rect 2770 1327 2800 1413
rect 70 1097 100 1183
rect 170 1097 200 1183
rect 270 1097 300 1183
rect 370 1097 400 1183
rect 470 1097 500 1183
rect 570 1097 600 1183
rect 670 1097 700 1183
rect 770 1097 800 1183
rect 870 1097 900 1183
rect 970 1097 1000 1183
rect 1070 1097 1100 1183
rect 1170 1097 1200 1183
rect 1270 1097 1300 1183
rect 1370 1097 1400 1183
rect 1470 1097 1500 1183
rect 1570 1097 1600 1183
rect 1670 1097 1700 1183
rect 70 957 100 1043
rect 70 817 100 903
rect 270 957 300 1043
rect 370 957 400 1043
rect 470 957 500 1043
rect 570 957 600 1043
rect 770 957 800 1043
rect 870 957 900 1043
rect 970 957 1000 1043
rect 1070 957 1100 1043
rect 1170 957 1200 1043
rect 1870 1097 1900 1183
rect 1970 1097 2000 1183
rect 3270 1467 3300 1553
rect 3370 1467 3400 1553
rect 3470 1467 3500 1553
rect 3870 1607 3900 1693
rect 4070 1747 4100 1833
rect 4070 1607 4100 1693
rect 3670 1467 3700 1553
rect 3770 1467 3800 1553
rect 3870 1467 3900 1553
rect 3970 1467 4000 1553
rect 4370 1887 4400 1973
rect 4570 1887 4600 1973
rect 4770 2027 4800 2113
rect 4870 2027 4900 2113
rect 5070 2027 5100 2113
rect 5170 2027 5200 2113
rect 5270 2027 5300 2113
rect 5370 2027 5400 2113
rect 5470 2027 5500 2113
rect 5570 2027 5600 2113
rect 5670 2027 5700 2113
rect 4770 1887 4800 1973
rect 4870 1887 4900 1973
rect 4970 1887 5000 1973
rect 5070 1887 5100 1973
rect 4270 1747 4300 1833
rect 4370 1747 4400 1833
rect 4470 1747 4500 1833
rect 4570 1747 4600 1833
rect 4670 1747 4700 1833
rect 4770 1747 4800 1833
rect 4270 1607 4300 1693
rect 4370 1607 4400 1693
rect 5270 1887 5300 1973
rect 5370 1887 5400 1973
rect 5470 1887 5500 1973
rect 5570 1887 5600 1973
rect 5670 1887 5700 1973
rect 6270 2167 6300 2253
rect 6370 2167 6400 2253
rect 6570 2167 6600 2253
rect 6670 2167 6700 2253
rect 5870 2027 5900 2113
rect 5970 2027 6000 2113
rect 6070 2027 6100 2113
rect 6170 2027 6200 2113
rect 6270 2027 6300 2113
rect 6370 2027 6400 2113
rect 6470 2027 6500 2113
rect 6570 2027 6600 2113
rect 6870 2167 6900 2253
rect 6770 2027 6800 2113
rect 5870 1887 5900 1973
rect 5970 1887 6000 1973
rect 6070 1887 6100 1973
rect 6170 1887 6200 1973
rect 6270 1887 6300 1973
rect 6370 1887 6400 1973
rect 6470 1887 6500 1973
rect 6570 1887 6600 1973
rect 6670 1887 6700 1973
rect 4970 1747 5000 1833
rect 5070 1747 5100 1833
rect 5170 1747 5200 1833
rect 5270 1747 5300 1833
rect 5370 1747 5400 1833
rect 5470 1747 5500 1833
rect 5570 1747 5600 1833
rect 5670 1747 5700 1833
rect 5770 1747 5800 1833
rect 5870 1747 5900 1833
rect 5970 1747 6000 1833
rect 6070 1747 6100 1833
rect 6170 1747 6200 1833
rect 6270 1747 6300 1833
rect 4570 1607 4600 1693
rect 4670 1607 4700 1693
rect 4770 1607 4800 1693
rect 4870 1607 4900 1693
rect 4170 1467 4200 1553
rect 4270 1467 4300 1553
rect 4370 1467 4400 1553
rect 4470 1467 4500 1553
rect 4570 1467 4600 1553
rect 4670 1467 4700 1553
rect 4770 1467 4800 1553
rect 2970 1327 3000 1413
rect 3070 1327 3100 1413
rect 3170 1327 3200 1413
rect 3270 1327 3300 1413
rect 3370 1327 3400 1413
rect 3470 1327 3500 1413
rect 3570 1327 3600 1413
rect 3670 1327 3700 1413
rect 3770 1327 3800 1413
rect 3870 1327 3900 1413
rect 3970 1327 4000 1413
rect 4070 1327 4100 1413
rect 4170 1327 4200 1413
rect 4270 1327 4300 1413
rect 4370 1327 4400 1413
rect 4470 1327 4500 1413
rect 4570 1327 4600 1413
rect 2170 1097 2200 1183
rect 2270 1097 2300 1183
rect 2370 1097 2400 1183
rect 2470 1097 2500 1183
rect 2570 1097 2600 1183
rect 2670 1097 2700 1183
rect 2770 1097 2800 1183
rect 2870 1097 2900 1183
rect 2970 1097 3000 1183
rect 1370 957 1400 1043
rect 1470 957 1500 1043
rect 1570 957 1600 1043
rect 1670 957 1700 1043
rect 1770 957 1800 1043
rect 1870 957 1900 1043
rect 1970 957 2000 1043
rect 2070 957 2100 1043
rect 2170 957 2200 1043
rect 2270 957 2300 1043
rect 2370 957 2400 1043
rect 2470 957 2500 1043
rect 2570 957 2600 1043
rect 2770 957 2800 1043
rect 3170 1097 3200 1183
rect 2970 957 3000 1043
rect 3070 957 3100 1043
rect 270 817 300 903
rect 370 817 400 903
rect 470 817 500 903
rect 570 817 600 903
rect 670 817 700 903
rect 770 817 800 903
rect 870 817 900 903
rect 970 817 1000 903
rect 1070 817 1100 903
rect 1170 817 1200 903
rect 1270 817 1300 903
rect 1370 817 1400 903
rect 1470 817 1500 903
rect 1570 817 1600 903
rect 1670 817 1700 903
rect 1770 817 1800 903
rect 1870 817 1900 903
rect 1970 817 2000 903
rect 2070 817 2100 903
rect 2170 817 2200 903
rect 2270 817 2300 903
rect 2370 817 2400 903
rect 2470 817 2500 903
rect 2570 817 2600 903
rect 2670 817 2700 903
rect 2770 817 2800 903
rect 2870 817 2900 903
rect 70 677 100 763
rect 170 677 200 763
rect 270 677 300 763
rect 370 677 400 763
rect 470 677 500 763
rect 670 677 700 763
rect 70 537 100 623
rect 170 537 200 623
rect 270 537 300 623
rect 370 537 400 623
rect 470 537 500 623
rect 570 537 600 623
rect 670 537 700 623
rect 70 397 100 483
rect 170 397 200 483
rect 270 397 300 483
rect 870 677 900 763
rect 970 677 1000 763
rect 1070 677 1100 763
rect 1170 677 1200 763
rect 870 537 900 623
rect 970 537 1000 623
rect 1070 537 1100 623
rect 1170 537 1200 623
rect 470 397 500 483
rect 570 397 600 483
rect 670 397 700 483
rect 770 397 800 483
rect 870 397 900 483
rect 970 397 1000 483
rect 1070 397 1100 483
rect 1370 677 1400 763
rect 1570 677 1600 763
rect 1670 677 1700 763
rect 1770 677 1800 763
rect 1870 677 1900 763
rect 1970 677 2000 763
rect 2170 677 2200 763
rect 2270 677 2300 763
rect 2370 677 2400 763
rect 1370 537 1400 623
rect 1470 537 1500 623
rect 1570 537 1600 623
rect 1670 537 1700 623
rect 1770 537 1800 623
rect 1870 537 1900 623
rect 1970 537 2000 623
rect 2070 537 2100 623
rect 1270 397 1300 483
rect 1370 397 1400 483
rect 1470 397 1500 483
rect 1570 397 1600 483
rect 1670 397 1700 483
rect 1770 397 1800 483
rect 70 257 100 343
rect 170 257 200 343
rect 270 257 300 343
rect 370 257 400 343
rect 470 257 500 343
rect 570 257 600 343
rect 670 257 700 343
rect 770 257 800 343
rect 870 257 900 343
rect 970 257 1000 343
rect 1070 257 1100 343
rect 1170 257 1200 343
rect 1270 257 1300 343
rect 1370 257 1400 343
rect 1470 257 1500 343
rect 1570 257 1600 343
rect 1670 257 1700 343
rect 70 117 100 203
rect 170 117 200 203
rect 270 117 300 203
rect 370 117 400 203
rect 470 117 500 203
rect 570 117 600 203
rect 670 117 700 203
rect 770 117 800 203
rect 870 117 900 203
rect 970 117 1000 203
rect 1070 117 1100 203
rect 1170 117 1200 203
rect 1270 117 1300 203
rect 1370 117 1400 203
rect 1470 117 1500 203
rect 1570 117 1600 203
rect 2570 677 2600 763
rect 2670 677 2700 763
rect 2770 677 2800 763
rect 2270 537 2300 623
rect 2370 537 2400 623
rect 2470 537 2500 623
rect 2570 537 2600 623
rect 2670 537 2700 623
rect 1970 397 2000 483
rect 2070 397 2100 483
rect 2170 397 2200 483
rect 2270 397 2300 483
rect 2470 397 2500 483
rect 2570 397 2600 483
rect 3370 1097 3400 1183
rect 3470 1097 3500 1183
rect 3570 1097 3600 1183
rect 3670 1097 3700 1183
rect 3270 957 3300 1043
rect 3470 957 3500 1043
rect 3570 957 3600 1043
rect 3870 1097 3900 1183
rect 3970 1097 4000 1183
rect 4070 1097 4100 1183
rect 4170 1097 4200 1183
rect 4270 1097 4300 1183
rect 4370 1097 4400 1183
rect 3770 957 3800 1043
rect 3070 817 3100 903
rect 3170 817 3200 903
rect 3270 817 3300 903
rect 3370 817 3400 903
rect 3470 817 3500 903
rect 3570 817 3600 903
rect 3670 817 3700 903
rect 3770 817 3800 903
rect 2970 677 3000 763
rect 3170 677 3200 763
rect 3270 677 3300 763
rect 3470 677 3500 763
rect 3570 677 3600 763
rect 4770 1327 4800 1413
rect 4570 1097 4600 1183
rect 5070 1607 5100 1693
rect 5170 1607 5200 1693
rect 5370 1607 5400 1693
rect 5470 1607 5500 1693
rect 5570 1607 5600 1693
rect 5770 1607 5800 1693
rect 5870 1607 5900 1693
rect 4970 1467 5000 1553
rect 5070 1467 5100 1553
rect 5170 1467 5200 1553
rect 5270 1467 5300 1553
rect 5370 1467 5400 1553
rect 5470 1467 5500 1553
rect 5570 1467 5600 1553
rect 5670 1467 5700 1553
rect 5770 1467 5800 1553
rect 4970 1327 5000 1413
rect 5070 1327 5100 1413
rect 6070 1607 6100 1693
rect 5970 1467 6000 1553
rect 7070 2307 7100 2393
rect 7170 2307 7200 2393
rect 8370 2677 8400 2763
rect 8470 2677 8500 2763
rect 8570 2677 8600 2763
rect 8670 2677 8700 2763
rect 8370 2537 8400 2623
rect 8570 2537 8600 2623
rect 8670 2537 8700 2623
rect 7370 2307 7400 2393
rect 7470 2307 7500 2393
rect 7570 2307 7600 2393
rect 7670 2307 7700 2393
rect 7770 2307 7800 2393
rect 7870 2307 7900 2393
rect 7970 2307 8000 2393
rect 8070 2307 8100 2393
rect 8170 2307 8200 2393
rect 8270 2307 8300 2393
rect 8370 2307 8400 2393
rect 8470 2307 8500 2393
rect 7070 2167 7100 2253
rect 7170 2167 7200 2253
rect 7270 2167 7300 2253
rect 7370 2167 7400 2253
rect 7470 2167 7500 2253
rect 7670 2167 7700 2253
rect 10170 3517 10200 3603
rect 10270 3517 10300 3603
rect 10370 3517 10400 3603
rect 10470 3517 10500 3603
rect 10570 3517 10600 3603
rect 11270 3747 11300 3833
rect 11370 3747 11400 3833
rect 11470 3747 11500 3833
rect 11670 3747 11700 3833
rect 11770 3747 11800 3833
rect 11870 3747 11900 3833
rect 11970 3747 12000 3833
rect 12070 3747 12100 3833
rect 10770 3517 10800 3603
rect 10870 3517 10900 3603
rect 10970 3517 11000 3603
rect 11070 3517 11100 3603
rect 11170 3517 11200 3603
rect 11270 3517 11300 3603
rect 11370 3517 11400 3603
rect 9870 3377 9900 3463
rect 9970 3377 10000 3463
rect 10070 3377 10100 3463
rect 10170 3377 10200 3463
rect 10270 3377 10300 3463
rect 10370 3377 10400 3463
rect 10470 3377 10500 3463
rect 10570 3377 10600 3463
rect 10670 3377 10700 3463
rect 10770 3377 10800 3463
rect 10870 3377 10900 3463
rect 10970 3377 11000 3463
rect 11070 3377 11100 3463
rect 11170 3377 11200 3463
rect 11270 3377 11300 3463
rect 11370 3377 11400 3463
rect 9670 3237 9700 3323
rect 9770 3237 9800 3323
rect 9870 3237 9900 3323
rect 9970 3237 10000 3323
rect 10070 3237 10100 3323
rect 10170 3237 10200 3323
rect 10270 3237 10300 3323
rect 8970 3097 9000 3183
rect 9070 3097 9100 3183
rect 9170 3097 9200 3183
rect 9270 3097 9300 3183
rect 9370 3097 9400 3183
rect 9470 3097 9500 3183
rect 9570 3097 9600 3183
rect 9670 3097 9700 3183
rect 9770 3097 9800 3183
rect 9870 3097 9900 3183
rect 8970 2957 9000 3043
rect 9070 2957 9100 3043
rect 9270 2957 9300 3043
rect 9370 2957 9400 3043
rect 10070 3097 10100 3183
rect 10270 3097 10300 3183
rect 10470 3237 10500 3323
rect 12270 3747 12300 3833
rect 12370 3747 12400 3833
rect 12470 3747 12500 3833
rect 12570 3747 12600 3833
rect 12670 3747 12700 3833
rect 12770 3747 12800 3833
rect 12970 3747 13000 3833
rect 13070 3747 13100 3833
rect 13280 3747 13310 3833
rect 13380 3747 13410 3833
rect 13480 3747 13510 3833
rect 13580 3747 13610 3833
rect 11570 3517 11600 3603
rect 11670 3517 11700 3603
rect 11770 3517 11800 3603
rect 11870 3517 11900 3603
rect 11970 3517 12000 3603
rect 12070 3517 12100 3603
rect 12170 3517 12200 3603
rect 12270 3517 12300 3603
rect 12370 3517 12400 3603
rect 12470 3517 12500 3603
rect 12570 3517 12600 3603
rect 12670 3517 12700 3603
rect 12770 3517 12800 3603
rect 12970 3517 13000 3603
rect 13070 3517 13100 3603
rect 13280 3517 13310 3603
rect 13380 3517 13410 3603
rect 13480 3517 13510 3603
rect 13580 3517 13610 3603
rect 11570 3377 11600 3463
rect 11670 3377 11700 3463
rect 11770 3377 11800 3463
rect 11870 3377 11900 3463
rect 11970 3377 12000 3463
rect 12070 3377 12100 3463
rect 12270 3377 12300 3463
rect 12370 3377 12400 3463
rect 12470 3377 12500 3463
rect 12570 3377 12600 3463
rect 12670 3377 12700 3463
rect 12770 3377 12800 3463
rect 12970 3377 13000 3463
rect 13070 3377 13100 3463
rect 13280 3377 13310 3463
rect 13380 3377 13410 3463
rect 13480 3377 13510 3463
rect 13580 3377 13610 3463
rect 10670 3237 10700 3323
rect 10770 3237 10800 3323
rect 10870 3237 10900 3323
rect 10970 3237 11000 3323
rect 11070 3237 11100 3323
rect 11170 3237 11200 3323
rect 11270 3237 11300 3323
rect 11370 3237 11400 3323
rect 11470 3237 11500 3323
rect 11570 3237 11600 3323
rect 11670 3237 11700 3323
rect 11770 3237 11800 3323
rect 11870 3237 11900 3323
rect 11970 3237 12000 3323
rect 12070 3237 12100 3323
rect 12170 3237 12200 3323
rect 12270 3237 12300 3323
rect 12370 3237 12400 3323
rect 10470 3097 10500 3183
rect 10570 3097 10600 3183
rect 10670 3097 10700 3183
rect 10770 3097 10800 3183
rect 10970 3097 11000 3183
rect 11070 3097 11100 3183
rect 11170 3097 11200 3183
rect 11270 3097 11300 3183
rect 11370 3097 11400 3183
rect 11470 3097 11500 3183
rect 9570 2957 9600 3043
rect 9670 2957 9700 3043
rect 9770 2957 9800 3043
rect 9870 2957 9900 3043
rect 9970 2957 10000 3043
rect 10070 2957 10100 3043
rect 10170 2957 10200 3043
rect 10270 2957 10300 3043
rect 10370 2957 10400 3043
rect 10470 2957 10500 3043
rect 10570 2957 10600 3043
rect 10670 2957 10700 3043
rect 10770 2957 10800 3043
rect 10870 2957 10900 3043
rect 10970 2957 11000 3043
rect 11070 2957 11100 3043
rect 11170 2957 11200 3043
rect 11270 2957 11300 3043
rect 11370 2957 11400 3043
rect 11470 2957 11500 3043
rect 8870 2817 8900 2903
rect 8970 2817 9000 2903
rect 9070 2817 9100 2903
rect 9170 2817 9200 2903
rect 9270 2817 9300 2903
rect 9370 2817 9400 2903
rect 9470 2817 9500 2903
rect 9570 2817 9600 2903
rect 9670 2817 9700 2903
rect 9770 2817 9800 2903
rect 9870 2817 9900 2903
rect 9970 2817 10000 2903
rect 10070 2817 10100 2903
rect 10170 2817 10200 2903
rect 10270 2817 10300 2903
rect 10370 2817 10400 2903
rect 10470 2817 10500 2903
rect 8870 2677 8900 2763
rect 9070 2677 9100 2763
rect 8870 2537 8900 2623
rect 8970 2537 9000 2623
rect 9270 2677 9300 2763
rect 9170 2537 9200 2623
rect 9470 2677 9500 2763
rect 9370 2537 9400 2623
rect 9470 2537 9500 2623
rect 9670 2677 9700 2763
rect 9770 2677 9800 2763
rect 9870 2677 9900 2763
rect 9670 2537 9700 2623
rect 9770 2537 9800 2623
rect 9870 2537 9900 2623
rect 8670 2307 8700 2393
rect 8770 2307 8800 2393
rect 8870 2307 8900 2393
rect 8970 2307 9000 2393
rect 9070 2307 9100 2393
rect 9170 2307 9200 2393
rect 9270 2307 9300 2393
rect 9370 2307 9400 2393
rect 9470 2307 9500 2393
rect 9570 2307 9600 2393
rect 7870 2167 7900 2253
rect 7970 2167 8000 2253
rect 8070 2167 8100 2253
rect 8170 2167 8200 2253
rect 8270 2167 8300 2253
rect 8370 2167 8400 2253
rect 8470 2167 8500 2253
rect 8570 2167 8600 2253
rect 8670 2167 8700 2253
rect 8770 2167 8800 2253
rect 6970 2027 7000 2113
rect 7070 2027 7100 2113
rect 7170 2027 7200 2113
rect 7270 2027 7300 2113
rect 7370 2027 7400 2113
rect 7470 2027 7500 2113
rect 7570 2027 7600 2113
rect 7670 2027 7700 2113
rect 7770 2027 7800 2113
rect 7870 2027 7900 2113
rect 7970 2027 8000 2113
rect 8070 2027 8100 2113
rect 6870 1887 6900 1973
rect 8270 2027 8300 2113
rect 8470 2027 8500 2113
rect 8570 2027 8600 2113
rect 8670 2027 8700 2113
rect 8970 2167 9000 2253
rect 8870 2027 8900 2113
rect 9170 2167 9200 2253
rect 9070 2027 9100 2113
rect 9170 2027 9200 2113
rect 9370 2167 9400 2253
rect 9470 2167 9500 2253
rect 10070 2677 10100 2763
rect 10170 2677 10200 2763
rect 10270 2677 10300 2763
rect 10370 2677 10400 2763
rect 10670 2817 10700 2903
rect 10770 2817 10800 2903
rect 10870 2817 10900 2903
rect 10970 2817 11000 2903
rect 11070 2817 11100 2903
rect 11170 2817 11200 2903
rect 11270 2817 11300 2903
rect 10570 2677 10600 2763
rect 12570 3237 12600 3323
rect 12670 3237 12700 3323
rect 12770 3237 12800 3323
rect 12970 3237 13000 3323
rect 13070 3237 13100 3323
rect 13280 3237 13310 3323
rect 13380 3237 13410 3323
rect 13480 3237 13510 3323
rect 13580 3237 13610 3323
rect 11670 3097 11700 3183
rect 11770 3097 11800 3183
rect 11870 3097 11900 3183
rect 11970 3097 12000 3183
rect 12070 3097 12100 3183
rect 12170 3097 12200 3183
rect 12270 3097 12300 3183
rect 12370 3097 12400 3183
rect 12470 3097 12500 3183
rect 12570 3097 12600 3183
rect 12670 3097 12700 3183
rect 12770 3097 12800 3183
rect 12970 3097 13000 3183
rect 13070 3097 13100 3183
rect 13280 3097 13310 3183
rect 13380 3097 13410 3183
rect 13480 3097 13510 3183
rect 13580 3097 13610 3183
rect 11670 2957 11700 3043
rect 11770 2957 11800 3043
rect 11870 2957 11900 3043
rect 11970 2957 12000 3043
rect 12070 2957 12100 3043
rect 12170 2957 12200 3043
rect 12270 2957 12300 3043
rect 12370 2957 12400 3043
rect 12470 2957 12500 3043
rect 12570 2957 12600 3043
rect 12670 2957 12700 3043
rect 12770 2957 12800 3043
rect 12970 2957 13000 3043
rect 13070 2957 13100 3043
rect 13280 2957 13310 3043
rect 13380 2957 13410 3043
rect 13480 2957 13510 3043
rect 13580 2957 13610 3043
rect 11470 2817 11500 2903
rect 11570 2817 11600 2903
rect 11670 2817 11700 2903
rect 11770 2817 11800 2903
rect 10770 2677 10800 2763
rect 10870 2677 10900 2763
rect 10970 2677 11000 2763
rect 11070 2677 11100 2763
rect 11170 2677 11200 2763
rect 11270 2677 11300 2763
rect 11370 2677 11400 2763
rect 11470 2677 11500 2763
rect 11570 2677 11600 2763
rect 10070 2537 10100 2623
rect 10170 2537 10200 2623
rect 10270 2537 10300 2623
rect 10370 2537 10400 2623
rect 10470 2537 10500 2623
rect 10570 2537 10600 2623
rect 10670 2537 10700 2623
rect 10770 2537 10800 2623
rect 10870 2537 10900 2623
rect 11070 2537 11100 2623
rect 11270 2537 11300 2623
rect 11470 2537 11500 2623
rect 11570 2537 11600 2623
rect 11970 2817 12000 2903
rect 12070 2817 12100 2903
rect 12170 2817 12200 2903
rect 12270 2817 12300 2903
rect 12370 2817 12400 2903
rect 12470 2817 12500 2903
rect 12570 2817 12600 2903
rect 12670 2817 12700 2903
rect 12770 2817 12800 2903
rect 12970 2817 13000 2903
rect 13070 2817 13100 2903
rect 13280 2817 13310 2903
rect 13380 2817 13410 2903
rect 13480 2817 13510 2903
rect 13580 2817 13610 2903
rect 11770 2677 11800 2763
rect 11870 2677 11900 2763
rect 11970 2677 12000 2763
rect 12070 2677 12100 2763
rect 12170 2677 12200 2763
rect 12270 2677 12300 2763
rect 12370 2677 12400 2763
rect 12470 2677 12500 2763
rect 12570 2677 12600 2763
rect 12670 2677 12700 2763
rect 12770 2677 12800 2763
rect 12970 2677 13000 2763
rect 13070 2677 13100 2763
rect 13280 2677 13310 2763
rect 13380 2677 13410 2763
rect 13480 2677 13510 2763
rect 13580 2677 13610 2763
rect 11770 2537 11800 2623
rect 11870 2537 11900 2623
rect 11970 2537 12000 2623
rect 12070 2537 12100 2623
rect 12170 2537 12200 2623
rect 12270 2537 12300 2623
rect 12370 2537 12400 2623
rect 12470 2537 12500 2623
rect 12570 2537 12600 2623
rect 12670 2537 12700 2623
rect 12770 2537 12800 2623
rect 12970 2537 13000 2623
rect 13070 2537 13100 2623
rect 13280 2537 13310 2623
rect 13380 2537 13410 2623
rect 13480 2537 13510 2623
rect 13580 2537 13610 2623
rect 9770 2307 9800 2393
rect 9870 2307 9900 2393
rect 9970 2307 10000 2393
rect 10070 2307 10100 2393
rect 10170 2307 10200 2393
rect 10270 2307 10300 2393
rect 10370 2307 10400 2393
rect 10470 2307 10500 2393
rect 10570 2307 10600 2393
rect 10670 2307 10700 2393
rect 10770 2307 10800 2393
rect 10870 2307 10900 2393
rect 10970 2307 11000 2393
rect 11070 2307 11100 2393
rect 11170 2307 11200 2393
rect 11270 2307 11300 2393
rect 11370 2307 11400 2393
rect 11470 2307 11500 2393
rect 11570 2307 11600 2393
rect 11670 2307 11700 2393
rect 9670 2167 9700 2253
rect 9770 2167 9800 2253
rect 9870 2167 9900 2253
rect 9970 2167 10000 2253
rect 10070 2167 10100 2253
rect 10170 2167 10200 2253
rect 10270 2167 10300 2253
rect 10370 2167 10400 2253
rect 10470 2167 10500 2253
rect 11870 2307 11900 2393
rect 12070 2307 12100 2393
rect 12170 2307 12200 2393
rect 12270 2307 12300 2393
rect 12370 2307 12400 2393
rect 12470 2307 12500 2393
rect 10670 2167 10700 2253
rect 10770 2167 10800 2253
rect 10870 2167 10900 2253
rect 10970 2167 11000 2253
rect 11070 2167 11100 2253
rect 11170 2167 11200 2253
rect 11270 2167 11300 2253
rect 11370 2167 11400 2253
rect 11470 2167 11500 2253
rect 11570 2167 11600 2253
rect 11670 2167 11700 2253
rect 11770 2167 11800 2253
rect 11870 2167 11900 2253
rect 11970 2167 12000 2253
rect 9370 2027 9400 2113
rect 9470 2027 9500 2113
rect 9570 2027 9600 2113
rect 9670 2027 9700 2113
rect 9770 2027 9800 2113
rect 9870 2027 9900 2113
rect 9970 2027 10000 2113
rect 10070 2027 10100 2113
rect 10170 2027 10200 2113
rect 10270 2027 10300 2113
rect 10370 2027 10400 2113
rect 10470 2027 10500 2113
rect 10570 2027 10600 2113
rect 10670 2027 10700 2113
rect 10770 2027 10800 2113
rect 10870 2027 10900 2113
rect 10970 2027 11000 2113
rect 11070 2027 11100 2113
rect 11170 2027 11200 2113
rect 7070 1887 7100 1973
rect 7170 1887 7200 1973
rect 7270 1887 7300 1973
rect 7370 1887 7400 1973
rect 7470 1887 7500 1973
rect 7570 1887 7600 1973
rect 7670 1887 7700 1973
rect 7770 1887 7800 1973
rect 7870 1887 7900 1973
rect 7970 1887 8000 1973
rect 8070 1887 8100 1973
rect 8170 1887 8200 1973
rect 8270 1887 8300 1973
rect 8370 1887 8400 1973
rect 8470 1887 8500 1973
rect 8570 1887 8600 1973
rect 8670 1887 8700 1973
rect 8770 1887 8800 1973
rect 8870 1887 8900 1973
rect 8970 1887 9000 1973
rect 9070 1887 9100 1973
rect 9170 1887 9200 1973
rect 9270 1887 9300 1973
rect 9370 1887 9400 1973
rect 9470 1887 9500 1973
rect 9570 1887 9600 1973
rect 9670 1887 9700 1973
rect 9770 1887 9800 1973
rect 9870 1887 9900 1973
rect 9970 1887 10000 1973
rect 10070 1887 10100 1973
rect 10170 1887 10200 1973
rect 10270 1887 10300 1973
rect 10370 1887 10400 1973
rect 10470 1887 10500 1973
rect 10570 1887 10600 1973
rect 10670 1887 10700 1973
rect 10770 1887 10800 1973
rect 10870 1887 10900 1973
rect 10970 1887 11000 1973
rect 6470 1747 6500 1833
rect 6570 1747 6600 1833
rect 6670 1747 6700 1833
rect 6770 1747 6800 1833
rect 6870 1747 6900 1833
rect 6970 1747 7000 1833
rect 7070 1747 7100 1833
rect 6270 1607 6300 1693
rect 6370 1607 6400 1693
rect 6470 1607 6500 1693
rect 6170 1467 6200 1553
rect 6270 1467 6300 1553
rect 5270 1327 5300 1413
rect 5370 1327 5400 1413
rect 5470 1327 5500 1413
rect 5570 1327 5600 1413
rect 5670 1327 5700 1413
rect 5770 1327 5800 1413
rect 5870 1327 5900 1413
rect 5970 1327 6000 1413
rect 6070 1327 6100 1413
rect 6170 1327 6200 1413
rect 4770 1097 4800 1183
rect 4870 1097 4900 1183
rect 4970 1097 5000 1183
rect 5070 1097 5100 1183
rect 5170 1097 5200 1183
rect 5270 1097 5300 1183
rect 5370 1097 5400 1183
rect 3970 957 4000 1043
rect 4070 957 4100 1043
rect 4170 957 4200 1043
rect 4270 957 4300 1043
rect 4370 957 4400 1043
rect 4470 957 4500 1043
rect 4570 957 4600 1043
rect 4670 957 4700 1043
rect 4770 957 4800 1043
rect 4970 957 5000 1043
rect 5070 957 5100 1043
rect 5170 957 5200 1043
rect 5270 957 5300 1043
rect 7270 1747 7300 1833
rect 7370 1747 7400 1833
rect 7570 1747 7600 1833
rect 7670 1747 7700 1833
rect 7870 1747 7900 1833
rect 7970 1747 8000 1833
rect 8170 1747 8200 1833
rect 8270 1747 8300 1833
rect 8370 1747 8400 1833
rect 8470 1747 8500 1833
rect 8570 1747 8600 1833
rect 8770 1747 8800 1833
rect 8870 1747 8900 1833
rect 8970 1747 9000 1833
rect 9070 1747 9100 1833
rect 9170 1747 9200 1833
rect 9270 1747 9300 1833
rect 9370 1747 9400 1833
rect 9470 1747 9500 1833
rect 9570 1747 9600 1833
rect 9670 1747 9700 1833
rect 9770 1747 9800 1833
rect 6670 1607 6700 1693
rect 6770 1607 6800 1693
rect 6870 1607 6900 1693
rect 6970 1607 7000 1693
rect 7070 1607 7100 1693
rect 7170 1607 7200 1693
rect 7270 1607 7300 1693
rect 7370 1607 7400 1693
rect 7470 1607 7500 1693
rect 7570 1607 7600 1693
rect 7670 1607 7700 1693
rect 7770 1607 7800 1693
rect 7870 1607 7900 1693
rect 7970 1607 8000 1693
rect 8070 1607 8100 1693
rect 8170 1607 8200 1693
rect 8270 1607 8300 1693
rect 8370 1607 8400 1693
rect 8470 1607 8500 1693
rect 8570 1607 8600 1693
rect 8670 1607 8700 1693
rect 8770 1607 8800 1693
rect 8870 1607 8900 1693
rect 8970 1607 9000 1693
rect 9070 1607 9100 1693
rect 9170 1607 9200 1693
rect 9270 1607 9300 1693
rect 9370 1607 9400 1693
rect 9470 1607 9500 1693
rect 6470 1467 6500 1553
rect 6570 1467 6600 1553
rect 6670 1467 6700 1553
rect 6770 1467 6800 1553
rect 6870 1467 6900 1553
rect 6970 1467 7000 1553
rect 7070 1467 7100 1553
rect 7170 1467 7200 1553
rect 7270 1467 7300 1553
rect 7370 1467 7400 1553
rect 7470 1467 7500 1553
rect 7570 1467 7600 1553
rect 7670 1467 7700 1553
rect 6370 1327 6400 1413
rect 6570 1327 6600 1413
rect 6670 1327 6700 1413
rect 6870 1327 6900 1413
rect 5570 1097 5600 1183
rect 5670 1097 5700 1183
rect 5770 1097 5800 1183
rect 5870 1097 5900 1183
rect 5970 1097 6000 1183
rect 6070 1097 6100 1183
rect 6170 1097 6200 1183
rect 6270 1097 6300 1183
rect 6370 1097 6400 1183
rect 6470 1097 6500 1183
rect 6570 1097 6600 1183
rect 6670 1097 6700 1183
rect 5470 957 5500 1043
rect 5570 957 5600 1043
rect 5670 957 5700 1043
rect 5770 957 5800 1043
rect 5870 957 5900 1043
rect 5970 957 6000 1043
rect 6070 957 6100 1043
rect 6170 957 6200 1043
rect 6270 957 6300 1043
rect 6370 957 6400 1043
rect 7870 1467 7900 1553
rect 7070 1327 7100 1413
rect 7170 1327 7200 1413
rect 7270 1327 7300 1413
rect 7370 1327 7400 1413
rect 7470 1327 7500 1413
rect 7570 1327 7600 1413
rect 7670 1327 7700 1413
rect 7770 1327 7800 1413
rect 7870 1327 7900 1413
rect 8070 1467 8100 1553
rect 8170 1467 8200 1553
rect 8270 1467 8300 1553
rect 8370 1467 8400 1553
rect 8470 1467 8500 1553
rect 8670 1467 8700 1553
rect 8770 1467 8800 1553
rect 8870 1467 8900 1553
rect 8970 1467 9000 1553
rect 9070 1467 9100 1553
rect 9170 1467 9200 1553
rect 9270 1467 9300 1553
rect 8070 1327 8100 1413
rect 8170 1327 8200 1413
rect 8270 1327 8300 1413
rect 8370 1327 8400 1413
rect 8470 1327 8500 1413
rect 8570 1327 8600 1413
rect 8670 1327 8700 1413
rect 8770 1327 8800 1413
rect 8870 1327 8900 1413
rect 8970 1327 9000 1413
rect 9070 1327 9100 1413
rect 9170 1327 9200 1413
rect 9270 1327 9300 1413
rect 9970 1747 10000 1833
rect 10170 1747 10200 1833
rect 10370 1747 10400 1833
rect 10570 1747 10600 1833
rect 10670 1747 10700 1833
rect 11170 1887 11200 1973
rect 11370 2027 11400 2113
rect 12170 2167 12200 2253
rect 12270 2167 12300 2253
rect 12670 2307 12700 2393
rect 12770 2307 12800 2393
rect 12970 2307 13000 2393
rect 13070 2307 13100 2393
rect 13280 2307 13310 2393
rect 13380 2307 13410 2393
rect 13480 2307 13510 2393
rect 13580 2307 13610 2393
rect 12470 2167 12500 2253
rect 12570 2167 12600 2253
rect 11570 2027 11600 2113
rect 11670 2027 11700 2113
rect 11770 2027 11800 2113
rect 11870 2027 11900 2113
rect 11970 2027 12000 2113
rect 12070 2027 12100 2113
rect 12170 2027 12200 2113
rect 12270 2027 12300 2113
rect 12370 2027 12400 2113
rect 12470 2027 12500 2113
rect 12570 2027 12600 2113
rect 11370 1887 11400 1973
rect 11470 1887 11500 1973
rect 11570 1887 11600 1973
rect 11670 1887 11700 1973
rect 11770 1887 11800 1973
rect 11870 1887 11900 1973
rect 11970 1887 12000 1973
rect 12070 1887 12100 1973
rect 12170 1887 12200 1973
rect 12270 1887 12300 1973
rect 12370 1887 12400 1973
rect 12470 1887 12500 1973
rect 12570 1887 12600 1973
rect 10870 1747 10900 1833
rect 10970 1747 11000 1833
rect 11070 1747 11100 1833
rect 11170 1747 11200 1833
rect 11270 1747 11300 1833
rect 11370 1747 11400 1833
rect 11470 1747 11500 1833
rect 11570 1747 11600 1833
rect 9670 1607 9700 1693
rect 9770 1607 9800 1693
rect 9870 1607 9900 1693
rect 9970 1607 10000 1693
rect 10070 1607 10100 1693
rect 10170 1607 10200 1693
rect 10270 1607 10300 1693
rect 10370 1607 10400 1693
rect 10470 1607 10500 1693
rect 10570 1607 10600 1693
rect 10670 1607 10700 1693
rect 10770 1607 10800 1693
rect 10870 1607 10900 1693
rect 9470 1467 9500 1553
rect 9570 1467 9600 1553
rect 9670 1467 9700 1553
rect 9770 1467 9800 1553
rect 9870 1467 9900 1553
rect 9970 1467 10000 1553
rect 10070 1467 10100 1553
rect 10170 1467 10200 1553
rect 10270 1467 10300 1553
rect 10370 1467 10400 1553
rect 10470 1467 10500 1553
rect 10570 1467 10600 1553
rect 10670 1467 10700 1553
rect 10770 1467 10800 1553
rect 10870 1467 10900 1553
rect 9470 1327 9500 1413
rect 9570 1327 9600 1413
rect 9670 1327 9700 1413
rect 9770 1327 9800 1413
rect 9870 1327 9900 1413
rect 9970 1327 10000 1413
rect 10070 1327 10100 1413
rect 10170 1327 10200 1413
rect 6870 1097 6900 1183
rect 6970 1097 7000 1183
rect 7070 1097 7100 1183
rect 7170 1097 7200 1183
rect 7270 1097 7300 1183
rect 7370 1097 7400 1183
rect 7470 1097 7500 1183
rect 7570 1097 7600 1183
rect 7670 1097 7700 1183
rect 7770 1097 7800 1183
rect 7870 1097 7900 1183
rect 7970 1097 8000 1183
rect 8070 1097 8100 1183
rect 8170 1097 8200 1183
rect 8270 1097 8300 1183
rect 8370 1097 8400 1183
rect 8470 1097 8500 1183
rect 8570 1097 8600 1183
rect 8670 1097 8700 1183
rect 8770 1097 8800 1183
rect 8870 1097 8900 1183
rect 8970 1097 9000 1183
rect 9070 1097 9100 1183
rect 9170 1097 9200 1183
rect 9270 1097 9300 1183
rect 9370 1097 9400 1183
rect 9470 1097 9500 1183
rect 9570 1097 9600 1183
rect 6570 957 6600 1043
rect 6670 957 6700 1043
rect 6770 957 6800 1043
rect 6870 957 6900 1043
rect 3970 817 4000 903
rect 4070 817 4100 903
rect 4170 817 4200 903
rect 4270 817 4300 903
rect 4370 817 4400 903
rect 4470 817 4500 903
rect 4570 817 4600 903
rect 4670 817 4700 903
rect 4770 817 4800 903
rect 4870 817 4900 903
rect 4970 817 5000 903
rect 5070 817 5100 903
rect 5170 817 5200 903
rect 5270 817 5300 903
rect 5370 817 5400 903
rect 5470 817 5500 903
rect 5570 817 5600 903
rect 5670 817 5700 903
rect 5770 817 5800 903
rect 5870 817 5900 903
rect 5970 817 6000 903
rect 6070 817 6100 903
rect 6170 817 6200 903
rect 6270 817 6300 903
rect 6370 817 6400 903
rect 6470 817 6500 903
rect 6570 817 6600 903
rect 3770 677 3800 763
rect 3870 677 3900 763
rect 3970 677 4000 763
rect 4070 677 4100 763
rect 4170 677 4200 763
rect 4270 677 4300 763
rect 4370 677 4400 763
rect 4470 677 4500 763
rect 4570 677 4600 763
rect 2870 537 2900 623
rect 2970 537 3000 623
rect 3070 537 3100 623
rect 3170 537 3200 623
rect 3270 537 3300 623
rect 3370 537 3400 623
rect 3470 537 3500 623
rect 3570 537 3600 623
rect 3670 537 3700 623
rect 3770 537 3800 623
rect 3870 537 3900 623
rect 4070 537 4100 623
rect 4770 677 4800 763
rect 4870 677 4900 763
rect 4970 677 5000 763
rect 5070 677 5100 763
rect 4270 537 4300 623
rect 4370 537 4400 623
rect 4470 537 4500 623
rect 4570 537 4600 623
rect 4670 537 4700 623
rect 4770 537 4800 623
rect 2770 397 2800 483
rect 2870 397 2900 483
rect 2970 397 3000 483
rect 3070 397 3100 483
rect 3170 397 3200 483
rect 3270 397 3300 483
rect 3370 397 3400 483
rect 3470 397 3500 483
rect 3570 397 3600 483
rect 3670 397 3700 483
rect 3770 397 3800 483
rect 3870 397 3900 483
rect 3970 397 4000 483
rect 4070 397 4100 483
rect 4170 397 4200 483
rect 4270 397 4300 483
rect 4370 397 4400 483
rect 1870 257 1900 343
rect 1970 257 2000 343
rect 2070 257 2100 343
rect 2170 257 2200 343
rect 2270 257 2300 343
rect 2370 257 2400 343
rect 2470 257 2500 343
rect 2570 257 2600 343
rect 2670 257 2700 343
rect 2770 257 2800 343
rect 1770 117 1800 203
rect 2970 257 3000 343
rect 4970 537 5000 623
rect 5270 677 5300 763
rect 5370 677 5400 763
rect 5470 677 5500 763
rect 5570 677 5600 763
rect 5670 677 5700 763
rect 5170 537 5200 623
rect 4570 397 4600 483
rect 4670 397 4700 483
rect 4770 397 4800 483
rect 4870 397 4900 483
rect 4970 397 5000 483
rect 5070 397 5100 483
rect 3170 257 3200 343
rect 3270 257 3300 343
rect 3370 257 3400 343
rect 3470 257 3500 343
rect 3570 257 3600 343
rect 3670 257 3700 343
rect 3770 257 3800 343
rect 3870 257 3900 343
rect 3970 257 4000 343
rect 4070 257 4100 343
rect 4170 257 4200 343
rect 4270 257 4300 343
rect 4370 257 4400 343
rect 4470 257 4500 343
rect 4670 257 4700 343
rect 4770 257 4800 343
rect 4970 257 5000 343
rect 5870 677 5900 763
rect 5970 677 6000 763
rect 6070 677 6100 763
rect 6170 677 6200 763
rect 6370 677 6400 763
rect 7070 957 7100 1043
rect 7270 957 7300 1043
rect 6770 817 6800 903
rect 6870 817 6900 903
rect 6970 817 7000 903
rect 7070 817 7100 903
rect 7170 817 7200 903
rect 7270 817 7300 903
rect 6570 677 6600 763
rect 6670 677 6700 763
rect 6770 677 6800 763
rect 6870 677 6900 763
rect 6970 677 7000 763
rect 7470 957 7500 1043
rect 7570 957 7600 1043
rect 7670 957 7700 1043
rect 7770 957 7800 1043
rect 7870 957 7900 1043
rect 7970 957 8000 1043
rect 8070 957 8100 1043
rect 8170 957 8200 1043
rect 8270 957 8300 1043
rect 8370 957 8400 1043
rect 8470 957 8500 1043
rect 8570 957 8600 1043
rect 7470 817 7500 903
rect 7670 817 7700 903
rect 7870 817 7900 903
rect 8070 817 8100 903
rect 8170 817 8200 903
rect 8270 817 8300 903
rect 8370 817 8400 903
rect 8470 817 8500 903
rect 8570 817 8600 903
rect 8770 957 8800 1043
rect 8770 817 8800 903
rect 8970 957 9000 1043
rect 9070 957 9100 1043
rect 9170 957 9200 1043
rect 9270 957 9300 1043
rect 9370 957 9400 1043
rect 9470 957 9500 1043
rect 11770 1747 11800 1833
rect 11870 1747 11900 1833
rect 11070 1607 11100 1693
rect 11170 1607 11200 1693
rect 11270 1607 11300 1693
rect 11370 1607 11400 1693
rect 11470 1607 11500 1693
rect 11570 1607 11600 1693
rect 11670 1607 11700 1693
rect 11070 1467 11100 1553
rect 10370 1327 10400 1413
rect 10470 1327 10500 1413
rect 10570 1327 10600 1413
rect 10670 1327 10700 1413
rect 10770 1327 10800 1413
rect 10870 1327 10900 1413
rect 10970 1327 11000 1413
rect 11070 1327 11100 1413
rect 12770 2167 12800 2253
rect 12970 2167 13000 2253
rect 13070 2167 13100 2253
rect 13280 2167 13310 2253
rect 13380 2167 13410 2253
rect 13480 2167 13510 2253
rect 13580 2167 13610 2253
rect 12770 2027 12800 2113
rect 12970 2027 13000 2113
rect 13070 2027 13100 2113
rect 13280 2027 13310 2113
rect 13380 2027 13410 2113
rect 13480 2027 13510 2113
rect 13580 2027 13610 2113
rect 12770 1887 12800 1973
rect 12970 1887 13000 1973
rect 13070 1887 13100 1973
rect 13280 1887 13310 1973
rect 13380 1887 13410 1973
rect 13480 1887 13510 1973
rect 13580 1887 13610 1973
rect 12070 1747 12100 1833
rect 12170 1747 12200 1833
rect 12270 1747 12300 1833
rect 12370 1747 12400 1833
rect 12470 1747 12500 1833
rect 12570 1747 12600 1833
rect 12670 1747 12700 1833
rect 12770 1747 12800 1833
rect 12970 1747 13000 1833
rect 13070 1747 13100 1833
rect 13280 1747 13310 1833
rect 13380 1747 13410 1833
rect 13480 1747 13510 1833
rect 13580 1747 13610 1833
rect 11870 1607 11900 1693
rect 11970 1607 12000 1693
rect 12070 1607 12100 1693
rect 12170 1607 12200 1693
rect 12270 1607 12300 1693
rect 12370 1607 12400 1693
rect 12470 1607 12500 1693
rect 12570 1607 12600 1693
rect 12670 1607 12700 1693
rect 12770 1607 12800 1693
rect 12970 1607 13000 1693
rect 13070 1607 13100 1693
rect 13280 1607 13310 1693
rect 13380 1607 13410 1693
rect 13480 1607 13510 1693
rect 13580 1607 13610 1693
rect 11270 1467 11300 1553
rect 11370 1467 11400 1553
rect 11470 1467 11500 1553
rect 11570 1467 11600 1553
rect 11670 1467 11700 1553
rect 11770 1467 11800 1553
rect 11870 1467 11900 1553
rect 11970 1467 12000 1553
rect 11270 1327 11300 1413
rect 11370 1327 11400 1413
rect 11470 1327 11500 1413
rect 11570 1327 11600 1413
rect 11670 1327 11700 1413
rect 9770 1097 9800 1183
rect 9870 1097 9900 1183
rect 9970 1097 10000 1183
rect 10070 1097 10100 1183
rect 10170 1097 10200 1183
rect 10270 1097 10300 1183
rect 10370 1097 10400 1183
rect 10470 1097 10500 1183
rect 10570 1097 10600 1183
rect 10670 1097 10700 1183
rect 10770 1097 10800 1183
rect 10870 1097 10900 1183
rect 10970 1097 11000 1183
rect 9670 957 9700 1043
rect 9770 957 9800 1043
rect 9870 957 9900 1043
rect 8970 817 9000 903
rect 9070 817 9100 903
rect 9170 817 9200 903
rect 9270 817 9300 903
rect 9370 817 9400 903
rect 9470 817 9500 903
rect 9570 817 9600 903
rect 9670 817 9700 903
rect 9770 817 9800 903
rect 9870 817 9900 903
rect 7170 677 7200 763
rect 7270 677 7300 763
rect 7370 677 7400 763
rect 7470 677 7500 763
rect 7570 677 7600 763
rect 7670 677 7700 763
rect 7770 677 7800 763
rect 7870 677 7900 763
rect 7970 677 8000 763
rect 8070 677 8100 763
rect 8170 677 8200 763
rect 8270 677 8300 763
rect 8370 677 8400 763
rect 8470 677 8500 763
rect 8570 677 8600 763
rect 8670 677 8700 763
rect 8770 677 8800 763
rect 8870 677 8900 763
rect 8970 677 9000 763
rect 9070 677 9100 763
rect 5370 537 5400 623
rect 5470 537 5500 623
rect 5570 537 5600 623
rect 5670 537 5700 623
rect 5770 537 5800 623
rect 5870 537 5900 623
rect 5970 537 6000 623
rect 6070 537 6100 623
rect 6170 537 6200 623
rect 6270 537 6300 623
rect 6370 537 6400 623
rect 6470 537 6500 623
rect 6570 537 6600 623
rect 6670 537 6700 623
rect 6770 537 6800 623
rect 6870 537 6900 623
rect 6970 537 7000 623
rect 7070 537 7100 623
rect 7170 537 7200 623
rect 7270 537 7300 623
rect 7370 537 7400 623
rect 7470 537 7500 623
rect 7570 537 7600 623
rect 7670 537 7700 623
rect 7770 537 7800 623
rect 7870 537 7900 623
rect 7970 537 8000 623
rect 8070 537 8100 623
rect 8170 537 8200 623
rect 8270 537 8300 623
rect 5270 397 5300 483
rect 5470 397 5500 483
rect 5570 397 5600 483
rect 5670 397 5700 483
rect 5770 397 5800 483
rect 5870 397 5900 483
rect 5970 397 6000 483
rect 6070 397 6100 483
rect 5170 257 5200 343
rect 5270 257 5300 343
rect 5370 257 5400 343
rect 5470 257 5500 343
rect 5570 257 5600 343
rect 5670 257 5700 343
rect 5770 257 5800 343
rect 5970 257 6000 343
rect 6270 397 6300 483
rect 6370 397 6400 483
rect 6170 257 6200 343
rect 6370 257 6400 343
rect 6570 397 6600 483
rect 6670 397 6700 483
rect 6770 397 6800 483
rect 6870 397 6900 483
rect 6970 397 7000 483
rect 7070 397 7100 483
rect 6570 257 6600 343
rect 6770 257 6800 343
rect 7270 397 7300 483
rect 7470 397 7500 483
rect 7670 397 7700 483
rect 7770 397 7800 483
rect 7870 397 7900 483
rect 7970 397 8000 483
rect 8070 397 8100 483
rect 8170 397 8200 483
rect 8270 397 8300 483
rect 6970 257 7000 343
rect 7070 257 7100 343
rect 7170 257 7200 343
rect 7270 257 7300 343
rect 7370 257 7400 343
rect 7470 257 7500 343
rect 7570 257 7600 343
rect 7670 257 7700 343
rect 7770 257 7800 343
rect 1970 117 2000 203
rect 2070 117 2100 203
rect 2170 117 2200 203
rect 2270 117 2300 203
rect 2370 117 2400 203
rect 2470 117 2500 203
rect 2570 117 2600 203
rect 2670 117 2700 203
rect 2770 117 2800 203
rect 2870 117 2900 203
rect 2970 117 3000 203
rect 3070 117 3100 203
rect 3170 117 3200 203
rect 3270 117 3300 203
rect 3370 117 3400 203
rect 3470 117 3500 203
rect 3570 117 3600 203
rect 3670 117 3700 203
rect 3770 117 3800 203
rect 3870 117 3900 203
rect 3970 117 4000 203
rect 4070 117 4100 203
rect 4170 117 4200 203
rect 4270 117 4300 203
rect 4370 117 4400 203
rect 4470 117 4500 203
rect 4570 117 4600 203
rect 4670 117 4700 203
rect 4770 117 4800 203
rect 4870 117 4900 203
rect 4970 117 5000 203
rect 5070 117 5100 203
rect 5170 117 5200 203
rect 5270 117 5300 203
rect 5370 117 5400 203
rect 5470 117 5500 203
rect 5570 117 5600 203
rect 5670 117 5700 203
rect 5770 117 5800 203
rect 5870 117 5900 203
rect 5970 117 6000 203
rect 6070 117 6100 203
rect 6170 117 6200 203
rect 6270 117 6300 203
rect 6370 117 6400 203
rect 6470 117 6500 203
rect 6570 117 6600 203
rect 6670 117 6700 203
rect 6770 117 6800 203
rect 6870 117 6900 203
rect 6970 117 7000 203
rect 7970 257 8000 343
rect 9270 677 9300 763
rect 9470 677 9500 763
rect 9570 677 9600 763
rect 9770 677 9800 763
rect 10070 957 10100 1043
rect 10170 957 10200 1043
rect 10270 957 10300 1043
rect 11170 1097 11200 1183
rect 11370 1097 11400 1183
rect 10470 957 10500 1043
rect 10570 957 10600 1043
rect 10670 957 10700 1043
rect 10770 957 10800 1043
rect 10870 957 10900 1043
rect 10970 957 11000 1043
rect 11070 957 11100 1043
rect 11170 957 11200 1043
rect 11270 957 11300 1043
rect 10070 817 10100 903
rect 10170 817 10200 903
rect 10270 817 10300 903
rect 10370 817 10400 903
rect 10470 817 10500 903
rect 10570 817 10600 903
rect 10670 817 10700 903
rect 9970 677 10000 763
rect 10070 677 10100 763
rect 10870 817 10900 903
rect 10270 677 10300 763
rect 10370 677 10400 763
rect 10470 677 10500 763
rect 10570 677 10600 763
rect 10670 677 10700 763
rect 10770 677 10800 763
rect 10870 677 10900 763
rect 8470 537 8500 623
rect 8570 537 8600 623
rect 8670 537 8700 623
rect 8770 537 8800 623
rect 8870 537 8900 623
rect 8970 537 9000 623
rect 9070 537 9100 623
rect 9170 537 9200 623
rect 9270 537 9300 623
rect 9370 537 9400 623
rect 9470 537 9500 623
rect 9570 537 9600 623
rect 9670 537 9700 623
rect 9770 537 9800 623
rect 9870 537 9900 623
rect 9970 537 10000 623
rect 10070 537 10100 623
rect 10170 537 10200 623
rect 8470 397 8500 483
rect 8570 397 8600 483
rect 8670 397 8700 483
rect 8770 397 8800 483
rect 8870 397 8900 483
rect 8970 397 9000 483
rect 9070 397 9100 483
rect 9170 397 9200 483
rect 9270 397 9300 483
rect 9370 397 9400 483
rect 9470 397 9500 483
rect 9570 397 9600 483
rect 9670 397 9700 483
rect 9770 397 9800 483
rect 9870 397 9900 483
rect 8170 257 8200 343
rect 8270 257 8300 343
rect 8370 257 8400 343
rect 8470 257 8500 343
rect 8570 257 8600 343
rect 8670 257 8700 343
rect 8870 257 8900 343
rect 8970 257 9000 343
rect 9170 257 9200 343
rect 10070 397 10100 483
rect 10170 397 10200 483
rect 9370 257 9400 343
rect 9470 257 9500 343
rect 9570 257 9600 343
rect 9670 257 9700 343
rect 9770 257 9800 343
rect 9870 257 9900 343
rect 9970 257 10000 343
rect 10070 257 10100 343
rect 10370 537 10400 623
rect 12170 1467 12200 1553
rect 12270 1467 12300 1553
rect 12370 1467 12400 1553
rect 11870 1327 11900 1413
rect 11970 1327 12000 1413
rect 12070 1327 12100 1413
rect 12170 1327 12200 1413
rect 12270 1327 12300 1413
rect 12370 1327 12400 1413
rect 11570 1097 11600 1183
rect 11670 1097 11700 1183
rect 11770 1097 11800 1183
rect 11870 1097 11900 1183
rect 11970 1097 12000 1183
rect 11470 957 11500 1043
rect 11570 957 11600 1043
rect 11770 957 11800 1043
rect 11870 957 11900 1043
rect 11070 817 11100 903
rect 11170 817 11200 903
rect 11270 817 11300 903
rect 11370 817 11400 903
rect 11470 817 11500 903
rect 11570 817 11600 903
rect 11670 817 11700 903
rect 11770 817 11800 903
rect 11870 817 11900 903
rect 11070 677 11100 763
rect 11170 677 11200 763
rect 11270 677 11300 763
rect 11370 677 11400 763
rect 11470 677 11500 763
rect 11570 677 11600 763
rect 11670 677 11700 763
rect 10570 537 10600 623
rect 10670 537 10700 623
rect 10770 537 10800 623
rect 10870 537 10900 623
rect 10970 537 11000 623
rect 11070 537 11100 623
rect 11170 537 11200 623
rect 10370 397 10400 483
rect 10470 397 10500 483
rect 10570 397 10600 483
rect 10670 397 10700 483
rect 10770 397 10800 483
rect 10970 397 11000 483
rect 11070 397 11100 483
rect 12570 1467 12600 1553
rect 12670 1467 12700 1553
rect 12770 1467 12800 1553
rect 12970 1467 13000 1553
rect 13070 1467 13100 1553
rect 13280 1467 13310 1553
rect 13380 1467 13410 1553
rect 13480 1467 13510 1553
rect 13580 1467 13610 1553
rect 12570 1327 12600 1413
rect 12670 1327 12700 1413
rect 12770 1327 12800 1413
rect 12970 1327 13000 1413
rect 13070 1327 13100 1413
rect 13280 1327 13310 1413
rect 13380 1327 13410 1413
rect 13480 1327 13510 1413
rect 13580 1327 13610 1413
rect 12170 1097 12200 1183
rect 12270 1097 12300 1183
rect 12370 1097 12400 1183
rect 12470 1097 12500 1183
rect 12570 1097 12600 1183
rect 12770 1097 12800 1183
rect 12970 1097 13000 1183
rect 13070 1097 13100 1183
rect 13280 1097 13310 1183
rect 13380 1097 13410 1183
rect 13480 1097 13510 1183
rect 13580 1097 13610 1183
rect 12070 957 12100 1043
rect 12170 957 12200 1043
rect 12270 957 12300 1043
rect 12370 957 12400 1043
rect 12470 957 12500 1043
rect 12570 957 12600 1043
rect 12670 957 12700 1043
rect 12770 957 12800 1043
rect 12970 957 13000 1043
rect 13070 957 13100 1043
rect 13280 957 13310 1043
rect 13380 957 13410 1043
rect 13480 957 13510 1043
rect 13580 957 13610 1043
rect 12070 817 12100 903
rect 12170 817 12200 903
rect 12270 817 12300 903
rect 11870 677 11900 763
rect 11970 677 12000 763
rect 12070 677 12100 763
rect 12470 817 12500 903
rect 12670 817 12700 903
rect 12770 817 12800 903
rect 12970 817 13000 903
rect 13070 817 13100 903
rect 13280 817 13310 903
rect 13380 817 13410 903
rect 13480 817 13510 903
rect 13580 817 13610 903
rect 12270 677 12300 763
rect 12370 677 12400 763
rect 12470 677 12500 763
rect 12570 677 12600 763
rect 12670 677 12700 763
rect 12770 677 12800 763
rect 12970 677 13000 763
rect 13070 677 13100 763
rect 13280 677 13310 763
rect 13380 677 13410 763
rect 13480 677 13510 763
rect 13580 677 13610 763
rect 11370 537 11400 623
rect 11470 537 11500 623
rect 11570 537 11600 623
rect 11670 537 11700 623
rect 11770 537 11800 623
rect 11870 537 11900 623
rect 11970 537 12000 623
rect 12070 537 12100 623
rect 12170 537 12200 623
rect 12270 537 12300 623
rect 12370 537 12400 623
rect 12470 537 12500 623
rect 12570 537 12600 623
rect 12670 537 12700 623
rect 12770 537 12800 623
rect 12970 537 13000 623
rect 13070 537 13100 623
rect 13280 537 13310 623
rect 13380 537 13410 623
rect 13480 537 13510 623
rect 13580 537 13610 623
rect 11270 397 11300 483
rect 11470 397 11500 483
rect 11570 397 11600 483
rect 11670 397 11700 483
rect 11770 397 11800 483
rect 11870 397 11900 483
rect 11970 397 12000 483
rect 12070 397 12100 483
rect 12170 397 12200 483
rect 12270 397 12300 483
rect 10270 257 10300 343
rect 10370 257 10400 343
rect 10470 257 10500 343
rect 10570 257 10600 343
rect 10670 257 10700 343
rect 10770 257 10800 343
rect 10870 257 10900 343
rect 10970 257 11000 343
rect 11070 257 11100 343
rect 11170 257 11200 343
rect 11270 257 11300 343
rect 11370 257 11400 343
rect 7170 117 7200 203
rect 7270 117 7300 203
rect 7370 117 7400 203
rect 7470 117 7500 203
rect 7570 117 7600 203
rect 7670 117 7700 203
rect 7770 117 7800 203
rect 7870 117 7900 203
rect 7970 117 8000 203
rect 8070 117 8100 203
rect 8170 117 8200 203
rect 8270 117 8300 203
rect 8370 117 8400 203
rect 8470 117 8500 203
rect 8570 117 8600 203
rect 8670 117 8700 203
rect 8770 117 8800 203
rect 8870 117 8900 203
rect 8970 117 9000 203
rect 9070 117 9100 203
rect 9170 117 9200 203
rect 9270 117 9300 203
rect 9370 117 9400 203
rect 9470 117 9500 203
rect 9570 117 9600 203
rect 9670 117 9700 203
rect 9770 117 9800 203
rect 9870 117 9900 203
rect 9970 117 10000 203
rect 10070 117 10100 203
rect 10170 117 10200 203
rect 10270 117 10300 203
rect 10370 117 10400 203
rect 10470 117 10500 203
rect 10570 117 10600 203
rect 10670 117 10700 203
rect 10770 117 10800 203
rect 10870 117 10900 203
rect 10970 117 11000 203
rect 11070 117 11100 203
rect 11170 117 11200 203
rect 11270 117 11300 203
rect 11370 117 11400 203
rect 11570 257 11600 343
rect 11670 257 11700 343
rect 11770 257 11800 343
rect 11870 257 11900 343
rect 11970 257 12000 343
rect 12070 257 12100 343
rect 12170 257 12200 343
rect 12470 397 12500 483
rect 12570 397 12600 483
rect 12670 397 12700 483
rect 12770 397 12800 483
rect 12970 397 13000 483
rect 13070 397 13100 483
rect 13280 397 13310 483
rect 13380 397 13410 483
rect 13480 397 13510 483
rect 13580 397 13610 483
rect 12370 257 12400 343
rect 12470 257 12500 343
rect 12570 257 12600 343
rect 12670 257 12700 343
rect 12770 257 12800 343
rect 12970 257 13000 343
rect 13070 257 13100 343
rect 13280 257 13310 343
rect 13380 257 13410 343
rect 13480 257 13510 343
rect 13580 257 13610 343
rect 11570 117 11600 203
rect 11670 117 11700 203
rect 11770 117 11800 203
rect 11870 117 11900 203
rect 11970 117 12000 203
rect 12070 117 12100 203
rect 12170 117 12200 203
rect 12270 117 12300 203
rect 12370 117 12400 203
rect 12470 117 12500 203
rect 12570 117 12600 203
rect 12670 117 12700 203
rect 12770 117 12800 203
rect 12970 117 13000 203
rect 13070 117 13100 203
rect 13280 117 13310 203
rect 13380 117 13410 203
rect 13480 117 13510 203
rect 13580 117 13610 203
rect -10 -940 108 -910
rect 162 -940 280 -910
rect 390 -940 508 -910
rect 562 -940 680 -910
rect 790 -940 908 -910
rect 962 -940 1080 -910
rect 1190 -940 1308 -910
rect 1362 -940 1480 -910
rect -10 -1040 108 -1010
rect 162 -1040 280 -1010
rect 390 -1040 508 -1010
rect 562 -1040 680 -1010
rect 1590 -940 1708 -910
rect 1762 -940 1880 -910
rect 1990 -940 2108 -910
rect 2162 -940 2280 -910
rect 790 -1040 908 -1010
rect 962 -1040 1080 -1010
rect 1190 -1040 1308 -1010
rect 1362 -1040 1480 -1010
rect -10 -1140 108 -1110
rect 162 -1140 280 -1110
rect 390 -1140 508 -1110
rect 562 -1140 680 -1110
rect 2390 -940 2508 -910
rect 2562 -940 2680 -910
rect 2790 -940 2908 -910
rect 2962 -940 3080 -910
rect 1590 -1040 1708 -1010
rect 1762 -1040 1880 -1010
rect 1990 -1040 2108 -1010
rect 2162 -1040 2280 -1010
rect 790 -1140 908 -1110
rect 962 -1140 1080 -1110
rect 1190 -1140 1308 -1110
rect 1362 -1140 1480 -1110
rect -10 -1240 108 -1210
rect 162 -1240 280 -1210
rect 390 -1240 508 -1210
rect 562 -1240 680 -1210
rect 3190 -940 3308 -910
rect 3362 -940 3480 -910
rect 3590 -940 3708 -910
rect 3762 -940 3880 -910
rect 2390 -1040 2508 -1010
rect 2562 -1040 2680 -1010
rect 2790 -1040 2908 -1010
rect 2962 -1040 3080 -1010
rect 1590 -1140 1708 -1110
rect 1762 -1140 1880 -1110
rect 1990 -1140 2108 -1110
rect 2162 -1140 2280 -1110
rect 790 -1240 908 -1210
rect 962 -1240 1080 -1210
rect 1190 -1240 1308 -1210
rect 1362 -1240 1480 -1210
rect -10 -1340 108 -1310
rect 162 -1340 280 -1310
rect 390 -1340 508 -1310
rect 562 -1340 680 -1310
rect 3990 -940 4108 -910
rect 4162 -940 4280 -910
rect 4390 -940 4508 -910
rect 4562 -940 4680 -910
rect 3190 -1040 3308 -1010
rect 3362 -1040 3480 -1010
rect 3590 -1040 3708 -1010
rect 3762 -1040 3880 -1010
rect 2390 -1140 2508 -1110
rect 2562 -1140 2680 -1110
rect 2790 -1140 2908 -1110
rect 2962 -1140 3080 -1110
rect 1590 -1240 1708 -1210
rect 1762 -1240 1880 -1210
rect 1990 -1240 2108 -1210
rect 2162 -1240 2280 -1210
rect 790 -1340 908 -1310
rect 962 -1340 1080 -1310
rect 1190 -1340 1308 -1310
rect 1362 -1340 1480 -1310
rect -10 -1440 108 -1410
rect 162 -1440 280 -1410
rect 390 -1440 508 -1410
rect 562 -1440 680 -1410
rect 4790 -940 4908 -910
rect 4962 -940 5080 -910
rect 5190 -940 5308 -910
rect 5362 -940 5480 -910
rect 3990 -1040 4108 -1010
rect 4162 -1040 4280 -1010
rect 4390 -1040 4508 -1010
rect 4562 -1040 4680 -1010
rect 3190 -1140 3308 -1110
rect 3362 -1140 3480 -1110
rect 3590 -1140 3708 -1110
rect 3762 -1140 3880 -1110
rect 2390 -1240 2508 -1210
rect 2562 -1240 2680 -1210
rect 2790 -1240 2908 -1210
rect 2962 -1240 3080 -1210
rect 1590 -1340 1708 -1310
rect 1762 -1340 1880 -1310
rect 1990 -1340 2108 -1310
rect 2162 -1340 2280 -1310
rect 790 -1440 908 -1410
rect 962 -1440 1080 -1410
rect 1190 -1440 1308 -1410
rect 1362 -1440 1480 -1410
rect -10 -1540 108 -1510
rect 162 -1540 280 -1510
rect 390 -1540 508 -1510
rect 562 -1540 680 -1510
rect 5590 -940 5708 -910
rect 5762 -940 5880 -910
rect 5990 -940 6108 -910
rect 6162 -940 6280 -910
rect 4790 -1040 4908 -1010
rect 4962 -1040 5080 -1010
rect 5190 -1040 5308 -1010
rect 5362 -1040 5480 -1010
rect 3990 -1140 4108 -1110
rect 4162 -1140 4280 -1110
rect 4390 -1140 4508 -1110
rect 4562 -1140 4680 -1110
rect 3190 -1240 3308 -1210
rect 3362 -1240 3480 -1210
rect 3590 -1240 3708 -1210
rect 3762 -1240 3880 -1210
rect 2390 -1340 2508 -1310
rect 2562 -1340 2680 -1310
rect 2790 -1340 2908 -1310
rect 2962 -1340 3080 -1310
rect 1590 -1440 1708 -1410
rect 1762 -1440 1880 -1410
rect 1990 -1440 2108 -1410
rect 2162 -1440 2280 -1410
rect 790 -1540 908 -1510
rect 962 -1540 1080 -1510
rect 1190 -1540 1308 -1510
rect 1362 -1540 1480 -1510
rect -10 -1640 108 -1610
rect 162 -1640 280 -1610
rect 390 -1640 508 -1610
rect 562 -1640 680 -1610
rect 6390 -940 6508 -910
rect 6562 -940 6680 -910
rect 6790 -940 6908 -910
rect 6962 -940 7080 -910
rect 5590 -1040 5708 -1010
rect 5762 -1040 5880 -1010
rect 5990 -1040 6108 -1010
rect 6162 -1040 6280 -1010
rect 4790 -1140 4908 -1110
rect 4962 -1140 5080 -1110
rect 5190 -1140 5308 -1110
rect 5362 -1140 5480 -1110
rect 3990 -1240 4108 -1210
rect 4162 -1240 4280 -1210
rect 4390 -1240 4508 -1210
rect 4562 -1240 4680 -1210
rect 3190 -1340 3308 -1310
rect 3362 -1340 3480 -1310
rect 3590 -1340 3708 -1310
rect 3762 -1340 3880 -1310
rect 2390 -1440 2508 -1410
rect 2562 -1440 2680 -1410
rect 2790 -1440 2908 -1410
rect 2962 -1440 3080 -1410
rect 1590 -1540 1708 -1510
rect 1762 -1540 1880 -1510
rect 1990 -1540 2108 -1510
rect 2162 -1540 2280 -1510
rect 790 -1640 908 -1610
rect 962 -1640 1080 -1610
rect 1190 -1640 1308 -1610
rect 1362 -1640 1480 -1610
rect -10 -1740 108 -1710
rect 162 -1740 280 -1710
rect 390 -1740 508 -1710
rect 562 -1740 680 -1710
rect 7190 -940 7308 -910
rect 7362 -940 7480 -910
rect 7590 -940 7708 -910
rect 7762 -940 7880 -910
rect 6390 -1040 6508 -1010
rect 6562 -1040 6680 -1010
rect 6790 -1040 6908 -1010
rect 6962 -1040 7080 -1010
rect 5590 -1140 5708 -1110
rect 5762 -1140 5880 -1110
rect 5990 -1140 6108 -1110
rect 6162 -1140 6280 -1110
rect 4790 -1240 4908 -1210
rect 4962 -1240 5080 -1210
rect 5190 -1240 5308 -1210
rect 5362 -1240 5480 -1210
rect 3990 -1340 4108 -1310
rect 4162 -1340 4280 -1310
rect 4390 -1340 4508 -1310
rect 4562 -1340 4680 -1310
rect 3190 -1440 3308 -1410
rect 3362 -1440 3480 -1410
rect 3590 -1440 3708 -1410
rect 3762 -1440 3880 -1410
rect 2390 -1540 2508 -1510
rect 2562 -1540 2680 -1510
rect 2790 -1540 2908 -1510
rect 2962 -1540 3080 -1510
rect 1590 -1640 1708 -1610
rect 1762 -1640 1880 -1610
rect 1990 -1640 2108 -1610
rect 2162 -1640 2280 -1610
rect 790 -1740 908 -1710
rect 962 -1740 1080 -1710
rect 1190 -1740 1308 -1710
rect 1362 -1740 1480 -1710
rect -10 -1840 108 -1810
rect 162 -1840 280 -1810
rect 390 -1840 508 -1810
rect 562 -1840 680 -1810
rect 7990 -940 8108 -910
rect 8162 -940 8280 -910
rect 8390 -940 8508 -910
rect 8562 -940 8680 -910
rect 7190 -1040 7308 -1010
rect 7362 -1040 7480 -1010
rect 7590 -1040 7708 -1010
rect 7762 -1040 7880 -1010
rect 6390 -1140 6508 -1110
rect 6562 -1140 6680 -1110
rect 6790 -1140 6908 -1110
rect 6962 -1140 7080 -1110
rect 5590 -1240 5708 -1210
rect 5762 -1240 5880 -1210
rect 5990 -1240 6108 -1210
rect 6162 -1240 6280 -1210
rect 4790 -1340 4908 -1310
rect 4962 -1340 5080 -1310
rect 5190 -1340 5308 -1310
rect 5362 -1340 5480 -1310
rect 3990 -1440 4108 -1410
rect 4162 -1440 4280 -1410
rect 4390 -1440 4508 -1410
rect 4562 -1440 4680 -1410
rect 3190 -1540 3308 -1510
rect 3362 -1540 3480 -1510
rect 3590 -1540 3708 -1510
rect 3762 -1540 3880 -1510
rect 2390 -1640 2508 -1610
rect 2562 -1640 2680 -1610
rect 2790 -1640 2908 -1610
rect 2962 -1640 3080 -1610
rect 1590 -1740 1708 -1710
rect 1762 -1740 1880 -1710
rect 1990 -1740 2108 -1710
rect 2162 -1740 2280 -1710
rect 790 -1840 908 -1810
rect 962 -1840 1080 -1810
rect 1190 -1840 1308 -1810
rect 1362 -1840 1480 -1810
rect -10 -1940 108 -1910
rect 162 -1940 280 -1910
rect 390 -1940 508 -1910
rect 562 -1940 680 -1910
rect 8790 -940 8908 -910
rect 8962 -940 9080 -910
rect 9190 -940 9308 -910
rect 9362 -940 9480 -910
rect 7990 -1040 8108 -1010
rect 8162 -1040 8280 -1010
rect 8390 -1040 8508 -1010
rect 8562 -1040 8680 -1010
rect 7190 -1140 7308 -1110
rect 7362 -1140 7480 -1110
rect 7590 -1140 7708 -1110
rect 7762 -1140 7880 -1110
rect 6390 -1240 6508 -1210
rect 6562 -1240 6680 -1210
rect 6790 -1240 6908 -1210
rect 6962 -1240 7080 -1210
rect 5590 -1340 5708 -1310
rect 5762 -1340 5880 -1310
rect 5990 -1340 6108 -1310
rect 6162 -1340 6280 -1310
rect 4790 -1440 4908 -1410
rect 4962 -1440 5080 -1410
rect 5190 -1440 5308 -1410
rect 5362 -1440 5480 -1410
rect 3990 -1540 4108 -1510
rect 4162 -1540 4280 -1510
rect 4390 -1540 4508 -1510
rect 4562 -1540 4680 -1510
rect 3190 -1640 3308 -1610
rect 3362 -1640 3480 -1610
rect 3590 -1640 3708 -1610
rect 3762 -1640 3880 -1610
rect 2390 -1740 2508 -1710
rect 2562 -1740 2680 -1710
rect 2790 -1740 2908 -1710
rect 2962 -1740 3080 -1710
rect 1590 -1840 1708 -1810
rect 1762 -1840 1880 -1810
rect 1990 -1840 2108 -1810
rect 2162 -1840 2280 -1810
rect 790 -1940 908 -1910
rect 962 -1940 1080 -1910
rect 1190 -1940 1308 -1910
rect 1362 -1940 1480 -1910
rect -10 -2040 108 -2010
rect 162 -2040 280 -2010
rect 390 -2040 508 -2010
rect 562 -2040 680 -2010
rect 9590 -940 9708 -910
rect 9762 -940 9880 -910
rect 9990 -940 10108 -910
rect 10162 -940 10280 -910
rect 8790 -1040 8908 -1010
rect 8962 -1040 9080 -1010
rect 9190 -1040 9308 -1010
rect 9362 -1040 9480 -1010
rect 7990 -1140 8108 -1110
rect 8162 -1140 8280 -1110
rect 8390 -1140 8508 -1110
rect 8562 -1140 8680 -1110
rect 7190 -1240 7308 -1210
rect 7362 -1240 7480 -1210
rect 7590 -1240 7708 -1210
rect 7762 -1240 7880 -1210
rect 6390 -1340 6508 -1310
rect 6562 -1340 6680 -1310
rect 6790 -1340 6908 -1310
rect 6962 -1340 7080 -1310
rect 5590 -1440 5708 -1410
rect 5762 -1440 5880 -1410
rect 5990 -1440 6108 -1410
rect 6162 -1440 6280 -1410
rect 4790 -1540 4908 -1510
rect 4962 -1540 5080 -1510
rect 5190 -1540 5308 -1510
rect 5362 -1540 5480 -1510
rect 3990 -1640 4108 -1610
rect 4162 -1640 4280 -1610
rect 4390 -1640 4508 -1610
rect 4562 -1640 4680 -1610
rect 3190 -1740 3308 -1710
rect 3362 -1740 3480 -1710
rect 3590 -1740 3708 -1710
rect 3762 -1740 3880 -1710
rect 2390 -1840 2508 -1810
rect 2562 -1840 2680 -1810
rect 2790 -1840 2908 -1810
rect 2962 -1840 3080 -1810
rect 1590 -1940 1708 -1910
rect 1762 -1940 1880 -1910
rect 1990 -1940 2108 -1910
rect 2162 -1940 2280 -1910
rect 790 -2040 908 -2010
rect 962 -2040 1080 -2010
rect 1190 -2040 1308 -2010
rect 1362 -2040 1480 -2010
rect 10390 -940 10508 -910
rect 10562 -940 10680 -910
rect 10790 -940 10908 -910
rect 10962 -940 11080 -910
rect 9590 -1040 9708 -1010
rect 9762 -1040 9880 -1010
rect 9990 -1040 10108 -1010
rect 10162 -1040 10280 -1010
rect 8790 -1140 8908 -1110
rect 8962 -1140 9080 -1110
rect 9190 -1140 9308 -1110
rect 9362 -1140 9480 -1110
rect 7990 -1240 8108 -1210
rect 8162 -1240 8280 -1210
rect 8390 -1240 8508 -1210
rect 8562 -1240 8680 -1210
rect 7190 -1340 7308 -1310
rect 7362 -1340 7480 -1310
rect 7590 -1340 7708 -1310
rect 7762 -1340 7880 -1310
rect 6390 -1440 6508 -1410
rect 6562 -1440 6680 -1410
rect 6790 -1440 6908 -1410
rect 6962 -1440 7080 -1410
rect 5590 -1540 5708 -1510
rect 5762 -1540 5880 -1510
rect 5990 -1540 6108 -1510
rect 6162 -1540 6280 -1510
rect 4790 -1640 4908 -1610
rect 4962 -1640 5080 -1610
rect 5190 -1640 5308 -1610
rect 5362 -1640 5480 -1610
rect 3990 -1740 4108 -1710
rect 4162 -1740 4280 -1710
rect 4390 -1740 4508 -1710
rect 4562 -1740 4680 -1710
rect 3190 -1840 3308 -1810
rect 3362 -1840 3480 -1810
rect 3590 -1840 3708 -1810
rect 3762 -1840 3880 -1810
rect 2390 -1940 2508 -1910
rect 2562 -1940 2680 -1910
rect 2790 -1940 2908 -1910
rect 2962 -1940 3080 -1910
rect 1590 -2040 1708 -2010
rect 1762 -2040 1880 -2010
rect 1990 -2040 2108 -2010
rect 2162 -2040 2280 -2010
rect 11190 -940 11308 -910
rect 11362 -940 11480 -910
rect 11590 -940 11708 -910
rect 11762 -940 11880 -910
rect 10390 -1040 10508 -1010
rect 10562 -1040 10680 -1010
rect 10790 -1040 10908 -1010
rect 10962 -1040 11080 -1010
rect 9590 -1140 9708 -1110
rect 9762 -1140 9880 -1110
rect 9990 -1140 10108 -1110
rect 10162 -1140 10280 -1110
rect 8790 -1240 8908 -1210
rect 8962 -1240 9080 -1210
rect 9190 -1240 9308 -1210
rect 9362 -1240 9480 -1210
rect 7990 -1340 8108 -1310
rect 8162 -1340 8280 -1310
rect 8390 -1340 8508 -1310
rect 8562 -1340 8680 -1310
rect 7190 -1440 7308 -1410
rect 7362 -1440 7480 -1410
rect 7590 -1440 7708 -1410
rect 7762 -1440 7880 -1410
rect 6390 -1540 6508 -1510
rect 6562 -1540 6680 -1510
rect 6790 -1540 6908 -1510
rect 6962 -1540 7080 -1510
rect 5590 -1640 5708 -1610
rect 5762 -1640 5880 -1610
rect 5990 -1640 6108 -1610
rect 6162 -1640 6280 -1610
rect 4790 -1740 4908 -1710
rect 4962 -1740 5080 -1710
rect 5190 -1740 5308 -1710
rect 5362 -1740 5480 -1710
rect 3990 -1840 4108 -1810
rect 4162 -1840 4280 -1810
rect 4390 -1840 4508 -1810
rect 4562 -1840 4680 -1810
rect 3190 -1940 3308 -1910
rect 3362 -1940 3480 -1910
rect 3590 -1940 3708 -1910
rect 3762 -1940 3880 -1910
rect 2390 -2040 2508 -2010
rect 2562 -2040 2680 -2010
rect 2790 -2040 2908 -2010
rect 2962 -2040 3080 -2010
rect 11990 -940 12108 -910
rect 12162 -940 12280 -910
rect 12390 -940 12508 -910
rect 12562 -940 12680 -910
rect 11190 -1040 11308 -1010
rect 11362 -1040 11480 -1010
rect 11590 -1040 11708 -1010
rect 11762 -1040 11880 -1010
rect 10390 -1140 10508 -1110
rect 10562 -1140 10680 -1110
rect 10790 -1140 10908 -1110
rect 10962 -1140 11080 -1110
rect 9590 -1240 9708 -1210
rect 9762 -1240 9880 -1210
rect 9990 -1240 10108 -1210
rect 10162 -1240 10280 -1210
rect 8790 -1340 8908 -1310
rect 8962 -1340 9080 -1310
rect 9190 -1340 9308 -1310
rect 9362 -1340 9480 -1310
rect 7990 -1440 8108 -1410
rect 8162 -1440 8280 -1410
rect 8390 -1440 8508 -1410
rect 8562 -1440 8680 -1410
rect 7190 -1540 7308 -1510
rect 7362 -1540 7480 -1510
rect 7590 -1540 7708 -1510
rect 7762 -1540 7880 -1510
rect 6390 -1640 6508 -1610
rect 6562 -1640 6680 -1610
rect 6790 -1640 6908 -1610
rect 6962 -1640 7080 -1610
rect 5590 -1740 5708 -1710
rect 5762 -1740 5880 -1710
rect 5990 -1740 6108 -1710
rect 6162 -1740 6280 -1710
rect 4790 -1840 4908 -1810
rect 4962 -1840 5080 -1810
rect 5190 -1840 5308 -1810
rect 5362 -1840 5480 -1810
rect 3990 -1940 4108 -1910
rect 4162 -1940 4280 -1910
rect 4390 -1940 4508 -1910
rect 4562 -1940 4680 -1910
rect 3190 -2040 3308 -2010
rect 3362 -2040 3480 -2010
rect 3590 -2040 3708 -2010
rect 3762 -2040 3880 -2010
rect 11990 -1040 12108 -1010
rect 12162 -1040 12280 -1010
rect 12390 -1040 12508 -1010
rect 12562 -1040 12680 -1010
rect 11190 -1140 11308 -1110
rect 11362 -1140 11480 -1110
rect 11590 -1140 11708 -1110
rect 11762 -1140 11880 -1110
rect 10390 -1240 10508 -1210
rect 10562 -1240 10680 -1210
rect 10790 -1240 10908 -1210
rect 10962 -1240 11080 -1210
rect 9590 -1340 9708 -1310
rect 9762 -1340 9880 -1310
rect 9990 -1340 10108 -1310
rect 10162 -1340 10280 -1310
rect 8790 -1440 8908 -1410
rect 8962 -1440 9080 -1410
rect 9190 -1440 9308 -1410
rect 9362 -1440 9480 -1410
rect 7990 -1540 8108 -1510
rect 8162 -1540 8280 -1510
rect 8390 -1540 8508 -1510
rect 8562 -1540 8680 -1510
rect 7190 -1640 7308 -1610
rect 7362 -1640 7480 -1610
rect 7590 -1640 7708 -1610
rect 7762 -1640 7880 -1610
rect 6390 -1740 6508 -1710
rect 6562 -1740 6680 -1710
rect 6790 -1740 6908 -1710
rect 6962 -1740 7080 -1710
rect 5590 -1840 5708 -1810
rect 5762 -1840 5880 -1810
rect 5990 -1840 6108 -1810
rect 6162 -1840 6280 -1810
rect 4790 -1940 4908 -1910
rect 4962 -1940 5080 -1910
rect 5190 -1940 5308 -1910
rect 5362 -1940 5480 -1910
rect 3990 -2040 4108 -2010
rect 4162 -2040 4280 -2010
rect 4390 -2040 4508 -2010
rect 4562 -2040 4680 -2010
rect 11990 -1140 12108 -1110
rect 12162 -1140 12280 -1110
rect 12390 -1140 12508 -1110
rect 12562 -1140 12680 -1110
rect 11190 -1240 11308 -1210
rect 11362 -1240 11480 -1210
rect 11590 -1240 11708 -1210
rect 11762 -1240 11880 -1210
rect 10390 -1340 10508 -1310
rect 10562 -1340 10680 -1310
rect 10790 -1340 10908 -1310
rect 10962 -1340 11080 -1310
rect 9590 -1440 9708 -1410
rect 9762 -1440 9880 -1410
rect 9990 -1440 10108 -1410
rect 10162 -1440 10280 -1410
rect 8790 -1540 8908 -1510
rect 8962 -1540 9080 -1510
rect 9190 -1540 9308 -1510
rect 9362 -1540 9480 -1510
rect 7990 -1640 8108 -1610
rect 8162 -1640 8280 -1610
rect 8390 -1640 8508 -1610
rect 8562 -1640 8680 -1610
rect 7190 -1740 7308 -1710
rect 7362 -1740 7480 -1710
rect 7590 -1740 7708 -1710
rect 7762 -1740 7880 -1710
rect 6390 -1840 6508 -1810
rect 6562 -1840 6680 -1810
rect 6790 -1840 6908 -1810
rect 6962 -1840 7080 -1810
rect 5590 -1940 5708 -1910
rect 5762 -1940 5880 -1910
rect 5990 -1940 6108 -1910
rect 6162 -1940 6280 -1910
rect 4790 -2040 4908 -2010
rect 4962 -2040 5080 -2010
rect 5190 -2040 5308 -2010
rect 5362 -2040 5480 -2010
rect 11990 -1240 12108 -1210
rect 12162 -1240 12280 -1210
rect 12390 -1240 12508 -1210
rect 12562 -1240 12680 -1210
rect 11190 -1340 11308 -1310
rect 11362 -1340 11480 -1310
rect 11590 -1340 11708 -1310
rect 11762 -1340 11880 -1310
rect 10390 -1440 10508 -1410
rect 10562 -1440 10680 -1410
rect 10790 -1440 10908 -1410
rect 10962 -1440 11080 -1410
rect 9590 -1540 9708 -1510
rect 9762 -1540 9880 -1510
rect 9990 -1540 10108 -1510
rect 10162 -1540 10280 -1510
rect 8790 -1640 8908 -1610
rect 8962 -1640 9080 -1610
rect 9190 -1640 9308 -1610
rect 9362 -1640 9480 -1610
rect 7990 -1740 8108 -1710
rect 8162 -1740 8280 -1710
rect 8390 -1740 8508 -1710
rect 8562 -1740 8680 -1710
rect 7190 -1840 7308 -1810
rect 7362 -1840 7480 -1810
rect 7590 -1840 7708 -1810
rect 7762 -1840 7880 -1810
rect 6390 -1940 6508 -1910
rect 6562 -1940 6680 -1910
rect 6790 -1940 6908 -1910
rect 6962 -1940 7080 -1910
rect 5590 -2040 5708 -2010
rect 5762 -2040 5880 -2010
rect 5990 -2040 6108 -2010
rect 6162 -2040 6280 -2010
rect 11990 -1340 12108 -1310
rect 12162 -1340 12280 -1310
rect 12390 -1340 12508 -1310
rect 12562 -1340 12680 -1310
rect 11190 -1440 11308 -1410
rect 11362 -1440 11480 -1410
rect 11590 -1440 11708 -1410
rect 11762 -1440 11880 -1410
rect 10390 -1540 10508 -1510
rect 10562 -1540 10680 -1510
rect 10790 -1540 10908 -1510
rect 10962 -1540 11080 -1510
rect 9590 -1640 9708 -1610
rect 9762 -1640 9880 -1610
rect 9990 -1640 10108 -1610
rect 10162 -1640 10280 -1610
rect 8790 -1740 8908 -1710
rect 8962 -1740 9080 -1710
rect 9190 -1740 9308 -1710
rect 9362 -1740 9480 -1710
rect 7990 -1840 8108 -1810
rect 8162 -1840 8280 -1810
rect 8390 -1840 8508 -1810
rect 8562 -1840 8680 -1810
rect 7190 -1940 7308 -1910
rect 7362 -1940 7480 -1910
rect 7590 -1940 7708 -1910
rect 7762 -1940 7880 -1910
rect 6390 -2040 6508 -2010
rect 6562 -2040 6680 -2010
rect 6790 -2040 6908 -2010
rect 6962 -2040 7080 -2010
rect 11990 -1440 12108 -1410
rect 12162 -1440 12280 -1410
rect 12390 -1440 12508 -1410
rect 12562 -1440 12680 -1410
rect 11190 -1540 11308 -1510
rect 11362 -1540 11480 -1510
rect 11590 -1540 11708 -1510
rect 11762 -1540 11880 -1510
rect 10390 -1640 10508 -1610
rect 10562 -1640 10680 -1610
rect 10790 -1640 10908 -1610
rect 10962 -1640 11080 -1610
rect 9590 -1740 9708 -1710
rect 9762 -1740 9880 -1710
rect 9990 -1740 10108 -1710
rect 10162 -1740 10280 -1710
rect 8790 -1840 8908 -1810
rect 8962 -1840 9080 -1810
rect 9190 -1840 9308 -1810
rect 9362 -1840 9480 -1810
rect 7990 -1940 8108 -1910
rect 8162 -1940 8280 -1910
rect 8390 -1940 8508 -1910
rect 8562 -1940 8680 -1910
rect 7190 -2040 7308 -2010
rect 7362 -2040 7480 -2010
rect 7590 -2040 7708 -2010
rect 7762 -2040 7880 -2010
rect 11990 -1540 12108 -1510
rect 12162 -1540 12280 -1510
rect 12390 -1540 12508 -1510
rect 12562 -1540 12680 -1510
rect 11190 -1640 11308 -1610
rect 11362 -1640 11480 -1610
rect 11590 -1640 11708 -1610
rect 11762 -1640 11880 -1610
rect 10390 -1740 10508 -1710
rect 10562 -1740 10680 -1710
rect 10790 -1740 10908 -1710
rect 10962 -1740 11080 -1710
rect 9590 -1840 9708 -1810
rect 9762 -1840 9880 -1810
rect 9990 -1840 10108 -1810
rect 10162 -1840 10280 -1810
rect 8790 -1940 8908 -1910
rect 8962 -1940 9080 -1910
rect 9190 -1940 9308 -1910
rect 9362 -1940 9480 -1910
rect 7990 -2040 8108 -2010
rect 8162 -2040 8280 -2010
rect 8390 -2040 8508 -2010
rect 8562 -2040 8680 -2010
rect 11990 -1640 12108 -1610
rect 12162 -1640 12280 -1610
rect 12390 -1640 12508 -1610
rect 12562 -1640 12680 -1610
rect 11190 -1740 11308 -1710
rect 11362 -1740 11480 -1710
rect 11590 -1740 11708 -1710
rect 11762 -1740 11880 -1710
rect 10390 -1840 10508 -1810
rect 10562 -1840 10680 -1810
rect 10790 -1840 10908 -1810
rect 10962 -1840 11080 -1810
rect 9590 -1940 9708 -1910
rect 9762 -1940 9880 -1910
rect 9990 -1940 10108 -1910
rect 10162 -1940 10280 -1910
rect 8790 -2040 8908 -2010
rect 8962 -2040 9080 -2010
rect 9190 -2040 9308 -2010
rect 9362 -2040 9480 -2010
rect 11990 -1740 12108 -1710
rect 12162 -1740 12280 -1710
rect 12390 -1740 12508 -1710
rect 12562 -1740 12680 -1710
rect 11190 -1840 11308 -1810
rect 11362 -1840 11480 -1810
rect 11590 -1840 11708 -1810
rect 11762 -1840 11880 -1810
rect 10390 -1940 10508 -1910
rect 10562 -1940 10680 -1910
rect 10790 -1940 10908 -1910
rect 10962 -1940 11080 -1910
rect 9590 -2040 9708 -2010
rect 9762 -2040 9880 -2010
rect 9990 -2040 10108 -2010
rect 10162 -2040 10280 -2010
rect 11990 -1840 12108 -1810
rect 12162 -1840 12280 -1810
rect 12390 -1840 12508 -1810
rect 12562 -1840 12680 -1810
rect 11190 -1940 11308 -1910
rect 11362 -1940 11480 -1910
rect 11590 -1940 11708 -1910
rect 11762 -1940 11880 -1910
rect 10390 -2040 10508 -2010
rect 10562 -2040 10680 -2010
rect 10790 -2040 10908 -2010
rect 10962 -2040 11080 -2010
rect 11990 -1940 12108 -1910
rect 12162 -1940 12280 -1910
rect 12390 -1940 12508 -1910
rect 12562 -1940 12680 -1910
rect 11190 -2040 11308 -2010
rect 11362 -2040 11480 -2010
rect 11590 -2040 11708 -2010
rect 11762 -2040 11880 -2010
rect 11990 -2040 12108 -2010
rect 12162 -2040 12280 -2010
rect 12390 -2040 12508 -2010
rect 12562 -2040 12680 -2010
<< ndiff >>
rect 16 4787 70 4813
rect 16 4753 24 4787
rect 58 4753 70 4787
rect 16 4727 70 4753
rect 100 4787 170 4813
rect 100 4753 118 4787
rect 152 4753 170 4787
rect 100 4727 170 4753
rect 200 4787 270 4813
rect 200 4753 218 4787
rect 252 4753 270 4787
rect 200 4727 270 4753
rect 300 4787 354 4813
rect 300 4753 312 4787
rect 346 4753 354 4787
rect 300 4727 354 4753
rect 416 4787 470 4813
rect 416 4753 424 4787
rect 458 4753 470 4787
rect 416 4727 470 4753
rect 500 4787 570 4813
rect 500 4753 518 4787
rect 552 4753 570 4787
rect 500 4727 570 4753
rect 600 4787 670 4813
rect 600 4753 618 4787
rect 652 4753 670 4787
rect 600 4727 670 4753
rect 700 4727 770 4813
rect 800 4727 870 4813
rect 900 4727 970 4813
rect 1000 4787 1070 4813
rect 1000 4753 1018 4787
rect 1052 4753 1070 4787
rect 1000 4727 1070 4753
rect 1100 4787 1154 4813
rect 1100 4753 1112 4787
rect 1146 4753 1154 4787
rect 1100 4727 1154 4753
rect 16 4587 70 4673
rect 100 4647 170 4673
rect 100 4613 118 4647
rect 152 4613 170 4647
rect 100 4587 170 4613
rect 200 4647 270 4673
rect 200 4613 218 4647
rect 252 4613 270 4647
rect 200 4587 270 4613
rect 300 4587 370 4673
rect 400 4587 470 4673
rect 500 4587 570 4673
rect 600 4647 670 4673
rect 600 4613 618 4647
rect 652 4613 670 4647
rect 600 4587 670 4613
rect 700 4647 770 4673
rect 700 4613 718 4647
rect 752 4613 770 4647
rect 700 4587 770 4613
rect 800 4587 870 4673
rect 900 4647 970 4673
rect 900 4613 918 4647
rect 952 4613 970 4647
rect 900 4587 970 4613
rect 1000 4647 1070 4673
rect 1000 4613 1018 4647
rect 1052 4613 1070 4647
rect 1000 4587 1070 4613
rect 1100 4647 1154 4673
rect 1100 4613 1112 4647
rect 1146 4613 1154 4647
rect 1100 4587 1154 4613
rect 16 4447 70 4533
rect 100 4447 170 4533
rect 200 4507 270 4533
rect 200 4473 218 4507
rect 252 4473 270 4507
rect 200 4447 270 4473
rect 300 4507 354 4533
rect 300 4473 312 4507
rect 346 4473 354 4507
rect 300 4447 354 4473
rect 1216 4787 1270 4813
rect 1216 4753 1224 4787
rect 1258 4753 1270 4787
rect 1216 4727 1270 4753
rect 1300 4787 1370 4813
rect 1300 4753 1318 4787
rect 1352 4753 1370 4787
rect 1300 4727 1370 4753
rect 1400 4787 1470 4813
rect 1400 4753 1418 4787
rect 1452 4753 1470 4787
rect 1400 4727 1470 4753
rect 1500 4727 1570 4813
rect 1600 4787 1670 4813
rect 1600 4753 1618 4787
rect 1652 4753 1670 4787
rect 1600 4727 1670 4753
rect 1700 4787 1770 4813
rect 1700 4753 1718 4787
rect 1752 4753 1770 4787
rect 1700 4727 1770 4753
rect 1800 4787 1870 4813
rect 1800 4753 1818 4787
rect 1852 4753 1870 4787
rect 1800 4727 1870 4753
rect 1900 4787 1970 4813
rect 1900 4753 1918 4787
rect 1952 4753 1970 4787
rect 1900 4727 1970 4753
rect 2000 4727 2070 4813
rect 2100 4727 2170 4813
rect 2200 4787 2270 4813
rect 2200 4753 2218 4787
rect 2252 4753 2270 4787
rect 2200 4727 2270 4753
rect 2300 4787 2354 4813
rect 2300 4753 2312 4787
rect 2346 4753 2354 4787
rect 2300 4727 2354 4753
rect 2416 4787 2470 4813
rect 2416 4753 2424 4787
rect 2458 4753 2470 4787
rect 2416 4727 2470 4753
rect 2500 4787 2570 4813
rect 2500 4753 2518 4787
rect 2552 4753 2570 4787
rect 2500 4727 2570 4753
rect 2600 4787 2670 4813
rect 2600 4753 2618 4787
rect 2652 4753 2670 4787
rect 2600 4727 2670 4753
rect 2700 4727 2770 4813
rect 2800 4727 2870 4813
rect 2900 4787 2970 4813
rect 2900 4753 2918 4787
rect 2952 4753 2970 4787
rect 2900 4727 2970 4753
rect 3000 4787 3070 4813
rect 3000 4753 3018 4787
rect 3052 4753 3070 4787
rect 3000 4727 3070 4753
rect 3100 4787 3154 4813
rect 3100 4753 3112 4787
rect 3146 4753 3154 4787
rect 3100 4727 3154 4753
rect 1216 4647 1270 4673
rect 1216 4613 1224 4647
rect 1258 4613 1270 4647
rect 1216 4587 1270 4613
rect 1300 4647 1370 4673
rect 1300 4613 1318 4647
rect 1352 4613 1370 4647
rect 1300 4587 1370 4613
rect 1400 4587 1470 4673
rect 1500 4647 1570 4673
rect 1500 4613 1518 4647
rect 1552 4613 1570 4647
rect 1500 4587 1570 4613
rect 1600 4647 1670 4673
rect 1600 4613 1618 4647
rect 1652 4613 1670 4647
rect 1600 4587 1670 4613
rect 1700 4647 1770 4673
rect 1700 4613 1718 4647
rect 1752 4613 1770 4647
rect 1700 4587 1770 4613
rect 1800 4587 1870 4673
rect 1900 4587 1970 4673
rect 2000 4647 2070 4673
rect 2000 4613 2018 4647
rect 2052 4613 2070 4647
rect 2000 4587 2070 4613
rect 2100 4647 2170 4673
rect 2100 4613 2118 4647
rect 2152 4613 2170 4647
rect 2100 4587 2170 4613
rect 2200 4587 2270 4673
rect 2300 4587 2370 4673
rect 2400 4587 2470 4673
rect 2500 4587 2570 4673
rect 2600 4647 2670 4673
rect 2600 4613 2618 4647
rect 2652 4613 2670 4647
rect 2600 4587 2670 4613
rect 2700 4647 2770 4673
rect 2700 4613 2718 4647
rect 2752 4613 2770 4647
rect 2700 4587 2770 4613
rect 2800 4647 2870 4673
rect 2800 4613 2818 4647
rect 2852 4613 2870 4647
rect 2800 4587 2870 4613
rect 2900 4647 2954 4673
rect 2900 4613 2912 4647
rect 2946 4613 2954 4647
rect 2900 4587 2954 4613
rect 416 4507 470 4533
rect 416 4473 424 4507
rect 458 4473 470 4507
rect 416 4447 470 4473
rect 500 4507 570 4533
rect 500 4473 518 4507
rect 552 4473 570 4507
rect 500 4447 570 4473
rect 600 4507 670 4533
rect 600 4473 618 4507
rect 652 4473 670 4507
rect 600 4447 670 4473
rect 700 4507 770 4533
rect 700 4473 718 4507
rect 752 4473 770 4507
rect 700 4447 770 4473
rect 800 4507 870 4533
rect 800 4473 818 4507
rect 852 4473 870 4507
rect 800 4447 870 4473
rect 900 4447 970 4533
rect 1000 4507 1070 4533
rect 1000 4473 1018 4507
rect 1052 4473 1070 4507
rect 1000 4447 1070 4473
rect 1100 4507 1170 4533
rect 1100 4473 1118 4507
rect 1152 4473 1170 4507
rect 1100 4447 1170 4473
rect 1200 4447 1270 4533
rect 1300 4447 1370 4533
rect 1400 4507 1470 4533
rect 1400 4473 1418 4507
rect 1452 4473 1470 4507
rect 1400 4447 1470 4473
rect 1500 4507 1570 4533
rect 1500 4473 1518 4507
rect 1552 4473 1570 4507
rect 1500 4447 1570 4473
rect 1600 4507 1654 4533
rect 1600 4473 1612 4507
rect 1646 4473 1654 4507
rect 1600 4447 1654 4473
rect 16 4367 70 4393
rect 16 4333 24 4367
rect 58 4333 70 4367
rect 16 4307 70 4333
rect 100 4367 170 4393
rect 100 4333 118 4367
rect 152 4333 170 4367
rect 100 4307 170 4333
rect 200 4367 270 4393
rect 200 4333 218 4367
rect 252 4333 270 4367
rect 200 4307 270 4333
rect 300 4307 370 4393
rect 400 4367 470 4393
rect 400 4333 418 4367
rect 452 4333 470 4367
rect 400 4307 470 4333
rect 500 4367 570 4393
rect 500 4333 518 4367
rect 552 4333 570 4367
rect 500 4307 570 4333
rect 600 4307 670 4393
rect 700 4307 770 4393
rect 800 4307 870 4393
rect 900 4307 970 4393
rect 1000 4367 1070 4393
rect 1000 4333 1018 4367
rect 1052 4333 1070 4367
rect 1000 4307 1070 4333
rect 1100 4367 1170 4393
rect 1100 4333 1118 4367
rect 1152 4333 1170 4367
rect 1100 4307 1170 4333
rect 1200 4367 1254 4393
rect 1200 4333 1212 4367
rect 1246 4333 1254 4367
rect 1200 4307 1254 4333
rect 16 4167 70 4253
rect 100 4227 170 4253
rect 100 4193 118 4227
rect 152 4193 170 4227
rect 100 4167 170 4193
rect 200 4227 270 4253
rect 200 4193 218 4227
rect 252 4193 270 4227
rect 200 4167 270 4193
rect 300 4167 370 4253
rect 400 4227 470 4253
rect 400 4193 418 4227
rect 452 4193 470 4227
rect 400 4167 470 4193
rect 500 4227 554 4253
rect 500 4193 512 4227
rect 546 4193 554 4227
rect 500 4167 554 4193
rect 16 4087 70 4113
rect 16 4053 24 4087
rect 58 4053 70 4087
rect 16 4027 70 4053
rect 100 4087 170 4113
rect 100 4053 118 4087
rect 152 4053 170 4087
rect 100 4027 170 4053
rect 200 4087 254 4113
rect 200 4053 212 4087
rect 246 4053 254 4087
rect 200 4027 254 4053
rect 316 4087 370 4113
rect 316 4053 324 4087
rect 358 4053 370 4087
rect 316 4027 370 4053
rect 400 4087 454 4113
rect 400 4053 412 4087
rect 446 4053 454 4087
rect 400 4027 454 4053
rect 616 4227 670 4253
rect 616 4193 624 4227
rect 658 4193 670 4227
rect 616 4167 670 4193
rect 700 4227 770 4253
rect 700 4193 718 4227
rect 752 4193 770 4227
rect 700 4167 770 4193
rect 800 4167 870 4253
rect 900 4167 970 4253
rect 1000 4227 1070 4253
rect 1000 4193 1018 4227
rect 1052 4193 1070 4227
rect 1000 4167 1070 4193
rect 1100 4227 1154 4253
rect 1100 4193 1112 4227
rect 1146 4193 1154 4227
rect 1100 4167 1154 4193
rect 1716 4507 1770 4533
rect 1716 4473 1724 4507
rect 1758 4473 1770 4507
rect 1716 4447 1770 4473
rect 1800 4507 1854 4533
rect 1800 4473 1812 4507
rect 1846 4473 1854 4507
rect 1800 4447 1854 4473
rect 1916 4507 1970 4533
rect 1916 4473 1924 4507
rect 1958 4473 1970 4507
rect 1916 4447 1970 4473
rect 2000 4507 2070 4533
rect 2000 4473 2018 4507
rect 2052 4473 2070 4507
rect 2000 4447 2070 4473
rect 2100 4507 2170 4533
rect 2100 4473 2118 4507
rect 2152 4473 2170 4507
rect 2100 4447 2170 4473
rect 2200 4507 2270 4533
rect 2200 4473 2218 4507
rect 2252 4473 2270 4507
rect 2200 4447 2270 4473
rect 2300 4507 2354 4533
rect 2300 4473 2312 4507
rect 2346 4473 2354 4507
rect 2300 4447 2354 4473
rect 1316 4367 1370 4393
rect 1316 4333 1324 4367
rect 1358 4333 1370 4367
rect 1316 4307 1370 4333
rect 1400 4367 1470 4393
rect 1400 4333 1418 4367
rect 1452 4333 1470 4367
rect 1400 4307 1470 4333
rect 1500 4367 1570 4393
rect 1500 4333 1518 4367
rect 1552 4333 1570 4367
rect 1500 4307 1570 4333
rect 1600 4307 1670 4393
rect 1700 4367 1770 4393
rect 1700 4333 1718 4367
rect 1752 4333 1770 4367
rect 1700 4307 1770 4333
rect 1800 4367 1870 4393
rect 1800 4333 1818 4367
rect 1852 4333 1870 4367
rect 1800 4307 1870 4333
rect 1900 4367 1954 4393
rect 1900 4333 1912 4367
rect 1946 4333 1954 4367
rect 1900 4307 1954 4333
rect 1216 4227 1270 4253
rect 1216 4193 1224 4227
rect 1258 4193 1270 4227
rect 1216 4167 1270 4193
rect 1300 4227 1370 4253
rect 1300 4193 1318 4227
rect 1352 4193 1370 4227
rect 1300 4167 1370 4193
rect 1400 4227 1470 4253
rect 1400 4193 1418 4227
rect 1452 4193 1470 4227
rect 1400 4167 1470 4193
rect 1500 4227 1570 4253
rect 1500 4193 1518 4227
rect 1552 4193 1570 4227
rect 1500 4167 1570 4193
rect 1600 4227 1670 4253
rect 1600 4193 1618 4227
rect 1652 4193 1670 4227
rect 1600 4167 1670 4193
rect 1700 4227 1770 4253
rect 1700 4193 1718 4227
rect 1752 4193 1770 4227
rect 1700 4167 1770 4193
rect 1800 4227 1870 4253
rect 1800 4193 1818 4227
rect 1852 4193 1870 4227
rect 1800 4167 1870 4193
rect 1900 4227 1954 4253
rect 1900 4193 1912 4227
rect 1946 4193 1954 4227
rect 1900 4167 1954 4193
rect 516 4087 570 4113
rect 516 4053 524 4087
rect 558 4053 570 4087
rect 516 4027 570 4053
rect 600 4087 670 4113
rect 600 4053 618 4087
rect 652 4053 670 4087
rect 600 4027 670 4053
rect 700 4027 770 4113
rect 800 4027 870 4113
rect 900 4087 970 4113
rect 900 4053 918 4087
rect 952 4053 970 4087
rect 900 4027 970 4053
rect 1000 4087 1070 4113
rect 1000 4053 1018 4087
rect 1052 4053 1070 4087
rect 1000 4027 1070 4053
rect 1100 4087 1170 4113
rect 1100 4053 1118 4087
rect 1152 4053 1170 4087
rect 1100 4027 1170 4053
rect 1200 4087 1270 4113
rect 1200 4053 1218 4087
rect 1252 4053 1270 4087
rect 1200 4027 1270 4053
rect 1300 4087 1354 4113
rect 1300 4053 1312 4087
rect 1346 4053 1354 4087
rect 1300 4027 1354 4053
rect 1416 4087 1470 4113
rect 1416 4053 1424 4087
rect 1458 4053 1470 4087
rect 1416 4027 1470 4053
rect 1500 4087 1570 4113
rect 1500 4053 1518 4087
rect 1552 4053 1570 4087
rect 1500 4027 1570 4053
rect 1600 4087 1654 4113
rect 1600 4053 1612 4087
rect 1646 4053 1654 4087
rect 1600 4027 1654 4053
rect 2416 4507 2470 4533
rect 2416 4473 2424 4507
rect 2458 4473 2470 4507
rect 2416 4447 2470 4473
rect 2500 4507 2570 4533
rect 2500 4473 2518 4507
rect 2552 4473 2570 4507
rect 2500 4447 2570 4473
rect 2600 4507 2654 4533
rect 2600 4473 2612 4507
rect 2646 4473 2654 4507
rect 2600 4447 2654 4473
rect 2716 4507 2770 4533
rect 2716 4473 2724 4507
rect 2758 4473 2770 4507
rect 2716 4447 2770 4473
rect 2800 4507 2854 4533
rect 2800 4473 2812 4507
rect 2846 4473 2854 4507
rect 2800 4447 2854 4473
rect 3216 4787 3270 4813
rect 3216 4753 3224 4787
rect 3258 4753 3270 4787
rect 3216 4727 3270 4753
rect 3300 4787 3370 4813
rect 3300 4753 3318 4787
rect 3352 4753 3370 4787
rect 3300 4727 3370 4753
rect 3400 4787 3454 4813
rect 3400 4753 3412 4787
rect 3446 4753 3454 4787
rect 3400 4727 3454 4753
rect 3516 4787 3570 4813
rect 3516 4753 3524 4787
rect 3558 4753 3570 4787
rect 3516 4727 3570 4753
rect 3600 4787 3670 4813
rect 3600 4753 3618 4787
rect 3652 4753 3670 4787
rect 3600 4727 3670 4753
rect 3700 4727 3770 4813
rect 3800 4727 3870 4813
rect 3900 4787 3970 4813
rect 3900 4753 3918 4787
rect 3952 4753 3970 4787
rect 3900 4727 3970 4753
rect 4000 4787 4070 4813
rect 4000 4753 4018 4787
rect 4052 4753 4070 4787
rect 4000 4727 4070 4753
rect 4100 4787 4170 4813
rect 4100 4753 4118 4787
rect 4152 4753 4170 4787
rect 4100 4727 4170 4753
rect 4200 4787 4254 4813
rect 4200 4753 4212 4787
rect 4246 4753 4254 4787
rect 4200 4727 4254 4753
rect 3016 4647 3070 4673
rect 3016 4613 3024 4647
rect 3058 4613 3070 4647
rect 3016 4587 3070 4613
rect 3100 4647 3170 4673
rect 3100 4613 3118 4647
rect 3152 4613 3170 4647
rect 3100 4587 3170 4613
rect 3200 4647 3270 4673
rect 3200 4613 3218 4647
rect 3252 4613 3270 4647
rect 3200 4587 3270 4613
rect 3300 4647 3370 4673
rect 3300 4613 3318 4647
rect 3352 4613 3370 4647
rect 3300 4587 3370 4613
rect 3400 4587 3470 4673
rect 3500 4647 3570 4673
rect 3500 4613 3518 4647
rect 3552 4613 3570 4647
rect 3500 4587 3570 4613
rect 3600 4647 3654 4673
rect 3600 4613 3612 4647
rect 3646 4613 3654 4647
rect 3600 4587 3654 4613
rect 4316 4787 4370 4813
rect 4316 4753 4324 4787
rect 4358 4753 4370 4787
rect 4316 4727 4370 4753
rect 4400 4787 4470 4813
rect 4400 4753 4418 4787
rect 4452 4753 4470 4787
rect 4400 4727 4470 4753
rect 4500 4787 4570 4813
rect 4500 4753 4518 4787
rect 4552 4753 4570 4787
rect 4500 4727 4570 4753
rect 4600 4787 4670 4813
rect 4600 4753 4618 4787
rect 4652 4753 4670 4787
rect 4600 4727 4670 4753
rect 4700 4787 4770 4813
rect 4700 4753 4718 4787
rect 4752 4753 4770 4787
rect 4700 4727 4770 4753
rect 4800 4727 4870 4813
rect 4900 4787 4970 4813
rect 4900 4753 4918 4787
rect 4952 4753 4970 4787
rect 4900 4727 4970 4753
rect 5000 4787 5070 4813
rect 5000 4753 5018 4787
rect 5052 4753 5070 4787
rect 5000 4727 5070 4753
rect 5100 4727 5170 4813
rect 5200 4727 5270 4813
rect 5300 4787 5370 4813
rect 5300 4753 5318 4787
rect 5352 4753 5370 4787
rect 5300 4727 5370 4753
rect 5400 4787 5470 4813
rect 5400 4753 5418 4787
rect 5452 4753 5470 4787
rect 5400 4727 5470 4753
rect 5500 4787 5570 4813
rect 5500 4753 5518 4787
rect 5552 4753 5570 4787
rect 5500 4727 5570 4753
rect 5600 4727 5670 4813
rect 5700 4727 5770 4813
rect 5800 4727 5870 4813
rect 5900 4787 5970 4813
rect 5900 4753 5918 4787
rect 5952 4753 5970 4787
rect 5900 4727 5970 4753
rect 6000 4787 6070 4813
rect 6000 4753 6018 4787
rect 6052 4753 6070 4787
rect 6000 4727 6070 4753
rect 6100 4727 6170 4813
rect 6200 4727 6270 4813
rect 6300 4787 6370 4813
rect 6300 4753 6318 4787
rect 6352 4753 6370 4787
rect 6300 4727 6370 4753
rect 6400 4787 6454 4813
rect 6400 4753 6412 4787
rect 6446 4753 6454 4787
rect 6400 4727 6454 4753
rect 3716 4647 3770 4673
rect 3716 4613 3724 4647
rect 3758 4613 3770 4647
rect 3716 4587 3770 4613
rect 3800 4647 3870 4673
rect 3800 4613 3818 4647
rect 3852 4613 3870 4647
rect 3800 4587 3870 4613
rect 3900 4587 3970 4673
rect 4000 4647 4070 4673
rect 4000 4613 4018 4647
rect 4052 4613 4070 4647
rect 4000 4587 4070 4613
rect 4100 4647 4170 4673
rect 4100 4613 4118 4647
rect 4152 4613 4170 4647
rect 4100 4587 4170 4613
rect 4200 4587 4270 4673
rect 4300 4647 4370 4673
rect 4300 4613 4318 4647
rect 4352 4613 4370 4647
rect 4300 4587 4370 4613
rect 4400 4647 4470 4673
rect 4400 4613 4418 4647
rect 4452 4613 4470 4647
rect 4400 4587 4470 4613
rect 4500 4587 4570 4673
rect 4600 4647 4670 4673
rect 4600 4613 4618 4647
rect 4652 4613 4670 4647
rect 4600 4587 4670 4613
rect 4700 4647 4754 4673
rect 4700 4613 4712 4647
rect 4746 4613 4754 4647
rect 4700 4587 4754 4613
rect 2916 4507 2970 4533
rect 2916 4473 2924 4507
rect 2958 4473 2970 4507
rect 2916 4447 2970 4473
rect 3000 4507 3070 4533
rect 3000 4473 3018 4507
rect 3052 4473 3070 4507
rect 3000 4447 3070 4473
rect 3100 4447 3170 4533
rect 3200 4447 3270 4533
rect 3300 4447 3370 4533
rect 3400 4447 3470 4533
rect 3500 4507 3570 4533
rect 3500 4473 3518 4507
rect 3552 4473 3570 4507
rect 3500 4447 3570 4473
rect 3600 4507 3670 4533
rect 3600 4473 3618 4507
rect 3652 4473 3670 4507
rect 3600 4447 3670 4473
rect 3700 4507 3754 4533
rect 3700 4473 3712 4507
rect 3746 4473 3754 4507
rect 3700 4447 3754 4473
rect 2016 4367 2070 4393
rect 2016 4333 2024 4367
rect 2058 4333 2070 4367
rect 2016 4307 2070 4333
rect 2100 4367 2170 4393
rect 2100 4333 2118 4367
rect 2152 4333 2170 4367
rect 2100 4307 2170 4333
rect 2200 4367 2270 4393
rect 2200 4333 2218 4367
rect 2252 4333 2270 4367
rect 2200 4307 2270 4333
rect 2300 4367 2370 4393
rect 2300 4333 2318 4367
rect 2352 4333 2370 4367
rect 2300 4307 2370 4333
rect 2400 4367 2470 4393
rect 2400 4333 2418 4367
rect 2452 4333 2470 4367
rect 2400 4307 2470 4333
rect 2500 4367 2570 4393
rect 2500 4333 2518 4367
rect 2552 4333 2570 4367
rect 2500 4307 2570 4333
rect 2600 4307 2670 4393
rect 2700 4307 2770 4393
rect 2800 4367 2870 4393
rect 2800 4333 2818 4367
rect 2852 4333 2870 4367
rect 2800 4307 2870 4333
rect 2900 4367 2970 4393
rect 2900 4333 2918 4367
rect 2952 4333 2970 4367
rect 2900 4307 2970 4333
rect 3000 4307 3070 4393
rect 3100 4367 3170 4393
rect 3100 4333 3118 4367
rect 3152 4333 3170 4367
rect 3100 4307 3170 4333
rect 3200 4367 3270 4393
rect 3200 4333 3218 4367
rect 3252 4333 3270 4367
rect 3200 4307 3270 4333
rect 3300 4367 3370 4393
rect 3300 4333 3318 4367
rect 3352 4333 3370 4367
rect 3300 4307 3370 4333
rect 3400 4307 3470 4393
rect 3500 4367 3570 4393
rect 3500 4333 3518 4367
rect 3552 4333 3570 4367
rect 3500 4307 3570 4333
rect 3600 4367 3670 4393
rect 3600 4333 3618 4367
rect 3652 4333 3670 4367
rect 3600 4307 3670 4333
rect 3700 4367 3754 4393
rect 3700 4333 3712 4367
rect 3746 4333 3754 4367
rect 3700 4307 3754 4333
rect 4816 4647 4870 4673
rect 4816 4613 4824 4647
rect 4858 4613 4870 4647
rect 4816 4587 4870 4613
rect 4900 4647 4970 4673
rect 4900 4613 4918 4647
rect 4952 4613 4970 4647
rect 4900 4587 4970 4613
rect 5000 4647 5054 4673
rect 5000 4613 5012 4647
rect 5046 4613 5054 4647
rect 5000 4587 5054 4613
rect 3816 4507 3870 4533
rect 3816 4473 3824 4507
rect 3858 4473 3870 4507
rect 3816 4447 3870 4473
rect 3900 4507 3970 4533
rect 3900 4473 3918 4507
rect 3952 4473 3970 4507
rect 3900 4447 3970 4473
rect 4000 4507 4070 4533
rect 4000 4473 4018 4507
rect 4052 4473 4070 4507
rect 4000 4447 4070 4473
rect 4100 4507 4170 4533
rect 4100 4473 4118 4507
rect 4152 4473 4170 4507
rect 4100 4447 4170 4473
rect 4200 4507 4270 4533
rect 4200 4473 4218 4507
rect 4252 4473 4270 4507
rect 4200 4447 4270 4473
rect 4300 4507 4370 4533
rect 4300 4473 4318 4507
rect 4352 4473 4370 4507
rect 4300 4447 4370 4473
rect 4400 4447 4470 4533
rect 4500 4447 4570 4533
rect 4600 4507 4670 4533
rect 4600 4473 4618 4507
rect 4652 4473 4670 4507
rect 4600 4447 4670 4473
rect 4700 4507 4770 4533
rect 4700 4473 4718 4507
rect 4752 4473 4770 4507
rect 4700 4447 4770 4473
rect 4800 4447 4870 4533
rect 4900 4507 4970 4533
rect 4900 4473 4918 4507
rect 4952 4473 4970 4507
rect 4900 4447 4970 4473
rect 5000 4507 5054 4533
rect 5000 4473 5012 4507
rect 5046 4473 5054 4507
rect 5000 4447 5054 4473
rect 5116 4647 5170 4673
rect 5116 4613 5124 4647
rect 5158 4613 5170 4647
rect 5116 4587 5170 4613
rect 5200 4647 5270 4673
rect 5200 4613 5218 4647
rect 5252 4613 5270 4647
rect 5200 4587 5270 4613
rect 5300 4647 5370 4673
rect 5300 4613 5318 4647
rect 5352 4613 5370 4647
rect 5300 4587 5370 4613
rect 5400 4587 5470 4673
rect 5500 4587 5570 4673
rect 5600 4587 5670 4673
rect 5700 4647 5770 4673
rect 5700 4613 5718 4647
rect 5752 4613 5770 4647
rect 5700 4587 5770 4613
rect 5800 4647 5854 4673
rect 5800 4613 5812 4647
rect 5846 4613 5854 4647
rect 5800 4587 5854 4613
rect 5116 4507 5170 4533
rect 5116 4473 5124 4507
rect 5158 4473 5170 4507
rect 5116 4447 5170 4473
rect 5200 4507 5270 4533
rect 5200 4473 5218 4507
rect 5252 4473 5270 4507
rect 5200 4447 5270 4473
rect 5300 4507 5354 4533
rect 5300 4473 5312 4507
rect 5346 4473 5354 4507
rect 5300 4447 5354 4473
rect 5916 4647 5970 4673
rect 5916 4613 5924 4647
rect 5958 4613 5970 4647
rect 5916 4587 5970 4613
rect 6000 4647 6070 4673
rect 6000 4613 6018 4647
rect 6052 4613 6070 4647
rect 6000 4587 6070 4613
rect 6100 4647 6170 4673
rect 6100 4613 6118 4647
rect 6152 4613 6170 4647
rect 6100 4587 6170 4613
rect 6200 4647 6270 4673
rect 6200 4613 6218 4647
rect 6252 4613 6270 4647
rect 6200 4587 6270 4613
rect 6300 4647 6370 4673
rect 6300 4613 6318 4647
rect 6352 4613 6370 4647
rect 6300 4587 6370 4613
rect 6400 4647 6454 4673
rect 6400 4613 6412 4647
rect 6446 4613 6454 4647
rect 6400 4587 6454 4613
rect 5416 4507 5470 4533
rect 5416 4473 5424 4507
rect 5458 4473 5470 4507
rect 5416 4447 5470 4473
rect 5500 4507 5570 4533
rect 5500 4473 5518 4507
rect 5552 4473 5570 4507
rect 5500 4447 5570 4473
rect 5600 4447 5670 4533
rect 5700 4447 5770 4533
rect 5800 4447 5870 4533
rect 5900 4507 5970 4533
rect 5900 4473 5918 4507
rect 5952 4473 5970 4507
rect 5900 4447 5970 4473
rect 6000 4507 6054 4533
rect 6000 4473 6012 4507
rect 6046 4473 6054 4507
rect 6000 4447 6054 4473
rect 3816 4367 3870 4393
rect 3816 4333 3824 4367
rect 3858 4333 3870 4367
rect 3816 4307 3870 4333
rect 3900 4367 3970 4393
rect 3900 4333 3918 4367
rect 3952 4333 3970 4367
rect 3900 4307 3970 4333
rect 4000 4367 4070 4393
rect 4000 4333 4018 4367
rect 4052 4333 4070 4367
rect 4000 4307 4070 4333
rect 4100 4367 4170 4393
rect 4100 4333 4118 4367
rect 4152 4333 4170 4367
rect 4100 4307 4170 4333
rect 4200 4367 4270 4393
rect 4200 4333 4218 4367
rect 4252 4333 4270 4367
rect 4200 4307 4270 4333
rect 4300 4307 4370 4393
rect 4400 4367 4470 4393
rect 4400 4333 4418 4367
rect 4452 4333 4470 4367
rect 4400 4307 4470 4333
rect 4500 4367 4570 4393
rect 4500 4333 4518 4367
rect 4552 4333 4570 4367
rect 4500 4307 4570 4333
rect 4600 4367 4670 4393
rect 4600 4333 4618 4367
rect 4652 4333 4670 4367
rect 4600 4307 4670 4333
rect 4700 4307 4770 4393
rect 4800 4367 4870 4393
rect 4800 4333 4818 4367
rect 4852 4333 4870 4367
rect 4800 4307 4870 4333
rect 4900 4367 4970 4393
rect 4900 4333 4918 4367
rect 4952 4333 4970 4367
rect 4900 4307 4970 4333
rect 5000 4367 5070 4393
rect 5000 4333 5018 4367
rect 5052 4333 5070 4367
rect 5000 4307 5070 4333
rect 5100 4307 5170 4393
rect 5200 4367 5270 4393
rect 5200 4333 5218 4367
rect 5252 4333 5270 4367
rect 5200 4307 5270 4333
rect 5300 4367 5370 4393
rect 5300 4333 5318 4367
rect 5352 4333 5370 4367
rect 5300 4307 5370 4333
rect 5400 4307 5470 4393
rect 5500 4367 5570 4393
rect 5500 4333 5518 4367
rect 5552 4333 5570 4367
rect 5500 4307 5570 4333
rect 5600 4367 5670 4393
rect 5600 4333 5618 4367
rect 5652 4333 5670 4367
rect 5600 4307 5670 4333
rect 5700 4307 5770 4393
rect 5800 4307 5870 4393
rect 5900 4367 5970 4393
rect 5900 4333 5918 4367
rect 5952 4333 5970 4367
rect 5900 4307 5970 4333
rect 6000 4367 6054 4393
rect 6000 4333 6012 4367
rect 6046 4333 6054 4367
rect 6000 4307 6054 4333
rect 2016 4227 2070 4253
rect 2016 4193 2024 4227
rect 2058 4193 2070 4227
rect 2016 4167 2070 4193
rect 2100 4227 2170 4253
rect 2100 4193 2118 4227
rect 2152 4193 2170 4227
rect 2100 4167 2170 4193
rect 2200 4167 2270 4253
rect 2300 4227 2370 4253
rect 2300 4193 2318 4227
rect 2352 4193 2370 4227
rect 2300 4167 2370 4193
rect 2400 4227 2470 4253
rect 2400 4193 2418 4227
rect 2452 4193 2470 4227
rect 2400 4167 2470 4193
rect 2500 4227 2570 4253
rect 2500 4193 2518 4227
rect 2552 4193 2570 4227
rect 2500 4167 2570 4193
rect 2600 4167 2670 4253
rect 2700 4167 2770 4253
rect 2800 4227 2870 4253
rect 2800 4193 2818 4227
rect 2852 4193 2870 4227
rect 2800 4167 2870 4193
rect 2900 4227 2970 4253
rect 2900 4193 2918 4227
rect 2952 4193 2970 4227
rect 2900 4167 2970 4193
rect 3000 4227 3070 4253
rect 3000 4193 3018 4227
rect 3052 4193 3070 4227
rect 3000 4167 3070 4193
rect 3100 4167 3170 4253
rect 3200 4227 3270 4253
rect 3200 4193 3218 4227
rect 3252 4193 3270 4227
rect 3200 4167 3270 4193
rect 3300 4227 3370 4253
rect 3300 4193 3318 4227
rect 3352 4193 3370 4227
rect 3300 4167 3370 4193
rect 3400 4167 3470 4253
rect 3500 4167 3570 4253
rect 3600 4227 3670 4253
rect 3600 4193 3618 4227
rect 3652 4193 3670 4227
rect 3600 4167 3670 4193
rect 3700 4227 3770 4253
rect 3700 4193 3718 4227
rect 3752 4193 3770 4227
rect 3700 4167 3770 4193
rect 3800 4227 3870 4253
rect 3800 4193 3818 4227
rect 3852 4193 3870 4227
rect 3800 4167 3870 4193
rect 3900 4227 3970 4253
rect 3900 4193 3918 4227
rect 3952 4193 3970 4227
rect 3900 4167 3970 4193
rect 4000 4227 4054 4253
rect 4000 4193 4012 4227
rect 4046 4193 4054 4227
rect 4000 4167 4054 4193
rect 1716 4087 1770 4113
rect 1716 4053 1724 4087
rect 1758 4053 1770 4087
rect 1716 4027 1770 4053
rect 1800 4087 1870 4113
rect 1800 4053 1818 4087
rect 1852 4053 1870 4087
rect 1800 4027 1870 4053
rect 1900 4027 1970 4113
rect 2000 4087 2070 4113
rect 2000 4053 2018 4087
rect 2052 4053 2070 4087
rect 2000 4027 2070 4053
rect 2100 4087 2170 4113
rect 2100 4053 2118 4087
rect 2152 4053 2170 4087
rect 2100 4027 2170 4053
rect 2200 4087 2254 4113
rect 2200 4053 2212 4087
rect 2246 4053 2254 4087
rect 2200 4027 2254 4053
rect 16 3947 70 3973
rect 16 3913 24 3947
rect 58 3913 70 3947
rect 16 3887 70 3913
rect 100 3947 170 3973
rect 100 3913 118 3947
rect 152 3913 170 3947
rect 100 3887 170 3913
rect 200 3947 270 3973
rect 200 3913 218 3947
rect 252 3913 270 3947
rect 200 3887 270 3913
rect 300 3947 370 3973
rect 300 3913 318 3947
rect 352 3913 370 3947
rect 300 3887 370 3913
rect 400 3887 470 3973
rect 500 3887 570 3973
rect 600 3947 670 3973
rect 600 3913 618 3947
rect 652 3913 670 3947
rect 600 3887 670 3913
rect 700 3947 770 3973
rect 700 3913 718 3947
rect 752 3913 770 3947
rect 700 3887 770 3913
rect 800 3887 870 3973
rect 900 3947 970 3973
rect 900 3913 918 3947
rect 952 3913 970 3947
rect 900 3887 970 3913
rect 1000 3947 1070 3973
rect 1000 3913 1018 3947
rect 1052 3913 1070 3947
rect 1000 3887 1070 3913
rect 1100 3947 1170 3973
rect 1100 3913 1118 3947
rect 1152 3913 1170 3947
rect 1100 3887 1170 3913
rect 1200 3887 1270 3973
rect 1300 3887 1370 3973
rect 1400 3887 1470 3973
rect 1500 3947 1570 3973
rect 1500 3913 1518 3947
rect 1552 3913 1570 3947
rect 1500 3887 1570 3913
rect 1600 3947 1670 3973
rect 1600 3913 1618 3947
rect 1652 3913 1670 3947
rect 1600 3887 1670 3913
rect 1700 3887 1770 3973
rect 1800 3947 1870 3973
rect 1800 3913 1818 3947
rect 1852 3913 1870 3947
rect 1800 3887 1870 3913
rect 1900 3947 1954 3973
rect 1900 3913 1912 3947
rect 1946 3913 1954 3947
rect 1900 3887 1954 3913
rect 2316 4087 2370 4113
rect 2316 4053 2324 4087
rect 2358 4053 2370 4087
rect 2316 4027 2370 4053
rect 2400 4087 2470 4113
rect 2400 4053 2418 4087
rect 2452 4053 2470 4087
rect 2400 4027 2470 4053
rect 2500 4087 2570 4113
rect 2500 4053 2518 4087
rect 2552 4053 2570 4087
rect 2500 4027 2570 4053
rect 2600 4087 2654 4113
rect 2600 4053 2612 4087
rect 2646 4053 2654 4087
rect 2600 4027 2654 4053
rect 2716 4087 2770 4113
rect 2716 4053 2724 4087
rect 2758 4053 2770 4087
rect 2716 4027 2770 4053
rect 2800 4087 2870 4113
rect 2800 4053 2818 4087
rect 2852 4053 2870 4087
rect 2800 4027 2870 4053
rect 2900 4087 2954 4113
rect 2900 4053 2912 4087
rect 2946 4053 2954 4087
rect 2900 4027 2954 4053
rect 3016 4087 3070 4113
rect 3016 4053 3024 4087
rect 3058 4053 3070 4087
rect 3016 4027 3070 4053
rect 3100 4087 3170 4113
rect 3100 4053 3118 4087
rect 3152 4053 3170 4087
rect 3100 4027 3170 4053
rect 3200 4087 3254 4113
rect 3200 4053 3212 4087
rect 3246 4053 3254 4087
rect 3200 4027 3254 4053
rect 4116 4227 4170 4253
rect 4116 4193 4124 4227
rect 4158 4193 4170 4227
rect 4116 4167 4170 4193
rect 4200 4227 4254 4253
rect 4200 4193 4212 4227
rect 4246 4193 4254 4227
rect 4200 4167 4254 4193
rect 3316 4087 3370 4113
rect 3316 4053 3324 4087
rect 3358 4053 3370 4087
rect 3316 4027 3370 4053
rect 3400 4087 3470 4113
rect 3400 4053 3418 4087
rect 3452 4053 3470 4087
rect 3400 4027 3470 4053
rect 3500 4087 3570 4113
rect 3500 4053 3518 4087
rect 3552 4053 3570 4087
rect 3500 4027 3570 4053
rect 3600 4087 3670 4113
rect 3600 4053 3618 4087
rect 3652 4053 3670 4087
rect 3600 4027 3670 4053
rect 3700 4027 3770 4113
rect 3800 4027 3870 4113
rect 3900 4087 3970 4113
rect 3900 4053 3918 4087
rect 3952 4053 3970 4087
rect 3900 4027 3970 4053
rect 4000 4087 4070 4113
rect 4000 4053 4018 4087
rect 4052 4053 4070 4087
rect 4000 4027 4070 4053
rect 4100 4087 4154 4113
rect 4100 4053 4112 4087
rect 4146 4053 4154 4087
rect 4100 4027 4154 4053
rect 2016 3947 2070 3973
rect 2016 3913 2024 3947
rect 2058 3913 2070 3947
rect 2016 3887 2070 3913
rect 2100 3947 2170 3973
rect 2100 3913 2118 3947
rect 2152 3913 2170 3947
rect 2100 3887 2170 3913
rect 2200 3887 2270 3973
rect 2300 3887 2370 3973
rect 2400 3887 2470 3973
rect 2500 3887 2570 3973
rect 2600 3887 2670 3973
rect 2700 3887 2770 3973
rect 2800 3887 2870 3973
rect 2900 3947 2970 3973
rect 2900 3913 2918 3947
rect 2952 3913 2970 3947
rect 2900 3887 2970 3913
rect 3000 3947 3070 3973
rect 3000 3913 3018 3947
rect 3052 3913 3070 3947
rect 3000 3887 3070 3913
rect 3100 3947 3170 3973
rect 3100 3913 3118 3947
rect 3152 3913 3170 3947
rect 3100 3887 3170 3913
rect 3200 3947 3270 3973
rect 3200 3913 3218 3947
rect 3252 3913 3270 3947
rect 3200 3887 3270 3913
rect 3300 3947 3370 3973
rect 3300 3913 3318 3947
rect 3352 3913 3370 3947
rect 3300 3887 3370 3913
rect 3400 3887 3470 3973
rect 3500 3887 3570 3973
rect 3600 3947 3670 3973
rect 3600 3913 3618 3947
rect 3652 3913 3670 3947
rect 3600 3887 3670 3913
rect 3700 3947 3770 3973
rect 3700 3913 3718 3947
rect 3752 3913 3770 3947
rect 3700 3887 3770 3913
rect 3800 3947 3870 3973
rect 3800 3913 3818 3947
rect 3852 3913 3870 3947
rect 3800 3887 3870 3913
rect 3900 3947 3954 3973
rect 3900 3913 3912 3947
rect 3946 3913 3954 3947
rect 3900 3887 3954 3913
rect 16 3807 70 3833
rect 16 3773 24 3807
rect 58 3773 70 3807
rect 16 3747 70 3773
rect 100 3807 170 3833
rect 100 3773 118 3807
rect 152 3773 170 3807
rect 100 3747 170 3773
rect 200 3807 270 3833
rect 200 3773 218 3807
rect 252 3773 270 3807
rect 200 3747 270 3773
rect 300 3747 370 3833
rect 400 3747 470 3833
rect 500 3747 570 3833
rect 600 3807 670 3833
rect 600 3773 618 3807
rect 652 3773 670 3807
rect 600 3747 670 3773
rect 700 3807 770 3833
rect 700 3773 718 3807
rect 752 3773 770 3807
rect 700 3747 770 3773
rect 800 3747 870 3833
rect 900 3747 970 3833
rect 1000 3807 1070 3833
rect 1000 3773 1018 3807
rect 1052 3773 1070 3807
rect 1000 3747 1070 3773
rect 1100 3807 1170 3833
rect 1100 3773 1118 3807
rect 1152 3773 1170 3807
rect 1100 3747 1170 3773
rect 1200 3747 1270 3833
rect 1300 3747 1370 3833
rect 1400 3747 1470 3833
rect 1500 3747 1570 3833
rect 1600 3747 1670 3833
rect 1700 3807 1770 3833
rect 1700 3773 1718 3807
rect 1752 3773 1770 3807
rect 1700 3747 1770 3773
rect 1800 3807 1870 3833
rect 1800 3773 1818 3807
rect 1852 3773 1870 3807
rect 1800 3747 1870 3773
rect 1900 3747 1970 3833
rect 2000 3807 2070 3833
rect 2000 3773 2018 3807
rect 2052 3773 2070 3807
rect 2000 3747 2070 3773
rect 2100 3807 2154 3833
rect 2100 3773 2112 3807
rect 2146 3773 2154 3807
rect 2100 3747 2154 3773
rect 16 3517 70 3603
rect 100 3517 170 3603
rect 200 3517 270 3603
rect 300 3517 370 3603
rect 400 3517 470 3603
rect 500 3577 570 3603
rect 500 3543 518 3577
rect 552 3543 570 3577
rect 500 3517 570 3543
rect 600 3577 670 3603
rect 600 3543 618 3577
rect 652 3543 670 3577
rect 600 3517 670 3543
rect 700 3577 770 3603
rect 700 3543 718 3577
rect 752 3543 770 3577
rect 700 3517 770 3543
rect 800 3577 854 3603
rect 800 3543 812 3577
rect 846 3543 854 3577
rect 800 3517 854 3543
rect 16 3437 70 3463
rect 16 3403 24 3437
rect 58 3403 70 3437
rect 16 3377 70 3403
rect 100 3437 170 3463
rect 100 3403 118 3437
rect 152 3403 170 3437
rect 100 3377 170 3403
rect 200 3437 270 3463
rect 200 3403 218 3437
rect 252 3403 270 3437
rect 200 3377 270 3403
rect 300 3437 354 3463
rect 300 3403 312 3437
rect 346 3403 354 3437
rect 300 3377 354 3403
rect 416 3437 470 3463
rect 416 3403 424 3437
rect 458 3403 470 3437
rect 416 3377 470 3403
rect 500 3437 554 3463
rect 500 3403 512 3437
rect 546 3403 554 3437
rect 500 3377 554 3403
rect 616 3437 670 3463
rect 616 3403 624 3437
rect 658 3403 670 3437
rect 616 3377 670 3403
rect 700 3437 754 3463
rect 700 3403 712 3437
rect 746 3403 754 3437
rect 700 3377 754 3403
rect 16 3237 70 3323
rect 100 3297 170 3323
rect 100 3263 118 3297
rect 152 3263 170 3297
rect 100 3237 170 3263
rect 200 3297 270 3323
rect 200 3263 218 3297
rect 252 3263 270 3297
rect 200 3237 270 3263
rect 300 3297 370 3323
rect 300 3263 318 3297
rect 352 3263 370 3297
rect 300 3237 370 3263
rect 400 3297 470 3323
rect 400 3263 418 3297
rect 452 3263 470 3297
rect 400 3237 470 3263
rect 500 3297 570 3323
rect 500 3263 518 3297
rect 552 3263 570 3297
rect 500 3237 570 3263
rect 600 3297 670 3323
rect 600 3263 618 3297
rect 652 3263 670 3297
rect 600 3237 670 3263
rect 700 3297 754 3323
rect 700 3263 712 3297
rect 746 3263 754 3297
rect 700 3237 754 3263
rect 16 3157 70 3183
rect 16 3123 24 3157
rect 58 3123 70 3157
rect 16 3097 70 3123
rect 100 3157 154 3183
rect 100 3123 112 3157
rect 146 3123 154 3157
rect 100 3097 154 3123
rect 916 3577 970 3603
rect 916 3543 924 3577
rect 958 3543 970 3577
rect 916 3517 970 3543
rect 1000 3577 1054 3603
rect 1000 3543 1012 3577
rect 1046 3543 1054 3577
rect 1000 3517 1054 3543
rect 816 3437 870 3463
rect 816 3403 824 3437
rect 858 3403 870 3437
rect 816 3377 870 3403
rect 900 3437 954 3463
rect 900 3403 912 3437
rect 946 3403 954 3437
rect 900 3377 954 3403
rect 816 3297 870 3323
rect 816 3263 824 3297
rect 858 3263 870 3297
rect 816 3237 870 3263
rect 900 3297 954 3323
rect 900 3263 912 3297
rect 946 3263 954 3297
rect 900 3237 954 3263
rect 2216 3807 2270 3833
rect 2216 3773 2224 3807
rect 2258 3773 2270 3807
rect 2216 3747 2270 3773
rect 2300 3807 2370 3833
rect 2300 3773 2318 3807
rect 2352 3773 2370 3807
rect 2300 3747 2370 3773
rect 2400 3807 2470 3833
rect 2400 3773 2418 3807
rect 2452 3773 2470 3807
rect 2400 3747 2470 3773
rect 2500 3807 2554 3833
rect 2500 3773 2512 3807
rect 2546 3773 2554 3807
rect 2500 3747 2554 3773
rect 2616 3807 2670 3833
rect 2616 3773 2624 3807
rect 2658 3773 2670 3807
rect 2616 3747 2670 3773
rect 2700 3807 2754 3833
rect 2700 3773 2712 3807
rect 2746 3773 2754 3807
rect 2700 3747 2754 3773
rect 1116 3577 1170 3603
rect 1116 3543 1124 3577
rect 1158 3543 1170 3577
rect 1116 3517 1170 3543
rect 1200 3577 1270 3603
rect 1200 3543 1218 3577
rect 1252 3543 1270 3577
rect 1200 3517 1270 3543
rect 1300 3577 1370 3603
rect 1300 3543 1318 3577
rect 1352 3543 1370 3577
rect 1300 3517 1370 3543
rect 1400 3577 1470 3603
rect 1400 3543 1418 3577
rect 1452 3543 1470 3577
rect 1400 3517 1470 3543
rect 1500 3517 1570 3603
rect 1600 3577 1670 3603
rect 1600 3543 1618 3577
rect 1652 3543 1670 3577
rect 1600 3517 1670 3543
rect 1700 3577 1770 3603
rect 1700 3543 1718 3577
rect 1752 3543 1770 3577
rect 1700 3517 1770 3543
rect 1800 3577 1870 3603
rect 1800 3543 1818 3577
rect 1852 3543 1870 3577
rect 1800 3517 1870 3543
rect 1900 3577 1970 3603
rect 1900 3543 1918 3577
rect 1952 3543 1970 3577
rect 1900 3517 1970 3543
rect 2000 3577 2070 3603
rect 2000 3543 2018 3577
rect 2052 3543 2070 3577
rect 2000 3517 2070 3543
rect 2100 3577 2170 3603
rect 2100 3543 2118 3577
rect 2152 3543 2170 3577
rect 2100 3517 2170 3543
rect 2200 3577 2270 3603
rect 2200 3543 2218 3577
rect 2252 3543 2270 3577
rect 2200 3517 2270 3543
rect 2300 3577 2370 3603
rect 2300 3543 2318 3577
rect 2352 3543 2370 3577
rect 2300 3517 2370 3543
rect 2400 3577 2470 3603
rect 2400 3543 2418 3577
rect 2452 3543 2470 3577
rect 2400 3517 2470 3543
rect 2500 3577 2554 3603
rect 2500 3543 2512 3577
rect 2546 3543 2554 3577
rect 2500 3517 2554 3543
rect 2816 3807 2870 3833
rect 2816 3773 2824 3807
rect 2858 3773 2870 3807
rect 2816 3747 2870 3773
rect 2900 3807 2970 3833
rect 2900 3773 2918 3807
rect 2952 3773 2970 3807
rect 2900 3747 2970 3773
rect 3000 3807 3070 3833
rect 3000 3773 3018 3807
rect 3052 3773 3070 3807
rect 3000 3747 3070 3773
rect 3100 3807 3154 3833
rect 3100 3773 3112 3807
rect 3146 3773 3154 3807
rect 3100 3747 3154 3773
rect 4016 3947 4070 3973
rect 4016 3913 4024 3947
rect 4058 3913 4070 3947
rect 4016 3887 4070 3913
rect 4100 3947 4154 3973
rect 4100 3913 4112 3947
rect 4146 3913 4154 3947
rect 4100 3887 4154 3913
rect 4316 4227 4370 4253
rect 4316 4193 4324 4227
rect 4358 4193 4370 4227
rect 4316 4167 4370 4193
rect 4400 4227 4454 4253
rect 4400 4193 4412 4227
rect 4446 4193 4454 4227
rect 4400 4167 4454 4193
rect 4216 4087 4270 4113
rect 4216 4053 4224 4087
rect 4258 4053 4270 4087
rect 4216 4027 4270 4053
rect 4300 4087 4354 4113
rect 4300 4053 4312 4087
rect 4346 4053 4354 4087
rect 4300 4027 4354 4053
rect 4516 4227 4570 4253
rect 4516 4193 4524 4227
rect 4558 4193 4570 4227
rect 4516 4167 4570 4193
rect 4600 4227 4654 4253
rect 4600 4193 4612 4227
rect 4646 4193 4654 4227
rect 4600 4167 4654 4193
rect 4416 4087 4470 4113
rect 4416 4053 4424 4087
rect 4458 4053 4470 4087
rect 4416 4027 4470 4053
rect 4500 4087 4554 4113
rect 4500 4053 4512 4087
rect 4546 4053 4554 4087
rect 4500 4027 4554 4053
rect 4716 4227 4770 4253
rect 4716 4193 4724 4227
rect 4758 4193 4770 4227
rect 4716 4167 4770 4193
rect 4800 4227 4854 4253
rect 4800 4193 4812 4227
rect 4846 4193 4854 4227
rect 4800 4167 4854 4193
rect 4616 4087 4670 4113
rect 4616 4053 4624 4087
rect 4658 4053 4670 4087
rect 4616 4027 4670 4053
rect 4700 4087 4754 4113
rect 4700 4053 4712 4087
rect 4746 4053 4754 4087
rect 4700 4027 4754 4053
rect 4916 4227 4970 4253
rect 4916 4193 4924 4227
rect 4958 4193 4970 4227
rect 4916 4167 4970 4193
rect 5000 4227 5070 4253
rect 5000 4193 5018 4227
rect 5052 4193 5070 4227
rect 5000 4167 5070 4193
rect 5100 4167 5170 4253
rect 5200 4167 5270 4253
rect 5300 4227 5370 4253
rect 5300 4193 5318 4227
rect 5352 4193 5370 4227
rect 5300 4167 5370 4193
rect 5400 4227 5470 4253
rect 5400 4193 5418 4227
rect 5452 4193 5470 4227
rect 5400 4167 5470 4193
rect 5500 4227 5554 4253
rect 5500 4193 5512 4227
rect 5546 4193 5554 4227
rect 5500 4167 5554 4193
rect 4816 4087 4870 4113
rect 4816 4053 4824 4087
rect 4858 4053 4870 4087
rect 4816 4027 4870 4053
rect 4900 4087 4954 4113
rect 4900 4053 4912 4087
rect 4946 4053 4954 4087
rect 4900 4027 4954 4053
rect 5016 4087 5070 4113
rect 5016 4053 5024 4087
rect 5058 4053 5070 4087
rect 5016 4027 5070 4053
rect 5100 4087 5170 4113
rect 5100 4053 5118 4087
rect 5152 4053 5170 4087
rect 5100 4027 5170 4053
rect 5200 4087 5254 4113
rect 5200 4053 5212 4087
rect 5246 4053 5254 4087
rect 5200 4027 5254 4053
rect 4216 3947 4270 3973
rect 4216 3913 4224 3947
rect 4258 3913 4270 3947
rect 4216 3887 4270 3913
rect 4300 3947 4370 3973
rect 4300 3913 4318 3947
rect 4352 3913 4370 3947
rect 4300 3887 4370 3913
rect 4400 3947 4470 3973
rect 4400 3913 4418 3947
rect 4452 3913 4470 3947
rect 4400 3887 4470 3913
rect 4500 3887 4570 3973
rect 4600 3947 4670 3973
rect 4600 3913 4618 3947
rect 4652 3913 4670 3947
rect 4600 3887 4670 3913
rect 4700 3947 4770 3973
rect 4700 3913 4718 3947
rect 4752 3913 4770 3947
rect 4700 3887 4770 3913
rect 4800 3887 4870 3973
rect 4900 3947 4970 3973
rect 4900 3913 4918 3947
rect 4952 3913 4970 3947
rect 4900 3887 4970 3913
rect 5000 3947 5054 3973
rect 5000 3913 5012 3947
rect 5046 3913 5054 3947
rect 5000 3887 5054 3913
rect 3216 3807 3270 3833
rect 3216 3773 3224 3807
rect 3258 3773 3270 3807
rect 3216 3747 3270 3773
rect 3300 3807 3370 3833
rect 3300 3773 3318 3807
rect 3352 3773 3370 3807
rect 3300 3747 3370 3773
rect 3400 3747 3470 3833
rect 3500 3747 3570 3833
rect 3600 3807 3670 3833
rect 3600 3773 3618 3807
rect 3652 3773 3670 3807
rect 3600 3747 3670 3773
rect 3700 3807 3770 3833
rect 3700 3773 3718 3807
rect 3752 3773 3770 3807
rect 3700 3747 3770 3773
rect 3800 3747 3870 3833
rect 3900 3807 3970 3833
rect 3900 3773 3918 3807
rect 3952 3773 3970 3807
rect 3900 3747 3970 3773
rect 4000 3807 4070 3833
rect 4000 3773 4018 3807
rect 4052 3773 4070 3807
rect 4000 3747 4070 3773
rect 4100 3747 4170 3833
rect 4200 3807 4270 3833
rect 4200 3773 4218 3807
rect 4252 3773 4270 3807
rect 4200 3747 4270 3773
rect 4300 3807 4370 3833
rect 4300 3773 4318 3807
rect 4352 3773 4370 3807
rect 4300 3747 4370 3773
rect 4400 3807 4470 3833
rect 4400 3773 4418 3807
rect 4452 3773 4470 3807
rect 4400 3747 4470 3773
rect 4500 3807 4554 3833
rect 4500 3773 4512 3807
rect 4546 3773 4554 3807
rect 4500 3747 4554 3773
rect 2616 3577 2670 3603
rect 2616 3543 2624 3577
rect 2658 3543 2670 3577
rect 2616 3517 2670 3543
rect 2700 3577 2770 3603
rect 2700 3543 2718 3577
rect 2752 3543 2770 3577
rect 2700 3517 2770 3543
rect 2800 3517 2870 3603
rect 2900 3577 2970 3603
rect 2900 3543 2918 3577
rect 2952 3543 2970 3577
rect 2900 3517 2970 3543
rect 3000 3577 3070 3603
rect 3000 3543 3018 3577
rect 3052 3543 3070 3577
rect 3000 3517 3070 3543
rect 3100 3577 3154 3603
rect 3100 3543 3112 3577
rect 3146 3543 3154 3577
rect 3100 3517 3154 3543
rect 5116 3947 5170 3973
rect 5116 3913 5124 3947
rect 5158 3913 5170 3947
rect 5116 3887 5170 3913
rect 5200 3947 5254 3973
rect 5200 3913 5212 3947
rect 5246 3913 5254 3947
rect 5200 3887 5254 3913
rect 5616 4227 5670 4253
rect 5616 4193 5624 4227
rect 5658 4193 5670 4227
rect 5616 4167 5670 4193
rect 5700 4227 5770 4253
rect 5700 4193 5718 4227
rect 5752 4193 5770 4227
rect 5700 4167 5770 4193
rect 5800 4167 5870 4253
rect 5900 4227 5970 4253
rect 5900 4193 5918 4227
rect 5952 4193 5970 4227
rect 5900 4167 5970 4193
rect 6000 4227 6054 4253
rect 6000 4193 6012 4227
rect 6046 4193 6054 4227
rect 6000 4167 6054 4193
rect 5316 4087 5370 4113
rect 5316 4053 5324 4087
rect 5358 4053 5370 4087
rect 5316 4027 5370 4053
rect 5400 4087 5470 4113
rect 5400 4053 5418 4087
rect 5452 4053 5470 4087
rect 5400 4027 5470 4053
rect 5500 4087 5570 4113
rect 5500 4053 5518 4087
rect 5552 4053 5570 4087
rect 5500 4027 5570 4053
rect 5600 4087 5654 4113
rect 5600 4053 5612 4087
rect 5646 4053 5654 4087
rect 5600 4027 5654 4053
rect 5316 3947 5370 3973
rect 5316 3913 5324 3947
rect 5358 3913 5370 3947
rect 5316 3887 5370 3913
rect 5400 3947 5470 3973
rect 5400 3913 5418 3947
rect 5452 3913 5470 3947
rect 5400 3887 5470 3913
rect 5500 3947 5554 3973
rect 5500 3913 5512 3947
rect 5546 3913 5554 3947
rect 5500 3887 5554 3913
rect 4616 3807 4670 3833
rect 4616 3773 4624 3807
rect 4658 3773 4670 3807
rect 4616 3747 4670 3773
rect 4700 3807 4770 3833
rect 4700 3773 4718 3807
rect 4752 3773 4770 3807
rect 4700 3747 4770 3773
rect 4800 3747 4870 3833
rect 4900 3747 4970 3833
rect 5000 3807 5070 3833
rect 5000 3773 5018 3807
rect 5052 3773 5070 3807
rect 5000 3747 5070 3773
rect 5100 3807 5170 3833
rect 5100 3773 5118 3807
rect 5152 3773 5170 3807
rect 5100 3747 5170 3773
rect 5200 3747 5270 3833
rect 5300 3807 5370 3833
rect 5300 3773 5318 3807
rect 5352 3773 5370 3807
rect 5300 3747 5370 3773
rect 5400 3807 5454 3833
rect 5400 3773 5412 3807
rect 5446 3773 5454 3807
rect 5400 3747 5454 3773
rect 3216 3577 3270 3603
rect 3216 3543 3224 3577
rect 3258 3543 3270 3577
rect 3216 3517 3270 3543
rect 3300 3577 3370 3603
rect 3300 3543 3318 3577
rect 3352 3543 3370 3577
rect 3300 3517 3370 3543
rect 3400 3517 3470 3603
rect 3500 3577 3570 3603
rect 3500 3543 3518 3577
rect 3552 3543 3570 3577
rect 3500 3517 3570 3543
rect 3600 3577 3670 3603
rect 3600 3543 3618 3577
rect 3652 3543 3670 3577
rect 3600 3517 3670 3543
rect 3700 3577 3770 3603
rect 3700 3543 3718 3577
rect 3752 3543 3770 3577
rect 3700 3517 3770 3543
rect 3800 3517 3870 3603
rect 3900 3517 3970 3603
rect 4000 3577 4070 3603
rect 4000 3543 4018 3577
rect 4052 3543 4070 3577
rect 4000 3517 4070 3543
rect 4100 3577 4170 3603
rect 4100 3543 4118 3577
rect 4152 3543 4170 3577
rect 4100 3517 4170 3543
rect 4200 3517 4270 3603
rect 4300 3577 4370 3603
rect 4300 3543 4318 3577
rect 4352 3543 4370 3577
rect 4300 3517 4370 3543
rect 4400 3577 4454 3603
rect 4400 3543 4412 3577
rect 4446 3543 4454 3577
rect 4400 3517 4454 3543
rect 1016 3437 1070 3463
rect 1016 3403 1024 3437
rect 1058 3403 1070 3437
rect 1016 3377 1070 3403
rect 1100 3437 1170 3463
rect 1100 3403 1118 3437
rect 1152 3403 1170 3437
rect 1100 3377 1170 3403
rect 1200 3437 1270 3463
rect 1200 3403 1218 3437
rect 1252 3403 1270 3437
rect 1200 3377 1270 3403
rect 1300 3377 1370 3463
rect 1400 3437 1470 3463
rect 1400 3403 1418 3437
rect 1452 3403 1470 3437
rect 1400 3377 1470 3403
rect 1500 3437 1570 3463
rect 1500 3403 1518 3437
rect 1552 3403 1570 3437
rect 1500 3377 1570 3403
rect 1600 3437 1670 3463
rect 1600 3403 1618 3437
rect 1652 3403 1670 3437
rect 1600 3377 1670 3403
rect 1700 3437 1770 3463
rect 1700 3403 1718 3437
rect 1752 3403 1770 3437
rect 1700 3377 1770 3403
rect 1800 3437 1870 3463
rect 1800 3403 1818 3437
rect 1852 3403 1870 3437
rect 1800 3377 1870 3403
rect 1900 3437 1970 3463
rect 1900 3403 1918 3437
rect 1952 3403 1970 3437
rect 1900 3377 1970 3403
rect 2000 3437 2070 3463
rect 2000 3403 2018 3437
rect 2052 3403 2070 3437
rect 2000 3377 2070 3403
rect 2100 3437 2170 3463
rect 2100 3403 2118 3437
rect 2152 3403 2170 3437
rect 2100 3377 2170 3403
rect 2200 3377 2270 3463
rect 2300 3377 2370 3463
rect 2400 3377 2470 3463
rect 2500 3437 2570 3463
rect 2500 3403 2518 3437
rect 2552 3403 2570 3437
rect 2500 3377 2570 3403
rect 2600 3437 2670 3463
rect 2600 3403 2618 3437
rect 2652 3403 2670 3437
rect 2600 3377 2670 3403
rect 2700 3437 2770 3463
rect 2700 3403 2718 3437
rect 2752 3403 2770 3437
rect 2700 3377 2770 3403
rect 2800 3377 2870 3463
rect 2900 3377 2970 3463
rect 3000 3437 3070 3463
rect 3000 3403 3018 3437
rect 3052 3403 3070 3437
rect 3000 3377 3070 3403
rect 3100 3437 3170 3463
rect 3100 3403 3118 3437
rect 3152 3403 3170 3437
rect 3100 3377 3170 3403
rect 3200 3377 3270 3463
rect 3300 3377 3370 3463
rect 3400 3377 3470 3463
rect 3500 3377 3570 3463
rect 3600 3437 3670 3463
rect 3600 3403 3618 3437
rect 3652 3403 3670 3437
rect 3600 3377 3670 3403
rect 3700 3437 3770 3463
rect 3700 3403 3718 3437
rect 3752 3403 3770 3437
rect 3700 3377 3770 3403
rect 3800 3437 3854 3463
rect 3800 3403 3812 3437
rect 3846 3403 3854 3437
rect 3800 3377 3854 3403
rect 1016 3297 1070 3323
rect 1016 3263 1024 3297
rect 1058 3263 1070 3297
rect 1016 3237 1070 3263
rect 1100 3297 1170 3323
rect 1100 3263 1118 3297
rect 1152 3263 1170 3297
rect 1100 3237 1170 3263
rect 1200 3297 1270 3323
rect 1200 3263 1218 3297
rect 1252 3263 1270 3297
rect 1200 3237 1270 3263
rect 1300 3297 1370 3323
rect 1300 3263 1318 3297
rect 1352 3263 1370 3297
rect 1300 3237 1370 3263
rect 1400 3297 1470 3323
rect 1400 3263 1418 3297
rect 1452 3263 1470 3297
rect 1400 3237 1470 3263
rect 1500 3297 1570 3323
rect 1500 3263 1518 3297
rect 1552 3263 1570 3297
rect 1500 3237 1570 3263
rect 1600 3297 1670 3323
rect 1600 3263 1618 3297
rect 1652 3263 1670 3297
rect 1600 3237 1670 3263
rect 1700 3297 1770 3323
rect 1700 3263 1718 3297
rect 1752 3263 1770 3297
rect 1700 3237 1770 3263
rect 1800 3297 1870 3323
rect 1800 3263 1818 3297
rect 1852 3263 1870 3297
rect 1800 3237 1870 3263
rect 1900 3297 1970 3323
rect 1900 3263 1918 3297
rect 1952 3263 1970 3297
rect 1900 3237 1970 3263
rect 2000 3297 2070 3323
rect 2000 3263 2018 3297
rect 2052 3263 2070 3297
rect 2000 3237 2070 3263
rect 2100 3297 2170 3323
rect 2100 3263 2118 3297
rect 2152 3263 2170 3297
rect 2100 3237 2170 3263
rect 2200 3297 2270 3323
rect 2200 3263 2218 3297
rect 2252 3263 2270 3297
rect 2200 3237 2270 3263
rect 2300 3297 2370 3323
rect 2300 3263 2318 3297
rect 2352 3263 2370 3297
rect 2300 3237 2370 3263
rect 2400 3297 2470 3323
rect 2400 3263 2418 3297
rect 2452 3263 2470 3297
rect 2400 3237 2470 3263
rect 2500 3237 2570 3323
rect 2600 3297 2670 3323
rect 2600 3263 2618 3297
rect 2652 3263 2670 3297
rect 2600 3237 2670 3263
rect 2700 3297 2754 3323
rect 2700 3263 2712 3297
rect 2746 3263 2754 3297
rect 2700 3237 2754 3263
rect 216 3157 270 3183
rect 216 3123 224 3157
rect 258 3123 270 3157
rect 216 3097 270 3123
rect 300 3157 370 3183
rect 300 3123 318 3157
rect 352 3123 370 3157
rect 300 3097 370 3123
rect 400 3157 470 3183
rect 400 3123 418 3157
rect 452 3123 470 3157
rect 400 3097 470 3123
rect 500 3157 570 3183
rect 500 3123 518 3157
rect 552 3123 570 3157
rect 500 3097 570 3123
rect 600 3157 670 3183
rect 600 3123 618 3157
rect 652 3123 670 3157
rect 600 3097 670 3123
rect 700 3097 770 3183
rect 800 3157 870 3183
rect 800 3123 818 3157
rect 852 3123 870 3157
rect 800 3097 870 3123
rect 900 3157 970 3183
rect 900 3123 918 3157
rect 952 3123 970 3157
rect 900 3097 970 3123
rect 1000 3097 1070 3183
rect 1100 3097 1170 3183
rect 1200 3157 1270 3183
rect 1200 3123 1218 3157
rect 1252 3123 1270 3157
rect 1200 3097 1270 3123
rect 1300 3157 1354 3183
rect 1300 3123 1312 3157
rect 1346 3123 1354 3157
rect 1300 3097 1354 3123
rect 16 2957 70 3043
rect 100 3017 170 3043
rect 100 2983 118 3017
rect 152 2983 170 3017
rect 100 2957 170 2983
rect 200 3017 270 3043
rect 200 2983 218 3017
rect 252 2983 270 3017
rect 200 2957 270 2983
rect 300 2957 370 3043
rect 400 3017 470 3043
rect 400 2983 418 3017
rect 452 2983 470 3017
rect 400 2957 470 2983
rect 500 3017 570 3043
rect 500 2983 518 3017
rect 552 2983 570 3017
rect 500 2957 570 2983
rect 600 3017 654 3043
rect 600 2983 612 3017
rect 646 2983 654 3017
rect 600 2957 654 2983
rect 1416 3157 1470 3183
rect 1416 3123 1424 3157
rect 1458 3123 1470 3157
rect 1416 3097 1470 3123
rect 1500 3157 1570 3183
rect 1500 3123 1518 3157
rect 1552 3123 1570 3157
rect 1500 3097 1570 3123
rect 1600 3097 1670 3183
rect 1700 3157 1770 3183
rect 1700 3123 1718 3157
rect 1752 3123 1770 3157
rect 1700 3097 1770 3123
rect 1800 3157 1870 3183
rect 1800 3123 1818 3157
rect 1852 3123 1870 3157
rect 1800 3097 1870 3123
rect 1900 3097 1970 3183
rect 2000 3157 2070 3183
rect 2000 3123 2018 3157
rect 2052 3123 2070 3157
rect 2000 3097 2070 3123
rect 2100 3157 2170 3183
rect 2100 3123 2118 3157
rect 2152 3123 2170 3157
rect 2100 3097 2170 3123
rect 2200 3097 2270 3183
rect 2300 3157 2370 3183
rect 2300 3123 2318 3157
rect 2352 3123 2370 3157
rect 2300 3097 2370 3123
rect 2400 3157 2470 3183
rect 2400 3123 2418 3157
rect 2452 3123 2470 3157
rect 2400 3097 2470 3123
rect 2500 3157 2554 3183
rect 2500 3123 2512 3157
rect 2546 3123 2554 3157
rect 2500 3097 2554 3123
rect 716 3017 770 3043
rect 716 2983 724 3017
rect 758 2983 770 3017
rect 716 2957 770 2983
rect 800 3017 870 3043
rect 800 2983 818 3017
rect 852 2983 870 3017
rect 800 2957 870 2983
rect 900 3017 970 3043
rect 900 2983 918 3017
rect 952 2983 970 3017
rect 900 2957 970 2983
rect 1000 2957 1070 3043
rect 1100 2957 1170 3043
rect 1200 3017 1270 3043
rect 1200 2983 1218 3017
rect 1252 2983 1270 3017
rect 1200 2957 1270 2983
rect 1300 3017 1370 3043
rect 1300 2983 1318 3017
rect 1352 2983 1370 3017
rect 1300 2957 1370 2983
rect 1400 2957 1470 3043
rect 1500 2957 1570 3043
rect 1600 2957 1670 3043
rect 1700 2957 1770 3043
rect 1800 3017 1870 3043
rect 1800 2983 1818 3017
rect 1852 2983 1870 3017
rect 1800 2957 1870 2983
rect 1900 3017 1970 3043
rect 1900 2983 1918 3017
rect 1952 2983 1970 3017
rect 1900 2957 1970 2983
rect 2000 3017 2054 3043
rect 2000 2983 2012 3017
rect 2046 2983 2054 3017
rect 2000 2957 2054 2983
rect 16 2877 70 2903
rect 16 2843 24 2877
rect 58 2843 70 2877
rect 16 2817 70 2843
rect 100 2877 170 2903
rect 100 2843 118 2877
rect 152 2843 170 2877
rect 100 2817 170 2843
rect 200 2877 270 2903
rect 200 2843 218 2877
rect 252 2843 270 2877
rect 200 2817 270 2843
rect 300 2817 370 2903
rect 400 2877 470 2903
rect 400 2843 418 2877
rect 452 2843 470 2877
rect 400 2817 470 2843
rect 500 2877 570 2903
rect 500 2843 518 2877
rect 552 2843 570 2877
rect 500 2817 570 2843
rect 600 2877 670 2903
rect 600 2843 618 2877
rect 652 2843 670 2877
rect 600 2817 670 2843
rect 700 2877 770 2903
rect 700 2843 718 2877
rect 752 2843 770 2877
rect 700 2817 770 2843
rect 800 2877 854 2903
rect 800 2843 812 2877
rect 846 2843 854 2877
rect 800 2817 854 2843
rect 2816 3297 2870 3323
rect 2816 3263 2824 3297
rect 2858 3263 2870 3297
rect 2816 3237 2870 3263
rect 2900 3297 2970 3323
rect 2900 3263 2918 3297
rect 2952 3263 2970 3297
rect 2900 3237 2970 3263
rect 3000 3297 3070 3323
rect 3000 3263 3018 3297
rect 3052 3263 3070 3297
rect 3000 3237 3070 3263
rect 3100 3297 3170 3323
rect 3100 3263 3118 3297
rect 3152 3263 3170 3297
rect 3100 3237 3170 3263
rect 3200 3297 3254 3323
rect 3200 3263 3212 3297
rect 3246 3263 3254 3297
rect 3200 3237 3254 3263
rect 2616 3157 2670 3183
rect 2616 3123 2624 3157
rect 2658 3123 2670 3157
rect 2616 3097 2670 3123
rect 2700 3157 2770 3183
rect 2700 3123 2718 3157
rect 2752 3123 2770 3157
rect 2700 3097 2770 3123
rect 2800 3157 2870 3183
rect 2800 3123 2818 3157
rect 2852 3123 2870 3157
rect 2800 3097 2870 3123
rect 2900 3157 2970 3183
rect 2900 3123 2918 3157
rect 2952 3123 2970 3157
rect 2900 3097 2970 3123
rect 3000 3097 3070 3183
rect 3100 3157 3170 3183
rect 3100 3123 3118 3157
rect 3152 3123 3170 3157
rect 3100 3097 3170 3123
rect 3200 3157 3254 3183
rect 3200 3123 3212 3157
rect 3246 3123 3254 3157
rect 3200 3097 3254 3123
rect 2116 3017 2170 3043
rect 2116 2983 2124 3017
rect 2158 2983 2170 3017
rect 2116 2957 2170 2983
rect 2200 3017 2270 3043
rect 2200 2983 2218 3017
rect 2252 2983 2270 3017
rect 2200 2957 2270 2983
rect 2300 2957 2370 3043
rect 2400 3017 2470 3043
rect 2400 2983 2418 3017
rect 2452 2983 2470 3017
rect 2400 2957 2470 2983
rect 2500 3017 2570 3043
rect 2500 2983 2518 3017
rect 2552 2983 2570 3017
rect 2500 2957 2570 2983
rect 2600 2957 2670 3043
rect 2700 3017 2770 3043
rect 2700 2983 2718 3017
rect 2752 2983 2770 3017
rect 2700 2957 2770 2983
rect 2800 3017 2870 3043
rect 2800 2983 2818 3017
rect 2852 2983 2870 3017
rect 2800 2957 2870 2983
rect 2900 3017 2970 3043
rect 2900 2983 2918 3017
rect 2952 2983 2970 3017
rect 2900 2957 2970 2983
rect 3000 3017 3054 3043
rect 3000 2983 3012 3017
rect 3046 2983 3054 3017
rect 3000 2957 3054 2983
rect 916 2877 970 2903
rect 916 2843 924 2877
rect 958 2843 970 2877
rect 916 2817 970 2843
rect 1000 2877 1070 2903
rect 1000 2843 1018 2877
rect 1052 2843 1070 2877
rect 1000 2817 1070 2843
rect 1100 2877 1170 2903
rect 1100 2843 1118 2877
rect 1152 2843 1170 2877
rect 1100 2817 1170 2843
rect 1200 2817 1270 2903
rect 1300 2877 1370 2903
rect 1300 2843 1318 2877
rect 1352 2843 1370 2877
rect 1300 2817 1370 2843
rect 1400 2877 1470 2903
rect 1400 2843 1418 2877
rect 1452 2843 1470 2877
rect 1400 2817 1470 2843
rect 1500 2817 1570 2903
rect 1600 2817 1670 2903
rect 1700 2817 1770 2903
rect 1800 2877 1870 2903
rect 1800 2843 1818 2877
rect 1852 2843 1870 2877
rect 1800 2817 1870 2843
rect 1900 2877 1970 2903
rect 1900 2843 1918 2877
rect 1952 2843 1970 2877
rect 1900 2817 1970 2843
rect 2000 2877 2070 2903
rect 2000 2843 2018 2877
rect 2052 2843 2070 2877
rect 2000 2817 2070 2843
rect 2100 2817 2170 2903
rect 2200 2817 2270 2903
rect 2300 2817 2370 2903
rect 2400 2817 2470 2903
rect 2500 2877 2570 2903
rect 2500 2843 2518 2877
rect 2552 2843 2570 2877
rect 2500 2817 2570 2843
rect 2600 2877 2654 2903
rect 2600 2843 2612 2877
rect 2646 2843 2654 2877
rect 2600 2817 2654 2843
rect 16 2677 70 2763
rect 100 2677 170 2763
rect 200 2737 270 2763
rect 200 2703 218 2737
rect 252 2703 270 2737
rect 200 2677 270 2703
rect 300 2737 370 2763
rect 300 2703 318 2737
rect 352 2703 370 2737
rect 300 2677 370 2703
rect 400 2737 470 2763
rect 400 2703 418 2737
rect 452 2703 470 2737
rect 400 2677 470 2703
rect 500 2737 570 2763
rect 500 2703 518 2737
rect 552 2703 570 2737
rect 500 2677 570 2703
rect 600 2677 670 2763
rect 700 2677 770 2763
rect 800 2677 870 2763
rect 900 2677 970 2763
rect 1000 2737 1070 2763
rect 1000 2703 1018 2737
rect 1052 2703 1070 2737
rect 1000 2677 1070 2703
rect 1100 2737 1154 2763
rect 1100 2703 1112 2737
rect 1146 2703 1154 2737
rect 1100 2677 1154 2703
rect 1216 2737 1270 2763
rect 1216 2703 1224 2737
rect 1258 2703 1270 2737
rect 1216 2677 1270 2703
rect 1300 2737 1370 2763
rect 1300 2703 1318 2737
rect 1352 2703 1370 2737
rect 1300 2677 1370 2703
rect 1400 2677 1470 2763
rect 1500 2677 1570 2763
rect 1600 2677 1670 2763
rect 1700 2677 1770 2763
rect 1800 2737 1870 2763
rect 1800 2703 1818 2737
rect 1852 2703 1870 2737
rect 1800 2677 1870 2703
rect 1900 2737 1970 2763
rect 1900 2703 1918 2737
rect 1952 2703 1970 2737
rect 1900 2677 1970 2703
rect 2000 2677 2070 2763
rect 2100 2677 2170 2763
rect 2200 2737 2270 2763
rect 2200 2703 2218 2737
rect 2252 2703 2270 2737
rect 2200 2677 2270 2703
rect 2300 2737 2354 2763
rect 2300 2703 2312 2737
rect 2346 2703 2354 2737
rect 2300 2677 2354 2703
rect 2716 2877 2770 2903
rect 2716 2843 2724 2877
rect 2758 2843 2770 2877
rect 2716 2817 2770 2843
rect 2800 2877 2870 2903
rect 2800 2843 2818 2877
rect 2852 2843 2870 2877
rect 2800 2817 2870 2843
rect 2900 2877 2954 2903
rect 2900 2843 2912 2877
rect 2946 2843 2954 2877
rect 2900 2817 2954 2843
rect 3316 3297 3370 3323
rect 3316 3263 3324 3297
rect 3358 3263 3370 3297
rect 3316 3237 3370 3263
rect 3400 3297 3454 3323
rect 3400 3263 3412 3297
rect 3446 3263 3454 3297
rect 3400 3237 3454 3263
rect 3916 3437 3970 3463
rect 3916 3403 3924 3437
rect 3958 3403 3970 3437
rect 3916 3377 3970 3403
rect 4000 3437 4070 3463
rect 4000 3403 4018 3437
rect 4052 3403 4070 3437
rect 4000 3377 4070 3403
rect 4100 3437 4170 3463
rect 4100 3403 4118 3437
rect 4152 3403 4170 3437
rect 4100 3377 4170 3403
rect 4200 3437 4270 3463
rect 4200 3403 4218 3437
rect 4252 3403 4270 3437
rect 4200 3377 4270 3403
rect 4300 3437 4370 3463
rect 4300 3403 4318 3437
rect 4352 3403 4370 3437
rect 4300 3377 4370 3403
rect 4400 3437 4454 3463
rect 4400 3403 4412 3437
rect 4446 3403 4454 3437
rect 4400 3377 4454 3403
rect 6516 4787 6570 4813
rect 6516 4753 6524 4787
rect 6558 4753 6570 4787
rect 6516 4727 6570 4753
rect 6600 4787 6670 4813
rect 6600 4753 6618 4787
rect 6652 4753 6670 4787
rect 6600 4727 6670 4753
rect 6700 4787 6770 4813
rect 6700 4753 6718 4787
rect 6752 4753 6770 4787
rect 6700 4727 6770 4753
rect 6800 4727 6870 4813
rect 6900 4727 6970 4813
rect 7000 4787 7070 4813
rect 7000 4753 7018 4787
rect 7052 4753 7070 4787
rect 7000 4727 7070 4753
rect 7100 4787 7170 4813
rect 7100 4753 7118 4787
rect 7152 4753 7170 4787
rect 7100 4727 7170 4753
rect 7200 4727 7270 4813
rect 7300 4787 7370 4813
rect 7300 4753 7318 4787
rect 7352 4753 7370 4787
rect 7300 4727 7370 4753
rect 7400 4787 7470 4813
rect 7400 4753 7418 4787
rect 7452 4753 7470 4787
rect 7400 4727 7470 4753
rect 7500 4787 7570 4813
rect 7500 4753 7518 4787
rect 7552 4753 7570 4787
rect 7500 4727 7570 4753
rect 7600 4787 7670 4813
rect 7600 4753 7618 4787
rect 7652 4753 7670 4787
rect 7600 4727 7670 4753
rect 7700 4787 7770 4813
rect 7700 4753 7718 4787
rect 7752 4753 7770 4787
rect 7700 4727 7770 4753
rect 7800 4787 7870 4813
rect 7800 4753 7818 4787
rect 7852 4753 7870 4787
rect 7800 4727 7870 4753
rect 7900 4727 7970 4813
rect 8000 4727 8070 4813
rect 8100 4787 8170 4813
rect 8100 4753 8118 4787
rect 8152 4753 8170 4787
rect 8100 4727 8170 4753
rect 8200 4787 8270 4813
rect 8200 4753 8218 4787
rect 8252 4753 8270 4787
rect 8200 4727 8270 4753
rect 8300 4787 8370 4813
rect 8300 4753 8318 4787
rect 8352 4753 8370 4787
rect 8300 4727 8370 4753
rect 8400 4787 8470 4813
rect 8400 4753 8418 4787
rect 8452 4753 8470 4787
rect 8400 4727 8470 4753
rect 8500 4727 8570 4813
rect 8600 4727 8670 4813
rect 8700 4727 8770 4813
rect 8800 4787 8870 4813
rect 8800 4753 8818 4787
rect 8852 4753 8870 4787
rect 8800 4727 8870 4753
rect 8900 4787 8970 4813
rect 8900 4753 8918 4787
rect 8952 4753 8970 4787
rect 8900 4727 8970 4753
rect 9000 4727 9070 4813
rect 9100 4727 9170 4813
rect 9200 4727 9270 4813
rect 9300 4727 9370 4813
rect 9400 4727 9470 4813
rect 9500 4727 9570 4813
rect 9600 4727 9670 4813
rect 9700 4787 9770 4813
rect 9700 4753 9718 4787
rect 9752 4753 9770 4787
rect 9700 4727 9770 4753
rect 9800 4787 9854 4813
rect 9800 4753 9812 4787
rect 9846 4753 9854 4787
rect 9800 4727 9854 4753
rect 6516 4647 6570 4673
rect 6516 4613 6524 4647
rect 6558 4613 6570 4647
rect 6516 4587 6570 4613
rect 6600 4647 6670 4673
rect 6600 4613 6618 4647
rect 6652 4613 6670 4647
rect 6600 4587 6670 4613
rect 6700 4647 6770 4673
rect 6700 4613 6718 4647
rect 6752 4613 6770 4647
rect 6700 4587 6770 4613
rect 6800 4647 6870 4673
rect 6800 4613 6818 4647
rect 6852 4613 6870 4647
rect 6800 4587 6870 4613
rect 6900 4647 6970 4673
rect 6900 4613 6918 4647
rect 6952 4613 6970 4647
rect 6900 4587 6970 4613
rect 7000 4647 7070 4673
rect 7000 4613 7018 4647
rect 7052 4613 7070 4647
rect 7000 4587 7070 4613
rect 7100 4647 7170 4673
rect 7100 4613 7118 4647
rect 7152 4613 7170 4647
rect 7100 4587 7170 4613
rect 7200 4647 7270 4673
rect 7200 4613 7218 4647
rect 7252 4613 7270 4647
rect 7200 4587 7270 4613
rect 7300 4587 7370 4673
rect 7400 4587 7470 4673
rect 7500 4587 7570 4673
rect 7600 4587 7670 4673
rect 7700 4587 7770 4673
rect 7800 4587 7870 4673
rect 7900 4647 7970 4673
rect 7900 4613 7918 4647
rect 7952 4613 7970 4647
rect 7900 4587 7970 4613
rect 8000 4647 8070 4673
rect 8000 4613 8018 4647
rect 8052 4613 8070 4647
rect 8000 4587 8070 4613
rect 8100 4647 8170 4673
rect 8100 4613 8118 4647
rect 8152 4613 8170 4647
rect 8100 4587 8170 4613
rect 8200 4647 8270 4673
rect 8200 4613 8218 4647
rect 8252 4613 8270 4647
rect 8200 4587 8270 4613
rect 8300 4647 8370 4673
rect 8300 4613 8318 4647
rect 8352 4613 8370 4647
rect 8300 4587 8370 4613
rect 8400 4587 8470 4673
rect 8500 4587 8570 4673
rect 8600 4647 8670 4673
rect 8600 4613 8618 4647
rect 8652 4613 8670 4647
rect 8600 4587 8670 4613
rect 8700 4647 8754 4673
rect 8700 4613 8712 4647
rect 8746 4613 8754 4647
rect 8700 4587 8754 4613
rect 6116 4507 6170 4533
rect 6116 4473 6124 4507
rect 6158 4473 6170 4507
rect 6116 4447 6170 4473
rect 6200 4507 6270 4533
rect 6200 4473 6218 4507
rect 6252 4473 6270 4507
rect 6200 4447 6270 4473
rect 6300 4447 6370 4533
rect 6400 4447 6470 4533
rect 6500 4447 6570 4533
rect 6600 4447 6670 4533
rect 6700 4447 6770 4533
rect 6800 4447 6870 4533
rect 6900 4447 6970 4533
rect 7000 4507 7070 4533
rect 7000 4473 7018 4507
rect 7052 4473 7070 4507
rect 7000 4447 7070 4473
rect 7100 4507 7170 4533
rect 7100 4473 7118 4507
rect 7152 4473 7170 4507
rect 7100 4447 7170 4473
rect 7200 4507 7270 4533
rect 7200 4473 7218 4507
rect 7252 4473 7270 4507
rect 7200 4447 7270 4473
rect 7300 4447 7370 4533
rect 7400 4447 7470 4533
rect 7500 4447 7570 4533
rect 7600 4447 7670 4533
rect 7700 4507 7770 4533
rect 7700 4473 7718 4507
rect 7752 4473 7770 4507
rect 7700 4447 7770 4473
rect 7800 4507 7870 4533
rect 7800 4473 7818 4507
rect 7852 4473 7870 4507
rect 7800 4447 7870 4473
rect 7900 4507 7970 4533
rect 7900 4473 7918 4507
rect 7952 4473 7970 4507
rect 7900 4447 7970 4473
rect 8000 4507 8054 4533
rect 8000 4473 8012 4507
rect 8046 4473 8054 4507
rect 8000 4447 8054 4473
rect 6116 4367 6170 4393
rect 6116 4333 6124 4367
rect 6158 4333 6170 4367
rect 6116 4307 6170 4333
rect 6200 4367 6270 4393
rect 6200 4333 6218 4367
rect 6252 4333 6270 4367
rect 6200 4307 6270 4333
rect 6300 4307 6370 4393
rect 6400 4367 6470 4393
rect 6400 4333 6418 4367
rect 6452 4333 6470 4367
rect 6400 4307 6470 4333
rect 6500 4367 6570 4393
rect 6500 4333 6518 4367
rect 6552 4333 6570 4367
rect 6500 4307 6570 4333
rect 6600 4367 6654 4393
rect 6600 4333 6612 4367
rect 6646 4333 6654 4367
rect 6600 4307 6654 4333
rect 6116 4227 6170 4253
rect 6116 4193 6124 4227
rect 6158 4193 6170 4227
rect 6116 4167 6170 4193
rect 6200 4227 6254 4253
rect 6200 4193 6212 4227
rect 6246 4193 6254 4227
rect 6200 4167 6254 4193
rect 6316 4227 6370 4253
rect 6316 4193 6324 4227
rect 6358 4193 6370 4227
rect 6316 4167 6370 4193
rect 6400 4227 6454 4253
rect 6400 4193 6412 4227
rect 6446 4193 6454 4227
rect 6400 4167 6454 4193
rect 6516 4227 6570 4253
rect 6516 4193 6524 4227
rect 6558 4193 6570 4227
rect 6516 4167 6570 4193
rect 6600 4227 6654 4253
rect 6600 4193 6612 4227
rect 6646 4193 6654 4227
rect 6600 4167 6654 4193
rect 6716 4367 6770 4393
rect 6716 4333 6724 4367
rect 6758 4333 6770 4367
rect 6716 4307 6770 4333
rect 6800 4367 6870 4393
rect 6800 4333 6818 4367
rect 6852 4333 6870 4367
rect 6800 4307 6870 4333
rect 6900 4307 6970 4393
rect 7000 4307 7070 4393
rect 7100 4367 7170 4393
rect 7100 4333 7118 4367
rect 7152 4333 7170 4367
rect 7100 4307 7170 4333
rect 7200 4367 7270 4393
rect 7200 4333 7218 4367
rect 7252 4333 7270 4367
rect 7200 4307 7270 4333
rect 7300 4367 7354 4393
rect 7300 4333 7312 4367
rect 7346 4333 7354 4367
rect 7300 4307 7354 4333
rect 6716 4227 6770 4253
rect 6716 4193 6724 4227
rect 6758 4193 6770 4227
rect 6716 4167 6770 4193
rect 6800 4227 6870 4253
rect 6800 4193 6818 4227
rect 6852 4193 6870 4227
rect 6800 4167 6870 4193
rect 6900 4167 6970 4253
rect 7000 4227 7070 4253
rect 7000 4193 7018 4227
rect 7052 4193 7070 4227
rect 7000 4167 7070 4193
rect 7100 4227 7154 4253
rect 7100 4193 7112 4227
rect 7146 4193 7154 4227
rect 7100 4167 7154 4193
rect 8116 4507 8170 4533
rect 8116 4473 8124 4507
rect 8158 4473 8170 4507
rect 8116 4447 8170 4473
rect 8200 4507 8270 4533
rect 8200 4473 8218 4507
rect 8252 4473 8270 4507
rect 8200 4447 8270 4473
rect 8300 4507 8354 4533
rect 8300 4473 8312 4507
rect 8346 4473 8354 4507
rect 8300 4447 8354 4473
rect 9916 4787 9970 4813
rect 9916 4753 9924 4787
rect 9958 4753 9970 4787
rect 9916 4727 9970 4753
rect 10000 4787 10070 4813
rect 10000 4753 10018 4787
rect 10052 4753 10070 4787
rect 10000 4727 10070 4753
rect 10100 4787 10170 4813
rect 10100 4753 10118 4787
rect 10152 4753 10170 4787
rect 10100 4727 10170 4753
rect 10200 4727 10270 4813
rect 10300 4727 10370 4813
rect 10400 4787 10470 4813
rect 10400 4753 10418 4787
rect 10452 4753 10470 4787
rect 10400 4727 10470 4753
rect 10500 4787 10570 4813
rect 10500 4753 10518 4787
rect 10552 4753 10570 4787
rect 10500 4727 10570 4753
rect 10600 4787 10670 4813
rect 10600 4753 10618 4787
rect 10652 4753 10670 4787
rect 10600 4727 10670 4753
rect 10700 4787 10754 4813
rect 10700 4753 10712 4787
rect 10746 4753 10754 4787
rect 10700 4727 10754 4753
rect 10816 4787 10870 4813
rect 10816 4753 10824 4787
rect 10858 4753 10870 4787
rect 10816 4727 10870 4753
rect 10900 4787 10970 4813
rect 10900 4753 10918 4787
rect 10952 4753 10970 4787
rect 10900 4727 10970 4753
rect 11000 4727 11070 4813
rect 11100 4787 11170 4813
rect 11100 4753 11118 4787
rect 11152 4753 11170 4787
rect 11100 4727 11170 4753
rect 11200 4787 11270 4813
rect 11200 4753 11218 4787
rect 11252 4753 11270 4787
rect 11200 4727 11270 4753
rect 11300 4787 11370 4813
rect 11300 4753 11318 4787
rect 11352 4753 11370 4787
rect 11300 4727 11370 4753
rect 11400 4727 11470 4813
rect 11500 4787 11570 4813
rect 11500 4753 11518 4787
rect 11552 4753 11570 4787
rect 11500 4727 11570 4753
rect 11600 4787 11654 4813
rect 11600 4753 11612 4787
rect 11646 4753 11654 4787
rect 11600 4727 11654 4753
rect 11716 4787 11770 4813
rect 11716 4753 11724 4787
rect 11758 4753 11770 4787
rect 11716 4727 11770 4753
rect 11800 4787 11870 4813
rect 11800 4753 11818 4787
rect 11852 4753 11870 4787
rect 11800 4727 11870 4753
rect 11900 4787 11970 4813
rect 11900 4753 11918 4787
rect 11952 4753 11970 4787
rect 11900 4727 11970 4753
rect 12000 4727 12070 4813
rect 12100 4787 12170 4813
rect 12100 4753 12118 4787
rect 12152 4753 12170 4787
rect 12100 4727 12170 4753
rect 12200 4787 12270 4813
rect 12200 4753 12218 4787
rect 12252 4753 12270 4787
rect 12200 4727 12270 4753
rect 12300 4787 12370 4813
rect 12300 4753 12318 4787
rect 12352 4753 12370 4787
rect 12300 4727 12370 4753
rect 12400 4787 12454 4813
rect 12400 4753 12412 4787
rect 12446 4753 12454 4787
rect 12400 4727 12454 4753
rect 12516 4787 12570 4813
rect 12516 4753 12524 4787
rect 12558 4753 12570 4787
rect 12516 4727 12570 4753
rect 12600 4787 12670 4813
rect 12600 4753 12618 4787
rect 12652 4753 12670 4787
rect 12600 4727 12670 4753
rect 12700 4787 12770 4813
rect 12700 4753 12718 4787
rect 12752 4753 12770 4787
rect 12700 4727 12770 4753
rect 12800 4787 12854 4813
rect 12800 4753 12812 4787
rect 12846 4753 12854 4787
rect 12800 4727 12854 4753
rect 12912 4802 12970 4813
rect 12912 4768 12924 4802
rect 12958 4768 12970 4802
rect 12912 4727 12970 4768
rect 13000 4787 13070 4813
rect 13000 4753 13018 4787
rect 13052 4753 13070 4787
rect 13000 4727 13070 4753
rect 13100 4772 13158 4813
rect 13100 4738 13112 4772
rect 13146 4738 13158 4772
rect 13100 4727 13158 4738
rect 13220 4787 13280 4813
rect 13220 4753 13228 4787
rect 13262 4753 13280 4787
rect 13220 4727 13280 4753
rect 13310 4787 13380 4813
rect 13310 4753 13328 4787
rect 13362 4753 13380 4787
rect 13310 4727 13380 4753
rect 13410 4787 13480 4813
rect 13410 4753 13428 4787
rect 13462 4753 13480 4787
rect 13410 4727 13480 4753
rect 13510 4787 13580 4813
rect 13510 4753 13528 4787
rect 13562 4753 13580 4787
rect 13510 4727 13580 4753
rect 13610 4787 13670 4813
rect 13610 4753 13628 4787
rect 13662 4753 13670 4787
rect 13610 4727 13670 4753
rect 8816 4647 8870 4673
rect 8816 4613 8824 4647
rect 8858 4613 8870 4647
rect 8816 4587 8870 4613
rect 8900 4647 8970 4673
rect 8900 4613 8918 4647
rect 8952 4613 8970 4647
rect 8900 4587 8970 4613
rect 9000 4587 9070 4673
rect 9100 4587 9170 4673
rect 9200 4587 9270 4673
rect 9300 4647 9370 4673
rect 9300 4613 9318 4647
rect 9352 4613 9370 4647
rect 9300 4587 9370 4613
rect 9400 4647 9470 4673
rect 9400 4613 9418 4647
rect 9452 4613 9470 4647
rect 9400 4587 9470 4613
rect 9500 4647 9570 4673
rect 9500 4613 9518 4647
rect 9552 4613 9570 4647
rect 9500 4587 9570 4613
rect 9600 4647 9670 4673
rect 9600 4613 9618 4647
rect 9652 4613 9670 4647
rect 9600 4587 9670 4613
rect 9700 4647 9770 4673
rect 9700 4613 9718 4647
rect 9752 4613 9770 4647
rect 9700 4587 9770 4613
rect 9800 4587 9870 4673
rect 9900 4647 9970 4673
rect 9900 4613 9918 4647
rect 9952 4613 9970 4647
rect 9900 4587 9970 4613
rect 10000 4647 10070 4673
rect 10000 4613 10018 4647
rect 10052 4613 10070 4647
rect 10000 4587 10070 4613
rect 10100 4647 10170 4673
rect 10100 4613 10118 4647
rect 10152 4613 10170 4647
rect 10100 4587 10170 4613
rect 10200 4587 10270 4673
rect 10300 4587 10370 4673
rect 10400 4587 10470 4673
rect 10500 4647 10570 4673
rect 10500 4613 10518 4647
rect 10552 4613 10570 4647
rect 10500 4587 10570 4613
rect 10600 4647 10670 4673
rect 10600 4613 10618 4647
rect 10652 4613 10670 4647
rect 10600 4587 10670 4613
rect 10700 4587 10770 4673
rect 10800 4587 10870 4673
rect 10900 4587 10970 4673
rect 11000 4587 11070 4673
rect 11100 4647 11170 4673
rect 11100 4613 11118 4647
rect 11152 4613 11170 4647
rect 11100 4587 11170 4613
rect 11200 4647 11270 4673
rect 11200 4613 11218 4647
rect 11252 4613 11270 4647
rect 11200 4587 11270 4613
rect 11300 4587 11370 4673
rect 11400 4647 11470 4673
rect 11400 4613 11418 4647
rect 11452 4613 11470 4647
rect 11400 4587 11470 4613
rect 11500 4647 11570 4673
rect 11500 4613 11518 4647
rect 11552 4613 11570 4647
rect 11500 4587 11570 4613
rect 11600 4647 11670 4673
rect 11600 4613 11618 4647
rect 11652 4613 11670 4647
rect 11600 4587 11670 4613
rect 11700 4647 11770 4673
rect 11700 4613 11718 4647
rect 11752 4613 11770 4647
rect 11700 4587 11770 4613
rect 11800 4647 11870 4673
rect 11800 4613 11818 4647
rect 11852 4613 11870 4647
rect 11800 4587 11870 4613
rect 11900 4647 11970 4673
rect 11900 4613 11918 4647
rect 11952 4613 11970 4647
rect 11900 4587 11970 4613
rect 12000 4587 12070 4673
rect 12100 4587 12170 4673
rect 12200 4587 12270 4673
rect 12300 4647 12370 4673
rect 12300 4613 12318 4647
rect 12352 4613 12370 4647
rect 12300 4587 12370 4613
rect 12400 4647 12470 4673
rect 12400 4613 12418 4647
rect 12452 4613 12470 4647
rect 12400 4587 12470 4613
rect 12500 4647 12570 4673
rect 12500 4613 12518 4647
rect 12552 4613 12570 4647
rect 12500 4587 12570 4613
rect 12600 4647 12654 4673
rect 12600 4613 12612 4647
rect 12646 4613 12654 4647
rect 12600 4587 12654 4613
rect 8416 4507 8470 4533
rect 8416 4473 8424 4507
rect 8458 4473 8470 4507
rect 8416 4447 8470 4473
rect 8500 4507 8570 4533
rect 8500 4473 8518 4507
rect 8552 4473 8570 4507
rect 8500 4447 8570 4473
rect 8600 4507 8670 4533
rect 8600 4473 8618 4507
rect 8652 4473 8670 4507
rect 8600 4447 8670 4473
rect 8700 4507 8770 4533
rect 8700 4473 8718 4507
rect 8752 4473 8770 4507
rect 8700 4447 8770 4473
rect 8800 4507 8854 4533
rect 8800 4473 8812 4507
rect 8846 4473 8854 4507
rect 8800 4447 8854 4473
rect 8916 4507 8970 4533
rect 8916 4473 8924 4507
rect 8958 4473 8970 4507
rect 8916 4447 8970 4473
rect 9000 4507 9054 4533
rect 9000 4473 9012 4507
rect 9046 4473 9054 4507
rect 9000 4447 9054 4473
rect 9116 4507 9170 4533
rect 9116 4473 9124 4507
rect 9158 4473 9170 4507
rect 9116 4447 9170 4473
rect 9200 4507 9270 4533
rect 9200 4473 9218 4507
rect 9252 4473 9270 4507
rect 9200 4447 9270 4473
rect 9300 4507 9354 4533
rect 9300 4473 9312 4507
rect 9346 4473 9354 4507
rect 9300 4447 9354 4473
rect 9416 4507 9470 4533
rect 9416 4473 9424 4507
rect 9458 4473 9470 4507
rect 9416 4447 9470 4473
rect 9500 4507 9570 4533
rect 9500 4473 9518 4507
rect 9552 4473 9570 4507
rect 9500 4447 9570 4473
rect 9600 4507 9654 4533
rect 9600 4473 9612 4507
rect 9646 4473 9654 4507
rect 9600 4447 9654 4473
rect 9716 4507 9770 4533
rect 9716 4473 9724 4507
rect 9758 4473 9770 4507
rect 9716 4447 9770 4473
rect 9800 4507 9870 4533
rect 9800 4473 9818 4507
rect 9852 4473 9870 4507
rect 9800 4447 9870 4473
rect 9900 4507 9954 4533
rect 9900 4473 9912 4507
rect 9946 4473 9954 4507
rect 9900 4447 9954 4473
rect 10016 4507 10070 4533
rect 10016 4473 10024 4507
rect 10058 4473 10070 4507
rect 10016 4447 10070 4473
rect 10100 4507 10170 4533
rect 10100 4473 10118 4507
rect 10152 4473 10170 4507
rect 10100 4447 10170 4473
rect 10200 4507 10254 4533
rect 10200 4473 10212 4507
rect 10246 4473 10254 4507
rect 10200 4447 10254 4473
rect 10316 4507 10370 4533
rect 10316 4473 10324 4507
rect 10358 4473 10370 4507
rect 10316 4447 10370 4473
rect 10400 4507 10470 4533
rect 10400 4473 10418 4507
rect 10452 4473 10470 4507
rect 10400 4447 10470 4473
rect 10500 4507 10554 4533
rect 10500 4473 10512 4507
rect 10546 4473 10554 4507
rect 10500 4447 10554 4473
rect 10616 4507 10670 4533
rect 10616 4473 10624 4507
rect 10658 4473 10670 4507
rect 10616 4447 10670 4473
rect 10700 4507 10754 4533
rect 10700 4473 10712 4507
rect 10746 4473 10754 4507
rect 10700 4447 10754 4473
rect 10816 4507 10870 4533
rect 10816 4473 10824 4507
rect 10858 4473 10870 4507
rect 10816 4447 10870 4473
rect 10900 4507 10954 4533
rect 10900 4473 10912 4507
rect 10946 4473 10954 4507
rect 10900 4447 10954 4473
rect 7416 4367 7470 4393
rect 7416 4333 7424 4367
rect 7458 4333 7470 4367
rect 7416 4307 7470 4333
rect 7500 4367 7570 4393
rect 7500 4333 7518 4367
rect 7552 4333 7570 4367
rect 7500 4307 7570 4333
rect 7600 4367 7670 4393
rect 7600 4333 7618 4367
rect 7652 4333 7670 4367
rect 7600 4307 7670 4333
rect 7700 4367 7770 4393
rect 7700 4333 7718 4367
rect 7752 4333 7770 4367
rect 7700 4307 7770 4333
rect 7800 4307 7870 4393
rect 7900 4307 7970 4393
rect 8000 4367 8070 4393
rect 8000 4333 8018 4367
rect 8052 4333 8070 4367
rect 8000 4307 8070 4333
rect 8100 4367 8170 4393
rect 8100 4333 8118 4367
rect 8152 4333 8170 4367
rect 8100 4307 8170 4333
rect 8200 4307 8270 4393
rect 8300 4367 8370 4393
rect 8300 4333 8318 4367
rect 8352 4333 8370 4367
rect 8300 4307 8370 4333
rect 8400 4367 8470 4393
rect 8400 4333 8418 4367
rect 8452 4333 8470 4367
rect 8400 4307 8470 4333
rect 8500 4307 8570 4393
rect 8600 4367 8670 4393
rect 8600 4333 8618 4367
rect 8652 4333 8670 4367
rect 8600 4307 8670 4333
rect 8700 4367 8770 4393
rect 8700 4333 8718 4367
rect 8752 4333 8770 4367
rect 8700 4307 8770 4333
rect 8800 4307 8870 4393
rect 8900 4367 8970 4393
rect 8900 4333 8918 4367
rect 8952 4333 8970 4367
rect 8900 4307 8970 4333
rect 9000 4367 9070 4393
rect 9000 4333 9018 4367
rect 9052 4333 9070 4367
rect 9000 4307 9070 4333
rect 9100 4367 9170 4393
rect 9100 4333 9118 4367
rect 9152 4333 9170 4367
rect 9100 4307 9170 4333
rect 9200 4307 9270 4393
rect 9300 4367 9370 4393
rect 9300 4333 9318 4367
rect 9352 4333 9370 4367
rect 9300 4307 9370 4333
rect 9400 4367 9470 4393
rect 9400 4333 9418 4367
rect 9452 4333 9470 4367
rect 9400 4307 9470 4333
rect 9500 4307 9570 4393
rect 9600 4307 9670 4393
rect 9700 4307 9770 4393
rect 9800 4307 9870 4393
rect 9900 4367 9970 4393
rect 9900 4333 9918 4367
rect 9952 4333 9970 4367
rect 9900 4307 9970 4333
rect 10000 4367 10070 4393
rect 10000 4333 10018 4367
rect 10052 4333 10070 4367
rect 10000 4307 10070 4333
rect 10100 4367 10170 4393
rect 10100 4333 10118 4367
rect 10152 4333 10170 4367
rect 10100 4307 10170 4333
rect 10200 4307 10270 4393
rect 10300 4367 10370 4393
rect 10300 4333 10318 4367
rect 10352 4333 10370 4367
rect 10300 4307 10370 4333
rect 10400 4367 10470 4393
rect 10400 4333 10418 4367
rect 10452 4333 10470 4367
rect 10400 4307 10470 4333
rect 10500 4307 10570 4393
rect 10600 4367 10670 4393
rect 10600 4333 10618 4367
rect 10652 4333 10670 4367
rect 10600 4307 10670 4333
rect 10700 4367 10770 4393
rect 10700 4333 10718 4367
rect 10752 4333 10770 4367
rect 10700 4307 10770 4333
rect 10800 4367 10854 4393
rect 10800 4333 10812 4367
rect 10846 4333 10854 4367
rect 10800 4307 10854 4333
rect 7216 4227 7270 4253
rect 7216 4193 7224 4227
rect 7258 4193 7270 4227
rect 7216 4167 7270 4193
rect 7300 4227 7370 4253
rect 7300 4193 7318 4227
rect 7352 4193 7370 4227
rect 7300 4167 7370 4193
rect 7400 4167 7470 4253
rect 7500 4227 7570 4253
rect 7500 4193 7518 4227
rect 7552 4193 7570 4227
rect 7500 4167 7570 4193
rect 7600 4227 7670 4253
rect 7600 4193 7618 4227
rect 7652 4193 7670 4227
rect 7600 4167 7670 4193
rect 7700 4227 7770 4253
rect 7700 4193 7718 4227
rect 7752 4193 7770 4227
rect 7700 4167 7770 4193
rect 7800 4167 7870 4253
rect 7900 4227 7970 4253
rect 7900 4193 7918 4227
rect 7952 4193 7970 4227
rect 7900 4167 7970 4193
rect 8000 4227 8070 4253
rect 8000 4193 8018 4227
rect 8052 4193 8070 4227
rect 8000 4167 8070 4193
rect 8100 4227 8154 4253
rect 8100 4193 8112 4227
rect 8146 4193 8154 4227
rect 8100 4167 8154 4193
rect 5716 4087 5770 4113
rect 5716 4053 5724 4087
rect 5758 4053 5770 4087
rect 5716 4027 5770 4053
rect 5800 4087 5870 4113
rect 5800 4053 5818 4087
rect 5852 4053 5870 4087
rect 5800 4027 5870 4053
rect 5900 4027 5970 4113
rect 6000 4027 6070 4113
rect 6100 4027 6170 4113
rect 6200 4087 6270 4113
rect 6200 4053 6218 4087
rect 6252 4053 6270 4087
rect 6200 4027 6270 4053
rect 6300 4087 6370 4113
rect 6300 4053 6318 4087
rect 6352 4053 6370 4087
rect 6300 4027 6370 4053
rect 6400 4087 6470 4113
rect 6400 4053 6418 4087
rect 6452 4053 6470 4087
rect 6400 4027 6470 4053
rect 6500 4087 6570 4113
rect 6500 4053 6518 4087
rect 6552 4053 6570 4087
rect 6500 4027 6570 4053
rect 6600 4027 6670 4113
rect 6700 4027 6770 4113
rect 6800 4087 6870 4113
rect 6800 4053 6818 4087
rect 6852 4053 6870 4087
rect 6800 4027 6870 4053
rect 6900 4087 6970 4113
rect 6900 4053 6918 4087
rect 6952 4053 6970 4087
rect 6900 4027 6970 4053
rect 7000 4087 7070 4113
rect 7000 4053 7018 4087
rect 7052 4053 7070 4087
rect 7000 4027 7070 4053
rect 7100 4087 7170 4113
rect 7100 4053 7118 4087
rect 7152 4053 7170 4087
rect 7100 4027 7170 4053
rect 7200 4087 7270 4113
rect 7200 4053 7218 4087
rect 7252 4053 7270 4087
rect 7200 4027 7270 4053
rect 7300 4087 7354 4113
rect 7300 4053 7312 4087
rect 7346 4053 7354 4087
rect 7300 4027 7354 4053
rect 5616 3947 5670 3973
rect 5616 3913 5624 3947
rect 5658 3913 5670 3947
rect 5616 3887 5670 3913
rect 5700 3947 5770 3973
rect 5700 3913 5718 3947
rect 5752 3913 5770 3947
rect 5700 3887 5770 3913
rect 5800 3947 5870 3973
rect 5800 3913 5818 3947
rect 5852 3913 5870 3947
rect 5800 3887 5870 3913
rect 5900 3947 5954 3973
rect 5900 3913 5912 3947
rect 5946 3913 5954 3947
rect 5900 3887 5954 3913
rect 5516 3807 5570 3833
rect 5516 3773 5524 3807
rect 5558 3773 5570 3807
rect 5516 3747 5570 3773
rect 5600 3807 5670 3833
rect 5600 3773 5618 3807
rect 5652 3773 5670 3807
rect 5600 3747 5670 3773
rect 5700 3807 5770 3833
rect 5700 3773 5718 3807
rect 5752 3773 5770 3807
rect 5700 3747 5770 3773
rect 5800 3807 5870 3833
rect 5800 3773 5818 3807
rect 5852 3773 5870 3807
rect 5800 3747 5870 3773
rect 5900 3807 5954 3833
rect 5900 3773 5912 3807
rect 5946 3773 5954 3807
rect 5900 3747 5954 3773
rect 4516 3577 4570 3603
rect 4516 3543 4524 3577
rect 4558 3543 4570 3577
rect 4516 3517 4570 3543
rect 4600 3577 4670 3603
rect 4600 3543 4618 3577
rect 4652 3543 4670 3577
rect 4600 3517 4670 3543
rect 4700 3577 4770 3603
rect 4700 3543 4718 3577
rect 4752 3543 4770 3577
rect 4700 3517 4770 3543
rect 4800 3517 4870 3603
rect 4900 3517 4970 3603
rect 5000 3517 5070 3603
rect 5100 3577 5170 3603
rect 5100 3543 5118 3577
rect 5152 3543 5170 3577
rect 5100 3517 5170 3543
rect 5200 3577 5270 3603
rect 5200 3543 5218 3577
rect 5252 3543 5270 3577
rect 5200 3517 5270 3543
rect 5300 3517 5370 3603
rect 5400 3577 5470 3603
rect 5400 3543 5418 3577
rect 5452 3543 5470 3577
rect 5400 3517 5470 3543
rect 5500 3577 5570 3603
rect 5500 3543 5518 3577
rect 5552 3543 5570 3577
rect 5500 3517 5570 3543
rect 5600 3577 5670 3603
rect 5600 3543 5618 3577
rect 5652 3543 5670 3577
rect 5600 3517 5670 3543
rect 5700 3577 5754 3603
rect 5700 3543 5712 3577
rect 5746 3543 5754 3577
rect 5700 3517 5754 3543
rect 4516 3437 4570 3463
rect 4516 3403 4524 3437
rect 4558 3403 4570 3437
rect 4516 3377 4570 3403
rect 4600 3437 4670 3463
rect 4600 3403 4618 3437
rect 4652 3403 4670 3437
rect 4600 3377 4670 3403
rect 4700 3437 4770 3463
rect 4700 3403 4718 3437
rect 4752 3403 4770 3437
rect 4700 3377 4770 3403
rect 4800 3437 4854 3463
rect 4800 3403 4812 3437
rect 4846 3403 4854 3437
rect 4800 3377 4854 3403
rect 4916 3437 4970 3463
rect 4916 3403 4924 3437
rect 4958 3403 4970 3437
rect 4916 3377 4970 3403
rect 5000 3437 5054 3463
rect 5000 3403 5012 3437
rect 5046 3403 5054 3437
rect 5000 3377 5054 3403
rect 6016 3947 6070 3973
rect 6016 3913 6024 3947
rect 6058 3913 6070 3947
rect 6016 3887 6070 3913
rect 6100 3947 6170 3973
rect 6100 3913 6118 3947
rect 6152 3913 6170 3947
rect 6100 3887 6170 3913
rect 6200 3947 6270 3973
rect 6200 3913 6218 3947
rect 6252 3913 6270 3947
rect 6200 3887 6270 3913
rect 6300 3947 6370 3973
rect 6300 3913 6318 3947
rect 6352 3913 6370 3947
rect 6300 3887 6370 3913
rect 6400 3887 6470 3973
rect 6500 3887 6570 3973
rect 6600 3947 6670 3973
rect 6600 3913 6618 3947
rect 6652 3913 6670 3947
rect 6600 3887 6670 3913
rect 6700 3947 6770 3973
rect 6700 3913 6718 3947
rect 6752 3913 6770 3947
rect 6700 3887 6770 3913
rect 6800 3947 6870 3973
rect 6800 3913 6818 3947
rect 6852 3913 6870 3947
rect 6800 3887 6870 3913
rect 6900 3947 6954 3973
rect 6900 3913 6912 3947
rect 6946 3913 6954 3947
rect 6900 3887 6954 3913
rect 7016 3947 7070 3973
rect 7016 3913 7024 3947
rect 7058 3913 7070 3947
rect 7016 3887 7070 3913
rect 7100 3947 7154 3973
rect 7100 3913 7112 3947
rect 7146 3913 7154 3947
rect 7100 3887 7154 3913
rect 7416 4087 7470 4113
rect 7416 4053 7424 4087
rect 7458 4053 7470 4087
rect 7416 4027 7470 4053
rect 7500 4087 7570 4113
rect 7500 4053 7518 4087
rect 7552 4053 7570 4087
rect 7500 4027 7570 4053
rect 7600 4087 7654 4113
rect 7600 4053 7612 4087
rect 7646 4053 7654 4087
rect 7600 4027 7654 4053
rect 7716 4087 7770 4113
rect 7716 4053 7724 4087
rect 7758 4053 7770 4087
rect 7716 4027 7770 4053
rect 7800 4087 7854 4113
rect 7800 4053 7812 4087
rect 7846 4053 7854 4087
rect 7800 4027 7854 4053
rect 8216 4227 8270 4253
rect 8216 4193 8224 4227
rect 8258 4193 8270 4227
rect 8216 4167 8270 4193
rect 8300 4227 8354 4253
rect 8300 4193 8312 4227
rect 8346 4193 8354 4227
rect 8300 4167 8354 4193
rect 8416 4227 8470 4253
rect 8416 4193 8424 4227
rect 8458 4193 8470 4227
rect 8416 4167 8470 4193
rect 8500 4227 8554 4253
rect 8500 4193 8512 4227
rect 8546 4193 8554 4227
rect 8500 4167 8554 4193
rect 8616 4227 8670 4253
rect 8616 4193 8624 4227
rect 8658 4193 8670 4227
rect 8616 4167 8670 4193
rect 8700 4227 8754 4253
rect 8700 4193 8712 4227
rect 8746 4193 8754 4227
rect 8700 4167 8754 4193
rect 7916 4087 7970 4113
rect 7916 4053 7924 4087
rect 7958 4053 7970 4087
rect 7916 4027 7970 4053
rect 8000 4087 8070 4113
rect 8000 4053 8018 4087
rect 8052 4053 8070 4087
rect 8000 4027 8070 4053
rect 8100 4087 8170 4113
rect 8100 4053 8118 4087
rect 8152 4053 8170 4087
rect 8100 4027 8170 4053
rect 8200 4027 8270 4113
rect 8300 4027 8370 4113
rect 8400 4087 8470 4113
rect 8400 4053 8418 4087
rect 8452 4053 8470 4087
rect 8400 4027 8470 4053
rect 8500 4087 8570 4113
rect 8500 4053 8518 4087
rect 8552 4053 8570 4087
rect 8500 4027 8570 4053
rect 8600 4087 8670 4113
rect 8600 4053 8618 4087
rect 8652 4053 8670 4087
rect 8600 4027 8670 4053
rect 8700 4087 8754 4113
rect 8700 4053 8712 4087
rect 8746 4053 8754 4087
rect 8700 4027 8754 4053
rect 7216 3947 7270 3973
rect 7216 3913 7224 3947
rect 7258 3913 7270 3947
rect 7216 3887 7270 3913
rect 7300 3947 7370 3973
rect 7300 3913 7318 3947
rect 7352 3913 7370 3947
rect 7300 3887 7370 3913
rect 7400 3947 7470 3973
rect 7400 3913 7418 3947
rect 7452 3913 7470 3947
rect 7400 3887 7470 3913
rect 7500 3947 7570 3973
rect 7500 3913 7518 3947
rect 7552 3913 7570 3947
rect 7500 3887 7570 3913
rect 7600 3947 7670 3973
rect 7600 3913 7618 3947
rect 7652 3913 7670 3947
rect 7600 3887 7670 3913
rect 7700 3887 7770 3973
rect 7800 3887 7870 3973
rect 7900 3887 7970 3973
rect 8000 3947 8070 3973
rect 8000 3913 8018 3947
rect 8052 3913 8070 3947
rect 8000 3887 8070 3913
rect 8100 3947 8170 3973
rect 8100 3913 8118 3947
rect 8152 3913 8170 3947
rect 8100 3887 8170 3913
rect 8200 3887 8270 3973
rect 8300 3887 8370 3973
rect 8400 3887 8470 3973
rect 8500 3947 8570 3973
rect 8500 3913 8518 3947
rect 8552 3913 8570 3947
rect 8500 3887 8570 3913
rect 8600 3947 8670 3973
rect 8600 3913 8618 3947
rect 8652 3913 8670 3947
rect 8600 3887 8670 3913
rect 8700 3947 8754 3973
rect 8700 3913 8712 3947
rect 8746 3913 8754 3947
rect 8700 3887 8754 3913
rect 6016 3807 6070 3833
rect 6016 3773 6024 3807
rect 6058 3773 6070 3807
rect 6016 3747 6070 3773
rect 6100 3807 6170 3833
rect 6100 3773 6118 3807
rect 6152 3773 6170 3807
rect 6100 3747 6170 3773
rect 6200 3747 6270 3833
rect 6300 3747 6370 3833
rect 6400 3747 6470 3833
rect 6500 3807 6570 3833
rect 6500 3773 6518 3807
rect 6552 3773 6570 3807
rect 6500 3747 6570 3773
rect 6600 3807 6670 3833
rect 6600 3773 6618 3807
rect 6652 3773 6670 3807
rect 6600 3747 6670 3773
rect 6700 3747 6770 3833
rect 6800 3747 6870 3833
rect 6900 3747 6970 3833
rect 7000 3747 7070 3833
rect 7100 3807 7170 3833
rect 7100 3773 7118 3807
rect 7152 3773 7170 3807
rect 7100 3747 7170 3773
rect 7200 3807 7270 3833
rect 7200 3773 7218 3807
rect 7252 3773 7270 3807
rect 7200 3747 7270 3773
rect 7300 3747 7370 3833
rect 7400 3747 7470 3833
rect 7500 3807 7570 3833
rect 7500 3773 7518 3807
rect 7552 3773 7570 3807
rect 7500 3747 7570 3773
rect 7600 3807 7654 3833
rect 7600 3773 7612 3807
rect 7646 3773 7654 3807
rect 7600 3747 7654 3773
rect 8816 4227 8870 4253
rect 8816 4193 8824 4227
rect 8858 4193 8870 4227
rect 8816 4167 8870 4193
rect 8900 4227 8954 4253
rect 8900 4193 8912 4227
rect 8946 4193 8954 4227
rect 8900 4167 8954 4193
rect 8816 4087 8870 4113
rect 8816 4053 8824 4087
rect 8858 4053 8870 4087
rect 8816 4027 8870 4053
rect 8900 4087 8954 4113
rect 8900 4053 8912 4087
rect 8946 4053 8954 4087
rect 8900 4027 8954 4053
rect 9016 4227 9070 4253
rect 9016 4193 9024 4227
rect 9058 4193 9070 4227
rect 9016 4167 9070 4193
rect 9100 4227 9170 4253
rect 9100 4193 9118 4227
rect 9152 4193 9170 4227
rect 9100 4167 9170 4193
rect 9200 4227 9270 4253
rect 9200 4193 9218 4227
rect 9252 4193 9270 4227
rect 9200 4167 9270 4193
rect 9300 4227 9354 4253
rect 9300 4193 9312 4227
rect 9346 4193 9354 4227
rect 9300 4167 9354 4193
rect 9416 4227 9470 4253
rect 9416 4193 9424 4227
rect 9458 4193 9470 4227
rect 9416 4167 9470 4193
rect 9500 4227 9554 4253
rect 9500 4193 9512 4227
rect 9546 4193 9554 4227
rect 9500 4167 9554 4193
rect 9016 4087 9070 4113
rect 9016 4053 9024 4087
rect 9058 4053 9070 4087
rect 9016 4027 9070 4053
rect 9100 4087 9170 4113
rect 9100 4053 9118 4087
rect 9152 4053 9170 4087
rect 9100 4027 9170 4053
rect 9200 4027 9270 4113
rect 9300 4087 9370 4113
rect 9300 4053 9318 4087
rect 9352 4053 9370 4087
rect 9300 4027 9370 4053
rect 9400 4087 9470 4113
rect 9400 4053 9418 4087
rect 9452 4053 9470 4087
rect 9400 4027 9470 4053
rect 9500 4087 9554 4113
rect 9500 4053 9512 4087
rect 9546 4053 9554 4087
rect 9500 4027 9554 4053
rect 8816 3947 8870 3973
rect 8816 3913 8824 3947
rect 8858 3913 8870 3947
rect 8816 3887 8870 3913
rect 8900 3947 8970 3973
rect 8900 3913 8918 3947
rect 8952 3913 8970 3947
rect 8900 3887 8970 3913
rect 9000 3887 9070 3973
rect 9100 3887 9170 3973
rect 9200 3887 9270 3973
rect 9300 3887 9370 3973
rect 9400 3947 9470 3973
rect 9400 3913 9418 3947
rect 9452 3913 9470 3947
rect 9400 3887 9470 3913
rect 9500 3947 9554 3973
rect 9500 3913 9512 3947
rect 9546 3913 9554 3947
rect 9500 3887 9554 3913
rect 7716 3807 7770 3833
rect 7716 3773 7724 3807
rect 7758 3773 7770 3807
rect 7716 3747 7770 3773
rect 7800 3807 7870 3833
rect 7800 3773 7818 3807
rect 7852 3773 7870 3807
rect 7800 3747 7870 3773
rect 7900 3807 7970 3833
rect 7900 3773 7918 3807
rect 7952 3773 7970 3807
rect 7900 3747 7970 3773
rect 8000 3807 8070 3833
rect 8000 3773 8018 3807
rect 8052 3773 8070 3807
rect 8000 3747 8070 3773
rect 8100 3807 8170 3833
rect 8100 3773 8118 3807
rect 8152 3773 8170 3807
rect 8100 3747 8170 3773
rect 8200 3807 8270 3833
rect 8200 3773 8218 3807
rect 8252 3773 8270 3807
rect 8200 3747 8270 3773
rect 8300 3807 8370 3833
rect 8300 3773 8318 3807
rect 8352 3773 8370 3807
rect 8300 3747 8370 3773
rect 8400 3807 8470 3833
rect 8400 3773 8418 3807
rect 8452 3773 8470 3807
rect 8400 3747 8470 3773
rect 8500 3747 8570 3833
rect 8600 3807 8670 3833
rect 8600 3773 8618 3807
rect 8652 3773 8670 3807
rect 8600 3747 8670 3773
rect 8700 3807 8770 3833
rect 8700 3773 8718 3807
rect 8752 3773 8770 3807
rect 8700 3747 8770 3773
rect 8800 3807 8870 3833
rect 8800 3773 8818 3807
rect 8852 3773 8870 3807
rect 8800 3747 8870 3773
rect 8900 3747 8970 3833
rect 9000 3747 9070 3833
rect 9100 3747 9170 3833
rect 9200 3807 9270 3833
rect 9200 3773 9218 3807
rect 9252 3773 9270 3807
rect 9200 3747 9270 3773
rect 9300 3807 9370 3833
rect 9300 3773 9318 3807
rect 9352 3773 9370 3807
rect 9300 3747 9370 3773
rect 9400 3807 9454 3833
rect 9400 3773 9412 3807
rect 9446 3773 9454 3807
rect 9400 3747 9454 3773
rect 5816 3577 5870 3603
rect 5816 3543 5824 3577
rect 5858 3543 5870 3577
rect 5816 3517 5870 3543
rect 5900 3577 5970 3603
rect 5900 3543 5918 3577
rect 5952 3543 5970 3577
rect 5900 3517 5970 3543
rect 6000 3577 6070 3603
rect 6000 3543 6018 3577
rect 6052 3543 6070 3577
rect 6000 3517 6070 3543
rect 6100 3517 6170 3603
rect 6200 3517 6270 3603
rect 6300 3517 6370 3603
rect 6400 3517 6470 3603
rect 6500 3517 6570 3603
rect 6600 3577 6670 3603
rect 6600 3543 6618 3577
rect 6652 3543 6670 3577
rect 6600 3517 6670 3543
rect 6700 3577 6770 3603
rect 6700 3543 6718 3577
rect 6752 3543 6770 3577
rect 6700 3517 6770 3543
rect 6800 3577 6870 3603
rect 6800 3543 6818 3577
rect 6852 3543 6870 3577
rect 6800 3517 6870 3543
rect 6900 3517 6970 3603
rect 7000 3517 7070 3603
rect 7100 3517 7170 3603
rect 7200 3517 7270 3603
rect 7300 3517 7370 3603
rect 7400 3577 7470 3603
rect 7400 3543 7418 3577
rect 7452 3543 7470 3577
rect 7400 3517 7470 3543
rect 7500 3577 7570 3603
rect 7500 3543 7518 3577
rect 7552 3543 7570 3577
rect 7500 3517 7570 3543
rect 7600 3577 7670 3603
rect 7600 3543 7618 3577
rect 7652 3543 7670 3577
rect 7600 3517 7670 3543
rect 7700 3517 7770 3603
rect 7800 3517 7870 3603
rect 7900 3517 7970 3603
rect 8000 3577 8070 3603
rect 8000 3543 8018 3577
rect 8052 3543 8070 3577
rect 8000 3517 8070 3543
rect 8100 3577 8170 3603
rect 8100 3543 8118 3577
rect 8152 3543 8170 3577
rect 8100 3517 8170 3543
rect 8200 3517 8270 3603
rect 8300 3577 8370 3603
rect 8300 3543 8318 3577
rect 8352 3543 8370 3577
rect 8300 3517 8370 3543
rect 8400 3577 8470 3603
rect 8400 3543 8418 3577
rect 8452 3543 8470 3577
rect 8400 3517 8470 3543
rect 8500 3577 8570 3603
rect 8500 3543 8518 3577
rect 8552 3543 8570 3577
rect 8500 3517 8570 3543
rect 8600 3517 8670 3603
rect 8700 3517 8770 3603
rect 8800 3577 8870 3603
rect 8800 3543 8818 3577
rect 8852 3543 8870 3577
rect 8800 3517 8870 3543
rect 8900 3577 8954 3603
rect 8900 3543 8912 3577
rect 8946 3543 8954 3577
rect 8900 3517 8954 3543
rect 5116 3437 5170 3463
rect 5116 3403 5124 3437
rect 5158 3403 5170 3437
rect 5116 3377 5170 3403
rect 5200 3437 5270 3463
rect 5200 3403 5218 3437
rect 5252 3403 5270 3437
rect 5200 3377 5270 3403
rect 5300 3377 5370 3463
rect 5400 3437 5470 3463
rect 5400 3403 5418 3437
rect 5452 3403 5470 3437
rect 5400 3377 5470 3403
rect 5500 3437 5570 3463
rect 5500 3403 5518 3437
rect 5552 3403 5570 3437
rect 5500 3377 5570 3403
rect 5600 3437 5670 3463
rect 5600 3403 5618 3437
rect 5652 3403 5670 3437
rect 5600 3377 5670 3403
rect 5700 3377 5770 3463
rect 5800 3377 5870 3463
rect 5900 3437 5970 3463
rect 5900 3403 5918 3437
rect 5952 3403 5970 3437
rect 5900 3377 5970 3403
rect 6000 3437 6054 3463
rect 6000 3403 6012 3437
rect 6046 3403 6054 3437
rect 6000 3377 6054 3403
rect 6116 3437 6170 3463
rect 6116 3403 6124 3437
rect 6158 3403 6170 3437
rect 6116 3377 6170 3403
rect 6200 3437 6270 3463
rect 6200 3403 6218 3437
rect 6252 3403 6270 3437
rect 6200 3377 6270 3403
rect 6300 3437 6370 3463
rect 6300 3403 6318 3437
rect 6352 3403 6370 3437
rect 6300 3377 6370 3403
rect 6400 3437 6454 3463
rect 6400 3403 6412 3437
rect 6446 3403 6454 3437
rect 6400 3377 6454 3403
rect 6516 3437 6570 3463
rect 6516 3403 6524 3437
rect 6558 3403 6570 3437
rect 6516 3377 6570 3403
rect 6600 3437 6670 3463
rect 6600 3403 6618 3437
rect 6652 3403 6670 3437
rect 6600 3377 6670 3403
rect 6700 3437 6754 3463
rect 6700 3403 6712 3437
rect 6746 3403 6754 3437
rect 6700 3377 6754 3403
rect 9016 3577 9070 3603
rect 9016 3543 9024 3577
rect 9058 3543 9070 3577
rect 9016 3517 9070 3543
rect 9100 3577 9154 3603
rect 9100 3543 9112 3577
rect 9146 3543 9154 3577
rect 9100 3517 9154 3543
rect 9216 3577 9270 3603
rect 9216 3543 9224 3577
rect 9258 3543 9270 3577
rect 9216 3517 9270 3543
rect 9300 3577 9354 3603
rect 9300 3543 9312 3577
rect 9346 3543 9354 3577
rect 9300 3517 9354 3543
rect 9616 4227 9670 4253
rect 9616 4193 9624 4227
rect 9658 4193 9670 4227
rect 9616 4167 9670 4193
rect 9700 4227 9754 4253
rect 9700 4193 9712 4227
rect 9746 4193 9754 4227
rect 9700 4167 9754 4193
rect 9816 4227 9870 4253
rect 9816 4193 9824 4227
rect 9858 4193 9870 4227
rect 9816 4167 9870 4193
rect 9900 4227 9970 4253
rect 9900 4193 9918 4227
rect 9952 4193 9970 4227
rect 9900 4167 9970 4193
rect 10000 4227 10054 4253
rect 10000 4193 10012 4227
rect 10046 4193 10054 4227
rect 10000 4167 10054 4193
rect 11016 4507 11070 4533
rect 11016 4473 11024 4507
rect 11058 4473 11070 4507
rect 11016 4447 11070 4473
rect 11100 4507 11170 4533
rect 11100 4473 11118 4507
rect 11152 4473 11170 4507
rect 11100 4447 11170 4473
rect 11200 4507 11254 4533
rect 11200 4473 11212 4507
rect 11246 4473 11254 4507
rect 11200 4447 11254 4473
rect 10916 4367 10970 4393
rect 10916 4333 10924 4367
rect 10958 4333 10970 4367
rect 10916 4307 10970 4333
rect 11000 4367 11070 4393
rect 11000 4333 11018 4367
rect 11052 4333 11070 4367
rect 11000 4307 11070 4333
rect 11100 4367 11154 4393
rect 11100 4333 11112 4367
rect 11146 4333 11154 4367
rect 11100 4307 11154 4333
rect 10116 4227 10170 4253
rect 10116 4193 10124 4227
rect 10158 4193 10170 4227
rect 10116 4167 10170 4193
rect 10200 4227 10270 4253
rect 10200 4193 10218 4227
rect 10252 4193 10270 4227
rect 10200 4167 10270 4193
rect 10300 4167 10370 4253
rect 10400 4167 10470 4253
rect 10500 4167 10570 4253
rect 10600 4227 10670 4253
rect 10600 4193 10618 4227
rect 10652 4193 10670 4227
rect 10600 4167 10670 4193
rect 10700 4227 10770 4253
rect 10700 4193 10718 4227
rect 10752 4193 10770 4227
rect 10700 4167 10770 4193
rect 10800 4227 10870 4253
rect 10800 4193 10818 4227
rect 10852 4193 10870 4227
rect 10800 4167 10870 4193
rect 10900 4227 10954 4253
rect 10900 4193 10912 4227
rect 10946 4193 10954 4227
rect 10900 4167 10954 4193
rect 9616 4087 9670 4113
rect 9616 4053 9624 4087
rect 9658 4053 9670 4087
rect 9616 4027 9670 4053
rect 9700 4087 9770 4113
rect 9700 4053 9718 4087
rect 9752 4053 9770 4087
rect 9700 4027 9770 4053
rect 9800 4027 9870 4113
rect 9900 4087 9970 4113
rect 9900 4053 9918 4087
rect 9952 4053 9970 4087
rect 9900 4027 9970 4053
rect 10000 4087 10070 4113
rect 10000 4053 10018 4087
rect 10052 4053 10070 4087
rect 10000 4027 10070 4053
rect 10100 4087 10170 4113
rect 10100 4053 10118 4087
rect 10152 4053 10170 4087
rect 10100 4027 10170 4053
rect 10200 4087 10270 4113
rect 10200 4053 10218 4087
rect 10252 4053 10270 4087
rect 10200 4027 10270 4053
rect 10300 4087 10370 4113
rect 10300 4053 10318 4087
rect 10352 4053 10370 4087
rect 10300 4027 10370 4053
rect 10400 4087 10470 4113
rect 10400 4053 10418 4087
rect 10452 4053 10470 4087
rect 10400 4027 10470 4053
rect 10500 4087 10570 4113
rect 10500 4053 10518 4087
rect 10552 4053 10570 4087
rect 10500 4027 10570 4053
rect 10600 4087 10654 4113
rect 10600 4053 10612 4087
rect 10646 4053 10654 4087
rect 10600 4027 10654 4053
rect 10716 4087 10770 4113
rect 10716 4053 10724 4087
rect 10758 4053 10770 4087
rect 10716 4027 10770 4053
rect 10800 4087 10854 4113
rect 10800 4053 10812 4087
rect 10846 4053 10854 4087
rect 10800 4027 10854 4053
rect 11316 4507 11370 4533
rect 11316 4473 11324 4507
rect 11358 4473 11370 4507
rect 11316 4447 11370 4473
rect 11400 4507 11470 4533
rect 11400 4473 11418 4507
rect 11452 4473 11470 4507
rect 11400 4447 11470 4473
rect 11500 4507 11570 4533
rect 11500 4473 11518 4507
rect 11552 4473 11570 4507
rect 11500 4447 11570 4473
rect 11600 4447 11670 4533
rect 11700 4447 11770 4533
rect 11800 4447 11870 4533
rect 11900 4507 11970 4533
rect 11900 4473 11918 4507
rect 11952 4473 11970 4507
rect 11900 4447 11970 4473
rect 12000 4507 12070 4533
rect 12000 4473 12018 4507
rect 12052 4473 12070 4507
rect 12000 4447 12070 4473
rect 12100 4507 12170 4533
rect 12100 4473 12118 4507
rect 12152 4473 12170 4507
rect 12100 4447 12170 4473
rect 12200 4447 12270 4533
rect 12300 4507 12370 4533
rect 12300 4473 12318 4507
rect 12352 4473 12370 4507
rect 12300 4447 12370 4473
rect 12400 4507 12454 4533
rect 12400 4473 12412 4507
rect 12446 4473 12454 4507
rect 12400 4447 12454 4473
rect 11216 4367 11270 4393
rect 11216 4333 11224 4367
rect 11258 4333 11270 4367
rect 11216 4307 11270 4333
rect 11300 4367 11370 4393
rect 11300 4333 11318 4367
rect 11352 4333 11370 4367
rect 11300 4307 11370 4333
rect 11400 4367 11470 4393
rect 11400 4333 11418 4367
rect 11452 4333 11470 4367
rect 11400 4307 11470 4333
rect 11500 4307 11570 4393
rect 11600 4307 11670 4393
rect 11700 4367 11770 4393
rect 11700 4333 11718 4367
rect 11752 4333 11770 4367
rect 11700 4307 11770 4333
rect 11800 4367 11870 4393
rect 11800 4333 11818 4367
rect 11852 4333 11870 4367
rect 11800 4307 11870 4333
rect 11900 4367 11954 4393
rect 11900 4333 11912 4367
rect 11946 4333 11954 4367
rect 11900 4307 11954 4333
rect 11016 4227 11070 4253
rect 11016 4193 11024 4227
rect 11058 4193 11070 4227
rect 11016 4167 11070 4193
rect 11100 4227 11170 4253
rect 11100 4193 11118 4227
rect 11152 4193 11170 4227
rect 11100 4167 11170 4193
rect 11200 4227 11270 4253
rect 11200 4193 11218 4227
rect 11252 4193 11270 4227
rect 11200 4167 11270 4193
rect 11300 4227 11354 4253
rect 11300 4193 11312 4227
rect 11346 4193 11354 4227
rect 11300 4167 11354 4193
rect 10916 4087 10970 4113
rect 10916 4053 10924 4087
rect 10958 4053 10970 4087
rect 10916 4027 10970 4053
rect 11000 4087 11070 4113
rect 11000 4053 11018 4087
rect 11052 4053 11070 4087
rect 11000 4027 11070 4053
rect 11100 4027 11170 4113
rect 11200 4087 11270 4113
rect 11200 4053 11218 4087
rect 11252 4053 11270 4087
rect 11200 4027 11270 4053
rect 11300 4087 11354 4113
rect 11300 4053 11312 4087
rect 11346 4053 11354 4087
rect 11300 4027 11354 4053
rect 9616 3947 9670 3973
rect 9616 3913 9624 3947
rect 9658 3913 9670 3947
rect 9616 3887 9670 3913
rect 9700 3947 9770 3973
rect 9700 3913 9718 3947
rect 9752 3913 9770 3947
rect 9700 3887 9770 3913
rect 9800 3947 9870 3973
rect 9800 3913 9818 3947
rect 9852 3913 9870 3947
rect 9800 3887 9870 3913
rect 9900 3887 9970 3973
rect 10000 3887 10070 3973
rect 10100 3947 10170 3973
rect 10100 3913 10118 3947
rect 10152 3913 10170 3947
rect 10100 3887 10170 3913
rect 10200 3947 10270 3973
rect 10200 3913 10218 3947
rect 10252 3913 10270 3947
rect 10200 3887 10270 3913
rect 10300 3947 10370 3973
rect 10300 3913 10318 3947
rect 10352 3913 10370 3947
rect 10300 3887 10370 3913
rect 10400 3947 10470 3973
rect 10400 3913 10418 3947
rect 10452 3913 10470 3947
rect 10400 3887 10470 3913
rect 10500 3887 10570 3973
rect 10600 3887 10670 3973
rect 10700 3887 10770 3973
rect 10800 3887 10870 3973
rect 10900 3947 10970 3973
rect 10900 3913 10918 3947
rect 10952 3913 10970 3947
rect 10900 3887 10970 3913
rect 11000 3947 11054 3973
rect 11000 3913 11012 3947
rect 11046 3913 11054 3947
rect 11000 3887 11054 3913
rect 9516 3807 9570 3833
rect 9516 3773 9524 3807
rect 9558 3773 9570 3807
rect 9516 3747 9570 3773
rect 9600 3807 9670 3833
rect 9600 3773 9618 3807
rect 9652 3773 9670 3807
rect 9600 3747 9670 3773
rect 9700 3807 9770 3833
rect 9700 3773 9718 3807
rect 9752 3773 9770 3807
rect 9700 3747 9770 3773
rect 9800 3747 9870 3833
rect 9900 3807 9970 3833
rect 9900 3773 9918 3807
rect 9952 3773 9970 3807
rect 9900 3747 9970 3773
rect 10000 3807 10054 3833
rect 10000 3773 10012 3807
rect 10046 3773 10054 3807
rect 10000 3747 10054 3773
rect 11416 4227 11470 4253
rect 11416 4193 11424 4227
rect 11458 4193 11470 4227
rect 11416 4167 11470 4193
rect 11500 4227 11554 4253
rect 11500 4193 11512 4227
rect 11546 4193 11554 4227
rect 11500 4167 11554 4193
rect 11416 4087 11470 4113
rect 11416 4053 11424 4087
rect 11458 4053 11470 4087
rect 11416 4027 11470 4053
rect 11500 4087 11554 4113
rect 11500 4053 11512 4087
rect 11546 4053 11554 4087
rect 11500 4027 11554 4053
rect 12716 4647 12770 4673
rect 12716 4613 12724 4647
rect 12758 4613 12770 4647
rect 12716 4587 12770 4613
rect 12800 4647 12854 4673
rect 12800 4613 12812 4647
rect 12846 4613 12854 4647
rect 12800 4587 12854 4613
rect 12912 4662 12970 4673
rect 12912 4628 12924 4662
rect 12958 4628 12970 4662
rect 12912 4587 12970 4628
rect 13000 4647 13070 4673
rect 13000 4613 13018 4647
rect 13052 4613 13070 4647
rect 13000 4587 13070 4613
rect 13100 4632 13158 4673
rect 13100 4598 13112 4632
rect 13146 4598 13158 4632
rect 13100 4587 13158 4598
rect 13220 4647 13280 4673
rect 13220 4613 13228 4647
rect 13262 4613 13280 4647
rect 13220 4587 13280 4613
rect 13310 4647 13380 4673
rect 13310 4613 13328 4647
rect 13362 4613 13380 4647
rect 13310 4587 13380 4613
rect 13410 4647 13480 4673
rect 13410 4613 13428 4647
rect 13462 4613 13480 4647
rect 13410 4587 13480 4613
rect 13510 4647 13580 4673
rect 13510 4613 13528 4647
rect 13562 4613 13580 4647
rect 13510 4587 13580 4613
rect 13610 4647 13670 4673
rect 13610 4613 13628 4647
rect 13662 4613 13670 4647
rect 13610 4587 13670 4613
rect 12516 4507 12570 4533
rect 12516 4473 12524 4507
rect 12558 4473 12570 4507
rect 12516 4447 12570 4473
rect 12600 4507 12670 4533
rect 12600 4473 12618 4507
rect 12652 4473 12670 4507
rect 12600 4447 12670 4473
rect 12700 4507 12770 4533
rect 12700 4473 12718 4507
rect 12752 4473 12770 4507
rect 12700 4447 12770 4473
rect 12800 4507 12854 4533
rect 12800 4473 12812 4507
rect 12846 4473 12854 4507
rect 12800 4447 12854 4473
rect 12912 4522 12970 4533
rect 12912 4488 12924 4522
rect 12958 4488 12970 4522
rect 12912 4447 12970 4488
rect 13000 4507 13070 4533
rect 13000 4473 13018 4507
rect 13052 4473 13070 4507
rect 13000 4447 13070 4473
rect 13100 4492 13158 4533
rect 13100 4458 13112 4492
rect 13146 4458 13158 4492
rect 13100 4447 13158 4458
rect 13220 4507 13280 4533
rect 13220 4473 13228 4507
rect 13262 4473 13280 4507
rect 13220 4447 13280 4473
rect 13310 4507 13380 4533
rect 13310 4473 13328 4507
rect 13362 4473 13380 4507
rect 13310 4447 13380 4473
rect 13410 4507 13480 4533
rect 13410 4473 13428 4507
rect 13462 4473 13480 4507
rect 13410 4447 13480 4473
rect 13510 4507 13580 4533
rect 13510 4473 13528 4507
rect 13562 4473 13580 4507
rect 13510 4447 13580 4473
rect 13610 4507 13670 4533
rect 13610 4473 13628 4507
rect 13662 4473 13670 4507
rect 13610 4447 13670 4473
rect 12016 4367 12070 4393
rect 12016 4333 12024 4367
rect 12058 4333 12070 4367
rect 12016 4307 12070 4333
rect 12100 4367 12170 4393
rect 12100 4333 12118 4367
rect 12152 4333 12170 4367
rect 12100 4307 12170 4333
rect 12200 4367 12270 4393
rect 12200 4333 12218 4367
rect 12252 4333 12270 4367
rect 12200 4307 12270 4333
rect 12300 4367 12370 4393
rect 12300 4333 12318 4367
rect 12352 4333 12370 4367
rect 12300 4307 12370 4333
rect 12400 4307 12470 4393
rect 12500 4367 12570 4393
rect 12500 4333 12518 4367
rect 12552 4333 12570 4367
rect 12500 4307 12570 4333
rect 12600 4367 12670 4393
rect 12600 4333 12618 4367
rect 12652 4333 12670 4367
rect 12600 4307 12670 4333
rect 12700 4367 12770 4393
rect 12700 4333 12718 4367
rect 12752 4333 12770 4367
rect 12700 4307 12770 4333
rect 12800 4367 12854 4393
rect 12800 4333 12812 4367
rect 12846 4333 12854 4367
rect 12800 4307 12854 4333
rect 12912 4382 12970 4393
rect 12912 4348 12924 4382
rect 12958 4348 12970 4382
rect 12912 4307 12970 4348
rect 13000 4367 13070 4393
rect 13000 4333 13018 4367
rect 13052 4333 13070 4367
rect 13000 4307 13070 4333
rect 13100 4352 13158 4393
rect 13100 4318 13112 4352
rect 13146 4318 13158 4352
rect 13100 4307 13158 4318
rect 13220 4367 13280 4393
rect 13220 4333 13228 4367
rect 13262 4333 13280 4367
rect 13220 4307 13280 4333
rect 13310 4367 13380 4393
rect 13310 4333 13328 4367
rect 13362 4333 13380 4367
rect 13310 4307 13380 4333
rect 13410 4367 13480 4393
rect 13410 4333 13428 4367
rect 13462 4333 13480 4367
rect 13410 4307 13480 4333
rect 13510 4367 13580 4393
rect 13510 4333 13528 4367
rect 13562 4333 13580 4367
rect 13510 4307 13580 4333
rect 13610 4367 13670 4393
rect 13610 4333 13628 4367
rect 13662 4333 13670 4367
rect 13610 4307 13670 4333
rect 11616 4227 11670 4253
rect 11616 4193 11624 4227
rect 11658 4193 11670 4227
rect 11616 4167 11670 4193
rect 11700 4227 11770 4253
rect 11700 4193 11718 4227
rect 11752 4193 11770 4227
rect 11700 4167 11770 4193
rect 11800 4167 11870 4253
rect 11900 4167 11970 4253
rect 12000 4167 12070 4253
rect 12100 4167 12170 4253
rect 12200 4167 12270 4253
rect 12300 4167 12370 4253
rect 12400 4167 12470 4253
rect 12500 4167 12570 4253
rect 12600 4227 12670 4253
rect 12600 4193 12618 4227
rect 12652 4193 12670 4227
rect 12600 4167 12670 4193
rect 12700 4227 12770 4253
rect 12700 4193 12718 4227
rect 12752 4193 12770 4227
rect 12700 4167 12770 4193
rect 12800 4167 12854 4253
rect 12912 4242 12970 4253
rect 12912 4208 12924 4242
rect 12958 4208 12970 4242
rect 12912 4167 12970 4208
rect 13000 4227 13070 4253
rect 13000 4193 13018 4227
rect 13052 4193 13070 4227
rect 13000 4167 13070 4193
rect 13100 4212 13158 4253
rect 13100 4178 13112 4212
rect 13146 4178 13158 4212
rect 13100 4167 13158 4178
rect 13220 4227 13280 4253
rect 13220 4193 13228 4227
rect 13262 4193 13280 4227
rect 13220 4167 13280 4193
rect 13310 4227 13380 4253
rect 13310 4193 13328 4227
rect 13362 4193 13380 4227
rect 13310 4167 13380 4193
rect 13410 4227 13480 4253
rect 13410 4193 13428 4227
rect 13462 4193 13480 4227
rect 13410 4167 13480 4193
rect 13510 4227 13580 4253
rect 13510 4193 13528 4227
rect 13562 4193 13580 4227
rect 13510 4167 13580 4193
rect 13610 4227 13670 4253
rect 13610 4193 13628 4227
rect 13662 4193 13670 4227
rect 13610 4167 13670 4193
rect 11616 4087 11670 4113
rect 11616 4053 11624 4087
rect 11658 4053 11670 4087
rect 11616 4027 11670 4053
rect 11700 4087 11770 4113
rect 11700 4053 11718 4087
rect 11752 4053 11770 4087
rect 11700 4027 11770 4053
rect 11800 4087 11854 4113
rect 11800 4053 11812 4087
rect 11846 4053 11854 4087
rect 11800 4027 11854 4053
rect 11916 4087 11970 4113
rect 11916 4053 11924 4087
rect 11958 4053 11970 4087
rect 11916 4027 11970 4053
rect 12000 4087 12070 4113
rect 12000 4053 12018 4087
rect 12052 4053 12070 4087
rect 12000 4027 12070 4053
rect 12100 4027 12170 4113
rect 12200 4027 12270 4113
rect 12300 4087 12370 4113
rect 12300 4053 12318 4087
rect 12352 4053 12370 4087
rect 12300 4027 12370 4053
rect 12400 4087 12470 4113
rect 12400 4053 12418 4087
rect 12452 4053 12470 4087
rect 12400 4027 12470 4053
rect 12500 4087 12570 4113
rect 12500 4053 12518 4087
rect 12552 4053 12570 4087
rect 12500 4027 12570 4053
rect 12600 4087 12654 4113
rect 12600 4053 12612 4087
rect 12646 4053 12654 4087
rect 12600 4027 12654 4053
rect 12716 4087 12770 4113
rect 12716 4053 12724 4087
rect 12758 4053 12770 4087
rect 12716 4027 12770 4053
rect 12800 4087 12854 4113
rect 12800 4053 12812 4087
rect 12846 4053 12854 4087
rect 12800 4027 12854 4053
rect 12912 4102 12970 4113
rect 12912 4068 12924 4102
rect 12958 4068 12970 4102
rect 12912 4027 12970 4068
rect 13000 4087 13070 4113
rect 13000 4053 13018 4087
rect 13052 4053 13070 4087
rect 13000 4027 13070 4053
rect 13100 4072 13158 4113
rect 13100 4038 13112 4072
rect 13146 4038 13158 4072
rect 13100 4027 13158 4038
rect 13220 4087 13280 4113
rect 13220 4053 13228 4087
rect 13262 4053 13280 4087
rect 13220 4027 13280 4053
rect 13310 4087 13380 4113
rect 13310 4053 13328 4087
rect 13362 4053 13380 4087
rect 13310 4027 13380 4053
rect 13410 4087 13480 4113
rect 13410 4053 13428 4087
rect 13462 4053 13480 4087
rect 13410 4027 13480 4053
rect 13510 4087 13580 4113
rect 13510 4053 13528 4087
rect 13562 4053 13580 4087
rect 13510 4027 13580 4053
rect 13610 4087 13670 4113
rect 13610 4053 13628 4087
rect 13662 4053 13670 4087
rect 13610 4027 13670 4053
rect 11116 3947 11170 3973
rect 11116 3913 11124 3947
rect 11158 3913 11170 3947
rect 11116 3887 11170 3913
rect 11200 3947 11270 3973
rect 11200 3913 11218 3947
rect 11252 3913 11270 3947
rect 11200 3887 11270 3913
rect 11300 3947 11370 3973
rect 11300 3913 11318 3947
rect 11352 3913 11370 3947
rect 11300 3887 11370 3913
rect 11400 3887 11470 3973
rect 11500 3887 11570 3973
rect 11600 3887 11670 3973
rect 11700 3947 11770 3973
rect 11700 3913 11718 3947
rect 11752 3913 11770 3947
rect 11700 3887 11770 3913
rect 11800 3947 11870 3973
rect 11800 3913 11818 3947
rect 11852 3913 11870 3947
rect 11800 3887 11870 3913
rect 11900 3887 11970 3973
rect 12000 3887 12070 3973
rect 12100 3947 12170 3973
rect 12100 3913 12118 3947
rect 12152 3913 12170 3947
rect 12100 3887 12170 3913
rect 12200 3947 12270 3973
rect 12200 3913 12218 3947
rect 12252 3913 12270 3947
rect 12200 3887 12270 3913
rect 12300 3947 12370 3973
rect 12300 3913 12318 3947
rect 12352 3913 12370 3947
rect 12300 3887 12370 3913
rect 12400 3887 12470 3973
rect 12500 3947 12570 3973
rect 12500 3913 12518 3947
rect 12552 3913 12570 3947
rect 12500 3887 12570 3913
rect 12600 3947 12670 3973
rect 12600 3913 12618 3947
rect 12652 3913 12670 3947
rect 12600 3887 12670 3913
rect 12700 3947 12770 3973
rect 12700 3913 12718 3947
rect 12752 3913 12770 3947
rect 12700 3887 12770 3913
rect 12800 3947 12854 3973
rect 12800 3913 12812 3947
rect 12846 3913 12854 3947
rect 12800 3887 12854 3913
rect 12912 3962 12970 3973
rect 12912 3928 12924 3962
rect 12958 3928 12970 3962
rect 12912 3887 12970 3928
rect 13000 3947 13070 3973
rect 13000 3913 13018 3947
rect 13052 3913 13070 3947
rect 13000 3887 13070 3913
rect 13100 3932 13158 3973
rect 13100 3898 13112 3932
rect 13146 3898 13158 3932
rect 13100 3887 13158 3898
rect 13220 3947 13280 3973
rect 13220 3913 13228 3947
rect 13262 3913 13280 3947
rect 13220 3887 13280 3913
rect 13310 3947 13380 3973
rect 13310 3913 13328 3947
rect 13362 3913 13380 3947
rect 13310 3887 13380 3913
rect 13410 3947 13480 3973
rect 13410 3913 13428 3947
rect 13462 3913 13480 3947
rect 13410 3887 13480 3913
rect 13510 3947 13580 3973
rect 13510 3913 13528 3947
rect 13562 3913 13580 3947
rect 13510 3887 13580 3913
rect 13610 3947 13670 3973
rect 13610 3913 13628 3947
rect 13662 3913 13670 3947
rect 13610 3887 13670 3913
rect 10116 3807 10170 3833
rect 10116 3773 10124 3807
rect 10158 3773 10170 3807
rect 10116 3747 10170 3773
rect 10200 3807 10270 3833
rect 10200 3773 10218 3807
rect 10252 3773 10270 3807
rect 10200 3747 10270 3773
rect 10300 3747 10370 3833
rect 10400 3807 10470 3833
rect 10400 3773 10418 3807
rect 10452 3773 10470 3807
rect 10400 3747 10470 3773
rect 10500 3807 10570 3833
rect 10500 3773 10518 3807
rect 10552 3773 10570 3807
rect 10500 3747 10570 3773
rect 10600 3807 10670 3833
rect 10600 3773 10618 3807
rect 10652 3773 10670 3807
rect 10600 3747 10670 3773
rect 10700 3807 10770 3833
rect 10700 3773 10718 3807
rect 10752 3773 10770 3807
rect 10700 3747 10770 3773
rect 10800 3807 10870 3833
rect 10800 3773 10818 3807
rect 10852 3773 10870 3807
rect 10800 3747 10870 3773
rect 10900 3807 10970 3833
rect 10900 3773 10918 3807
rect 10952 3773 10970 3807
rect 10900 3747 10970 3773
rect 11000 3807 11070 3833
rect 11000 3773 11018 3807
rect 11052 3773 11070 3807
rect 11000 3747 11070 3773
rect 11100 3807 11154 3833
rect 11100 3773 11112 3807
rect 11146 3773 11154 3807
rect 11100 3747 11154 3773
rect 9416 3577 9470 3603
rect 9416 3543 9424 3577
rect 9458 3543 9470 3577
rect 9416 3517 9470 3543
rect 9500 3577 9570 3603
rect 9500 3543 9518 3577
rect 9552 3543 9570 3577
rect 9500 3517 9570 3543
rect 9600 3577 9670 3603
rect 9600 3543 9618 3577
rect 9652 3543 9670 3577
rect 9600 3517 9670 3543
rect 9700 3577 9770 3603
rect 9700 3543 9718 3577
rect 9752 3543 9770 3577
rect 9700 3517 9770 3543
rect 9800 3577 9870 3603
rect 9800 3543 9818 3577
rect 9852 3543 9870 3577
rect 9800 3517 9870 3543
rect 9900 3577 9970 3603
rect 9900 3543 9918 3577
rect 9952 3543 9970 3577
rect 9900 3517 9970 3543
rect 10000 3577 10054 3603
rect 10000 3543 10012 3577
rect 10046 3543 10054 3577
rect 10000 3517 10054 3543
rect 6816 3437 6870 3463
rect 6816 3403 6824 3437
rect 6858 3403 6870 3437
rect 6816 3377 6870 3403
rect 6900 3437 6970 3463
rect 6900 3403 6918 3437
rect 6952 3403 6970 3437
rect 6900 3377 6970 3403
rect 7000 3377 7070 3463
rect 7100 3377 7170 3463
rect 7200 3377 7270 3463
rect 7300 3437 7370 3463
rect 7300 3403 7318 3437
rect 7352 3403 7370 3437
rect 7300 3377 7370 3403
rect 7400 3437 7470 3463
rect 7400 3403 7418 3437
rect 7452 3403 7470 3437
rect 7400 3377 7470 3403
rect 7500 3377 7570 3463
rect 7600 3377 7670 3463
rect 7700 3437 7770 3463
rect 7700 3403 7718 3437
rect 7752 3403 7770 3437
rect 7700 3377 7770 3403
rect 7800 3437 7870 3463
rect 7800 3403 7818 3437
rect 7852 3403 7870 3437
rect 7800 3377 7870 3403
rect 7900 3437 7970 3463
rect 7900 3403 7918 3437
rect 7952 3403 7970 3437
rect 7900 3377 7970 3403
rect 8000 3437 8070 3463
rect 8000 3403 8018 3437
rect 8052 3403 8070 3437
rect 8000 3377 8070 3403
rect 8100 3377 8170 3463
rect 8200 3377 8270 3463
rect 8300 3377 8370 3463
rect 8400 3437 8470 3463
rect 8400 3403 8418 3437
rect 8452 3403 8470 3437
rect 8400 3377 8470 3403
rect 8500 3437 8570 3463
rect 8500 3403 8518 3437
rect 8552 3403 8570 3437
rect 8500 3377 8570 3403
rect 8600 3437 8670 3463
rect 8600 3403 8618 3437
rect 8652 3403 8670 3437
rect 8600 3377 8670 3403
rect 8700 3437 8770 3463
rect 8700 3403 8718 3437
rect 8752 3403 8770 3437
rect 8700 3377 8770 3403
rect 8800 3377 8870 3463
rect 8900 3437 8970 3463
rect 8900 3403 8918 3437
rect 8952 3403 8970 3437
rect 8900 3377 8970 3403
rect 9000 3437 9070 3463
rect 9000 3403 9018 3437
rect 9052 3403 9070 3437
rect 9000 3377 9070 3403
rect 9100 3437 9170 3463
rect 9100 3403 9118 3437
rect 9152 3403 9170 3437
rect 9100 3377 9170 3403
rect 9200 3437 9270 3463
rect 9200 3403 9218 3437
rect 9252 3403 9270 3437
rect 9200 3377 9270 3403
rect 9300 3437 9370 3463
rect 9300 3403 9318 3437
rect 9352 3403 9370 3437
rect 9300 3377 9370 3403
rect 9400 3437 9454 3463
rect 9400 3403 9412 3437
rect 9446 3403 9454 3437
rect 9400 3377 9454 3403
rect 3516 3297 3570 3323
rect 3516 3263 3524 3297
rect 3558 3263 3570 3297
rect 3516 3237 3570 3263
rect 3600 3297 3670 3323
rect 3600 3263 3618 3297
rect 3652 3263 3670 3297
rect 3600 3237 3670 3263
rect 3700 3237 3770 3323
rect 3800 3237 3870 3323
rect 3900 3237 3970 3323
rect 4000 3237 4070 3323
rect 4100 3297 4170 3323
rect 4100 3263 4118 3297
rect 4152 3263 4170 3297
rect 4100 3237 4170 3263
rect 4200 3297 4270 3323
rect 4200 3263 4218 3297
rect 4252 3263 4270 3297
rect 4200 3237 4270 3263
rect 4300 3297 4370 3323
rect 4300 3263 4318 3297
rect 4352 3263 4370 3297
rect 4300 3237 4370 3263
rect 4400 3297 4470 3323
rect 4400 3263 4418 3297
rect 4452 3263 4470 3297
rect 4400 3237 4470 3263
rect 4500 3237 4570 3323
rect 4600 3237 4670 3323
rect 4700 3297 4770 3323
rect 4700 3263 4718 3297
rect 4752 3263 4770 3297
rect 4700 3237 4770 3263
rect 4800 3297 4870 3323
rect 4800 3263 4818 3297
rect 4852 3263 4870 3297
rect 4800 3237 4870 3263
rect 4900 3237 4970 3323
rect 5000 3297 5070 3323
rect 5000 3263 5018 3297
rect 5052 3263 5070 3297
rect 5000 3237 5070 3263
rect 5100 3297 5170 3323
rect 5100 3263 5118 3297
rect 5152 3263 5170 3297
rect 5100 3237 5170 3263
rect 5200 3297 5270 3323
rect 5200 3263 5218 3297
rect 5252 3263 5270 3297
rect 5200 3237 5270 3263
rect 5300 3237 5370 3323
rect 5400 3297 5470 3323
rect 5400 3263 5418 3297
rect 5452 3263 5470 3297
rect 5400 3237 5470 3263
rect 5500 3297 5570 3323
rect 5500 3263 5518 3297
rect 5552 3263 5570 3297
rect 5500 3237 5570 3263
rect 5600 3297 5670 3323
rect 5600 3263 5618 3297
rect 5652 3263 5670 3297
rect 5600 3237 5670 3263
rect 5700 3237 5770 3323
rect 5800 3297 5870 3323
rect 5800 3263 5818 3297
rect 5852 3263 5870 3297
rect 5800 3237 5870 3263
rect 5900 3297 5970 3323
rect 5900 3263 5918 3297
rect 5952 3263 5970 3297
rect 5900 3237 5970 3263
rect 6000 3297 6070 3323
rect 6000 3263 6018 3297
rect 6052 3263 6070 3297
rect 6000 3237 6070 3263
rect 6100 3237 6170 3323
rect 6200 3237 6270 3323
rect 6300 3297 6370 3323
rect 6300 3263 6318 3297
rect 6352 3263 6370 3297
rect 6300 3237 6370 3263
rect 6400 3297 6470 3323
rect 6400 3263 6418 3297
rect 6452 3263 6470 3297
rect 6400 3237 6470 3263
rect 6500 3297 6570 3323
rect 6500 3263 6518 3297
rect 6552 3263 6570 3297
rect 6500 3237 6570 3263
rect 6600 3297 6670 3323
rect 6600 3263 6618 3297
rect 6652 3263 6670 3297
rect 6600 3237 6670 3263
rect 6700 3297 6770 3323
rect 6700 3263 6718 3297
rect 6752 3263 6770 3297
rect 6700 3237 6770 3263
rect 6800 3297 6870 3323
rect 6800 3263 6818 3297
rect 6852 3263 6870 3297
rect 6800 3237 6870 3263
rect 6900 3237 6970 3323
rect 7000 3237 7070 3323
rect 7100 3297 7170 3323
rect 7100 3263 7118 3297
rect 7152 3263 7170 3297
rect 7100 3237 7170 3263
rect 7200 3297 7270 3323
rect 7200 3263 7218 3297
rect 7252 3263 7270 3297
rect 7200 3237 7270 3263
rect 7300 3297 7354 3323
rect 7300 3263 7312 3297
rect 7346 3263 7354 3297
rect 7300 3237 7354 3263
rect 3316 3157 3370 3183
rect 3316 3123 3324 3157
rect 3358 3123 3370 3157
rect 3316 3097 3370 3123
rect 3400 3157 3470 3183
rect 3400 3123 3418 3157
rect 3452 3123 3470 3157
rect 3400 3097 3470 3123
rect 3500 3157 3570 3183
rect 3500 3123 3518 3157
rect 3552 3123 3570 3157
rect 3500 3097 3570 3123
rect 3600 3157 3654 3183
rect 3600 3123 3612 3157
rect 3646 3123 3654 3157
rect 3600 3097 3654 3123
rect 3716 3157 3770 3183
rect 3716 3123 3724 3157
rect 3758 3123 3770 3157
rect 3716 3097 3770 3123
rect 3800 3157 3870 3183
rect 3800 3123 3818 3157
rect 3852 3123 3870 3157
rect 3800 3097 3870 3123
rect 3900 3157 3970 3183
rect 3900 3123 3918 3157
rect 3952 3123 3970 3157
rect 3900 3097 3970 3123
rect 4000 3157 4070 3183
rect 4000 3123 4018 3157
rect 4052 3123 4070 3157
rect 4000 3097 4070 3123
rect 4100 3157 4170 3183
rect 4100 3123 4118 3157
rect 4152 3123 4170 3157
rect 4100 3097 4170 3123
rect 4200 3157 4270 3183
rect 4200 3123 4218 3157
rect 4252 3123 4270 3157
rect 4200 3097 4270 3123
rect 4300 3157 4370 3183
rect 4300 3123 4318 3157
rect 4352 3123 4370 3157
rect 4300 3097 4370 3123
rect 4400 3097 4470 3183
rect 4500 3157 4570 3183
rect 4500 3123 4518 3157
rect 4552 3123 4570 3157
rect 4500 3097 4570 3123
rect 4600 3157 4670 3183
rect 4600 3123 4618 3157
rect 4652 3123 4670 3157
rect 4600 3097 4670 3123
rect 4700 3157 4770 3183
rect 4700 3123 4718 3157
rect 4752 3123 4770 3157
rect 4700 3097 4770 3123
rect 4800 3097 4870 3183
rect 4900 3097 4970 3183
rect 5000 3097 5070 3183
rect 5100 3097 5170 3183
rect 5200 3157 5270 3183
rect 5200 3123 5218 3157
rect 5252 3123 5270 3157
rect 5200 3097 5270 3123
rect 5300 3157 5370 3183
rect 5300 3123 5318 3157
rect 5352 3123 5370 3157
rect 5300 3097 5370 3123
rect 5400 3157 5454 3183
rect 5400 3123 5412 3157
rect 5446 3123 5454 3157
rect 5400 3097 5454 3123
rect 3116 3017 3170 3043
rect 3116 2983 3124 3017
rect 3158 2983 3170 3017
rect 3116 2957 3170 2983
rect 3200 3017 3270 3043
rect 3200 2983 3218 3017
rect 3252 2983 3270 3017
rect 3200 2957 3270 2983
rect 3300 3017 3370 3043
rect 3300 2983 3318 3017
rect 3352 2983 3370 3017
rect 3300 2957 3370 2983
rect 3400 3017 3470 3043
rect 3400 2983 3418 3017
rect 3452 2983 3470 3017
rect 3400 2957 3470 2983
rect 3500 2957 3570 3043
rect 3600 2957 3670 3043
rect 3700 3017 3770 3043
rect 3700 2983 3718 3017
rect 3752 2983 3770 3017
rect 3700 2957 3770 2983
rect 3800 3017 3854 3043
rect 3800 2983 3812 3017
rect 3846 2983 3854 3017
rect 3800 2957 3854 2983
rect 3016 2877 3070 2903
rect 3016 2843 3024 2877
rect 3058 2843 3070 2877
rect 3016 2817 3070 2843
rect 3100 2877 3170 2903
rect 3100 2843 3118 2877
rect 3152 2843 3170 2877
rect 3100 2817 3170 2843
rect 3200 2877 3270 2903
rect 3200 2843 3218 2877
rect 3252 2843 3270 2877
rect 3200 2817 3270 2843
rect 3300 2877 3354 2903
rect 3300 2843 3312 2877
rect 3346 2843 3354 2877
rect 3300 2817 3354 2843
rect 3916 3017 3970 3043
rect 3916 2983 3924 3017
rect 3958 2983 3970 3017
rect 3916 2957 3970 2983
rect 4000 3017 4070 3043
rect 4000 2983 4018 3017
rect 4052 2983 4070 3017
rect 4000 2957 4070 2983
rect 4100 3017 4170 3043
rect 4100 2983 4118 3017
rect 4152 2983 4170 3017
rect 4100 2957 4170 2983
rect 4200 3017 4270 3043
rect 4200 2983 4218 3017
rect 4252 2983 4270 3017
rect 4200 2957 4270 2983
rect 4300 2957 4370 3043
rect 4400 3017 4470 3043
rect 4400 2983 4418 3017
rect 4452 2983 4470 3017
rect 4400 2957 4470 2983
rect 4500 3017 4554 3043
rect 4500 2983 4512 3017
rect 4546 2983 4554 3017
rect 4500 2957 4554 2983
rect 3416 2877 3470 2903
rect 3416 2843 3424 2877
rect 3458 2843 3470 2877
rect 3416 2817 3470 2843
rect 3500 2877 3570 2903
rect 3500 2843 3518 2877
rect 3552 2843 3570 2877
rect 3500 2817 3570 2843
rect 3600 2877 3670 2903
rect 3600 2843 3618 2877
rect 3652 2843 3670 2877
rect 3600 2817 3670 2843
rect 3700 2877 3770 2903
rect 3700 2843 3718 2877
rect 3752 2843 3770 2877
rect 3700 2817 3770 2843
rect 3800 2877 3870 2903
rect 3800 2843 3818 2877
rect 3852 2843 3870 2877
rect 3800 2817 3870 2843
rect 3900 2877 3954 2903
rect 3900 2843 3912 2877
rect 3946 2843 3954 2877
rect 3900 2817 3954 2843
rect 4616 3017 4670 3043
rect 4616 2983 4624 3017
rect 4658 2983 4670 3017
rect 4616 2957 4670 2983
rect 4700 3017 4770 3043
rect 4700 2983 4718 3017
rect 4752 2983 4770 3017
rect 4700 2957 4770 2983
rect 4800 3017 4870 3043
rect 4800 2983 4818 3017
rect 4852 2983 4870 3017
rect 4800 2957 4870 2983
rect 4900 3017 4954 3043
rect 4900 2983 4912 3017
rect 4946 2983 4954 3017
rect 4900 2957 4954 2983
rect 5516 3157 5570 3183
rect 5516 3123 5524 3157
rect 5558 3123 5570 3157
rect 5516 3097 5570 3123
rect 5600 3157 5654 3183
rect 5600 3123 5612 3157
rect 5646 3123 5654 3157
rect 5600 3097 5654 3123
rect 5716 3157 5770 3183
rect 5716 3123 5724 3157
rect 5758 3123 5770 3157
rect 5716 3097 5770 3123
rect 5800 3157 5854 3183
rect 5800 3123 5812 3157
rect 5846 3123 5854 3157
rect 5800 3097 5854 3123
rect 5916 3157 5970 3183
rect 5916 3123 5924 3157
rect 5958 3123 5970 3157
rect 5916 3097 5970 3123
rect 6000 3157 6070 3183
rect 6000 3123 6018 3157
rect 6052 3123 6070 3157
rect 6000 3097 6070 3123
rect 6100 3097 6170 3183
rect 6200 3157 6270 3183
rect 6200 3123 6218 3157
rect 6252 3123 6270 3157
rect 6200 3097 6270 3123
rect 6300 3157 6354 3183
rect 6300 3123 6312 3157
rect 6346 3123 6354 3157
rect 6300 3097 6354 3123
rect 5016 3017 5070 3043
rect 5016 2983 5024 3017
rect 5058 2983 5070 3017
rect 5016 2957 5070 2983
rect 5100 3017 5170 3043
rect 5100 2983 5118 3017
rect 5152 2983 5170 3017
rect 5100 2957 5170 2983
rect 5200 2957 5270 3043
rect 5300 2957 5370 3043
rect 5400 3017 5470 3043
rect 5400 2983 5418 3017
rect 5452 2983 5470 3017
rect 5400 2957 5470 2983
rect 5500 3017 5570 3043
rect 5500 2983 5518 3017
rect 5552 2983 5570 3017
rect 5500 2957 5570 2983
rect 5600 2957 5670 3043
rect 5700 2957 5770 3043
rect 5800 3017 5870 3043
rect 5800 2983 5818 3017
rect 5852 2983 5870 3017
rect 5800 2957 5870 2983
rect 5900 3017 5954 3043
rect 5900 2983 5912 3017
rect 5946 2983 5954 3017
rect 5900 2957 5954 2983
rect 4016 2877 4070 2903
rect 4016 2843 4024 2877
rect 4058 2843 4070 2877
rect 4016 2817 4070 2843
rect 4100 2877 4170 2903
rect 4100 2843 4118 2877
rect 4152 2843 4170 2877
rect 4100 2817 4170 2843
rect 4200 2877 4270 2903
rect 4200 2843 4218 2877
rect 4252 2843 4270 2877
rect 4200 2817 4270 2843
rect 4300 2817 4370 2903
rect 4400 2877 4470 2903
rect 4400 2843 4418 2877
rect 4452 2843 4470 2877
rect 4400 2817 4470 2843
rect 4500 2877 4570 2903
rect 4500 2843 4518 2877
rect 4552 2843 4570 2877
rect 4500 2817 4570 2843
rect 4600 2817 4670 2903
rect 4700 2817 4770 2903
rect 4800 2817 4870 2903
rect 4900 2817 4970 2903
rect 5000 2817 5070 2903
rect 5100 2817 5170 2903
rect 5200 2877 5270 2903
rect 5200 2843 5218 2877
rect 5252 2843 5270 2877
rect 5200 2817 5270 2843
rect 5300 2877 5354 2903
rect 5300 2843 5312 2877
rect 5346 2843 5354 2877
rect 5300 2817 5354 2843
rect 2416 2737 2470 2763
rect 2416 2703 2424 2737
rect 2458 2703 2470 2737
rect 2416 2677 2470 2703
rect 2500 2737 2570 2763
rect 2500 2703 2518 2737
rect 2552 2703 2570 2737
rect 2500 2677 2570 2703
rect 2600 2737 2670 2763
rect 2600 2703 2618 2737
rect 2652 2703 2670 2737
rect 2600 2677 2670 2703
rect 2700 2737 2770 2763
rect 2700 2703 2718 2737
rect 2752 2703 2770 2737
rect 2700 2677 2770 2703
rect 2800 2677 2870 2763
rect 2900 2677 2970 2763
rect 3000 2737 3070 2763
rect 3000 2703 3018 2737
rect 3052 2703 3070 2737
rect 3000 2677 3070 2703
rect 3100 2737 3170 2763
rect 3100 2703 3118 2737
rect 3152 2703 3170 2737
rect 3100 2677 3170 2703
rect 3200 2737 3270 2763
rect 3200 2703 3218 2737
rect 3252 2703 3270 2737
rect 3200 2677 3270 2703
rect 3300 2737 3370 2763
rect 3300 2703 3318 2737
rect 3352 2703 3370 2737
rect 3300 2677 3370 2703
rect 3400 2677 3470 2763
rect 3500 2737 3570 2763
rect 3500 2703 3518 2737
rect 3552 2703 3570 2737
rect 3500 2677 3570 2703
rect 3600 2737 3670 2763
rect 3600 2703 3618 2737
rect 3652 2703 3670 2737
rect 3600 2677 3670 2703
rect 3700 2677 3770 2763
rect 3800 2677 3870 2763
rect 3900 2737 3970 2763
rect 3900 2703 3918 2737
rect 3952 2703 3970 2737
rect 3900 2677 3970 2703
rect 4000 2737 4070 2763
rect 4000 2703 4018 2737
rect 4052 2703 4070 2737
rect 4000 2677 4070 2703
rect 4100 2737 4154 2763
rect 4100 2703 4112 2737
rect 4146 2703 4154 2737
rect 4100 2677 4154 2703
rect 16 2537 70 2623
rect 100 2597 170 2623
rect 100 2563 118 2597
rect 152 2563 170 2597
rect 100 2537 170 2563
rect 200 2597 270 2623
rect 200 2563 218 2597
rect 252 2563 270 2597
rect 200 2537 270 2563
rect 300 2537 370 2623
rect 400 2597 470 2623
rect 400 2563 418 2597
rect 452 2563 470 2597
rect 400 2537 470 2563
rect 500 2597 570 2623
rect 500 2563 518 2597
rect 552 2563 570 2597
rect 500 2537 570 2563
rect 600 2597 670 2623
rect 600 2563 618 2597
rect 652 2563 670 2597
rect 600 2537 670 2563
rect 700 2597 770 2623
rect 700 2563 718 2597
rect 752 2563 770 2597
rect 700 2537 770 2563
rect 800 2537 870 2623
rect 900 2537 970 2623
rect 1000 2597 1070 2623
rect 1000 2563 1018 2597
rect 1052 2563 1070 2597
rect 1000 2537 1070 2563
rect 1100 2597 1170 2623
rect 1100 2563 1118 2597
rect 1152 2563 1170 2597
rect 1100 2537 1170 2563
rect 1200 2597 1270 2623
rect 1200 2563 1218 2597
rect 1252 2563 1270 2597
rect 1200 2537 1270 2563
rect 1300 2597 1370 2623
rect 1300 2563 1318 2597
rect 1352 2563 1370 2597
rect 1300 2537 1370 2563
rect 1400 2597 1470 2623
rect 1400 2563 1418 2597
rect 1452 2563 1470 2597
rect 1400 2537 1470 2563
rect 1500 2597 1570 2623
rect 1500 2563 1518 2597
rect 1552 2563 1570 2597
rect 1500 2537 1570 2563
rect 1600 2597 1670 2623
rect 1600 2563 1618 2597
rect 1652 2563 1670 2597
rect 1600 2537 1670 2563
rect 1700 2537 1770 2623
rect 1800 2597 1870 2623
rect 1800 2563 1818 2597
rect 1852 2563 1870 2597
rect 1800 2537 1870 2563
rect 1900 2597 1970 2623
rect 1900 2563 1918 2597
rect 1952 2563 1970 2597
rect 1900 2537 1970 2563
rect 2000 2597 2070 2623
rect 2000 2563 2018 2597
rect 2052 2563 2070 2597
rect 2000 2537 2070 2563
rect 2100 2537 2170 2623
rect 2200 2537 2270 2623
rect 2300 2597 2370 2623
rect 2300 2563 2318 2597
rect 2352 2563 2370 2597
rect 2300 2537 2370 2563
rect 2400 2597 2470 2623
rect 2400 2563 2418 2597
rect 2452 2563 2470 2597
rect 2400 2537 2470 2563
rect 2500 2597 2554 2623
rect 2500 2563 2512 2597
rect 2546 2563 2554 2597
rect 2500 2537 2554 2563
rect 16 2367 70 2393
rect 16 2333 24 2367
rect 58 2333 70 2367
rect 16 2307 70 2333
rect 100 2367 154 2393
rect 100 2333 112 2367
rect 146 2333 154 2367
rect 100 2307 154 2333
rect 216 2367 270 2393
rect 216 2333 224 2367
rect 258 2333 270 2367
rect 216 2307 270 2333
rect 300 2367 370 2393
rect 300 2333 318 2367
rect 352 2333 370 2367
rect 300 2307 370 2333
rect 400 2367 454 2393
rect 400 2333 412 2367
rect 446 2333 454 2367
rect 400 2307 454 2333
rect 516 2367 570 2393
rect 516 2333 524 2367
rect 558 2333 570 2367
rect 516 2307 570 2333
rect 600 2367 654 2393
rect 600 2333 612 2367
rect 646 2333 654 2367
rect 600 2307 654 2333
rect 716 2367 770 2393
rect 716 2333 724 2367
rect 758 2333 770 2367
rect 716 2307 770 2333
rect 800 2367 870 2393
rect 800 2333 818 2367
rect 852 2333 870 2367
rect 800 2307 870 2333
rect 900 2367 970 2393
rect 900 2333 918 2367
rect 952 2333 970 2367
rect 900 2307 970 2333
rect 1000 2307 1070 2393
rect 1100 2307 1170 2393
rect 1200 2307 1270 2393
rect 1300 2307 1370 2393
rect 1400 2367 1470 2393
rect 1400 2333 1418 2367
rect 1452 2333 1470 2367
rect 1400 2307 1470 2333
rect 1500 2367 1570 2393
rect 1500 2333 1518 2367
rect 1552 2333 1570 2367
rect 1500 2307 1570 2333
rect 1600 2307 1670 2393
rect 1700 2367 1770 2393
rect 1700 2333 1718 2367
rect 1752 2333 1770 2367
rect 1700 2307 1770 2333
rect 1800 2367 1870 2393
rect 1800 2333 1818 2367
rect 1852 2333 1870 2367
rect 1800 2307 1870 2333
rect 1900 2307 1970 2393
rect 2000 2367 2070 2393
rect 2000 2333 2018 2367
rect 2052 2333 2070 2367
rect 2000 2307 2070 2333
rect 2100 2367 2170 2393
rect 2100 2333 2118 2367
rect 2152 2333 2170 2367
rect 2100 2307 2170 2333
rect 2200 2367 2270 2393
rect 2200 2333 2218 2367
rect 2252 2333 2270 2367
rect 2200 2307 2270 2333
rect 2300 2367 2354 2393
rect 2300 2333 2312 2367
rect 2346 2333 2354 2367
rect 2300 2307 2354 2333
rect 16 2227 70 2253
rect 16 2193 24 2227
rect 58 2193 70 2227
rect 16 2167 70 2193
rect 100 2227 170 2253
rect 100 2193 118 2227
rect 152 2193 170 2227
rect 100 2167 170 2193
rect 200 2167 270 2253
rect 300 2227 370 2253
rect 300 2193 318 2227
rect 352 2193 370 2227
rect 300 2167 370 2193
rect 400 2227 470 2253
rect 400 2193 418 2227
rect 452 2193 470 2227
rect 400 2167 470 2193
rect 500 2227 570 2253
rect 500 2193 518 2227
rect 552 2193 570 2227
rect 500 2167 570 2193
rect 600 2167 670 2253
rect 700 2227 770 2253
rect 700 2193 718 2227
rect 752 2193 770 2227
rect 700 2167 770 2193
rect 800 2227 854 2253
rect 800 2193 812 2227
rect 846 2193 854 2227
rect 800 2167 854 2193
rect 16 2027 70 2113
rect 100 2027 170 2113
rect 200 2027 270 2113
rect 300 2087 370 2113
rect 300 2053 318 2087
rect 352 2053 370 2087
rect 300 2027 370 2053
rect 400 2087 470 2113
rect 400 2053 418 2087
rect 452 2053 470 2087
rect 400 2027 470 2053
rect 500 2087 570 2113
rect 500 2053 518 2087
rect 552 2053 570 2087
rect 500 2027 570 2053
rect 600 2087 670 2113
rect 600 2053 618 2087
rect 652 2053 670 2087
rect 600 2027 670 2053
rect 700 2087 754 2113
rect 700 2053 712 2087
rect 746 2053 754 2087
rect 700 2027 754 2053
rect 916 2227 970 2253
rect 916 2193 924 2227
rect 958 2193 970 2227
rect 916 2167 970 2193
rect 1000 2227 1054 2253
rect 1000 2193 1012 2227
rect 1046 2193 1054 2227
rect 1000 2167 1054 2193
rect 2616 2597 2670 2623
rect 2616 2563 2624 2597
rect 2658 2563 2670 2597
rect 2616 2537 2670 2563
rect 2700 2597 2770 2623
rect 2700 2563 2718 2597
rect 2752 2563 2770 2597
rect 2700 2537 2770 2563
rect 2800 2597 2870 2623
rect 2800 2563 2818 2597
rect 2852 2563 2870 2597
rect 2800 2537 2870 2563
rect 2900 2597 2970 2623
rect 2900 2563 2918 2597
rect 2952 2563 2970 2597
rect 2900 2537 2970 2563
rect 3000 2597 3070 2623
rect 3000 2563 3018 2597
rect 3052 2563 3070 2597
rect 3000 2537 3070 2563
rect 3100 2597 3170 2623
rect 3100 2563 3118 2597
rect 3152 2563 3170 2597
rect 3100 2537 3170 2563
rect 3200 2597 3270 2623
rect 3200 2563 3218 2597
rect 3252 2563 3270 2597
rect 3200 2537 3270 2563
rect 3300 2597 3354 2623
rect 3300 2563 3312 2597
rect 3346 2563 3354 2597
rect 3300 2537 3354 2563
rect 2416 2367 2470 2393
rect 2416 2333 2424 2367
rect 2458 2333 2470 2367
rect 2416 2307 2470 2333
rect 2500 2367 2570 2393
rect 2500 2333 2518 2367
rect 2552 2333 2570 2367
rect 2500 2307 2570 2333
rect 2600 2367 2654 2393
rect 2600 2333 2612 2367
rect 2646 2333 2654 2367
rect 2600 2307 2654 2333
rect 1116 2227 1170 2253
rect 1116 2193 1124 2227
rect 1158 2193 1170 2227
rect 1116 2167 1170 2193
rect 1200 2227 1270 2253
rect 1200 2193 1218 2227
rect 1252 2193 1270 2227
rect 1200 2167 1270 2193
rect 1300 2227 1370 2253
rect 1300 2193 1318 2227
rect 1352 2193 1370 2227
rect 1300 2167 1370 2193
rect 1400 2167 1470 2253
rect 1500 2167 1570 2253
rect 1600 2227 1670 2253
rect 1600 2193 1618 2227
rect 1652 2193 1670 2227
rect 1600 2167 1670 2193
rect 1700 2227 1770 2253
rect 1700 2193 1718 2227
rect 1752 2193 1770 2227
rect 1700 2167 1770 2193
rect 1800 2167 1870 2253
rect 1900 2227 1970 2253
rect 1900 2193 1918 2227
rect 1952 2193 1970 2227
rect 1900 2167 1970 2193
rect 2000 2227 2070 2253
rect 2000 2193 2018 2227
rect 2052 2193 2070 2227
rect 2000 2167 2070 2193
rect 2100 2167 2170 2253
rect 2200 2167 2270 2253
rect 2300 2167 2370 2253
rect 2400 2167 2470 2253
rect 2500 2227 2570 2253
rect 2500 2193 2518 2227
rect 2552 2193 2570 2227
rect 2500 2167 2570 2193
rect 2600 2227 2654 2253
rect 2600 2193 2612 2227
rect 2646 2193 2654 2227
rect 2600 2167 2654 2193
rect 816 2087 870 2113
rect 816 2053 824 2087
rect 858 2053 870 2087
rect 816 2027 870 2053
rect 900 2087 970 2113
rect 900 2053 918 2087
rect 952 2053 970 2087
rect 900 2027 970 2053
rect 1000 2027 1070 2113
rect 1100 2027 1170 2113
rect 1200 2027 1270 2113
rect 1300 2087 1370 2113
rect 1300 2053 1318 2087
rect 1352 2053 1370 2087
rect 1300 2027 1370 2053
rect 1400 2087 1454 2113
rect 1400 2053 1412 2087
rect 1446 2053 1454 2087
rect 1400 2027 1454 2053
rect 16 1887 70 1973
rect 100 1947 170 1973
rect 100 1913 118 1947
rect 152 1913 170 1947
rect 100 1887 170 1913
rect 200 1947 270 1973
rect 200 1913 218 1947
rect 252 1913 270 1947
rect 200 1887 270 1913
rect 300 1947 370 1973
rect 300 1913 318 1947
rect 352 1913 370 1947
rect 300 1887 370 1913
rect 400 1947 470 1973
rect 400 1913 418 1947
rect 452 1913 470 1947
rect 400 1887 470 1913
rect 500 1947 570 1973
rect 500 1913 518 1947
rect 552 1913 570 1947
rect 500 1887 570 1913
rect 600 1947 670 1973
rect 600 1913 618 1947
rect 652 1913 670 1947
rect 600 1887 670 1913
rect 700 1947 770 1973
rect 700 1913 718 1947
rect 752 1913 770 1947
rect 700 1887 770 1913
rect 800 1947 870 1973
rect 800 1913 818 1947
rect 852 1913 870 1947
rect 800 1887 870 1913
rect 900 1947 954 1973
rect 900 1913 912 1947
rect 946 1913 954 1947
rect 900 1887 954 1913
rect 3416 2597 3470 2623
rect 3416 2563 3424 2597
rect 3458 2563 3470 2597
rect 3416 2537 3470 2563
rect 3500 2597 3570 2623
rect 3500 2563 3518 2597
rect 3552 2563 3570 2597
rect 3500 2537 3570 2563
rect 3600 2597 3670 2623
rect 3600 2563 3618 2597
rect 3652 2563 3670 2597
rect 3600 2537 3670 2563
rect 3700 2537 3770 2623
rect 3800 2597 3870 2623
rect 3800 2563 3818 2597
rect 3852 2563 3870 2597
rect 3800 2537 3870 2563
rect 3900 2597 3954 2623
rect 3900 2563 3912 2597
rect 3946 2563 3954 2597
rect 3900 2537 3954 2563
rect 4016 2597 4070 2623
rect 4016 2563 4024 2597
rect 4058 2563 4070 2597
rect 4016 2537 4070 2563
rect 4100 2597 4154 2623
rect 4100 2563 4112 2597
rect 4146 2563 4154 2597
rect 4100 2537 4154 2563
rect 4216 2737 4270 2763
rect 4216 2703 4224 2737
rect 4258 2703 4270 2737
rect 4216 2677 4270 2703
rect 4300 2737 4370 2763
rect 4300 2703 4318 2737
rect 4352 2703 4370 2737
rect 4300 2677 4370 2703
rect 4400 2677 4470 2763
rect 4500 2737 4570 2763
rect 4500 2703 4518 2737
rect 4552 2703 4570 2737
rect 4500 2677 4570 2703
rect 4600 2737 4670 2763
rect 4600 2703 4618 2737
rect 4652 2703 4670 2737
rect 4600 2677 4670 2703
rect 4700 2737 4754 2763
rect 4700 2703 4712 2737
rect 4746 2703 4754 2737
rect 4700 2677 4754 2703
rect 4216 2597 4270 2623
rect 4216 2563 4224 2597
rect 4258 2563 4270 2597
rect 4216 2537 4270 2563
rect 4300 2597 4354 2623
rect 4300 2563 4312 2597
rect 4346 2563 4354 2597
rect 4300 2537 4354 2563
rect 4416 2597 4470 2623
rect 4416 2563 4424 2597
rect 4458 2563 4470 2597
rect 4416 2537 4470 2563
rect 4500 2597 4570 2623
rect 4500 2563 4518 2597
rect 4552 2563 4570 2597
rect 4500 2537 4570 2563
rect 4600 2597 4670 2623
rect 4600 2563 4618 2597
rect 4652 2563 4670 2597
rect 4600 2537 4670 2563
rect 4700 2597 4754 2623
rect 4700 2563 4712 2597
rect 4746 2563 4754 2597
rect 4700 2537 4754 2563
rect 4816 2737 4870 2763
rect 4816 2703 4824 2737
rect 4858 2703 4870 2737
rect 4816 2677 4870 2703
rect 4900 2737 4970 2763
rect 4900 2703 4918 2737
rect 4952 2703 4970 2737
rect 4900 2677 4970 2703
rect 5000 2737 5070 2763
rect 5000 2703 5018 2737
rect 5052 2703 5070 2737
rect 5000 2677 5070 2703
rect 5100 2737 5154 2763
rect 5100 2703 5112 2737
rect 5146 2703 5154 2737
rect 5100 2677 5154 2703
rect 5216 2737 5270 2763
rect 5216 2703 5224 2737
rect 5258 2703 5270 2737
rect 5216 2677 5270 2703
rect 5300 2737 5354 2763
rect 5300 2703 5312 2737
rect 5346 2703 5354 2737
rect 5300 2677 5354 2703
rect 6416 3157 6470 3183
rect 6416 3123 6424 3157
rect 6458 3123 6470 3157
rect 6416 3097 6470 3123
rect 6500 3157 6554 3183
rect 6500 3123 6512 3157
rect 6546 3123 6554 3157
rect 6500 3097 6554 3123
rect 6616 3157 6670 3183
rect 6616 3123 6624 3157
rect 6658 3123 6670 3157
rect 6616 3097 6670 3123
rect 6700 3157 6770 3183
rect 6700 3123 6718 3157
rect 6752 3123 6770 3157
rect 6700 3097 6770 3123
rect 6800 3157 6870 3183
rect 6800 3123 6818 3157
rect 6852 3123 6870 3157
rect 6800 3097 6870 3123
rect 6900 3157 6970 3183
rect 6900 3123 6918 3157
rect 6952 3123 6970 3157
rect 6900 3097 6970 3123
rect 7000 3157 7054 3183
rect 7000 3123 7012 3157
rect 7046 3123 7054 3157
rect 7000 3097 7054 3123
rect 9516 3437 9570 3463
rect 9516 3403 9524 3437
rect 9558 3403 9570 3437
rect 9516 3377 9570 3403
rect 9600 3437 9670 3463
rect 9600 3403 9618 3437
rect 9652 3403 9670 3437
rect 9600 3377 9670 3403
rect 9700 3437 9754 3463
rect 9700 3403 9712 3437
rect 9746 3403 9754 3437
rect 9700 3377 9754 3403
rect 7416 3297 7470 3323
rect 7416 3263 7424 3297
rect 7458 3263 7470 3297
rect 7416 3237 7470 3263
rect 7500 3297 7570 3323
rect 7500 3263 7518 3297
rect 7552 3263 7570 3297
rect 7500 3237 7570 3263
rect 7600 3297 7670 3323
rect 7600 3263 7618 3297
rect 7652 3263 7670 3297
rect 7600 3237 7670 3263
rect 7700 3297 7770 3323
rect 7700 3263 7718 3297
rect 7752 3263 7770 3297
rect 7700 3237 7770 3263
rect 7800 3297 7870 3323
rect 7800 3263 7818 3297
rect 7852 3263 7870 3297
rect 7800 3237 7870 3263
rect 7900 3297 7970 3323
rect 7900 3263 7918 3297
rect 7952 3263 7970 3297
rect 7900 3237 7970 3263
rect 8000 3297 8070 3323
rect 8000 3263 8018 3297
rect 8052 3263 8070 3297
rect 8000 3237 8070 3263
rect 8100 3297 8170 3323
rect 8100 3263 8118 3297
rect 8152 3263 8170 3297
rect 8100 3237 8170 3263
rect 8200 3297 8270 3323
rect 8200 3263 8218 3297
rect 8252 3263 8270 3297
rect 8200 3237 8270 3263
rect 8300 3297 8370 3323
rect 8300 3263 8318 3297
rect 8352 3263 8370 3297
rect 8300 3237 8370 3263
rect 8400 3237 8470 3323
rect 8500 3237 8570 3323
rect 8600 3297 8670 3323
rect 8600 3263 8618 3297
rect 8652 3263 8670 3297
rect 8600 3237 8670 3263
rect 8700 3297 8770 3323
rect 8700 3263 8718 3297
rect 8752 3263 8770 3297
rect 8700 3237 8770 3263
rect 8800 3237 8870 3323
rect 8900 3237 8970 3323
rect 9000 3237 9070 3323
rect 9100 3237 9170 3323
rect 9200 3297 9270 3323
rect 9200 3263 9218 3297
rect 9252 3263 9270 3297
rect 9200 3237 9270 3263
rect 9300 3297 9370 3323
rect 9300 3263 9318 3297
rect 9352 3263 9370 3297
rect 9300 3237 9370 3263
rect 9400 3297 9470 3323
rect 9400 3263 9418 3297
rect 9452 3263 9470 3297
rect 9400 3237 9470 3263
rect 9500 3297 9554 3323
rect 9500 3263 9512 3297
rect 9546 3263 9554 3297
rect 9500 3237 9554 3263
rect 7116 3157 7170 3183
rect 7116 3123 7124 3157
rect 7158 3123 7170 3157
rect 7116 3097 7170 3123
rect 7200 3157 7270 3183
rect 7200 3123 7218 3157
rect 7252 3123 7270 3157
rect 7200 3097 7270 3123
rect 7300 3097 7370 3183
rect 7400 3097 7470 3183
rect 7500 3097 7570 3183
rect 7600 3157 7670 3183
rect 7600 3123 7618 3157
rect 7652 3123 7670 3157
rect 7600 3097 7670 3123
rect 7700 3157 7770 3183
rect 7700 3123 7718 3157
rect 7752 3123 7770 3157
rect 7700 3097 7770 3123
rect 7800 3097 7870 3183
rect 7900 3157 7970 3183
rect 7900 3123 7918 3157
rect 7952 3123 7970 3157
rect 7900 3097 7970 3123
rect 8000 3157 8070 3183
rect 8000 3123 8018 3157
rect 8052 3123 8070 3157
rect 8000 3097 8070 3123
rect 8100 3157 8154 3183
rect 8100 3123 8112 3157
rect 8146 3123 8154 3157
rect 8100 3097 8154 3123
rect 6016 3017 6070 3043
rect 6016 2983 6024 3017
rect 6058 2983 6070 3017
rect 6016 2957 6070 2983
rect 6100 3017 6170 3043
rect 6100 2983 6118 3017
rect 6152 2983 6170 3017
rect 6100 2957 6170 2983
rect 6200 3017 6270 3043
rect 6200 2983 6218 3017
rect 6252 2983 6270 3017
rect 6200 2957 6270 2983
rect 6300 2957 6370 3043
rect 6400 3017 6470 3043
rect 6400 2983 6418 3017
rect 6452 2983 6470 3017
rect 6400 2957 6470 2983
rect 6500 3017 6570 3043
rect 6500 2983 6518 3017
rect 6552 2983 6570 3017
rect 6500 2957 6570 2983
rect 6600 3017 6670 3043
rect 6600 2983 6618 3017
rect 6652 2983 6670 3017
rect 6600 2957 6670 2983
rect 6700 3017 6770 3043
rect 6700 2983 6718 3017
rect 6752 2983 6770 3017
rect 6700 2957 6770 2983
rect 6800 3017 6870 3043
rect 6800 2983 6818 3017
rect 6852 2983 6870 3017
rect 6800 2957 6870 2983
rect 6900 3017 6970 3043
rect 6900 2983 6918 3017
rect 6952 2983 6970 3017
rect 6900 2957 6970 2983
rect 7000 3017 7070 3043
rect 7000 2983 7018 3017
rect 7052 2983 7070 3017
rect 7000 2957 7070 2983
rect 7100 2957 7170 3043
rect 7200 2957 7270 3043
rect 7300 2957 7370 3043
rect 7400 2957 7470 3043
rect 7500 3017 7570 3043
rect 7500 2983 7518 3017
rect 7552 2983 7570 3017
rect 7500 2957 7570 2983
rect 7600 3017 7670 3043
rect 7600 2983 7618 3017
rect 7652 2983 7670 3017
rect 7600 2957 7670 2983
rect 7700 3017 7770 3043
rect 7700 2983 7718 3017
rect 7752 2983 7770 3017
rect 7700 2957 7770 2983
rect 7800 3017 7870 3043
rect 7800 2983 7818 3017
rect 7852 2983 7870 3017
rect 7800 2957 7870 2983
rect 7900 3017 7970 3043
rect 7900 2983 7918 3017
rect 7952 2983 7970 3017
rect 7900 2957 7970 2983
rect 8000 3017 8054 3043
rect 8000 2983 8012 3017
rect 8046 2983 8054 3017
rect 8000 2957 8054 2983
rect 5416 2877 5470 2903
rect 5416 2843 5424 2877
rect 5458 2843 5470 2877
rect 5416 2817 5470 2843
rect 5500 2877 5570 2903
rect 5500 2843 5518 2877
rect 5552 2843 5570 2877
rect 5500 2817 5570 2843
rect 5600 2877 5670 2903
rect 5600 2843 5618 2877
rect 5652 2843 5670 2877
rect 5600 2817 5670 2843
rect 5700 2817 5770 2903
rect 5800 2817 5870 2903
rect 5900 2877 5970 2903
rect 5900 2843 5918 2877
rect 5952 2843 5970 2877
rect 5900 2817 5970 2843
rect 6000 2877 6054 2903
rect 6000 2843 6012 2877
rect 6046 2843 6054 2877
rect 6000 2817 6054 2843
rect 5416 2737 5470 2763
rect 5416 2703 5424 2737
rect 5458 2703 5470 2737
rect 5416 2677 5470 2703
rect 5500 2737 5570 2763
rect 5500 2703 5518 2737
rect 5552 2703 5570 2737
rect 5500 2677 5570 2703
rect 5600 2737 5670 2763
rect 5600 2703 5618 2737
rect 5652 2703 5670 2737
rect 5600 2677 5670 2703
rect 5700 2737 5770 2763
rect 5700 2703 5718 2737
rect 5752 2703 5770 2737
rect 5700 2677 5770 2703
rect 5800 2677 5870 2763
rect 5900 2737 5970 2763
rect 5900 2703 5918 2737
rect 5952 2703 5970 2737
rect 5900 2677 5970 2703
rect 6000 2737 6054 2763
rect 6000 2703 6012 2737
rect 6046 2703 6054 2737
rect 6000 2677 6054 2703
rect 6116 2877 6170 2903
rect 6116 2843 6124 2877
rect 6158 2843 6170 2877
rect 6116 2817 6170 2843
rect 6200 2877 6270 2903
rect 6200 2843 6218 2877
rect 6252 2843 6270 2877
rect 6200 2817 6270 2843
rect 6300 2817 6370 2903
rect 6400 2817 6470 2903
rect 6500 2817 6570 2903
rect 6600 2817 6670 2903
rect 6700 2877 6770 2903
rect 6700 2843 6718 2877
rect 6752 2843 6770 2877
rect 6700 2817 6770 2843
rect 6800 2877 6870 2903
rect 6800 2843 6818 2877
rect 6852 2843 6870 2877
rect 6800 2817 6870 2843
rect 6900 2877 6954 2903
rect 6900 2843 6912 2877
rect 6946 2843 6954 2877
rect 6900 2817 6954 2843
rect 6116 2737 6170 2763
rect 6116 2703 6124 2737
rect 6158 2703 6170 2737
rect 6116 2677 6170 2703
rect 6200 2737 6254 2763
rect 6200 2703 6212 2737
rect 6246 2703 6254 2737
rect 6200 2677 6254 2703
rect 4816 2597 4870 2623
rect 4816 2563 4824 2597
rect 4858 2563 4870 2597
rect 4816 2537 4870 2563
rect 4900 2597 4970 2623
rect 4900 2563 4918 2597
rect 4952 2563 4970 2597
rect 4900 2537 4970 2563
rect 5000 2537 5070 2623
rect 5100 2537 5170 2623
rect 5200 2537 5270 2623
rect 5300 2537 5370 2623
rect 5400 2537 5470 2623
rect 5500 2597 5570 2623
rect 5500 2563 5518 2597
rect 5552 2563 5570 2597
rect 5500 2537 5570 2563
rect 5600 2597 5670 2623
rect 5600 2563 5618 2597
rect 5652 2563 5670 2597
rect 5600 2537 5670 2563
rect 5700 2597 5770 2623
rect 5700 2563 5718 2597
rect 5752 2563 5770 2597
rect 5700 2537 5770 2563
rect 5800 2597 5870 2623
rect 5800 2563 5818 2597
rect 5852 2563 5870 2597
rect 5800 2537 5870 2563
rect 5900 2597 5970 2623
rect 5900 2563 5918 2597
rect 5952 2563 5970 2597
rect 5900 2537 5970 2563
rect 6000 2537 6070 2623
rect 6100 2597 6170 2623
rect 6100 2563 6118 2597
rect 6152 2563 6170 2597
rect 6100 2537 6170 2563
rect 6200 2597 6254 2623
rect 6200 2563 6212 2597
rect 6246 2563 6254 2597
rect 6200 2537 6254 2563
rect 6316 2737 6370 2763
rect 6316 2703 6324 2737
rect 6358 2703 6370 2737
rect 6316 2677 6370 2703
rect 6400 2737 6470 2763
rect 6400 2703 6418 2737
rect 6452 2703 6470 2737
rect 6400 2677 6470 2703
rect 6500 2737 6554 2763
rect 6500 2703 6512 2737
rect 6546 2703 6554 2737
rect 6500 2677 6554 2703
rect 7016 2877 7070 2903
rect 7016 2843 7024 2877
rect 7058 2843 7070 2877
rect 7016 2817 7070 2843
rect 7100 2877 7170 2903
rect 7100 2843 7118 2877
rect 7152 2843 7170 2877
rect 7100 2817 7170 2843
rect 7200 2877 7270 2903
rect 7200 2843 7218 2877
rect 7252 2843 7270 2877
rect 7200 2817 7270 2843
rect 7300 2877 7354 2903
rect 7300 2843 7312 2877
rect 7346 2843 7354 2877
rect 7300 2817 7354 2843
rect 7416 2877 7470 2903
rect 7416 2843 7424 2877
rect 7458 2843 7470 2877
rect 7416 2817 7470 2843
rect 7500 2877 7570 2903
rect 7500 2843 7518 2877
rect 7552 2843 7570 2877
rect 7500 2817 7570 2843
rect 7600 2877 7670 2903
rect 7600 2843 7618 2877
rect 7652 2843 7670 2877
rect 7600 2817 7670 2843
rect 7700 2877 7770 2903
rect 7700 2843 7718 2877
rect 7752 2843 7770 2877
rect 7700 2817 7770 2843
rect 7800 2877 7870 2903
rect 7800 2843 7818 2877
rect 7852 2843 7870 2877
rect 7800 2817 7870 2843
rect 7900 2877 7954 2903
rect 7900 2843 7912 2877
rect 7946 2843 7954 2877
rect 7900 2817 7954 2843
rect 8216 3157 8270 3183
rect 8216 3123 8224 3157
rect 8258 3123 8270 3157
rect 8216 3097 8270 3123
rect 8300 3157 8370 3183
rect 8300 3123 8318 3157
rect 8352 3123 8370 3157
rect 8300 3097 8370 3123
rect 8400 3157 8470 3183
rect 8400 3123 8418 3157
rect 8452 3123 8470 3157
rect 8400 3097 8470 3123
rect 8500 3097 8570 3183
rect 8600 3097 8670 3183
rect 8700 3157 8770 3183
rect 8700 3123 8718 3157
rect 8752 3123 8770 3157
rect 8700 3097 8770 3123
rect 8800 3157 8854 3183
rect 8800 3123 8812 3157
rect 8846 3123 8854 3157
rect 8800 3097 8854 3123
rect 8116 3017 8170 3043
rect 8116 2983 8124 3017
rect 8158 2983 8170 3017
rect 8116 2957 8170 2983
rect 8200 3017 8270 3043
rect 8200 2983 8218 3017
rect 8252 2983 8270 3017
rect 8200 2957 8270 2983
rect 8300 3017 8370 3043
rect 8300 2983 8318 3017
rect 8352 2983 8370 3017
rect 8300 2957 8370 2983
rect 8400 2957 8470 3043
rect 8500 2957 8570 3043
rect 8600 3017 8670 3043
rect 8600 2983 8618 3017
rect 8652 2983 8670 3017
rect 8600 2957 8670 2983
rect 8700 3017 8770 3043
rect 8700 2983 8718 3017
rect 8752 2983 8770 3017
rect 8700 2957 8770 2983
rect 8800 3017 8854 3043
rect 8800 2983 8812 3017
rect 8846 2983 8854 3017
rect 8800 2957 8854 2983
rect 8016 2877 8070 2903
rect 8016 2843 8024 2877
rect 8058 2843 8070 2877
rect 8016 2817 8070 2843
rect 8100 2877 8170 2903
rect 8100 2843 8118 2877
rect 8152 2843 8170 2877
rect 8100 2817 8170 2843
rect 8200 2877 8270 2903
rect 8200 2843 8218 2877
rect 8252 2843 8270 2877
rect 8200 2817 8270 2843
rect 8300 2817 8370 2903
rect 8400 2817 8470 2903
rect 8500 2817 8570 2903
rect 8600 2877 8670 2903
rect 8600 2843 8618 2877
rect 8652 2843 8670 2877
rect 8600 2817 8670 2843
rect 8700 2877 8754 2903
rect 8700 2843 8712 2877
rect 8746 2843 8754 2877
rect 8700 2817 8754 2843
rect 6616 2737 6670 2763
rect 6616 2703 6624 2737
rect 6658 2703 6670 2737
rect 6616 2677 6670 2703
rect 6700 2737 6770 2763
rect 6700 2703 6718 2737
rect 6752 2703 6770 2737
rect 6700 2677 6770 2703
rect 6800 2737 6870 2763
rect 6800 2703 6818 2737
rect 6852 2703 6870 2737
rect 6800 2677 6870 2703
rect 6900 2737 6970 2763
rect 6900 2703 6918 2737
rect 6952 2703 6970 2737
rect 6900 2677 6970 2703
rect 7000 2677 7070 2763
rect 7100 2737 7170 2763
rect 7100 2703 7118 2737
rect 7152 2703 7170 2737
rect 7100 2677 7170 2703
rect 7200 2737 7270 2763
rect 7200 2703 7218 2737
rect 7252 2703 7270 2737
rect 7200 2677 7270 2703
rect 7300 2677 7370 2763
rect 7400 2677 7470 2763
rect 7500 2737 7570 2763
rect 7500 2703 7518 2737
rect 7552 2703 7570 2737
rect 7500 2677 7570 2703
rect 7600 2737 7670 2763
rect 7600 2703 7618 2737
rect 7652 2703 7670 2737
rect 7600 2677 7670 2703
rect 7700 2677 7770 2763
rect 7800 2677 7870 2763
rect 7900 2677 7970 2763
rect 8000 2737 8070 2763
rect 8000 2703 8018 2737
rect 8052 2703 8070 2737
rect 8000 2677 8070 2703
rect 8100 2737 8170 2763
rect 8100 2703 8118 2737
rect 8152 2703 8170 2737
rect 8100 2677 8170 2703
rect 8200 2737 8254 2763
rect 8200 2703 8212 2737
rect 8246 2703 8254 2737
rect 8200 2677 8254 2703
rect 6316 2597 6370 2623
rect 6316 2563 6324 2597
rect 6358 2563 6370 2597
rect 6316 2537 6370 2563
rect 6400 2597 6470 2623
rect 6400 2563 6418 2597
rect 6452 2563 6470 2597
rect 6400 2537 6470 2563
rect 6500 2537 6570 2623
rect 6600 2597 6670 2623
rect 6600 2563 6618 2597
rect 6652 2563 6670 2597
rect 6600 2537 6670 2563
rect 6700 2597 6754 2623
rect 6700 2563 6712 2597
rect 6746 2563 6754 2597
rect 6700 2537 6754 2563
rect 6816 2597 6870 2623
rect 6816 2563 6824 2597
rect 6858 2563 6870 2597
rect 6816 2537 6870 2563
rect 6900 2597 6970 2623
rect 6900 2563 6918 2597
rect 6952 2563 6970 2597
rect 6900 2537 6970 2563
rect 7000 2537 7070 2623
rect 7100 2597 7170 2623
rect 7100 2563 7118 2597
rect 7152 2563 7170 2597
rect 7100 2537 7170 2563
rect 7200 2597 7270 2623
rect 7200 2563 7218 2597
rect 7252 2563 7270 2597
rect 7200 2537 7270 2563
rect 7300 2537 7370 2623
rect 7400 2597 7470 2623
rect 7400 2563 7418 2597
rect 7452 2563 7470 2597
rect 7400 2537 7470 2563
rect 7500 2597 7570 2623
rect 7500 2563 7518 2597
rect 7552 2563 7570 2597
rect 7500 2537 7570 2563
rect 7600 2537 7670 2623
rect 7700 2537 7770 2623
rect 7800 2537 7870 2623
rect 7900 2537 7970 2623
rect 8000 2597 8070 2623
rect 8000 2563 8018 2597
rect 8052 2563 8070 2597
rect 8000 2537 8070 2563
rect 8100 2597 8170 2623
rect 8100 2563 8118 2597
rect 8152 2563 8170 2597
rect 8100 2537 8170 2563
rect 8200 2597 8254 2623
rect 8200 2563 8212 2597
rect 8246 2563 8254 2597
rect 8200 2537 8254 2563
rect 2716 2367 2770 2393
rect 2716 2333 2724 2367
rect 2758 2333 2770 2367
rect 2716 2307 2770 2333
rect 2800 2367 2870 2393
rect 2800 2333 2818 2367
rect 2852 2333 2870 2367
rect 2800 2307 2870 2333
rect 2900 2367 2970 2393
rect 2900 2333 2918 2367
rect 2952 2333 2970 2367
rect 2900 2307 2970 2333
rect 3000 2307 3070 2393
rect 3100 2367 3170 2393
rect 3100 2333 3118 2367
rect 3152 2333 3170 2367
rect 3100 2307 3170 2333
rect 3200 2367 3270 2393
rect 3200 2333 3218 2367
rect 3252 2333 3270 2367
rect 3200 2307 3270 2333
rect 3300 2307 3370 2393
rect 3400 2307 3470 2393
rect 3500 2307 3570 2393
rect 3600 2367 3670 2393
rect 3600 2333 3618 2367
rect 3652 2333 3670 2367
rect 3600 2307 3670 2333
rect 3700 2367 3770 2393
rect 3700 2333 3718 2367
rect 3752 2333 3770 2367
rect 3700 2307 3770 2333
rect 3800 2307 3870 2393
rect 3900 2307 3970 2393
rect 4000 2367 4070 2393
rect 4000 2333 4018 2367
rect 4052 2333 4070 2367
rect 4000 2307 4070 2333
rect 4100 2367 4170 2393
rect 4100 2333 4118 2367
rect 4152 2333 4170 2367
rect 4100 2307 4170 2333
rect 4200 2367 4270 2393
rect 4200 2333 4218 2367
rect 4252 2333 4270 2367
rect 4200 2307 4270 2333
rect 4300 2367 4370 2393
rect 4300 2333 4318 2367
rect 4352 2333 4370 2367
rect 4300 2307 4370 2333
rect 4400 2367 4470 2393
rect 4400 2333 4418 2367
rect 4452 2333 4470 2367
rect 4400 2307 4470 2333
rect 4500 2307 4570 2393
rect 4600 2307 4670 2393
rect 4700 2307 4770 2393
rect 4800 2307 4870 2393
rect 4900 2367 4970 2393
rect 4900 2333 4918 2367
rect 4952 2333 4970 2367
rect 4900 2307 4970 2333
rect 5000 2367 5070 2393
rect 5000 2333 5018 2367
rect 5052 2333 5070 2367
rect 5000 2307 5070 2333
rect 5100 2307 5170 2393
rect 5200 2307 5270 2393
rect 5300 2307 5370 2393
rect 5400 2307 5470 2393
rect 5500 2367 5570 2393
rect 5500 2333 5518 2367
rect 5552 2333 5570 2367
rect 5500 2307 5570 2333
rect 5600 2367 5670 2393
rect 5600 2333 5618 2367
rect 5652 2333 5670 2367
rect 5600 2307 5670 2333
rect 5700 2367 5770 2393
rect 5700 2333 5718 2367
rect 5752 2333 5770 2367
rect 5700 2307 5770 2333
rect 5800 2367 5870 2393
rect 5800 2333 5818 2367
rect 5852 2333 5870 2367
rect 5800 2307 5870 2333
rect 5900 2367 5970 2393
rect 5900 2333 5918 2367
rect 5952 2333 5970 2367
rect 5900 2307 5970 2333
rect 6000 2307 6070 2393
rect 6100 2307 6170 2393
rect 6200 2307 6270 2393
rect 6300 2307 6370 2393
rect 6400 2367 6470 2393
rect 6400 2333 6418 2367
rect 6452 2333 6470 2367
rect 6400 2307 6470 2333
rect 6500 2367 6570 2393
rect 6500 2333 6518 2367
rect 6552 2333 6570 2367
rect 6500 2307 6570 2333
rect 6600 2367 6670 2393
rect 6600 2333 6618 2367
rect 6652 2333 6670 2367
rect 6600 2307 6670 2333
rect 6700 2307 6770 2393
rect 6800 2367 6870 2393
rect 6800 2333 6818 2367
rect 6852 2333 6870 2367
rect 6800 2307 6870 2333
rect 6900 2367 6954 2393
rect 6900 2333 6912 2367
rect 6946 2333 6954 2367
rect 6900 2307 6954 2333
rect 2716 2227 2770 2253
rect 2716 2193 2724 2227
rect 2758 2193 2770 2227
rect 2716 2167 2770 2193
rect 2800 2227 2854 2253
rect 2800 2193 2812 2227
rect 2846 2193 2854 2227
rect 2800 2167 2854 2193
rect 1516 2087 1570 2113
rect 1516 2053 1524 2087
rect 1558 2053 1570 2087
rect 1516 2027 1570 2053
rect 1600 2087 1670 2113
rect 1600 2053 1618 2087
rect 1652 2053 1670 2087
rect 1600 2027 1670 2053
rect 1700 2027 1770 2113
rect 1800 2027 1870 2113
rect 1900 2087 1970 2113
rect 1900 2053 1918 2087
rect 1952 2053 1970 2087
rect 1900 2027 1970 2053
rect 2000 2087 2070 2113
rect 2000 2053 2018 2087
rect 2052 2053 2070 2087
rect 2000 2027 2070 2053
rect 2100 2087 2170 2113
rect 2100 2053 2118 2087
rect 2152 2053 2170 2087
rect 2100 2027 2170 2053
rect 2200 2027 2270 2113
rect 2300 2027 2370 2113
rect 2400 2027 2470 2113
rect 2500 2027 2570 2113
rect 2600 2087 2670 2113
rect 2600 2053 2618 2087
rect 2652 2053 2670 2087
rect 2600 2027 2670 2053
rect 2700 2087 2754 2113
rect 2700 2053 2712 2087
rect 2746 2053 2754 2087
rect 2700 2027 2754 2053
rect 1016 1947 1070 1973
rect 1016 1913 1024 1947
rect 1058 1913 1070 1947
rect 1016 1887 1070 1913
rect 1100 1947 1170 1973
rect 1100 1913 1118 1947
rect 1152 1913 1170 1947
rect 1100 1887 1170 1913
rect 1200 1887 1270 1973
rect 1300 1887 1370 1973
rect 1400 1947 1470 1973
rect 1400 1913 1418 1947
rect 1452 1913 1470 1947
rect 1400 1887 1470 1913
rect 1500 1947 1554 1973
rect 1500 1913 1512 1947
rect 1546 1913 1554 1947
rect 1500 1887 1554 1913
rect 2916 2227 2970 2253
rect 2916 2193 2924 2227
rect 2958 2193 2970 2227
rect 2916 2167 2970 2193
rect 3000 2227 3054 2253
rect 3000 2193 3012 2227
rect 3046 2193 3054 2227
rect 3000 2167 3054 2193
rect 2816 2087 2870 2113
rect 2816 2053 2824 2087
rect 2858 2053 2870 2087
rect 2816 2027 2870 2053
rect 2900 2087 2954 2113
rect 2900 2053 2912 2087
rect 2946 2053 2954 2087
rect 2900 2027 2954 2053
rect 3116 2227 3170 2253
rect 3116 2193 3124 2227
rect 3158 2193 3170 2227
rect 3116 2167 3170 2193
rect 3200 2227 3270 2253
rect 3200 2193 3218 2227
rect 3252 2193 3270 2227
rect 3200 2167 3270 2193
rect 3300 2227 3354 2253
rect 3300 2193 3312 2227
rect 3346 2193 3354 2227
rect 3300 2167 3354 2193
rect 3416 2227 3470 2253
rect 3416 2193 3424 2227
rect 3458 2193 3470 2227
rect 3416 2167 3470 2193
rect 3500 2227 3570 2253
rect 3500 2193 3518 2227
rect 3552 2193 3570 2227
rect 3500 2167 3570 2193
rect 3600 2227 3654 2253
rect 3600 2193 3612 2227
rect 3646 2193 3654 2227
rect 3600 2167 3654 2193
rect 3016 2087 3070 2113
rect 3016 2053 3024 2087
rect 3058 2053 3070 2087
rect 3016 2027 3070 2053
rect 3100 2087 3170 2113
rect 3100 2053 3118 2087
rect 3152 2053 3170 2087
rect 3100 2027 3170 2053
rect 3200 2087 3270 2113
rect 3200 2053 3218 2087
rect 3252 2053 3270 2087
rect 3200 2027 3270 2053
rect 3300 2027 3370 2113
rect 3400 2087 3470 2113
rect 3400 2053 3418 2087
rect 3452 2053 3470 2087
rect 3400 2027 3470 2053
rect 3500 2087 3554 2113
rect 3500 2053 3512 2087
rect 3546 2053 3554 2087
rect 3500 2027 3554 2053
rect 3716 2227 3770 2253
rect 3716 2193 3724 2227
rect 3758 2193 3770 2227
rect 3716 2167 3770 2193
rect 3800 2227 3854 2253
rect 3800 2193 3812 2227
rect 3846 2193 3854 2227
rect 3800 2167 3854 2193
rect 3916 2227 3970 2253
rect 3916 2193 3924 2227
rect 3958 2193 3970 2227
rect 3916 2167 3970 2193
rect 4000 2227 4070 2253
rect 4000 2193 4018 2227
rect 4052 2193 4070 2227
rect 4000 2167 4070 2193
rect 4100 2227 4170 2253
rect 4100 2193 4118 2227
rect 4152 2193 4170 2227
rect 4100 2167 4170 2193
rect 4200 2227 4270 2253
rect 4200 2193 4218 2227
rect 4252 2193 4270 2227
rect 4200 2167 4270 2193
rect 4300 2227 4354 2253
rect 4300 2193 4312 2227
rect 4346 2193 4354 2227
rect 4300 2167 4354 2193
rect 4416 2227 4470 2253
rect 4416 2193 4424 2227
rect 4458 2193 4470 2227
rect 4416 2167 4470 2193
rect 4500 2227 4570 2253
rect 4500 2193 4518 2227
rect 4552 2193 4570 2227
rect 4500 2167 4570 2193
rect 4600 2167 4670 2253
rect 4700 2167 4770 2253
rect 4800 2167 4870 2253
rect 4900 2227 4970 2253
rect 4900 2193 4918 2227
rect 4952 2193 4970 2227
rect 4900 2167 4970 2193
rect 5000 2227 5070 2253
rect 5000 2193 5018 2227
rect 5052 2193 5070 2227
rect 5000 2167 5070 2193
rect 5100 2227 5170 2253
rect 5100 2193 5118 2227
rect 5152 2193 5170 2227
rect 5100 2167 5170 2193
rect 5200 2167 5270 2253
rect 5300 2167 5370 2253
rect 5400 2167 5470 2253
rect 5500 2167 5570 2253
rect 5600 2167 5670 2253
rect 5700 2167 5770 2253
rect 5800 2227 5870 2253
rect 5800 2193 5818 2227
rect 5852 2193 5870 2227
rect 5800 2167 5870 2193
rect 5900 2227 5970 2253
rect 5900 2193 5918 2227
rect 5952 2193 5970 2227
rect 5900 2167 5970 2193
rect 6000 2227 6070 2253
rect 6000 2193 6018 2227
rect 6052 2193 6070 2227
rect 6000 2167 6070 2193
rect 6100 2227 6154 2253
rect 6100 2193 6112 2227
rect 6146 2193 6154 2227
rect 6100 2167 6154 2193
rect 3616 2087 3670 2113
rect 3616 2053 3624 2087
rect 3658 2053 3670 2087
rect 3616 2027 3670 2053
rect 3700 2087 3770 2113
rect 3700 2053 3718 2087
rect 3752 2053 3770 2087
rect 3700 2027 3770 2053
rect 3800 2027 3870 2113
rect 3900 2027 3970 2113
rect 4000 2087 4070 2113
rect 4000 2053 4018 2087
rect 4052 2053 4070 2087
rect 4000 2027 4070 2053
rect 4100 2087 4170 2113
rect 4100 2053 4118 2087
rect 4152 2053 4170 2087
rect 4100 2027 4170 2053
rect 4200 2027 4270 2113
rect 4300 2087 4370 2113
rect 4300 2053 4318 2087
rect 4352 2053 4370 2087
rect 4300 2027 4370 2053
rect 4400 2087 4470 2113
rect 4400 2053 4418 2087
rect 4452 2053 4470 2087
rect 4400 2027 4470 2053
rect 4500 2087 4570 2113
rect 4500 2053 4518 2087
rect 4552 2053 4570 2087
rect 4500 2027 4570 2053
rect 4600 2087 4654 2113
rect 4600 2053 4612 2087
rect 4646 2053 4654 2087
rect 4600 2027 4654 2053
rect 1616 1947 1670 1973
rect 1616 1913 1624 1947
rect 1658 1913 1670 1947
rect 1616 1887 1670 1913
rect 1700 1947 1770 1973
rect 1700 1913 1718 1947
rect 1752 1913 1770 1947
rect 1700 1887 1770 1913
rect 1800 1947 1870 1973
rect 1800 1913 1818 1947
rect 1852 1913 1870 1947
rect 1800 1887 1870 1913
rect 1900 1947 1970 1973
rect 1900 1913 1918 1947
rect 1952 1913 1970 1947
rect 1900 1887 1970 1913
rect 2000 1947 2070 1973
rect 2000 1913 2018 1947
rect 2052 1913 2070 1947
rect 2000 1887 2070 1913
rect 2100 1947 2170 1973
rect 2100 1913 2118 1947
rect 2152 1913 2170 1947
rect 2100 1887 2170 1913
rect 2200 1947 2270 1973
rect 2200 1913 2218 1947
rect 2252 1913 2270 1947
rect 2200 1887 2270 1913
rect 2300 1887 2370 1973
rect 2400 1887 2470 1973
rect 2500 1947 2570 1973
rect 2500 1913 2518 1947
rect 2552 1913 2570 1947
rect 2500 1887 2570 1913
rect 2600 1947 2670 1973
rect 2600 1913 2618 1947
rect 2652 1913 2670 1947
rect 2600 1887 2670 1913
rect 2700 1887 2770 1973
rect 2800 1947 2870 1973
rect 2800 1913 2818 1947
rect 2852 1913 2870 1947
rect 2800 1887 2870 1913
rect 2900 1947 2970 1973
rect 2900 1913 2918 1947
rect 2952 1913 2970 1947
rect 2900 1887 2970 1913
rect 3000 1887 3070 1973
rect 3100 1887 3170 1973
rect 3200 1947 3270 1973
rect 3200 1913 3218 1947
rect 3252 1913 3270 1947
rect 3200 1887 3270 1913
rect 3300 1947 3370 1973
rect 3300 1913 3318 1947
rect 3352 1913 3370 1947
rect 3300 1887 3370 1913
rect 3400 1887 3470 1973
rect 3500 1947 3570 1973
rect 3500 1913 3518 1947
rect 3552 1913 3570 1947
rect 3500 1887 3570 1913
rect 3600 1947 3654 1973
rect 3600 1913 3612 1947
rect 3646 1913 3654 1947
rect 3600 1887 3654 1913
rect 16 1747 70 1833
rect 100 1807 170 1833
rect 100 1773 118 1807
rect 152 1773 170 1807
rect 100 1747 170 1773
rect 200 1807 270 1833
rect 200 1773 218 1807
rect 252 1773 270 1807
rect 200 1747 270 1773
rect 300 1807 370 1833
rect 300 1773 318 1807
rect 352 1773 370 1807
rect 300 1747 370 1773
rect 400 1747 470 1833
rect 500 1747 570 1833
rect 600 1747 670 1833
rect 700 1807 770 1833
rect 700 1773 718 1807
rect 752 1773 770 1807
rect 700 1747 770 1773
rect 800 1807 870 1833
rect 800 1773 818 1807
rect 852 1773 870 1807
rect 800 1747 870 1773
rect 900 1807 970 1833
rect 900 1773 918 1807
rect 952 1773 970 1807
rect 900 1747 970 1773
rect 1000 1807 1070 1833
rect 1000 1773 1018 1807
rect 1052 1773 1070 1807
rect 1000 1747 1070 1773
rect 1100 1807 1170 1833
rect 1100 1773 1118 1807
rect 1152 1773 1170 1807
rect 1100 1747 1170 1773
rect 1200 1807 1270 1833
rect 1200 1773 1218 1807
rect 1252 1773 1270 1807
rect 1200 1747 1270 1773
rect 1300 1807 1370 1833
rect 1300 1773 1318 1807
rect 1352 1773 1370 1807
rect 1300 1747 1370 1773
rect 1400 1807 1470 1833
rect 1400 1773 1418 1807
rect 1452 1773 1470 1807
rect 1400 1747 1470 1773
rect 1500 1807 1570 1833
rect 1500 1773 1518 1807
rect 1552 1773 1570 1807
rect 1500 1747 1570 1773
rect 1600 1807 1670 1833
rect 1600 1773 1618 1807
rect 1652 1773 1670 1807
rect 1600 1747 1670 1773
rect 1700 1747 1770 1833
rect 1800 1747 1870 1833
rect 1900 1747 1970 1833
rect 2000 1747 2070 1833
rect 2100 1807 2170 1833
rect 2100 1773 2118 1807
rect 2152 1773 2170 1807
rect 2100 1747 2170 1773
rect 2200 1807 2270 1833
rect 2200 1773 2218 1807
rect 2252 1773 2270 1807
rect 2200 1747 2270 1773
rect 2300 1807 2370 1833
rect 2300 1773 2318 1807
rect 2352 1773 2370 1807
rect 2300 1747 2370 1773
rect 2400 1807 2470 1833
rect 2400 1773 2418 1807
rect 2452 1773 2470 1807
rect 2400 1747 2470 1773
rect 2500 1747 2570 1833
rect 2600 1747 2670 1833
rect 2700 1807 2770 1833
rect 2700 1773 2718 1807
rect 2752 1773 2770 1807
rect 2700 1747 2770 1773
rect 2800 1807 2870 1833
rect 2800 1773 2818 1807
rect 2852 1773 2870 1807
rect 2800 1747 2870 1773
rect 2900 1747 2970 1833
rect 3000 1807 3070 1833
rect 3000 1773 3018 1807
rect 3052 1773 3070 1807
rect 3000 1747 3070 1773
rect 3100 1807 3154 1833
rect 3100 1773 3112 1807
rect 3146 1773 3154 1807
rect 3100 1747 3154 1773
rect 16 1607 70 1693
rect 100 1667 170 1693
rect 100 1633 118 1667
rect 152 1633 170 1667
rect 100 1607 170 1633
rect 200 1667 270 1693
rect 200 1633 218 1667
rect 252 1633 270 1667
rect 200 1607 270 1633
rect 300 1607 370 1693
rect 400 1607 470 1693
rect 500 1667 570 1693
rect 500 1633 518 1667
rect 552 1633 570 1667
rect 500 1607 570 1633
rect 600 1667 654 1693
rect 600 1633 612 1667
rect 646 1633 654 1667
rect 600 1607 654 1633
rect 16 1467 70 1553
rect 100 1527 170 1553
rect 100 1493 118 1527
rect 152 1493 170 1527
rect 100 1467 170 1493
rect 200 1527 270 1553
rect 200 1493 218 1527
rect 252 1493 270 1527
rect 200 1467 270 1493
rect 300 1527 370 1553
rect 300 1493 318 1527
rect 352 1493 370 1527
rect 300 1467 370 1493
rect 400 1527 454 1553
rect 400 1493 412 1527
rect 446 1493 454 1527
rect 400 1467 454 1493
rect 716 1667 770 1693
rect 716 1633 724 1667
rect 758 1633 770 1667
rect 716 1607 770 1633
rect 800 1667 870 1693
rect 800 1633 818 1667
rect 852 1633 870 1667
rect 800 1607 870 1633
rect 900 1667 970 1693
rect 900 1633 918 1667
rect 952 1633 970 1667
rect 900 1607 970 1633
rect 1000 1667 1054 1693
rect 1000 1633 1012 1667
rect 1046 1633 1054 1667
rect 1000 1607 1054 1633
rect 1116 1667 1170 1693
rect 1116 1633 1124 1667
rect 1158 1633 1170 1667
rect 1116 1607 1170 1633
rect 1200 1667 1254 1693
rect 1200 1633 1212 1667
rect 1246 1633 1254 1667
rect 1200 1607 1254 1633
rect 1316 1667 1370 1693
rect 1316 1633 1324 1667
rect 1358 1633 1370 1667
rect 1316 1607 1370 1633
rect 1400 1667 1470 1693
rect 1400 1633 1418 1667
rect 1452 1633 1470 1667
rect 1400 1607 1470 1633
rect 1500 1667 1554 1693
rect 1500 1633 1512 1667
rect 1546 1633 1554 1667
rect 1500 1607 1554 1633
rect 1616 1667 1670 1693
rect 1616 1633 1624 1667
rect 1658 1633 1670 1667
rect 1616 1607 1670 1633
rect 1700 1667 1770 1693
rect 1700 1633 1718 1667
rect 1752 1633 1770 1667
rect 1700 1607 1770 1633
rect 1800 1667 1870 1693
rect 1800 1633 1818 1667
rect 1852 1633 1870 1667
rect 1800 1607 1870 1633
rect 1900 1667 1970 1693
rect 1900 1633 1918 1667
rect 1952 1633 1970 1667
rect 1900 1607 1970 1633
rect 2000 1667 2070 1693
rect 2000 1633 2018 1667
rect 2052 1633 2070 1667
rect 2000 1607 2070 1633
rect 2100 1667 2170 1693
rect 2100 1633 2118 1667
rect 2152 1633 2170 1667
rect 2100 1607 2170 1633
rect 2200 1667 2270 1693
rect 2200 1633 2218 1667
rect 2252 1633 2270 1667
rect 2200 1607 2270 1633
rect 2300 1607 2370 1693
rect 2400 1667 2470 1693
rect 2400 1633 2418 1667
rect 2452 1633 2470 1667
rect 2400 1607 2470 1633
rect 2500 1667 2570 1693
rect 2500 1633 2518 1667
rect 2552 1633 2570 1667
rect 2500 1607 2570 1633
rect 2600 1667 2654 1693
rect 2600 1633 2612 1667
rect 2646 1633 2654 1667
rect 2600 1607 2654 1633
rect 516 1527 570 1553
rect 516 1493 524 1527
rect 558 1493 570 1527
rect 516 1467 570 1493
rect 600 1527 670 1553
rect 600 1493 618 1527
rect 652 1493 670 1527
rect 600 1467 670 1493
rect 700 1527 770 1553
rect 700 1493 718 1527
rect 752 1493 770 1527
rect 700 1467 770 1493
rect 800 1467 870 1553
rect 900 1527 970 1553
rect 900 1493 918 1527
rect 952 1493 970 1527
rect 900 1467 970 1493
rect 1000 1527 1070 1553
rect 1000 1493 1018 1527
rect 1052 1493 1070 1527
rect 1000 1467 1070 1493
rect 1100 1467 1170 1553
rect 1200 1467 1270 1553
rect 1300 1467 1370 1553
rect 1400 1467 1470 1553
rect 1500 1527 1570 1553
rect 1500 1493 1518 1527
rect 1552 1493 1570 1527
rect 1500 1467 1570 1493
rect 1600 1527 1670 1553
rect 1600 1493 1618 1527
rect 1652 1493 1670 1527
rect 1600 1467 1670 1493
rect 1700 1527 1770 1553
rect 1700 1493 1718 1527
rect 1752 1493 1770 1527
rect 1700 1467 1770 1493
rect 1800 1467 1870 1553
rect 1900 1527 1970 1553
rect 1900 1493 1918 1527
rect 1952 1493 1970 1527
rect 1900 1467 1970 1493
rect 2000 1527 2070 1553
rect 2000 1493 2018 1527
rect 2052 1493 2070 1527
rect 2000 1467 2070 1493
rect 2100 1527 2170 1553
rect 2100 1493 2118 1527
rect 2152 1493 2170 1527
rect 2100 1467 2170 1493
rect 2200 1467 2270 1553
rect 2300 1527 2370 1553
rect 2300 1493 2318 1527
rect 2352 1493 2370 1527
rect 2300 1467 2370 1493
rect 2400 1527 2470 1553
rect 2400 1493 2418 1527
rect 2452 1493 2470 1527
rect 2400 1467 2470 1493
rect 2500 1527 2554 1553
rect 2500 1493 2512 1527
rect 2546 1493 2554 1527
rect 2500 1467 2554 1493
rect 16 1327 70 1413
rect 100 1327 170 1413
rect 200 1327 270 1413
rect 300 1327 370 1413
rect 400 1327 470 1413
rect 500 1387 570 1413
rect 500 1353 518 1387
rect 552 1353 570 1387
rect 500 1327 570 1353
rect 600 1387 670 1413
rect 600 1353 618 1387
rect 652 1353 670 1387
rect 600 1327 670 1353
rect 700 1387 770 1413
rect 700 1353 718 1387
rect 752 1353 770 1387
rect 700 1327 770 1353
rect 800 1387 854 1413
rect 800 1353 812 1387
rect 846 1353 854 1387
rect 800 1327 854 1353
rect 3216 1807 3270 1833
rect 3216 1773 3224 1807
rect 3258 1773 3270 1807
rect 3216 1747 3270 1773
rect 3300 1807 3354 1833
rect 3300 1773 3312 1807
rect 3346 1773 3354 1807
rect 3300 1747 3354 1773
rect 3716 1947 3770 1973
rect 3716 1913 3724 1947
rect 3758 1913 3770 1947
rect 3716 1887 3770 1913
rect 3800 1947 3870 1973
rect 3800 1913 3818 1947
rect 3852 1913 3870 1947
rect 3800 1887 3870 1913
rect 3900 1887 3970 1973
rect 4000 1887 4070 1973
rect 4100 1947 4170 1973
rect 4100 1913 4118 1947
rect 4152 1913 4170 1947
rect 4100 1887 4170 1913
rect 4200 1947 4254 1973
rect 4200 1913 4212 1947
rect 4246 1913 4254 1947
rect 4200 1887 4254 1913
rect 3416 1807 3470 1833
rect 3416 1773 3424 1807
rect 3458 1773 3470 1807
rect 3416 1747 3470 1773
rect 3500 1807 3570 1833
rect 3500 1773 3518 1807
rect 3552 1773 3570 1807
rect 3500 1747 3570 1773
rect 3600 1807 3670 1833
rect 3600 1773 3618 1807
rect 3652 1773 3670 1807
rect 3600 1747 3670 1773
rect 3700 1747 3770 1833
rect 3800 1807 3870 1833
rect 3800 1773 3818 1807
rect 3852 1773 3870 1807
rect 3800 1747 3870 1773
rect 3900 1807 3954 1833
rect 3900 1773 3912 1807
rect 3946 1773 3954 1807
rect 3900 1747 3954 1773
rect 2716 1667 2770 1693
rect 2716 1633 2724 1667
rect 2758 1633 2770 1667
rect 2716 1607 2770 1633
rect 2800 1667 2870 1693
rect 2800 1633 2818 1667
rect 2852 1633 2870 1667
rect 2800 1607 2870 1633
rect 2900 1667 2970 1693
rect 2900 1633 2918 1667
rect 2952 1633 2970 1667
rect 2900 1607 2970 1633
rect 3000 1607 3070 1693
rect 3100 1667 3170 1693
rect 3100 1633 3118 1667
rect 3152 1633 3170 1667
rect 3100 1607 3170 1633
rect 3200 1667 3270 1693
rect 3200 1633 3218 1667
rect 3252 1633 3270 1667
rect 3200 1607 3270 1633
rect 3300 1607 3370 1693
rect 3400 1667 3470 1693
rect 3400 1633 3418 1667
rect 3452 1633 3470 1667
rect 3400 1607 3470 1633
rect 3500 1667 3570 1693
rect 3500 1633 3518 1667
rect 3552 1633 3570 1667
rect 3500 1607 3570 1633
rect 3600 1667 3670 1693
rect 3600 1633 3618 1667
rect 3652 1633 3670 1667
rect 3600 1607 3670 1633
rect 3700 1667 3754 1693
rect 3700 1633 3712 1667
rect 3746 1633 3754 1667
rect 3700 1607 3754 1633
rect 2616 1527 2670 1553
rect 2616 1493 2624 1527
rect 2658 1493 2670 1527
rect 2616 1467 2670 1493
rect 2700 1527 2770 1553
rect 2700 1493 2718 1527
rect 2752 1493 2770 1527
rect 2700 1467 2770 1493
rect 2800 1467 2870 1553
rect 2900 1527 2970 1553
rect 2900 1493 2918 1527
rect 2952 1493 2970 1527
rect 2900 1467 2970 1493
rect 3000 1527 3070 1553
rect 3000 1493 3018 1527
rect 3052 1493 3070 1527
rect 3000 1467 3070 1493
rect 3100 1527 3154 1553
rect 3100 1493 3112 1527
rect 3146 1493 3154 1527
rect 3100 1467 3154 1493
rect 916 1387 970 1413
rect 916 1353 924 1387
rect 958 1353 970 1387
rect 916 1327 970 1353
rect 1000 1387 1070 1413
rect 1000 1353 1018 1387
rect 1052 1353 1070 1387
rect 1000 1327 1070 1353
rect 1100 1387 1170 1413
rect 1100 1353 1118 1387
rect 1152 1353 1170 1387
rect 1100 1327 1170 1353
rect 1200 1327 1270 1413
rect 1300 1387 1370 1413
rect 1300 1353 1318 1387
rect 1352 1353 1370 1387
rect 1300 1327 1370 1353
rect 1400 1387 1470 1413
rect 1400 1353 1418 1387
rect 1452 1353 1470 1387
rect 1400 1327 1470 1353
rect 1500 1387 1570 1413
rect 1500 1353 1518 1387
rect 1552 1353 1570 1387
rect 1500 1327 1570 1353
rect 1600 1327 1670 1413
rect 1700 1327 1770 1413
rect 1800 1387 1870 1413
rect 1800 1353 1818 1387
rect 1852 1353 1870 1387
rect 1800 1327 1870 1353
rect 1900 1387 1970 1413
rect 1900 1353 1918 1387
rect 1952 1353 1970 1387
rect 1900 1327 1970 1353
rect 2000 1327 2070 1413
rect 2100 1387 2170 1413
rect 2100 1353 2118 1387
rect 2152 1353 2170 1387
rect 2100 1327 2170 1353
rect 2200 1387 2270 1413
rect 2200 1353 2218 1387
rect 2252 1353 2270 1387
rect 2200 1327 2270 1353
rect 2300 1387 2370 1413
rect 2300 1353 2318 1387
rect 2352 1353 2370 1387
rect 2300 1327 2370 1353
rect 2400 1327 2470 1413
rect 2500 1327 2570 1413
rect 2600 1327 2670 1413
rect 2700 1387 2770 1413
rect 2700 1353 2718 1387
rect 2752 1353 2770 1387
rect 2700 1327 2770 1353
rect 2800 1387 2854 1413
rect 2800 1353 2812 1387
rect 2846 1353 2854 1387
rect 2800 1327 2854 1353
rect 16 1097 70 1183
rect 100 1157 170 1183
rect 100 1123 118 1157
rect 152 1123 170 1157
rect 100 1097 170 1123
rect 200 1157 270 1183
rect 200 1123 218 1157
rect 252 1123 270 1157
rect 200 1097 270 1123
rect 300 1097 370 1183
rect 400 1097 470 1183
rect 500 1097 570 1183
rect 600 1097 670 1183
rect 700 1097 770 1183
rect 800 1097 870 1183
rect 900 1097 970 1183
rect 1000 1097 1070 1183
rect 1100 1157 1170 1183
rect 1100 1123 1118 1157
rect 1152 1123 1170 1157
rect 1100 1097 1170 1123
rect 1200 1157 1270 1183
rect 1200 1123 1218 1157
rect 1252 1123 1270 1157
rect 1200 1097 1270 1123
rect 1300 1157 1370 1183
rect 1300 1123 1318 1157
rect 1352 1123 1370 1157
rect 1300 1097 1370 1123
rect 1400 1097 1470 1183
rect 1500 1097 1570 1183
rect 1600 1157 1670 1183
rect 1600 1123 1618 1157
rect 1652 1123 1670 1157
rect 1600 1097 1670 1123
rect 1700 1157 1754 1183
rect 1700 1123 1712 1157
rect 1746 1123 1754 1157
rect 1700 1097 1754 1123
rect 16 1017 70 1043
rect 16 983 24 1017
rect 58 983 70 1017
rect 16 957 70 983
rect 100 1017 154 1043
rect 100 983 112 1017
rect 146 983 154 1017
rect 100 957 154 983
rect 16 877 70 903
rect 16 843 24 877
rect 58 843 70 877
rect 16 817 70 843
rect 100 877 154 903
rect 100 843 112 877
rect 146 843 154 877
rect 100 817 154 843
rect 216 1017 270 1043
rect 216 983 224 1017
rect 258 983 270 1017
rect 216 957 270 983
rect 300 1017 370 1043
rect 300 983 318 1017
rect 352 983 370 1017
rect 300 957 370 983
rect 400 1017 470 1043
rect 400 983 418 1017
rect 452 983 470 1017
rect 400 957 470 983
rect 500 1017 570 1043
rect 500 983 518 1017
rect 552 983 570 1017
rect 500 957 570 983
rect 600 1017 654 1043
rect 600 983 612 1017
rect 646 983 654 1017
rect 600 957 654 983
rect 716 1017 770 1043
rect 716 983 724 1017
rect 758 983 770 1017
rect 716 957 770 983
rect 800 1017 870 1043
rect 800 983 818 1017
rect 852 983 870 1017
rect 800 957 870 983
rect 900 957 970 1043
rect 1000 1017 1070 1043
rect 1000 983 1018 1017
rect 1052 983 1070 1017
rect 1000 957 1070 983
rect 1100 1017 1170 1043
rect 1100 983 1118 1017
rect 1152 983 1170 1017
rect 1100 957 1170 983
rect 1200 1017 1254 1043
rect 1200 983 1212 1017
rect 1246 983 1254 1017
rect 1200 957 1254 983
rect 1816 1157 1870 1183
rect 1816 1123 1824 1157
rect 1858 1123 1870 1157
rect 1816 1097 1870 1123
rect 1900 1157 1970 1183
rect 1900 1123 1918 1157
rect 1952 1123 1970 1157
rect 1900 1097 1970 1123
rect 2000 1157 2054 1183
rect 2000 1123 2012 1157
rect 2046 1123 2054 1157
rect 2000 1097 2054 1123
rect 3216 1527 3270 1553
rect 3216 1493 3224 1527
rect 3258 1493 3270 1527
rect 3216 1467 3270 1493
rect 3300 1527 3370 1553
rect 3300 1493 3318 1527
rect 3352 1493 3370 1527
rect 3300 1467 3370 1493
rect 3400 1527 3470 1553
rect 3400 1493 3418 1527
rect 3452 1493 3470 1527
rect 3400 1467 3470 1493
rect 3500 1527 3554 1553
rect 3500 1493 3512 1527
rect 3546 1493 3554 1527
rect 3500 1467 3554 1493
rect 3816 1667 3870 1693
rect 3816 1633 3824 1667
rect 3858 1633 3870 1667
rect 3816 1607 3870 1633
rect 3900 1667 3954 1693
rect 3900 1633 3912 1667
rect 3946 1633 3954 1667
rect 3900 1607 3954 1633
rect 4016 1807 4070 1833
rect 4016 1773 4024 1807
rect 4058 1773 4070 1807
rect 4016 1747 4070 1773
rect 4100 1807 4154 1833
rect 4100 1773 4112 1807
rect 4146 1773 4154 1807
rect 4100 1747 4154 1773
rect 4016 1667 4070 1693
rect 4016 1633 4024 1667
rect 4058 1633 4070 1667
rect 4016 1607 4070 1633
rect 4100 1667 4154 1693
rect 4100 1633 4112 1667
rect 4146 1633 4154 1667
rect 4100 1607 4154 1633
rect 3616 1527 3670 1553
rect 3616 1493 3624 1527
rect 3658 1493 3670 1527
rect 3616 1467 3670 1493
rect 3700 1527 3770 1553
rect 3700 1493 3718 1527
rect 3752 1493 3770 1527
rect 3700 1467 3770 1493
rect 3800 1527 3870 1553
rect 3800 1493 3818 1527
rect 3852 1493 3870 1527
rect 3800 1467 3870 1493
rect 3900 1527 3970 1553
rect 3900 1493 3918 1527
rect 3952 1493 3970 1527
rect 3900 1467 3970 1493
rect 4000 1527 4054 1553
rect 4000 1493 4012 1527
rect 4046 1493 4054 1527
rect 4000 1467 4054 1493
rect 4316 1947 4370 1973
rect 4316 1913 4324 1947
rect 4358 1913 4370 1947
rect 4316 1887 4370 1913
rect 4400 1947 4454 1973
rect 4400 1913 4412 1947
rect 4446 1913 4454 1947
rect 4400 1887 4454 1913
rect 4516 1947 4570 1973
rect 4516 1913 4524 1947
rect 4558 1913 4570 1947
rect 4516 1887 4570 1913
rect 4600 1947 4654 1973
rect 4600 1913 4612 1947
rect 4646 1913 4654 1947
rect 4600 1887 4654 1913
rect 4716 2087 4770 2113
rect 4716 2053 4724 2087
rect 4758 2053 4770 2087
rect 4716 2027 4770 2053
rect 4800 2087 4870 2113
rect 4800 2053 4818 2087
rect 4852 2053 4870 2087
rect 4800 2027 4870 2053
rect 4900 2087 4954 2113
rect 4900 2053 4912 2087
rect 4946 2053 4954 2087
rect 4900 2027 4954 2053
rect 5016 2087 5070 2113
rect 5016 2053 5024 2087
rect 5058 2053 5070 2087
rect 5016 2027 5070 2053
rect 5100 2087 5170 2113
rect 5100 2053 5118 2087
rect 5152 2053 5170 2087
rect 5100 2027 5170 2053
rect 5200 2027 5270 2113
rect 5300 2027 5370 2113
rect 5400 2027 5470 2113
rect 5500 2027 5570 2113
rect 5600 2087 5670 2113
rect 5600 2053 5618 2087
rect 5652 2053 5670 2087
rect 5600 2027 5670 2053
rect 5700 2087 5754 2113
rect 5700 2053 5712 2087
rect 5746 2053 5754 2087
rect 5700 2027 5754 2053
rect 4716 1947 4770 1973
rect 4716 1913 4724 1947
rect 4758 1913 4770 1947
rect 4716 1887 4770 1913
rect 4800 1947 4870 1973
rect 4800 1913 4818 1947
rect 4852 1913 4870 1947
rect 4800 1887 4870 1913
rect 4900 1887 4970 1973
rect 5000 1947 5070 1973
rect 5000 1913 5018 1947
rect 5052 1913 5070 1947
rect 5000 1887 5070 1913
rect 5100 1947 5154 1973
rect 5100 1913 5112 1947
rect 5146 1913 5154 1947
rect 5100 1887 5154 1913
rect 4216 1807 4270 1833
rect 4216 1773 4224 1807
rect 4258 1773 4270 1807
rect 4216 1747 4270 1773
rect 4300 1807 4370 1833
rect 4300 1773 4318 1807
rect 4352 1773 4370 1807
rect 4300 1747 4370 1773
rect 4400 1747 4470 1833
rect 4500 1747 4570 1833
rect 4600 1747 4670 1833
rect 4700 1807 4770 1833
rect 4700 1773 4718 1807
rect 4752 1773 4770 1807
rect 4700 1747 4770 1773
rect 4800 1807 4854 1833
rect 4800 1773 4812 1807
rect 4846 1773 4854 1807
rect 4800 1747 4854 1773
rect 4216 1667 4270 1693
rect 4216 1633 4224 1667
rect 4258 1633 4270 1667
rect 4216 1607 4270 1633
rect 4300 1667 4370 1693
rect 4300 1633 4318 1667
rect 4352 1633 4370 1667
rect 4300 1607 4370 1633
rect 4400 1667 4454 1693
rect 4400 1633 4412 1667
rect 4446 1633 4454 1667
rect 4400 1607 4454 1633
rect 5216 1947 5270 1973
rect 5216 1913 5224 1947
rect 5258 1913 5270 1947
rect 5216 1887 5270 1913
rect 5300 1947 5370 1973
rect 5300 1913 5318 1947
rect 5352 1913 5370 1947
rect 5300 1887 5370 1913
rect 5400 1947 5470 1973
rect 5400 1913 5418 1947
rect 5452 1913 5470 1947
rect 5400 1887 5470 1913
rect 5500 1947 5570 1973
rect 5500 1913 5518 1947
rect 5552 1913 5570 1947
rect 5500 1887 5570 1913
rect 5600 1947 5670 1973
rect 5600 1913 5618 1947
rect 5652 1913 5670 1947
rect 5600 1887 5670 1913
rect 5700 1947 5754 1973
rect 5700 1913 5712 1947
rect 5746 1913 5754 1947
rect 5700 1887 5754 1913
rect 6216 2227 6270 2253
rect 6216 2193 6224 2227
rect 6258 2193 6270 2227
rect 6216 2167 6270 2193
rect 6300 2227 6370 2253
rect 6300 2193 6318 2227
rect 6352 2193 6370 2227
rect 6300 2167 6370 2193
rect 6400 2227 6454 2253
rect 6400 2193 6412 2227
rect 6446 2193 6454 2227
rect 6400 2167 6454 2193
rect 6516 2227 6570 2253
rect 6516 2193 6524 2227
rect 6558 2193 6570 2227
rect 6516 2167 6570 2193
rect 6600 2227 6670 2253
rect 6600 2193 6618 2227
rect 6652 2193 6670 2227
rect 6600 2167 6670 2193
rect 6700 2227 6754 2253
rect 6700 2193 6712 2227
rect 6746 2193 6754 2227
rect 6700 2167 6754 2193
rect 5816 2087 5870 2113
rect 5816 2053 5824 2087
rect 5858 2053 5870 2087
rect 5816 2027 5870 2053
rect 5900 2087 5970 2113
rect 5900 2053 5918 2087
rect 5952 2053 5970 2087
rect 5900 2027 5970 2053
rect 6000 2087 6070 2113
rect 6000 2053 6018 2087
rect 6052 2053 6070 2087
rect 6000 2027 6070 2053
rect 6100 2087 6170 2113
rect 6100 2053 6118 2087
rect 6152 2053 6170 2087
rect 6100 2027 6170 2053
rect 6200 2027 6270 2113
rect 6300 2027 6370 2113
rect 6400 2027 6470 2113
rect 6500 2087 6570 2113
rect 6500 2053 6518 2087
rect 6552 2053 6570 2087
rect 6500 2027 6570 2053
rect 6600 2087 6654 2113
rect 6600 2053 6612 2087
rect 6646 2053 6654 2087
rect 6600 2027 6654 2053
rect 6816 2227 6870 2253
rect 6816 2193 6824 2227
rect 6858 2193 6870 2227
rect 6816 2167 6870 2193
rect 6900 2227 6954 2253
rect 6900 2193 6912 2227
rect 6946 2193 6954 2227
rect 6900 2167 6954 2193
rect 6716 2087 6770 2113
rect 6716 2053 6724 2087
rect 6758 2053 6770 2087
rect 6716 2027 6770 2053
rect 6800 2087 6854 2113
rect 6800 2053 6812 2087
rect 6846 2053 6854 2087
rect 6800 2027 6854 2053
rect 5816 1947 5870 1973
rect 5816 1913 5824 1947
rect 5858 1913 5870 1947
rect 5816 1887 5870 1913
rect 5900 1947 5970 1973
rect 5900 1913 5918 1947
rect 5952 1913 5970 1947
rect 5900 1887 5970 1913
rect 6000 1887 6070 1973
rect 6100 1887 6170 1973
rect 6200 1947 6270 1973
rect 6200 1913 6218 1947
rect 6252 1913 6270 1947
rect 6200 1887 6270 1913
rect 6300 1947 6370 1973
rect 6300 1913 6318 1947
rect 6352 1913 6370 1947
rect 6300 1887 6370 1913
rect 6400 1947 6470 1973
rect 6400 1913 6418 1947
rect 6452 1913 6470 1947
rect 6400 1887 6470 1913
rect 6500 1947 6570 1973
rect 6500 1913 6518 1947
rect 6552 1913 6570 1947
rect 6500 1887 6570 1913
rect 6600 1947 6670 1973
rect 6600 1913 6618 1947
rect 6652 1913 6670 1947
rect 6600 1887 6670 1913
rect 6700 1947 6754 1973
rect 6700 1913 6712 1947
rect 6746 1913 6754 1947
rect 6700 1887 6754 1913
rect 4916 1807 4970 1833
rect 4916 1773 4924 1807
rect 4958 1773 4970 1807
rect 4916 1747 4970 1773
rect 5000 1807 5070 1833
rect 5000 1773 5018 1807
rect 5052 1773 5070 1807
rect 5000 1747 5070 1773
rect 5100 1807 5170 1833
rect 5100 1773 5118 1807
rect 5152 1773 5170 1807
rect 5100 1747 5170 1773
rect 5200 1807 5270 1833
rect 5200 1773 5218 1807
rect 5252 1773 5270 1807
rect 5200 1747 5270 1773
rect 5300 1807 5370 1833
rect 5300 1773 5318 1807
rect 5352 1773 5370 1807
rect 5300 1747 5370 1773
rect 5400 1807 5470 1833
rect 5400 1773 5418 1807
rect 5452 1773 5470 1807
rect 5400 1747 5470 1773
rect 5500 1807 5570 1833
rect 5500 1773 5518 1807
rect 5552 1773 5570 1807
rect 5500 1747 5570 1773
rect 5600 1747 5670 1833
rect 5700 1747 5770 1833
rect 5800 1747 5870 1833
rect 5900 1747 5970 1833
rect 6000 1747 6070 1833
rect 6100 1747 6170 1833
rect 6200 1807 6270 1833
rect 6200 1773 6218 1807
rect 6252 1773 6270 1807
rect 6200 1747 6270 1773
rect 6300 1807 6354 1833
rect 6300 1773 6312 1807
rect 6346 1773 6354 1807
rect 6300 1747 6354 1773
rect 4516 1667 4570 1693
rect 4516 1633 4524 1667
rect 4558 1633 4570 1667
rect 4516 1607 4570 1633
rect 4600 1667 4670 1693
rect 4600 1633 4618 1667
rect 4652 1633 4670 1667
rect 4600 1607 4670 1633
rect 4700 1667 4770 1693
rect 4700 1633 4718 1667
rect 4752 1633 4770 1667
rect 4700 1607 4770 1633
rect 4800 1667 4870 1693
rect 4800 1633 4818 1667
rect 4852 1633 4870 1667
rect 4800 1607 4870 1633
rect 4900 1667 4954 1693
rect 4900 1633 4912 1667
rect 4946 1633 4954 1667
rect 4900 1607 4954 1633
rect 4116 1527 4170 1553
rect 4116 1493 4124 1527
rect 4158 1493 4170 1527
rect 4116 1467 4170 1493
rect 4200 1527 4270 1553
rect 4200 1493 4218 1527
rect 4252 1493 4270 1527
rect 4200 1467 4270 1493
rect 4300 1527 4370 1553
rect 4300 1493 4318 1527
rect 4352 1493 4370 1527
rect 4300 1467 4370 1493
rect 4400 1527 4470 1553
rect 4400 1493 4418 1527
rect 4452 1493 4470 1527
rect 4400 1467 4470 1493
rect 4500 1467 4570 1553
rect 4600 1527 4670 1553
rect 4600 1493 4618 1527
rect 4652 1493 4670 1527
rect 4600 1467 4670 1493
rect 4700 1527 4770 1553
rect 4700 1493 4718 1527
rect 4752 1493 4770 1527
rect 4700 1467 4770 1493
rect 4800 1527 4854 1553
rect 4800 1493 4812 1527
rect 4846 1493 4854 1527
rect 4800 1467 4854 1493
rect 2916 1387 2970 1413
rect 2916 1353 2924 1387
rect 2958 1353 2970 1387
rect 2916 1327 2970 1353
rect 3000 1387 3070 1413
rect 3000 1353 3018 1387
rect 3052 1353 3070 1387
rect 3000 1327 3070 1353
rect 3100 1327 3170 1413
rect 3200 1387 3270 1413
rect 3200 1353 3218 1387
rect 3252 1353 3270 1387
rect 3200 1327 3270 1353
rect 3300 1387 3370 1413
rect 3300 1353 3318 1387
rect 3352 1353 3370 1387
rect 3300 1327 3370 1353
rect 3400 1387 3470 1413
rect 3400 1353 3418 1387
rect 3452 1353 3470 1387
rect 3400 1327 3470 1353
rect 3500 1387 3570 1413
rect 3500 1353 3518 1387
rect 3552 1353 3570 1387
rect 3500 1327 3570 1353
rect 3600 1327 3670 1413
rect 3700 1327 3770 1413
rect 3800 1387 3870 1413
rect 3800 1353 3818 1387
rect 3852 1353 3870 1387
rect 3800 1327 3870 1353
rect 3900 1387 3970 1413
rect 3900 1353 3918 1387
rect 3952 1353 3970 1387
rect 3900 1327 3970 1353
rect 4000 1387 4070 1413
rect 4000 1353 4018 1387
rect 4052 1353 4070 1387
rect 4000 1327 4070 1353
rect 4100 1387 4170 1413
rect 4100 1353 4118 1387
rect 4152 1353 4170 1387
rect 4100 1327 4170 1353
rect 4200 1327 4270 1413
rect 4300 1387 4370 1413
rect 4300 1353 4318 1387
rect 4352 1353 4370 1387
rect 4300 1327 4370 1353
rect 4400 1387 4470 1413
rect 4400 1353 4418 1387
rect 4452 1353 4470 1387
rect 4400 1327 4470 1353
rect 4500 1387 4570 1413
rect 4500 1353 4518 1387
rect 4552 1353 4570 1387
rect 4500 1327 4570 1353
rect 4600 1387 4654 1413
rect 4600 1353 4612 1387
rect 4646 1353 4654 1387
rect 4600 1327 4654 1353
rect 2116 1157 2170 1183
rect 2116 1123 2124 1157
rect 2158 1123 2170 1157
rect 2116 1097 2170 1123
rect 2200 1157 2270 1183
rect 2200 1123 2218 1157
rect 2252 1123 2270 1157
rect 2200 1097 2270 1123
rect 2300 1097 2370 1183
rect 2400 1097 2470 1183
rect 2500 1097 2570 1183
rect 2600 1097 2670 1183
rect 2700 1097 2770 1183
rect 2800 1097 2870 1183
rect 2900 1157 2970 1183
rect 2900 1123 2918 1157
rect 2952 1123 2970 1157
rect 2900 1097 2970 1123
rect 3000 1157 3054 1183
rect 3000 1123 3012 1157
rect 3046 1123 3054 1157
rect 3000 1097 3054 1123
rect 1316 1017 1370 1043
rect 1316 983 1324 1017
rect 1358 983 1370 1017
rect 1316 957 1370 983
rect 1400 1017 1470 1043
rect 1400 983 1418 1017
rect 1452 983 1470 1017
rect 1400 957 1470 983
rect 1500 957 1570 1043
rect 1600 1017 1670 1043
rect 1600 983 1618 1017
rect 1652 983 1670 1017
rect 1600 957 1670 983
rect 1700 1017 1770 1043
rect 1700 983 1718 1017
rect 1752 983 1770 1017
rect 1700 957 1770 983
rect 1800 957 1870 1043
rect 1900 957 1970 1043
rect 2000 1017 2070 1043
rect 2000 983 2018 1017
rect 2052 983 2070 1017
rect 2000 957 2070 983
rect 2100 1017 2170 1043
rect 2100 983 2118 1017
rect 2152 983 2170 1017
rect 2100 957 2170 983
rect 2200 1017 2270 1043
rect 2200 983 2218 1017
rect 2252 983 2270 1017
rect 2200 957 2270 983
rect 2300 1017 2370 1043
rect 2300 983 2318 1017
rect 2352 983 2370 1017
rect 2300 957 2370 983
rect 2400 1017 2470 1043
rect 2400 983 2418 1017
rect 2452 983 2470 1017
rect 2400 957 2470 983
rect 2500 1017 2570 1043
rect 2500 983 2518 1017
rect 2552 983 2570 1017
rect 2500 957 2570 983
rect 2600 1017 2654 1043
rect 2600 983 2612 1017
rect 2646 983 2654 1017
rect 2600 957 2654 983
rect 2716 1017 2770 1043
rect 2716 983 2724 1017
rect 2758 983 2770 1017
rect 2716 957 2770 983
rect 2800 1017 2854 1043
rect 2800 983 2812 1017
rect 2846 983 2854 1017
rect 2800 957 2854 983
rect 3116 1157 3170 1183
rect 3116 1123 3124 1157
rect 3158 1123 3170 1157
rect 3116 1097 3170 1123
rect 3200 1157 3254 1183
rect 3200 1123 3212 1157
rect 3246 1123 3254 1157
rect 3200 1097 3254 1123
rect 2916 1017 2970 1043
rect 2916 983 2924 1017
rect 2958 983 2970 1017
rect 2916 957 2970 983
rect 3000 1017 3070 1043
rect 3000 983 3018 1017
rect 3052 983 3070 1017
rect 3000 957 3070 983
rect 3100 1017 3154 1043
rect 3100 983 3112 1017
rect 3146 983 3154 1017
rect 3100 957 3154 983
rect 216 877 270 903
rect 216 843 224 877
rect 258 843 270 877
rect 216 817 270 843
rect 300 877 370 903
rect 300 843 318 877
rect 352 843 370 877
rect 300 817 370 843
rect 400 877 470 903
rect 400 843 418 877
rect 452 843 470 877
rect 400 817 470 843
rect 500 877 570 903
rect 500 843 518 877
rect 552 843 570 877
rect 500 817 570 843
rect 600 877 670 903
rect 600 843 618 877
rect 652 843 670 877
rect 600 817 670 843
rect 700 877 770 903
rect 700 843 718 877
rect 752 843 770 877
rect 700 817 770 843
rect 800 817 870 903
rect 900 877 970 903
rect 900 843 918 877
rect 952 843 970 877
rect 900 817 970 843
rect 1000 877 1070 903
rect 1000 843 1018 877
rect 1052 843 1070 877
rect 1000 817 1070 843
rect 1100 877 1170 903
rect 1100 843 1118 877
rect 1152 843 1170 877
rect 1100 817 1170 843
rect 1200 877 1270 903
rect 1200 843 1218 877
rect 1252 843 1270 877
rect 1200 817 1270 843
rect 1300 817 1370 903
rect 1400 817 1470 903
rect 1500 817 1570 903
rect 1600 877 1670 903
rect 1600 843 1618 877
rect 1652 843 1670 877
rect 1600 817 1670 843
rect 1700 877 1770 903
rect 1700 843 1718 877
rect 1752 843 1770 877
rect 1700 817 1770 843
rect 1800 817 1870 903
rect 1900 877 1970 903
rect 1900 843 1918 877
rect 1952 843 1970 877
rect 1900 817 1970 843
rect 2000 877 2070 903
rect 2000 843 2018 877
rect 2052 843 2070 877
rect 2000 817 2070 843
rect 2100 877 2170 903
rect 2100 843 2118 877
rect 2152 843 2170 877
rect 2100 817 2170 843
rect 2200 817 2270 903
rect 2300 817 2370 903
rect 2400 877 2470 903
rect 2400 843 2418 877
rect 2452 843 2470 877
rect 2400 817 2470 843
rect 2500 877 2570 903
rect 2500 843 2518 877
rect 2552 843 2570 877
rect 2500 817 2570 843
rect 2600 817 2670 903
rect 2700 877 2770 903
rect 2700 843 2718 877
rect 2752 843 2770 877
rect 2700 817 2770 843
rect 2800 877 2870 903
rect 2800 843 2818 877
rect 2852 843 2870 877
rect 2800 817 2870 843
rect 2900 877 2954 903
rect 2900 843 2912 877
rect 2946 843 2954 877
rect 2900 817 2954 843
rect 16 677 70 763
rect 100 737 170 763
rect 100 703 118 737
rect 152 703 170 737
rect 100 677 170 703
rect 200 737 270 763
rect 200 703 218 737
rect 252 703 270 737
rect 200 677 270 703
rect 300 677 370 763
rect 400 737 470 763
rect 400 703 418 737
rect 452 703 470 737
rect 400 677 470 703
rect 500 737 554 763
rect 500 703 512 737
rect 546 703 554 737
rect 500 677 554 703
rect 616 737 670 763
rect 616 703 624 737
rect 658 703 670 737
rect 616 677 670 703
rect 700 737 754 763
rect 700 703 712 737
rect 746 703 754 737
rect 700 677 754 703
rect 16 537 70 623
rect 100 537 170 623
rect 200 537 270 623
rect 300 537 370 623
rect 400 597 470 623
rect 400 563 418 597
rect 452 563 470 597
rect 400 537 470 563
rect 500 597 570 623
rect 500 563 518 597
rect 552 563 570 597
rect 500 537 570 563
rect 600 597 670 623
rect 600 563 618 597
rect 652 563 670 597
rect 600 537 670 563
rect 700 597 754 623
rect 700 563 712 597
rect 746 563 754 597
rect 700 537 754 563
rect 16 397 70 483
rect 100 457 170 483
rect 100 423 118 457
rect 152 423 170 457
rect 100 397 170 423
rect 200 457 270 483
rect 200 423 218 457
rect 252 423 270 457
rect 200 397 270 423
rect 300 457 354 483
rect 300 423 312 457
rect 346 423 354 457
rect 300 397 354 423
rect 816 737 870 763
rect 816 703 824 737
rect 858 703 870 737
rect 816 677 870 703
rect 900 737 970 763
rect 900 703 918 737
rect 952 703 970 737
rect 900 677 970 703
rect 1000 677 1070 763
rect 1100 737 1170 763
rect 1100 703 1118 737
rect 1152 703 1170 737
rect 1100 677 1170 703
rect 1200 737 1254 763
rect 1200 703 1212 737
rect 1246 703 1254 737
rect 1200 677 1254 703
rect 816 597 870 623
rect 816 563 824 597
rect 858 563 870 597
rect 816 537 870 563
rect 900 597 970 623
rect 900 563 918 597
rect 952 563 970 597
rect 900 537 970 563
rect 1000 537 1070 623
rect 1100 597 1170 623
rect 1100 563 1118 597
rect 1152 563 1170 597
rect 1100 537 1170 563
rect 1200 597 1254 623
rect 1200 563 1212 597
rect 1246 563 1254 597
rect 1200 537 1254 563
rect 416 457 470 483
rect 416 423 424 457
rect 458 423 470 457
rect 416 397 470 423
rect 500 457 570 483
rect 500 423 518 457
rect 552 423 570 457
rect 500 397 570 423
rect 600 397 670 483
rect 700 397 770 483
rect 800 397 870 483
rect 900 457 970 483
rect 900 423 918 457
rect 952 423 970 457
rect 900 397 970 423
rect 1000 457 1070 483
rect 1000 423 1018 457
rect 1052 423 1070 457
rect 1000 397 1070 423
rect 1100 457 1154 483
rect 1100 423 1112 457
rect 1146 423 1154 457
rect 1100 397 1154 423
rect 1316 737 1370 763
rect 1316 703 1324 737
rect 1358 703 1370 737
rect 1316 677 1370 703
rect 1400 737 1454 763
rect 1400 703 1412 737
rect 1446 703 1454 737
rect 1400 677 1454 703
rect 1516 737 1570 763
rect 1516 703 1524 737
rect 1558 703 1570 737
rect 1516 677 1570 703
rect 1600 737 1670 763
rect 1600 703 1618 737
rect 1652 703 1670 737
rect 1600 677 1670 703
rect 1700 677 1770 763
rect 1800 737 1870 763
rect 1800 703 1818 737
rect 1852 703 1870 737
rect 1800 677 1870 703
rect 1900 737 1970 763
rect 1900 703 1918 737
rect 1952 703 1970 737
rect 1900 677 1970 703
rect 2000 737 2054 763
rect 2000 703 2012 737
rect 2046 703 2054 737
rect 2000 677 2054 703
rect 2116 737 2170 763
rect 2116 703 2124 737
rect 2158 703 2170 737
rect 2116 677 2170 703
rect 2200 737 2270 763
rect 2200 703 2218 737
rect 2252 703 2270 737
rect 2200 677 2270 703
rect 2300 737 2370 763
rect 2300 703 2318 737
rect 2352 703 2370 737
rect 2300 677 2370 703
rect 2400 737 2454 763
rect 2400 703 2412 737
rect 2446 703 2454 737
rect 2400 677 2454 703
rect 1316 597 1370 623
rect 1316 563 1324 597
rect 1358 563 1370 597
rect 1316 537 1370 563
rect 1400 597 1470 623
rect 1400 563 1418 597
rect 1452 563 1470 597
rect 1400 537 1470 563
rect 1500 597 1570 623
rect 1500 563 1518 597
rect 1552 563 1570 597
rect 1500 537 1570 563
rect 1600 537 1670 623
rect 1700 597 1770 623
rect 1700 563 1718 597
rect 1752 563 1770 597
rect 1700 537 1770 563
rect 1800 597 1870 623
rect 1800 563 1818 597
rect 1852 563 1870 597
rect 1800 537 1870 563
rect 1900 597 1970 623
rect 1900 563 1918 597
rect 1952 563 1970 597
rect 1900 537 1970 563
rect 2000 597 2070 623
rect 2000 563 2018 597
rect 2052 563 2070 597
rect 2000 537 2070 563
rect 2100 597 2154 623
rect 2100 563 2112 597
rect 2146 563 2154 597
rect 2100 537 2154 563
rect 1216 457 1270 483
rect 1216 423 1224 457
rect 1258 423 1270 457
rect 1216 397 1270 423
rect 1300 457 1370 483
rect 1300 423 1318 457
rect 1352 423 1370 457
rect 1300 397 1370 423
rect 1400 457 1470 483
rect 1400 423 1418 457
rect 1452 423 1470 457
rect 1400 397 1470 423
rect 1500 397 1570 483
rect 1600 457 1670 483
rect 1600 423 1618 457
rect 1652 423 1670 457
rect 1600 397 1670 423
rect 1700 457 1770 483
rect 1700 423 1718 457
rect 1752 423 1770 457
rect 1700 397 1770 423
rect 1800 457 1854 483
rect 1800 423 1812 457
rect 1846 423 1854 457
rect 1800 397 1854 423
rect 16 257 70 343
rect 100 317 170 343
rect 100 283 118 317
rect 152 283 170 317
rect 100 257 170 283
rect 200 317 270 343
rect 200 283 218 317
rect 252 283 270 317
rect 200 257 270 283
rect 300 257 370 343
rect 400 257 470 343
rect 500 257 570 343
rect 600 257 670 343
rect 700 257 770 343
rect 800 317 870 343
rect 800 283 818 317
rect 852 283 870 317
rect 800 257 870 283
rect 900 317 970 343
rect 900 283 918 317
rect 952 283 970 317
rect 900 257 970 283
rect 1000 317 1070 343
rect 1000 283 1018 317
rect 1052 283 1070 317
rect 1000 257 1070 283
rect 1100 257 1170 343
rect 1200 317 1270 343
rect 1200 283 1218 317
rect 1252 283 1270 317
rect 1200 257 1270 283
rect 1300 317 1370 343
rect 1300 283 1318 317
rect 1352 283 1370 317
rect 1300 257 1370 283
rect 1400 257 1470 343
rect 1500 257 1570 343
rect 1600 317 1670 343
rect 1600 283 1618 317
rect 1652 283 1670 317
rect 1600 257 1670 283
rect 1700 317 1754 343
rect 1700 283 1712 317
rect 1746 283 1754 317
rect 1700 257 1754 283
rect 16 177 70 203
rect 16 143 24 177
rect 58 143 70 177
rect 16 117 70 143
rect 100 177 170 203
rect 100 143 118 177
rect 152 143 170 177
rect 100 117 170 143
rect 200 177 270 203
rect 200 143 218 177
rect 252 143 270 177
rect 200 117 270 143
rect 300 177 370 203
rect 300 143 318 177
rect 352 143 370 177
rect 300 117 370 143
rect 400 177 470 203
rect 400 143 418 177
rect 452 143 470 177
rect 400 117 470 143
rect 500 177 570 203
rect 500 143 518 177
rect 552 143 570 177
rect 500 117 570 143
rect 600 177 670 203
rect 600 143 618 177
rect 652 143 670 177
rect 600 117 670 143
rect 700 177 770 203
rect 700 143 718 177
rect 752 143 770 177
rect 700 117 770 143
rect 800 117 870 203
rect 900 117 970 203
rect 1000 117 1070 203
rect 1100 117 1170 203
rect 1200 177 1270 203
rect 1200 143 1218 177
rect 1252 143 1270 177
rect 1200 117 1270 143
rect 1300 177 1370 203
rect 1300 143 1318 177
rect 1352 143 1370 177
rect 1300 117 1370 143
rect 1400 177 1470 203
rect 1400 143 1418 177
rect 1452 143 1470 177
rect 1400 117 1470 143
rect 1500 177 1570 203
rect 1500 143 1518 177
rect 1552 143 1570 177
rect 1500 117 1570 143
rect 1600 177 1654 203
rect 1600 143 1612 177
rect 1646 143 1654 177
rect 1600 117 1654 143
rect 2516 737 2570 763
rect 2516 703 2524 737
rect 2558 703 2570 737
rect 2516 677 2570 703
rect 2600 737 2670 763
rect 2600 703 2618 737
rect 2652 703 2670 737
rect 2600 677 2670 703
rect 2700 737 2770 763
rect 2700 703 2718 737
rect 2752 703 2770 737
rect 2700 677 2770 703
rect 2800 737 2854 763
rect 2800 703 2812 737
rect 2846 703 2854 737
rect 2800 677 2854 703
rect 2216 597 2270 623
rect 2216 563 2224 597
rect 2258 563 2270 597
rect 2216 537 2270 563
rect 2300 597 2370 623
rect 2300 563 2318 597
rect 2352 563 2370 597
rect 2300 537 2370 563
rect 2400 597 2470 623
rect 2400 563 2418 597
rect 2452 563 2470 597
rect 2400 537 2470 563
rect 2500 537 2570 623
rect 2600 597 2670 623
rect 2600 563 2618 597
rect 2652 563 2670 597
rect 2600 537 2670 563
rect 2700 597 2754 623
rect 2700 563 2712 597
rect 2746 563 2754 597
rect 2700 537 2754 563
rect 1916 457 1970 483
rect 1916 423 1924 457
rect 1958 423 1970 457
rect 1916 397 1970 423
rect 2000 457 2070 483
rect 2000 423 2018 457
rect 2052 423 2070 457
rect 2000 397 2070 423
rect 2100 397 2170 483
rect 2200 457 2270 483
rect 2200 423 2218 457
rect 2252 423 2270 457
rect 2200 397 2270 423
rect 2300 457 2354 483
rect 2300 423 2312 457
rect 2346 423 2354 457
rect 2300 397 2354 423
rect 2416 457 2470 483
rect 2416 423 2424 457
rect 2458 423 2470 457
rect 2416 397 2470 423
rect 2500 457 2570 483
rect 2500 423 2518 457
rect 2552 423 2570 457
rect 2500 397 2570 423
rect 2600 457 2654 483
rect 2600 423 2612 457
rect 2646 423 2654 457
rect 2600 397 2654 423
rect 3316 1157 3370 1183
rect 3316 1123 3324 1157
rect 3358 1123 3370 1157
rect 3316 1097 3370 1123
rect 3400 1157 3470 1183
rect 3400 1123 3418 1157
rect 3452 1123 3470 1157
rect 3400 1097 3470 1123
rect 3500 1097 3570 1183
rect 3600 1157 3670 1183
rect 3600 1123 3618 1157
rect 3652 1123 3670 1157
rect 3600 1097 3670 1123
rect 3700 1157 3754 1183
rect 3700 1123 3712 1157
rect 3746 1123 3754 1157
rect 3700 1097 3754 1123
rect 3216 1017 3270 1043
rect 3216 983 3224 1017
rect 3258 983 3270 1017
rect 3216 957 3270 983
rect 3300 1017 3354 1043
rect 3300 983 3312 1017
rect 3346 983 3354 1017
rect 3300 957 3354 983
rect 3416 1017 3470 1043
rect 3416 983 3424 1017
rect 3458 983 3470 1017
rect 3416 957 3470 983
rect 3500 1017 3570 1043
rect 3500 983 3518 1017
rect 3552 983 3570 1017
rect 3500 957 3570 983
rect 3600 1017 3654 1043
rect 3600 983 3612 1017
rect 3646 983 3654 1017
rect 3600 957 3654 983
rect 3816 1157 3870 1183
rect 3816 1123 3824 1157
rect 3858 1123 3870 1157
rect 3816 1097 3870 1123
rect 3900 1157 3970 1183
rect 3900 1123 3918 1157
rect 3952 1123 3970 1157
rect 3900 1097 3970 1123
rect 4000 1157 4070 1183
rect 4000 1123 4018 1157
rect 4052 1123 4070 1157
rect 4000 1097 4070 1123
rect 4100 1097 4170 1183
rect 4200 1097 4270 1183
rect 4300 1157 4370 1183
rect 4300 1123 4318 1157
rect 4352 1123 4370 1157
rect 4300 1097 4370 1123
rect 4400 1157 4454 1183
rect 4400 1123 4412 1157
rect 4446 1123 4454 1157
rect 4400 1097 4454 1123
rect 3716 1017 3770 1043
rect 3716 983 3724 1017
rect 3758 983 3770 1017
rect 3716 957 3770 983
rect 3800 1017 3854 1043
rect 3800 983 3812 1017
rect 3846 983 3854 1017
rect 3800 957 3854 983
rect 3016 877 3070 903
rect 3016 843 3024 877
rect 3058 843 3070 877
rect 3016 817 3070 843
rect 3100 877 3170 903
rect 3100 843 3118 877
rect 3152 843 3170 877
rect 3100 817 3170 843
rect 3200 817 3270 903
rect 3300 877 3370 903
rect 3300 843 3318 877
rect 3352 843 3370 877
rect 3300 817 3370 843
rect 3400 877 3470 903
rect 3400 843 3418 877
rect 3452 843 3470 877
rect 3400 817 3470 843
rect 3500 877 3570 903
rect 3500 843 3518 877
rect 3552 843 3570 877
rect 3500 817 3570 843
rect 3600 877 3670 903
rect 3600 843 3618 877
rect 3652 843 3670 877
rect 3600 817 3670 843
rect 3700 877 3770 903
rect 3700 843 3718 877
rect 3752 843 3770 877
rect 3700 817 3770 843
rect 3800 877 3854 903
rect 3800 843 3812 877
rect 3846 843 3854 877
rect 3800 817 3854 843
rect 2916 737 2970 763
rect 2916 703 2924 737
rect 2958 703 2970 737
rect 2916 677 2970 703
rect 3000 737 3054 763
rect 3000 703 3012 737
rect 3046 703 3054 737
rect 3000 677 3054 703
rect 3116 737 3170 763
rect 3116 703 3124 737
rect 3158 703 3170 737
rect 3116 677 3170 703
rect 3200 737 3270 763
rect 3200 703 3218 737
rect 3252 703 3270 737
rect 3200 677 3270 703
rect 3300 737 3354 763
rect 3300 703 3312 737
rect 3346 703 3354 737
rect 3300 677 3354 703
rect 3416 737 3470 763
rect 3416 703 3424 737
rect 3458 703 3470 737
rect 3416 677 3470 703
rect 3500 737 3570 763
rect 3500 703 3518 737
rect 3552 703 3570 737
rect 3500 677 3570 703
rect 3600 737 3654 763
rect 3600 703 3612 737
rect 3646 703 3654 737
rect 3600 677 3654 703
rect 4716 1387 4770 1413
rect 4716 1353 4724 1387
rect 4758 1353 4770 1387
rect 4716 1327 4770 1353
rect 4800 1387 4854 1413
rect 4800 1353 4812 1387
rect 4846 1353 4854 1387
rect 4800 1327 4854 1353
rect 4516 1157 4570 1183
rect 4516 1123 4524 1157
rect 4558 1123 4570 1157
rect 4516 1097 4570 1123
rect 4600 1157 4654 1183
rect 4600 1123 4612 1157
rect 4646 1123 4654 1157
rect 4600 1097 4654 1123
rect 5016 1667 5070 1693
rect 5016 1633 5024 1667
rect 5058 1633 5070 1667
rect 5016 1607 5070 1633
rect 5100 1667 5170 1693
rect 5100 1633 5118 1667
rect 5152 1633 5170 1667
rect 5100 1607 5170 1633
rect 5200 1667 5254 1693
rect 5200 1633 5212 1667
rect 5246 1633 5254 1667
rect 5200 1607 5254 1633
rect 5316 1667 5370 1693
rect 5316 1633 5324 1667
rect 5358 1633 5370 1667
rect 5316 1607 5370 1633
rect 5400 1667 5470 1693
rect 5400 1633 5418 1667
rect 5452 1633 5470 1667
rect 5400 1607 5470 1633
rect 5500 1667 5570 1693
rect 5500 1633 5518 1667
rect 5552 1633 5570 1667
rect 5500 1607 5570 1633
rect 5600 1667 5654 1693
rect 5600 1633 5612 1667
rect 5646 1633 5654 1667
rect 5600 1607 5654 1633
rect 5716 1667 5770 1693
rect 5716 1633 5724 1667
rect 5758 1633 5770 1667
rect 5716 1607 5770 1633
rect 5800 1667 5870 1693
rect 5800 1633 5818 1667
rect 5852 1633 5870 1667
rect 5800 1607 5870 1633
rect 5900 1667 5954 1693
rect 5900 1633 5912 1667
rect 5946 1633 5954 1667
rect 5900 1607 5954 1633
rect 4916 1527 4970 1553
rect 4916 1493 4924 1527
rect 4958 1493 4970 1527
rect 4916 1467 4970 1493
rect 5000 1527 5070 1553
rect 5000 1493 5018 1527
rect 5052 1493 5070 1527
rect 5000 1467 5070 1493
rect 5100 1527 5170 1553
rect 5100 1493 5118 1527
rect 5152 1493 5170 1527
rect 5100 1467 5170 1493
rect 5200 1527 5270 1553
rect 5200 1493 5218 1527
rect 5252 1493 5270 1527
rect 5200 1467 5270 1493
rect 5300 1527 5370 1553
rect 5300 1493 5318 1527
rect 5352 1493 5370 1527
rect 5300 1467 5370 1493
rect 5400 1527 5470 1553
rect 5400 1493 5418 1527
rect 5452 1493 5470 1527
rect 5400 1467 5470 1493
rect 5500 1527 5570 1553
rect 5500 1493 5518 1527
rect 5552 1493 5570 1527
rect 5500 1467 5570 1493
rect 5600 1467 5670 1553
rect 5700 1527 5770 1553
rect 5700 1493 5718 1527
rect 5752 1493 5770 1527
rect 5700 1467 5770 1493
rect 5800 1527 5854 1553
rect 5800 1493 5812 1527
rect 5846 1493 5854 1527
rect 5800 1467 5854 1493
rect 4916 1387 4970 1413
rect 4916 1353 4924 1387
rect 4958 1353 4970 1387
rect 4916 1327 4970 1353
rect 5000 1387 5070 1413
rect 5000 1353 5018 1387
rect 5052 1353 5070 1387
rect 5000 1327 5070 1353
rect 5100 1387 5154 1413
rect 5100 1353 5112 1387
rect 5146 1353 5154 1387
rect 5100 1327 5154 1353
rect 6016 1667 6070 1693
rect 6016 1633 6024 1667
rect 6058 1633 6070 1667
rect 6016 1607 6070 1633
rect 6100 1667 6154 1693
rect 6100 1633 6112 1667
rect 6146 1633 6154 1667
rect 6100 1607 6154 1633
rect 5916 1527 5970 1553
rect 5916 1493 5924 1527
rect 5958 1493 5970 1527
rect 5916 1467 5970 1493
rect 6000 1527 6054 1553
rect 6000 1493 6012 1527
rect 6046 1493 6054 1527
rect 6000 1467 6054 1493
rect 7016 2367 7070 2393
rect 7016 2333 7024 2367
rect 7058 2333 7070 2367
rect 7016 2307 7070 2333
rect 7100 2367 7170 2393
rect 7100 2333 7118 2367
rect 7152 2333 7170 2367
rect 7100 2307 7170 2333
rect 7200 2367 7254 2393
rect 7200 2333 7212 2367
rect 7246 2333 7254 2367
rect 7200 2307 7254 2333
rect 8316 2737 8370 2763
rect 8316 2703 8324 2737
rect 8358 2703 8370 2737
rect 8316 2677 8370 2703
rect 8400 2737 8470 2763
rect 8400 2703 8418 2737
rect 8452 2703 8470 2737
rect 8400 2677 8470 2703
rect 8500 2737 8570 2763
rect 8500 2703 8518 2737
rect 8552 2703 8570 2737
rect 8500 2677 8570 2703
rect 8600 2737 8670 2763
rect 8600 2703 8618 2737
rect 8652 2703 8670 2737
rect 8600 2677 8670 2703
rect 8700 2737 8754 2763
rect 8700 2703 8712 2737
rect 8746 2703 8754 2737
rect 8700 2677 8754 2703
rect 8316 2597 8370 2623
rect 8316 2563 8324 2597
rect 8358 2563 8370 2597
rect 8316 2537 8370 2563
rect 8400 2597 8454 2623
rect 8400 2563 8412 2597
rect 8446 2563 8454 2597
rect 8400 2537 8454 2563
rect 8516 2597 8570 2623
rect 8516 2563 8524 2597
rect 8558 2563 8570 2597
rect 8516 2537 8570 2563
rect 8600 2597 8670 2623
rect 8600 2563 8618 2597
rect 8652 2563 8670 2597
rect 8600 2537 8670 2563
rect 8700 2597 8754 2623
rect 8700 2563 8712 2597
rect 8746 2563 8754 2597
rect 8700 2537 8754 2563
rect 7316 2367 7370 2393
rect 7316 2333 7324 2367
rect 7358 2333 7370 2367
rect 7316 2307 7370 2333
rect 7400 2367 7470 2393
rect 7400 2333 7418 2367
rect 7452 2333 7470 2367
rect 7400 2307 7470 2333
rect 7500 2307 7570 2393
rect 7600 2307 7670 2393
rect 7700 2367 7770 2393
rect 7700 2333 7718 2367
rect 7752 2333 7770 2367
rect 7700 2307 7770 2333
rect 7800 2367 7870 2393
rect 7800 2333 7818 2367
rect 7852 2333 7870 2367
rect 7800 2307 7870 2333
rect 7900 2307 7970 2393
rect 8000 2307 8070 2393
rect 8100 2307 8170 2393
rect 8200 2307 8270 2393
rect 8300 2307 8370 2393
rect 8400 2367 8470 2393
rect 8400 2333 8418 2367
rect 8452 2333 8470 2367
rect 8400 2307 8470 2333
rect 8500 2367 8554 2393
rect 8500 2333 8512 2367
rect 8546 2333 8554 2367
rect 8500 2307 8554 2333
rect 7016 2227 7070 2253
rect 7016 2193 7024 2227
rect 7058 2193 7070 2227
rect 7016 2167 7070 2193
rect 7100 2227 7170 2253
rect 7100 2193 7118 2227
rect 7152 2193 7170 2227
rect 7100 2167 7170 2193
rect 7200 2167 7270 2253
rect 7300 2167 7370 2253
rect 7400 2227 7470 2253
rect 7400 2193 7418 2227
rect 7452 2193 7470 2227
rect 7400 2167 7470 2193
rect 7500 2227 7554 2253
rect 7500 2193 7512 2227
rect 7546 2193 7554 2227
rect 7500 2167 7554 2193
rect 7616 2227 7670 2253
rect 7616 2193 7624 2227
rect 7658 2193 7670 2227
rect 7616 2167 7670 2193
rect 7700 2227 7754 2253
rect 7700 2193 7712 2227
rect 7746 2193 7754 2227
rect 7700 2167 7754 2193
rect 10116 3577 10170 3603
rect 10116 3543 10124 3577
rect 10158 3543 10170 3577
rect 10116 3517 10170 3543
rect 10200 3577 10270 3603
rect 10200 3543 10218 3577
rect 10252 3543 10270 3577
rect 10200 3517 10270 3543
rect 10300 3517 10370 3603
rect 10400 3517 10470 3603
rect 10500 3577 10570 3603
rect 10500 3543 10518 3577
rect 10552 3543 10570 3577
rect 10500 3517 10570 3543
rect 10600 3577 10654 3603
rect 10600 3543 10612 3577
rect 10646 3543 10654 3577
rect 10600 3517 10654 3543
rect 11216 3807 11270 3833
rect 11216 3773 11224 3807
rect 11258 3773 11270 3807
rect 11216 3747 11270 3773
rect 11300 3807 11370 3833
rect 11300 3773 11318 3807
rect 11352 3773 11370 3807
rect 11300 3747 11370 3773
rect 11400 3807 11470 3833
rect 11400 3773 11418 3807
rect 11452 3773 11470 3807
rect 11400 3747 11470 3773
rect 11500 3807 11554 3833
rect 11500 3773 11512 3807
rect 11546 3773 11554 3807
rect 11500 3747 11554 3773
rect 11616 3807 11670 3833
rect 11616 3773 11624 3807
rect 11658 3773 11670 3807
rect 11616 3747 11670 3773
rect 11700 3807 11770 3833
rect 11700 3773 11718 3807
rect 11752 3773 11770 3807
rect 11700 3747 11770 3773
rect 11800 3807 11870 3833
rect 11800 3773 11818 3807
rect 11852 3773 11870 3807
rect 11800 3747 11870 3773
rect 11900 3807 11970 3833
rect 11900 3773 11918 3807
rect 11952 3773 11970 3807
rect 11900 3747 11970 3773
rect 12000 3807 12070 3833
rect 12000 3773 12018 3807
rect 12052 3773 12070 3807
rect 12000 3747 12070 3773
rect 12100 3807 12154 3833
rect 12100 3773 12112 3807
rect 12146 3773 12154 3807
rect 12100 3747 12154 3773
rect 10716 3577 10770 3603
rect 10716 3543 10724 3577
rect 10758 3543 10770 3577
rect 10716 3517 10770 3543
rect 10800 3577 10870 3603
rect 10800 3543 10818 3577
rect 10852 3543 10870 3577
rect 10800 3517 10870 3543
rect 10900 3577 10970 3603
rect 10900 3543 10918 3577
rect 10952 3543 10970 3577
rect 10900 3517 10970 3543
rect 11000 3517 11070 3603
rect 11100 3517 11170 3603
rect 11200 3517 11270 3603
rect 11300 3577 11370 3603
rect 11300 3543 11318 3577
rect 11352 3543 11370 3577
rect 11300 3517 11370 3543
rect 11400 3577 11454 3603
rect 11400 3543 11412 3577
rect 11446 3543 11454 3577
rect 11400 3517 11454 3543
rect 9816 3437 9870 3463
rect 9816 3403 9824 3437
rect 9858 3403 9870 3437
rect 9816 3377 9870 3403
rect 9900 3437 9970 3463
rect 9900 3403 9918 3437
rect 9952 3403 9970 3437
rect 9900 3377 9970 3403
rect 10000 3437 10070 3463
rect 10000 3403 10018 3437
rect 10052 3403 10070 3437
rect 10000 3377 10070 3403
rect 10100 3377 10170 3463
rect 10200 3377 10270 3463
rect 10300 3437 10370 3463
rect 10300 3403 10318 3437
rect 10352 3403 10370 3437
rect 10300 3377 10370 3403
rect 10400 3437 10470 3463
rect 10400 3403 10418 3437
rect 10452 3403 10470 3437
rect 10400 3377 10470 3403
rect 10500 3377 10570 3463
rect 10600 3377 10670 3463
rect 10700 3377 10770 3463
rect 10800 3377 10870 3463
rect 10900 3437 10970 3463
rect 10900 3403 10918 3437
rect 10952 3403 10970 3437
rect 10900 3377 10970 3403
rect 11000 3437 11070 3463
rect 11000 3403 11018 3437
rect 11052 3403 11070 3437
rect 11000 3377 11070 3403
rect 11100 3377 11170 3463
rect 11200 3377 11270 3463
rect 11300 3437 11370 3463
rect 11300 3403 11318 3437
rect 11352 3403 11370 3437
rect 11300 3377 11370 3403
rect 11400 3437 11454 3463
rect 11400 3403 11412 3437
rect 11446 3403 11454 3437
rect 11400 3377 11454 3403
rect 9616 3297 9670 3323
rect 9616 3263 9624 3297
rect 9658 3263 9670 3297
rect 9616 3237 9670 3263
rect 9700 3297 9770 3323
rect 9700 3263 9718 3297
rect 9752 3263 9770 3297
rect 9700 3237 9770 3263
rect 9800 3297 9870 3323
rect 9800 3263 9818 3297
rect 9852 3263 9870 3297
rect 9800 3237 9870 3263
rect 9900 3237 9970 3323
rect 10000 3237 10070 3323
rect 10100 3297 10170 3323
rect 10100 3263 10118 3297
rect 10152 3263 10170 3297
rect 10100 3237 10170 3263
rect 10200 3297 10270 3323
rect 10200 3263 10218 3297
rect 10252 3263 10270 3297
rect 10200 3237 10270 3263
rect 10300 3297 10354 3323
rect 10300 3263 10312 3297
rect 10346 3263 10354 3297
rect 10300 3237 10354 3263
rect 8916 3157 8970 3183
rect 8916 3123 8924 3157
rect 8958 3123 8970 3157
rect 8916 3097 8970 3123
rect 9000 3157 9070 3183
rect 9000 3123 9018 3157
rect 9052 3123 9070 3157
rect 9000 3097 9070 3123
rect 9100 3157 9170 3183
rect 9100 3123 9118 3157
rect 9152 3123 9170 3157
rect 9100 3097 9170 3123
rect 9200 3157 9270 3183
rect 9200 3123 9218 3157
rect 9252 3123 9270 3157
rect 9200 3097 9270 3123
rect 9300 3097 9370 3183
rect 9400 3157 9470 3183
rect 9400 3123 9418 3157
rect 9452 3123 9470 3157
rect 9400 3097 9470 3123
rect 9500 3157 9570 3183
rect 9500 3123 9518 3157
rect 9552 3123 9570 3157
rect 9500 3097 9570 3123
rect 9600 3157 9670 3183
rect 9600 3123 9618 3157
rect 9652 3123 9670 3157
rect 9600 3097 9670 3123
rect 9700 3157 9770 3183
rect 9700 3123 9718 3157
rect 9752 3123 9770 3157
rect 9700 3097 9770 3123
rect 9800 3157 9870 3183
rect 9800 3123 9818 3157
rect 9852 3123 9870 3157
rect 9800 3097 9870 3123
rect 9900 3157 9954 3183
rect 9900 3123 9912 3157
rect 9946 3123 9954 3157
rect 9900 3097 9954 3123
rect 8916 3017 8970 3043
rect 8916 2983 8924 3017
rect 8958 2983 8970 3017
rect 8916 2957 8970 2983
rect 9000 3017 9070 3043
rect 9000 2983 9018 3017
rect 9052 2983 9070 3017
rect 9000 2957 9070 2983
rect 9100 3017 9154 3043
rect 9100 2983 9112 3017
rect 9146 2983 9154 3017
rect 9100 2957 9154 2983
rect 9216 3017 9270 3043
rect 9216 2983 9224 3017
rect 9258 2983 9270 3017
rect 9216 2957 9270 2983
rect 9300 3017 9370 3043
rect 9300 2983 9318 3017
rect 9352 2983 9370 3017
rect 9300 2957 9370 2983
rect 9400 3017 9454 3043
rect 9400 2983 9412 3017
rect 9446 2983 9454 3017
rect 9400 2957 9454 2983
rect 10016 3157 10070 3183
rect 10016 3123 10024 3157
rect 10058 3123 10070 3157
rect 10016 3097 10070 3123
rect 10100 3157 10154 3183
rect 10100 3123 10112 3157
rect 10146 3123 10154 3157
rect 10100 3097 10154 3123
rect 10216 3157 10270 3183
rect 10216 3123 10224 3157
rect 10258 3123 10270 3157
rect 10216 3097 10270 3123
rect 10300 3157 10354 3183
rect 10300 3123 10312 3157
rect 10346 3123 10354 3157
rect 10300 3097 10354 3123
rect 10416 3297 10470 3323
rect 10416 3263 10424 3297
rect 10458 3263 10470 3297
rect 10416 3237 10470 3263
rect 10500 3297 10554 3323
rect 10500 3263 10512 3297
rect 10546 3263 10554 3297
rect 10500 3237 10554 3263
rect 12216 3807 12270 3833
rect 12216 3773 12224 3807
rect 12258 3773 12270 3807
rect 12216 3747 12270 3773
rect 12300 3807 12370 3833
rect 12300 3773 12318 3807
rect 12352 3773 12370 3807
rect 12300 3747 12370 3773
rect 12400 3807 12470 3833
rect 12400 3773 12418 3807
rect 12452 3773 12470 3807
rect 12400 3747 12470 3773
rect 12500 3807 12570 3833
rect 12500 3773 12518 3807
rect 12552 3773 12570 3807
rect 12500 3747 12570 3773
rect 12600 3747 12670 3833
rect 12700 3747 12770 3833
rect 12800 3747 12854 3833
rect 12912 3822 12970 3833
rect 12912 3788 12924 3822
rect 12958 3788 12970 3822
rect 12912 3747 12970 3788
rect 13000 3807 13070 3833
rect 13000 3773 13018 3807
rect 13052 3773 13070 3807
rect 13000 3747 13070 3773
rect 13100 3792 13158 3833
rect 13100 3758 13112 3792
rect 13146 3758 13158 3792
rect 13100 3747 13158 3758
rect 13220 3807 13280 3833
rect 13220 3773 13228 3807
rect 13262 3773 13280 3807
rect 13220 3747 13280 3773
rect 13310 3807 13380 3833
rect 13310 3773 13328 3807
rect 13362 3773 13380 3807
rect 13310 3747 13380 3773
rect 13410 3807 13480 3833
rect 13410 3773 13428 3807
rect 13462 3773 13480 3807
rect 13410 3747 13480 3773
rect 13510 3807 13580 3833
rect 13510 3773 13528 3807
rect 13562 3773 13580 3807
rect 13510 3747 13580 3773
rect 13610 3807 13670 3833
rect 13610 3773 13628 3807
rect 13662 3773 13670 3807
rect 13610 3747 13670 3773
rect 11516 3577 11570 3603
rect 11516 3543 11524 3577
rect 11558 3543 11570 3577
rect 11516 3517 11570 3543
rect 11600 3577 11670 3603
rect 11600 3543 11618 3577
rect 11652 3543 11670 3577
rect 11600 3517 11670 3543
rect 11700 3577 11770 3603
rect 11700 3543 11718 3577
rect 11752 3543 11770 3577
rect 11700 3517 11770 3543
rect 11800 3517 11870 3603
rect 11900 3517 11970 3603
rect 12000 3577 12070 3603
rect 12000 3543 12018 3577
rect 12052 3543 12070 3577
rect 12000 3517 12070 3543
rect 12100 3577 12170 3603
rect 12100 3543 12118 3577
rect 12152 3543 12170 3577
rect 12100 3517 12170 3543
rect 12200 3577 12270 3603
rect 12200 3543 12218 3577
rect 12252 3543 12270 3577
rect 12200 3517 12270 3543
rect 12300 3517 12370 3603
rect 12400 3517 12470 3603
rect 12500 3577 12570 3603
rect 12500 3543 12518 3577
rect 12552 3543 12570 3577
rect 12500 3517 12570 3543
rect 12600 3577 12670 3603
rect 12600 3543 12618 3577
rect 12652 3543 12670 3577
rect 12600 3517 12670 3543
rect 12700 3517 12770 3603
rect 12800 3517 12854 3603
rect 12912 3592 12970 3603
rect 12912 3558 12924 3592
rect 12958 3558 12970 3592
rect 12912 3517 12970 3558
rect 13000 3577 13070 3603
rect 13000 3543 13018 3577
rect 13052 3543 13070 3577
rect 13000 3517 13070 3543
rect 13100 3562 13158 3603
rect 13100 3528 13112 3562
rect 13146 3528 13158 3562
rect 13100 3517 13158 3528
rect 13220 3577 13280 3603
rect 13220 3543 13228 3577
rect 13262 3543 13280 3577
rect 13220 3517 13280 3543
rect 13310 3577 13380 3603
rect 13310 3543 13328 3577
rect 13362 3543 13380 3577
rect 13310 3517 13380 3543
rect 13410 3577 13480 3603
rect 13410 3543 13428 3577
rect 13462 3543 13480 3577
rect 13410 3517 13480 3543
rect 13510 3577 13580 3603
rect 13510 3543 13528 3577
rect 13562 3543 13580 3577
rect 13510 3517 13580 3543
rect 13610 3577 13670 3603
rect 13610 3543 13628 3577
rect 13662 3543 13670 3577
rect 13610 3517 13670 3543
rect 11516 3437 11570 3463
rect 11516 3403 11524 3437
rect 11558 3403 11570 3437
rect 11516 3377 11570 3403
rect 11600 3437 11670 3463
rect 11600 3403 11618 3437
rect 11652 3403 11670 3437
rect 11600 3377 11670 3403
rect 11700 3437 11770 3463
rect 11700 3403 11718 3437
rect 11752 3403 11770 3437
rect 11700 3377 11770 3403
rect 11800 3377 11870 3463
rect 11900 3437 11970 3463
rect 11900 3403 11918 3437
rect 11952 3403 11970 3437
rect 11900 3377 11970 3403
rect 12000 3437 12070 3463
rect 12000 3403 12018 3437
rect 12052 3403 12070 3437
rect 12000 3377 12070 3403
rect 12100 3437 12154 3463
rect 12100 3403 12112 3437
rect 12146 3403 12154 3437
rect 12100 3377 12154 3403
rect 12216 3437 12270 3463
rect 12216 3403 12224 3437
rect 12258 3403 12270 3437
rect 12216 3377 12270 3403
rect 12300 3437 12370 3463
rect 12300 3403 12318 3437
rect 12352 3403 12370 3437
rect 12300 3377 12370 3403
rect 12400 3377 12470 3463
rect 12500 3377 12570 3463
rect 12600 3437 12670 3463
rect 12600 3403 12618 3437
rect 12652 3403 12670 3437
rect 12600 3377 12670 3403
rect 12700 3437 12770 3463
rect 12700 3403 12718 3437
rect 12752 3403 12770 3437
rect 12700 3377 12770 3403
rect 12800 3437 12854 3463
rect 12800 3403 12812 3437
rect 12846 3403 12854 3437
rect 12800 3377 12854 3403
rect 12912 3452 12970 3463
rect 12912 3418 12924 3452
rect 12958 3418 12970 3452
rect 12912 3377 12970 3418
rect 13000 3437 13070 3463
rect 13000 3403 13018 3437
rect 13052 3403 13070 3437
rect 13000 3377 13070 3403
rect 13100 3422 13158 3463
rect 13100 3388 13112 3422
rect 13146 3388 13158 3422
rect 13100 3377 13158 3388
rect 13220 3437 13280 3463
rect 13220 3403 13228 3437
rect 13262 3403 13280 3437
rect 13220 3377 13280 3403
rect 13310 3437 13380 3463
rect 13310 3403 13328 3437
rect 13362 3403 13380 3437
rect 13310 3377 13380 3403
rect 13410 3437 13480 3463
rect 13410 3403 13428 3437
rect 13462 3403 13480 3437
rect 13410 3377 13480 3403
rect 13510 3437 13580 3463
rect 13510 3403 13528 3437
rect 13562 3403 13580 3437
rect 13510 3377 13580 3403
rect 13610 3437 13670 3463
rect 13610 3403 13628 3437
rect 13662 3403 13670 3437
rect 13610 3377 13670 3403
rect 10616 3297 10670 3323
rect 10616 3263 10624 3297
rect 10658 3263 10670 3297
rect 10616 3237 10670 3263
rect 10700 3297 10770 3323
rect 10700 3263 10718 3297
rect 10752 3263 10770 3297
rect 10700 3237 10770 3263
rect 10800 3297 10870 3323
rect 10800 3263 10818 3297
rect 10852 3263 10870 3297
rect 10800 3237 10870 3263
rect 10900 3297 10970 3323
rect 10900 3263 10918 3297
rect 10952 3263 10970 3297
rect 10900 3237 10970 3263
rect 11000 3297 11070 3323
rect 11000 3263 11018 3297
rect 11052 3263 11070 3297
rect 11000 3237 11070 3263
rect 11100 3297 11170 3323
rect 11100 3263 11118 3297
rect 11152 3263 11170 3297
rect 11100 3237 11170 3263
rect 11200 3297 11270 3323
rect 11200 3263 11218 3297
rect 11252 3263 11270 3297
rect 11200 3237 11270 3263
rect 11300 3297 11370 3323
rect 11300 3263 11318 3297
rect 11352 3263 11370 3297
rect 11300 3237 11370 3263
rect 11400 3297 11470 3323
rect 11400 3263 11418 3297
rect 11452 3263 11470 3297
rect 11400 3237 11470 3263
rect 11500 3297 11570 3323
rect 11500 3263 11518 3297
rect 11552 3263 11570 3297
rect 11500 3237 11570 3263
rect 11600 3297 11670 3323
rect 11600 3263 11618 3297
rect 11652 3263 11670 3297
rect 11600 3237 11670 3263
rect 11700 3297 11770 3323
rect 11700 3263 11718 3297
rect 11752 3263 11770 3297
rect 11700 3237 11770 3263
rect 11800 3297 11870 3323
rect 11800 3263 11818 3297
rect 11852 3263 11870 3297
rect 11800 3237 11870 3263
rect 11900 3237 11970 3323
rect 12000 3237 12070 3323
rect 12100 3237 12170 3323
rect 12200 3237 12270 3323
rect 12300 3297 12370 3323
rect 12300 3263 12318 3297
rect 12352 3263 12370 3297
rect 12300 3237 12370 3263
rect 12400 3297 12454 3323
rect 12400 3263 12412 3297
rect 12446 3263 12454 3297
rect 12400 3237 12454 3263
rect 10416 3157 10470 3183
rect 10416 3123 10424 3157
rect 10458 3123 10470 3157
rect 10416 3097 10470 3123
rect 10500 3157 10570 3183
rect 10500 3123 10518 3157
rect 10552 3123 10570 3157
rect 10500 3097 10570 3123
rect 10600 3097 10670 3183
rect 10700 3157 10770 3183
rect 10700 3123 10718 3157
rect 10752 3123 10770 3157
rect 10700 3097 10770 3123
rect 10800 3157 10854 3183
rect 10800 3123 10812 3157
rect 10846 3123 10854 3157
rect 10800 3097 10854 3123
rect 10916 3157 10970 3183
rect 10916 3123 10924 3157
rect 10958 3123 10970 3157
rect 10916 3097 10970 3123
rect 11000 3157 11070 3183
rect 11000 3123 11018 3157
rect 11052 3123 11070 3157
rect 11000 3097 11070 3123
rect 11100 3157 11170 3183
rect 11100 3123 11118 3157
rect 11152 3123 11170 3157
rect 11100 3097 11170 3123
rect 11200 3097 11270 3183
rect 11300 3097 11370 3183
rect 11400 3157 11470 3183
rect 11400 3123 11418 3157
rect 11452 3123 11470 3157
rect 11400 3097 11470 3123
rect 11500 3157 11554 3183
rect 11500 3123 11512 3157
rect 11546 3123 11554 3157
rect 11500 3097 11554 3123
rect 9516 3017 9570 3043
rect 9516 2983 9524 3017
rect 9558 2983 9570 3017
rect 9516 2957 9570 2983
rect 9600 3017 9670 3043
rect 9600 2983 9618 3017
rect 9652 2983 9670 3017
rect 9600 2957 9670 2983
rect 9700 2957 9770 3043
rect 9800 2957 9870 3043
rect 9900 3017 9970 3043
rect 9900 2983 9918 3017
rect 9952 2983 9970 3017
rect 9900 2957 9970 2983
rect 10000 3017 10070 3043
rect 10000 2983 10018 3017
rect 10052 2983 10070 3017
rect 10000 2957 10070 2983
rect 10100 3017 10170 3043
rect 10100 2983 10118 3017
rect 10152 2983 10170 3017
rect 10100 2957 10170 2983
rect 10200 2957 10270 3043
rect 10300 2957 10370 3043
rect 10400 3017 10470 3043
rect 10400 2983 10418 3017
rect 10452 2983 10470 3017
rect 10400 2957 10470 2983
rect 10500 3017 10570 3043
rect 10500 2983 10518 3017
rect 10552 2983 10570 3017
rect 10500 2957 10570 2983
rect 10600 3017 10670 3043
rect 10600 2983 10618 3017
rect 10652 2983 10670 3017
rect 10600 2957 10670 2983
rect 10700 2957 10770 3043
rect 10800 2957 10870 3043
rect 10900 2957 10970 3043
rect 11000 3017 11070 3043
rect 11000 2983 11018 3017
rect 11052 2983 11070 3017
rect 11000 2957 11070 2983
rect 11100 3017 11170 3043
rect 11100 2983 11118 3017
rect 11152 2983 11170 3017
rect 11100 2957 11170 2983
rect 11200 2957 11270 3043
rect 11300 3017 11370 3043
rect 11300 2983 11318 3017
rect 11352 2983 11370 3017
rect 11300 2957 11370 2983
rect 11400 3017 11470 3043
rect 11400 2983 11418 3017
rect 11452 2983 11470 3017
rect 11400 2957 11470 2983
rect 11500 3017 11554 3043
rect 11500 2983 11512 3017
rect 11546 2983 11554 3017
rect 11500 2957 11554 2983
rect 8816 2877 8870 2903
rect 8816 2843 8824 2877
rect 8858 2843 8870 2877
rect 8816 2817 8870 2843
rect 8900 2877 8970 2903
rect 8900 2843 8918 2877
rect 8952 2843 8970 2877
rect 8900 2817 8970 2843
rect 9000 2877 9070 2903
rect 9000 2843 9018 2877
rect 9052 2843 9070 2877
rect 9000 2817 9070 2843
rect 9100 2877 9170 2903
rect 9100 2843 9118 2877
rect 9152 2843 9170 2877
rect 9100 2817 9170 2843
rect 9200 2817 9270 2903
rect 9300 2877 9370 2903
rect 9300 2843 9318 2877
rect 9352 2843 9370 2877
rect 9300 2817 9370 2843
rect 9400 2877 9470 2903
rect 9400 2843 9418 2877
rect 9452 2843 9470 2877
rect 9400 2817 9470 2843
rect 9500 2817 9570 2903
rect 9600 2817 9670 2903
rect 9700 2817 9770 2903
rect 9800 2877 9870 2903
rect 9800 2843 9818 2877
rect 9852 2843 9870 2877
rect 9800 2817 9870 2843
rect 9900 2877 9970 2903
rect 9900 2843 9918 2877
rect 9952 2843 9970 2877
rect 9900 2817 9970 2843
rect 10000 2817 10070 2903
rect 10100 2877 10170 2903
rect 10100 2843 10118 2877
rect 10152 2843 10170 2877
rect 10100 2817 10170 2843
rect 10200 2877 10270 2903
rect 10200 2843 10218 2877
rect 10252 2843 10270 2877
rect 10200 2817 10270 2843
rect 10300 2877 10370 2903
rect 10300 2843 10318 2877
rect 10352 2843 10370 2877
rect 10300 2817 10370 2843
rect 10400 2877 10470 2903
rect 10400 2843 10418 2877
rect 10452 2843 10470 2877
rect 10400 2817 10470 2843
rect 10500 2877 10554 2903
rect 10500 2843 10512 2877
rect 10546 2843 10554 2877
rect 10500 2817 10554 2843
rect 8816 2737 8870 2763
rect 8816 2703 8824 2737
rect 8858 2703 8870 2737
rect 8816 2677 8870 2703
rect 8900 2737 8954 2763
rect 8900 2703 8912 2737
rect 8946 2703 8954 2737
rect 8900 2677 8954 2703
rect 9016 2737 9070 2763
rect 9016 2703 9024 2737
rect 9058 2703 9070 2737
rect 9016 2677 9070 2703
rect 9100 2737 9154 2763
rect 9100 2703 9112 2737
rect 9146 2703 9154 2737
rect 9100 2677 9154 2703
rect 8816 2597 8870 2623
rect 8816 2563 8824 2597
rect 8858 2563 8870 2597
rect 8816 2537 8870 2563
rect 8900 2597 8970 2623
rect 8900 2563 8918 2597
rect 8952 2563 8970 2597
rect 8900 2537 8970 2563
rect 9000 2597 9054 2623
rect 9000 2563 9012 2597
rect 9046 2563 9054 2597
rect 9000 2537 9054 2563
rect 9216 2737 9270 2763
rect 9216 2703 9224 2737
rect 9258 2703 9270 2737
rect 9216 2677 9270 2703
rect 9300 2737 9354 2763
rect 9300 2703 9312 2737
rect 9346 2703 9354 2737
rect 9300 2677 9354 2703
rect 9116 2597 9170 2623
rect 9116 2563 9124 2597
rect 9158 2563 9170 2597
rect 9116 2537 9170 2563
rect 9200 2597 9254 2623
rect 9200 2563 9212 2597
rect 9246 2563 9254 2597
rect 9200 2537 9254 2563
rect 9416 2737 9470 2763
rect 9416 2703 9424 2737
rect 9458 2703 9470 2737
rect 9416 2677 9470 2703
rect 9500 2737 9554 2763
rect 9500 2703 9512 2737
rect 9546 2703 9554 2737
rect 9500 2677 9554 2703
rect 9316 2597 9370 2623
rect 9316 2563 9324 2597
rect 9358 2563 9370 2597
rect 9316 2537 9370 2563
rect 9400 2597 9470 2623
rect 9400 2563 9418 2597
rect 9452 2563 9470 2597
rect 9400 2537 9470 2563
rect 9500 2597 9554 2623
rect 9500 2563 9512 2597
rect 9546 2563 9554 2597
rect 9500 2537 9554 2563
rect 9616 2737 9670 2763
rect 9616 2703 9624 2737
rect 9658 2703 9670 2737
rect 9616 2677 9670 2703
rect 9700 2737 9770 2763
rect 9700 2703 9718 2737
rect 9752 2703 9770 2737
rect 9700 2677 9770 2703
rect 9800 2737 9870 2763
rect 9800 2703 9818 2737
rect 9852 2703 9870 2737
rect 9800 2677 9870 2703
rect 9900 2737 9954 2763
rect 9900 2703 9912 2737
rect 9946 2703 9954 2737
rect 9900 2677 9954 2703
rect 9616 2597 9670 2623
rect 9616 2563 9624 2597
rect 9658 2563 9670 2597
rect 9616 2537 9670 2563
rect 9700 2597 9770 2623
rect 9700 2563 9718 2597
rect 9752 2563 9770 2597
rect 9700 2537 9770 2563
rect 9800 2597 9870 2623
rect 9800 2563 9818 2597
rect 9852 2563 9870 2597
rect 9800 2537 9870 2563
rect 9900 2597 9954 2623
rect 9900 2563 9912 2597
rect 9946 2563 9954 2597
rect 9900 2537 9954 2563
rect 8616 2367 8670 2393
rect 8616 2333 8624 2367
rect 8658 2333 8670 2367
rect 8616 2307 8670 2333
rect 8700 2367 8770 2393
rect 8700 2333 8718 2367
rect 8752 2333 8770 2367
rect 8700 2307 8770 2333
rect 8800 2307 8870 2393
rect 8900 2367 8970 2393
rect 8900 2333 8918 2367
rect 8952 2333 8970 2367
rect 8900 2307 8970 2333
rect 9000 2367 9070 2393
rect 9000 2333 9018 2367
rect 9052 2333 9070 2367
rect 9000 2307 9070 2333
rect 9100 2367 9170 2393
rect 9100 2333 9118 2367
rect 9152 2333 9170 2367
rect 9100 2307 9170 2333
rect 9200 2307 9270 2393
rect 9300 2307 9370 2393
rect 9400 2307 9470 2393
rect 9500 2367 9570 2393
rect 9500 2333 9518 2367
rect 9552 2333 9570 2367
rect 9500 2307 9570 2333
rect 9600 2367 9654 2393
rect 9600 2333 9612 2367
rect 9646 2333 9654 2367
rect 9600 2307 9654 2333
rect 7816 2227 7870 2253
rect 7816 2193 7824 2227
rect 7858 2193 7870 2227
rect 7816 2167 7870 2193
rect 7900 2227 7970 2253
rect 7900 2193 7918 2227
rect 7952 2193 7970 2227
rect 7900 2167 7970 2193
rect 8000 2167 8070 2253
rect 8100 2167 8170 2253
rect 8200 2227 8270 2253
rect 8200 2193 8218 2227
rect 8252 2193 8270 2227
rect 8200 2167 8270 2193
rect 8300 2227 8370 2253
rect 8300 2193 8318 2227
rect 8352 2193 8370 2227
rect 8300 2167 8370 2193
rect 8400 2167 8470 2253
rect 8500 2227 8570 2253
rect 8500 2193 8518 2227
rect 8552 2193 8570 2227
rect 8500 2167 8570 2193
rect 8600 2227 8670 2253
rect 8600 2193 8618 2227
rect 8652 2193 8670 2227
rect 8600 2167 8670 2193
rect 8700 2227 8770 2253
rect 8700 2193 8718 2227
rect 8752 2193 8770 2227
rect 8700 2167 8770 2193
rect 8800 2227 8854 2253
rect 8800 2193 8812 2227
rect 8846 2193 8854 2227
rect 8800 2167 8854 2193
rect 6916 2087 6970 2113
rect 6916 2053 6924 2087
rect 6958 2053 6970 2087
rect 6916 2027 6970 2053
rect 7000 2087 7070 2113
rect 7000 2053 7018 2087
rect 7052 2053 7070 2087
rect 7000 2027 7070 2053
rect 7100 2087 7170 2113
rect 7100 2053 7118 2087
rect 7152 2053 7170 2087
rect 7100 2027 7170 2053
rect 7200 2027 7270 2113
rect 7300 2027 7370 2113
rect 7400 2087 7470 2113
rect 7400 2053 7418 2087
rect 7452 2053 7470 2087
rect 7400 2027 7470 2053
rect 7500 2087 7570 2113
rect 7500 2053 7518 2087
rect 7552 2053 7570 2087
rect 7500 2027 7570 2053
rect 7600 2027 7670 2113
rect 7700 2027 7770 2113
rect 7800 2027 7870 2113
rect 7900 2027 7970 2113
rect 8000 2087 8070 2113
rect 8000 2053 8018 2087
rect 8052 2053 8070 2087
rect 8000 2027 8070 2053
rect 8100 2087 8154 2113
rect 8100 2053 8112 2087
rect 8146 2053 8154 2087
rect 8100 2027 8154 2053
rect 6816 1947 6870 1973
rect 6816 1913 6824 1947
rect 6858 1913 6870 1947
rect 6816 1887 6870 1913
rect 6900 1947 6954 1973
rect 6900 1913 6912 1947
rect 6946 1913 6954 1947
rect 6900 1887 6954 1913
rect 8216 2087 8270 2113
rect 8216 2053 8224 2087
rect 8258 2053 8270 2087
rect 8216 2027 8270 2053
rect 8300 2087 8354 2113
rect 8300 2053 8312 2087
rect 8346 2053 8354 2087
rect 8300 2027 8354 2053
rect 8416 2087 8470 2113
rect 8416 2053 8424 2087
rect 8458 2053 8470 2087
rect 8416 2027 8470 2053
rect 8500 2087 8570 2113
rect 8500 2053 8518 2087
rect 8552 2053 8570 2087
rect 8500 2027 8570 2053
rect 8600 2087 8670 2113
rect 8600 2053 8618 2087
rect 8652 2053 8670 2087
rect 8600 2027 8670 2053
rect 8700 2087 8754 2113
rect 8700 2053 8712 2087
rect 8746 2053 8754 2087
rect 8700 2027 8754 2053
rect 8916 2227 8970 2253
rect 8916 2193 8924 2227
rect 8958 2193 8970 2227
rect 8916 2167 8970 2193
rect 9000 2227 9054 2253
rect 9000 2193 9012 2227
rect 9046 2193 9054 2227
rect 9000 2167 9054 2193
rect 8816 2087 8870 2113
rect 8816 2053 8824 2087
rect 8858 2053 8870 2087
rect 8816 2027 8870 2053
rect 8900 2087 8954 2113
rect 8900 2053 8912 2087
rect 8946 2053 8954 2087
rect 8900 2027 8954 2053
rect 9116 2227 9170 2253
rect 9116 2193 9124 2227
rect 9158 2193 9170 2227
rect 9116 2167 9170 2193
rect 9200 2227 9254 2253
rect 9200 2193 9212 2227
rect 9246 2193 9254 2227
rect 9200 2167 9254 2193
rect 9016 2087 9070 2113
rect 9016 2053 9024 2087
rect 9058 2053 9070 2087
rect 9016 2027 9070 2053
rect 9100 2087 9170 2113
rect 9100 2053 9118 2087
rect 9152 2053 9170 2087
rect 9100 2027 9170 2053
rect 9200 2087 9254 2113
rect 9200 2053 9212 2087
rect 9246 2053 9254 2087
rect 9200 2027 9254 2053
rect 9316 2227 9370 2253
rect 9316 2193 9324 2227
rect 9358 2193 9370 2227
rect 9316 2167 9370 2193
rect 9400 2227 9470 2253
rect 9400 2193 9418 2227
rect 9452 2193 9470 2227
rect 9400 2167 9470 2193
rect 9500 2227 9554 2253
rect 9500 2193 9512 2227
rect 9546 2193 9554 2227
rect 9500 2167 9554 2193
rect 10016 2737 10070 2763
rect 10016 2703 10024 2737
rect 10058 2703 10070 2737
rect 10016 2677 10070 2703
rect 10100 2737 10170 2763
rect 10100 2703 10118 2737
rect 10152 2703 10170 2737
rect 10100 2677 10170 2703
rect 10200 2737 10270 2763
rect 10200 2703 10218 2737
rect 10252 2703 10270 2737
rect 10200 2677 10270 2703
rect 10300 2737 10370 2763
rect 10300 2703 10318 2737
rect 10352 2703 10370 2737
rect 10300 2677 10370 2703
rect 10400 2737 10454 2763
rect 10400 2703 10412 2737
rect 10446 2703 10454 2737
rect 10400 2677 10454 2703
rect 10616 2877 10670 2903
rect 10616 2843 10624 2877
rect 10658 2843 10670 2877
rect 10616 2817 10670 2843
rect 10700 2877 10770 2903
rect 10700 2843 10718 2877
rect 10752 2843 10770 2877
rect 10700 2817 10770 2843
rect 10800 2817 10870 2903
rect 10900 2877 10970 2903
rect 10900 2843 10918 2877
rect 10952 2843 10970 2877
rect 10900 2817 10970 2843
rect 11000 2877 11070 2903
rect 11000 2843 11018 2877
rect 11052 2843 11070 2877
rect 11000 2817 11070 2843
rect 11100 2877 11170 2903
rect 11100 2843 11118 2877
rect 11152 2843 11170 2877
rect 11100 2817 11170 2843
rect 11200 2877 11270 2903
rect 11200 2843 11218 2877
rect 11252 2843 11270 2877
rect 11200 2817 11270 2843
rect 11300 2877 11354 2903
rect 11300 2843 11312 2877
rect 11346 2843 11354 2877
rect 11300 2817 11354 2843
rect 10516 2737 10570 2763
rect 10516 2703 10524 2737
rect 10558 2703 10570 2737
rect 10516 2677 10570 2703
rect 10600 2737 10654 2763
rect 10600 2703 10612 2737
rect 10646 2703 10654 2737
rect 10600 2677 10654 2703
rect 12516 3297 12570 3323
rect 12516 3263 12524 3297
rect 12558 3263 12570 3297
rect 12516 3237 12570 3263
rect 12600 3297 12670 3323
rect 12600 3263 12618 3297
rect 12652 3263 12670 3297
rect 12600 3237 12670 3263
rect 12700 3297 12770 3323
rect 12700 3263 12718 3297
rect 12752 3263 12770 3297
rect 12700 3237 12770 3263
rect 12800 3237 12854 3323
rect 12912 3312 12970 3323
rect 12912 3278 12924 3312
rect 12958 3278 12970 3312
rect 12912 3237 12970 3278
rect 13000 3297 13070 3323
rect 13000 3263 13018 3297
rect 13052 3263 13070 3297
rect 13000 3237 13070 3263
rect 13100 3282 13158 3323
rect 13100 3248 13112 3282
rect 13146 3248 13158 3282
rect 13100 3237 13158 3248
rect 13220 3297 13280 3323
rect 13220 3263 13228 3297
rect 13262 3263 13280 3297
rect 13220 3237 13280 3263
rect 13310 3297 13380 3323
rect 13310 3263 13328 3297
rect 13362 3263 13380 3297
rect 13310 3237 13380 3263
rect 13410 3297 13480 3323
rect 13410 3263 13428 3297
rect 13462 3263 13480 3297
rect 13410 3237 13480 3263
rect 13510 3297 13580 3323
rect 13510 3263 13528 3297
rect 13562 3263 13580 3297
rect 13510 3237 13580 3263
rect 13610 3297 13670 3323
rect 13610 3263 13628 3297
rect 13662 3263 13670 3297
rect 13610 3237 13670 3263
rect 11616 3157 11670 3183
rect 11616 3123 11624 3157
rect 11658 3123 11670 3157
rect 11616 3097 11670 3123
rect 11700 3157 11770 3183
rect 11700 3123 11718 3157
rect 11752 3123 11770 3157
rect 11700 3097 11770 3123
rect 11800 3157 11870 3183
rect 11800 3123 11818 3157
rect 11852 3123 11870 3157
rect 11800 3097 11870 3123
rect 11900 3097 11970 3183
rect 12000 3157 12070 3183
rect 12000 3123 12018 3157
rect 12052 3123 12070 3157
rect 12000 3097 12070 3123
rect 12100 3157 12170 3183
rect 12100 3123 12118 3157
rect 12152 3123 12170 3157
rect 12100 3097 12170 3123
rect 12200 3097 12270 3183
rect 12300 3157 12370 3183
rect 12300 3123 12318 3157
rect 12352 3123 12370 3157
rect 12300 3097 12370 3123
rect 12400 3157 12470 3183
rect 12400 3123 12418 3157
rect 12452 3123 12470 3157
rect 12400 3097 12470 3123
rect 12500 3157 12570 3183
rect 12500 3123 12518 3157
rect 12552 3123 12570 3157
rect 12500 3097 12570 3123
rect 12600 3157 12670 3183
rect 12600 3123 12618 3157
rect 12652 3123 12670 3157
rect 12600 3097 12670 3123
rect 12700 3157 12770 3183
rect 12700 3123 12718 3157
rect 12752 3123 12770 3157
rect 12700 3097 12770 3123
rect 12800 3097 12854 3183
rect 12912 3172 12970 3183
rect 12912 3138 12924 3172
rect 12958 3138 12970 3172
rect 12912 3097 12970 3138
rect 13000 3157 13070 3183
rect 13000 3123 13018 3157
rect 13052 3123 13070 3157
rect 13000 3097 13070 3123
rect 13100 3142 13158 3183
rect 13100 3108 13112 3142
rect 13146 3108 13158 3142
rect 13100 3097 13158 3108
rect 13220 3157 13280 3183
rect 13220 3123 13228 3157
rect 13262 3123 13280 3157
rect 13220 3097 13280 3123
rect 13310 3157 13380 3183
rect 13310 3123 13328 3157
rect 13362 3123 13380 3157
rect 13310 3097 13380 3123
rect 13410 3157 13480 3183
rect 13410 3123 13428 3157
rect 13462 3123 13480 3157
rect 13410 3097 13480 3123
rect 13510 3157 13580 3183
rect 13510 3123 13528 3157
rect 13562 3123 13580 3157
rect 13510 3097 13580 3123
rect 13610 3157 13670 3183
rect 13610 3123 13628 3157
rect 13662 3123 13670 3157
rect 13610 3097 13670 3123
rect 11616 3017 11670 3043
rect 11616 2983 11624 3017
rect 11658 2983 11670 3017
rect 11616 2957 11670 2983
rect 11700 3017 11770 3043
rect 11700 2983 11718 3017
rect 11752 2983 11770 3017
rect 11700 2957 11770 2983
rect 11800 3017 11870 3043
rect 11800 2983 11818 3017
rect 11852 2983 11870 3017
rect 11800 2957 11870 2983
rect 11900 3017 11970 3043
rect 11900 2983 11918 3017
rect 11952 2983 11970 3017
rect 11900 2957 11970 2983
rect 12000 3017 12070 3043
rect 12000 2983 12018 3017
rect 12052 2983 12070 3017
rect 12000 2957 12070 2983
rect 12100 2957 12170 3043
rect 12200 3017 12270 3043
rect 12200 2983 12218 3017
rect 12252 2983 12270 3017
rect 12200 2957 12270 2983
rect 12300 3017 12370 3043
rect 12300 2983 12318 3017
rect 12352 2983 12370 3017
rect 12300 2957 12370 2983
rect 12400 2957 12470 3043
rect 12500 2957 12570 3043
rect 12600 2957 12670 3043
rect 12700 3017 12770 3043
rect 12700 2983 12718 3017
rect 12752 2983 12770 3017
rect 12700 2957 12770 2983
rect 12800 3017 12854 3043
rect 12800 2983 12812 3017
rect 12846 2983 12854 3017
rect 12800 2957 12854 2983
rect 12912 3032 12970 3043
rect 12912 2998 12924 3032
rect 12958 2998 12970 3032
rect 12912 2957 12970 2998
rect 13000 3017 13070 3043
rect 13000 2983 13018 3017
rect 13052 2983 13070 3017
rect 13000 2957 13070 2983
rect 13100 3002 13158 3043
rect 13100 2968 13112 3002
rect 13146 2968 13158 3002
rect 13100 2957 13158 2968
rect 13220 3017 13280 3043
rect 13220 2983 13228 3017
rect 13262 2983 13280 3017
rect 13220 2957 13280 2983
rect 13310 3017 13380 3043
rect 13310 2983 13328 3017
rect 13362 2983 13380 3017
rect 13310 2957 13380 2983
rect 13410 3017 13480 3043
rect 13410 2983 13428 3017
rect 13462 2983 13480 3017
rect 13410 2957 13480 2983
rect 13510 3017 13580 3043
rect 13510 2983 13528 3017
rect 13562 2983 13580 3017
rect 13510 2957 13580 2983
rect 13610 3017 13670 3043
rect 13610 2983 13628 3017
rect 13662 2983 13670 3017
rect 13610 2957 13670 2983
rect 11416 2877 11470 2903
rect 11416 2843 11424 2877
rect 11458 2843 11470 2877
rect 11416 2817 11470 2843
rect 11500 2877 11570 2903
rect 11500 2843 11518 2877
rect 11552 2843 11570 2877
rect 11500 2817 11570 2843
rect 11600 2877 11670 2903
rect 11600 2843 11618 2877
rect 11652 2843 11670 2877
rect 11600 2817 11670 2843
rect 11700 2877 11770 2903
rect 11700 2843 11718 2877
rect 11752 2843 11770 2877
rect 11700 2817 11770 2843
rect 11800 2877 11854 2903
rect 11800 2843 11812 2877
rect 11846 2843 11854 2877
rect 11800 2817 11854 2843
rect 10716 2737 10770 2763
rect 10716 2703 10724 2737
rect 10758 2703 10770 2737
rect 10716 2677 10770 2703
rect 10800 2737 10870 2763
rect 10800 2703 10818 2737
rect 10852 2703 10870 2737
rect 10800 2677 10870 2703
rect 10900 2737 10970 2763
rect 10900 2703 10918 2737
rect 10952 2703 10970 2737
rect 10900 2677 10970 2703
rect 11000 2677 11070 2763
rect 11100 2677 11170 2763
rect 11200 2677 11270 2763
rect 11300 2677 11370 2763
rect 11400 2677 11470 2763
rect 11500 2737 11570 2763
rect 11500 2703 11518 2737
rect 11552 2703 11570 2737
rect 11500 2677 11570 2703
rect 11600 2737 11654 2763
rect 11600 2703 11612 2737
rect 11646 2703 11654 2737
rect 11600 2677 11654 2703
rect 10016 2597 10070 2623
rect 10016 2563 10024 2597
rect 10058 2563 10070 2597
rect 10016 2537 10070 2563
rect 10100 2597 10170 2623
rect 10100 2563 10118 2597
rect 10152 2563 10170 2597
rect 10100 2537 10170 2563
rect 10200 2597 10270 2623
rect 10200 2563 10218 2597
rect 10252 2563 10270 2597
rect 10200 2537 10270 2563
rect 10300 2537 10370 2623
rect 10400 2537 10470 2623
rect 10500 2537 10570 2623
rect 10600 2597 10670 2623
rect 10600 2563 10618 2597
rect 10652 2563 10670 2597
rect 10600 2537 10670 2563
rect 10700 2597 10770 2623
rect 10700 2563 10718 2597
rect 10752 2563 10770 2597
rect 10700 2537 10770 2563
rect 10800 2597 10870 2623
rect 10800 2563 10818 2597
rect 10852 2563 10870 2597
rect 10800 2537 10870 2563
rect 10900 2597 10954 2623
rect 10900 2563 10912 2597
rect 10946 2563 10954 2597
rect 10900 2537 10954 2563
rect 11016 2597 11070 2623
rect 11016 2563 11024 2597
rect 11058 2563 11070 2597
rect 11016 2537 11070 2563
rect 11100 2597 11154 2623
rect 11100 2563 11112 2597
rect 11146 2563 11154 2597
rect 11100 2537 11154 2563
rect 11216 2597 11270 2623
rect 11216 2563 11224 2597
rect 11258 2563 11270 2597
rect 11216 2537 11270 2563
rect 11300 2597 11354 2623
rect 11300 2563 11312 2597
rect 11346 2563 11354 2597
rect 11300 2537 11354 2563
rect 11416 2597 11470 2623
rect 11416 2563 11424 2597
rect 11458 2563 11470 2597
rect 11416 2537 11470 2563
rect 11500 2597 11570 2623
rect 11500 2563 11518 2597
rect 11552 2563 11570 2597
rect 11500 2537 11570 2563
rect 11600 2597 11654 2623
rect 11600 2563 11612 2597
rect 11646 2563 11654 2597
rect 11600 2537 11654 2563
rect 11916 2877 11970 2903
rect 11916 2843 11924 2877
rect 11958 2843 11970 2877
rect 11916 2817 11970 2843
rect 12000 2877 12070 2903
rect 12000 2843 12018 2877
rect 12052 2843 12070 2877
rect 12000 2817 12070 2843
rect 12100 2817 12170 2903
rect 12200 2817 12270 2903
rect 12300 2817 12370 2903
rect 12400 2817 12470 2903
rect 12500 2817 12570 2903
rect 12600 2817 12670 2903
rect 12700 2877 12770 2903
rect 12700 2843 12718 2877
rect 12752 2843 12770 2877
rect 12700 2817 12770 2843
rect 12800 2877 12854 2903
rect 12800 2843 12812 2877
rect 12846 2843 12854 2877
rect 12800 2817 12854 2843
rect 12912 2892 12970 2903
rect 12912 2858 12924 2892
rect 12958 2858 12970 2892
rect 12912 2817 12970 2858
rect 13000 2877 13070 2903
rect 13000 2843 13018 2877
rect 13052 2843 13070 2877
rect 13000 2817 13070 2843
rect 13100 2862 13158 2903
rect 13100 2828 13112 2862
rect 13146 2828 13158 2862
rect 13100 2817 13158 2828
rect 13220 2877 13280 2903
rect 13220 2843 13228 2877
rect 13262 2843 13280 2877
rect 13220 2817 13280 2843
rect 13310 2877 13380 2903
rect 13310 2843 13328 2877
rect 13362 2843 13380 2877
rect 13310 2817 13380 2843
rect 13410 2877 13480 2903
rect 13410 2843 13428 2877
rect 13462 2843 13480 2877
rect 13410 2817 13480 2843
rect 13510 2877 13580 2903
rect 13510 2843 13528 2877
rect 13562 2843 13580 2877
rect 13510 2817 13580 2843
rect 13610 2877 13670 2903
rect 13610 2843 13628 2877
rect 13662 2843 13670 2877
rect 13610 2817 13670 2843
rect 11716 2737 11770 2763
rect 11716 2703 11724 2737
rect 11758 2703 11770 2737
rect 11716 2677 11770 2703
rect 11800 2737 11870 2763
rect 11800 2703 11818 2737
rect 11852 2703 11870 2737
rect 11800 2677 11870 2703
rect 11900 2737 11970 2763
rect 11900 2703 11918 2737
rect 11952 2703 11970 2737
rect 11900 2677 11970 2703
rect 12000 2677 12070 2763
rect 12100 2677 12170 2763
rect 12200 2737 12270 2763
rect 12200 2703 12218 2737
rect 12252 2703 12270 2737
rect 12200 2677 12270 2703
rect 12300 2737 12370 2763
rect 12300 2703 12318 2737
rect 12352 2703 12370 2737
rect 12300 2677 12370 2703
rect 12400 2737 12470 2763
rect 12400 2703 12418 2737
rect 12452 2703 12470 2737
rect 12400 2677 12470 2703
rect 12500 2737 12570 2763
rect 12500 2703 12518 2737
rect 12552 2703 12570 2737
rect 12500 2677 12570 2703
rect 12600 2737 12670 2763
rect 12600 2703 12618 2737
rect 12652 2703 12670 2737
rect 12600 2677 12670 2703
rect 12700 2737 12770 2763
rect 12700 2703 12718 2737
rect 12752 2703 12770 2737
rect 12700 2677 12770 2703
rect 12800 2677 12854 2763
rect 12912 2752 12970 2763
rect 12912 2718 12924 2752
rect 12958 2718 12970 2752
rect 12912 2677 12970 2718
rect 13000 2737 13070 2763
rect 13000 2703 13018 2737
rect 13052 2703 13070 2737
rect 13000 2677 13070 2703
rect 13100 2722 13158 2763
rect 13100 2688 13112 2722
rect 13146 2688 13158 2722
rect 13100 2677 13158 2688
rect 13220 2737 13280 2763
rect 13220 2703 13228 2737
rect 13262 2703 13280 2737
rect 13220 2677 13280 2703
rect 13310 2737 13380 2763
rect 13310 2703 13328 2737
rect 13362 2703 13380 2737
rect 13310 2677 13380 2703
rect 13410 2737 13480 2763
rect 13410 2703 13428 2737
rect 13462 2703 13480 2737
rect 13410 2677 13480 2703
rect 13510 2737 13580 2763
rect 13510 2703 13528 2737
rect 13562 2703 13580 2737
rect 13510 2677 13580 2703
rect 13610 2737 13670 2763
rect 13610 2703 13628 2737
rect 13662 2703 13670 2737
rect 13610 2677 13670 2703
rect 11716 2597 11770 2623
rect 11716 2563 11724 2597
rect 11758 2563 11770 2597
rect 11716 2537 11770 2563
rect 11800 2597 11870 2623
rect 11800 2563 11818 2597
rect 11852 2563 11870 2597
rect 11800 2537 11870 2563
rect 11900 2537 11970 2623
rect 12000 2537 12070 2623
rect 12100 2537 12170 2623
rect 12200 2597 12270 2623
rect 12200 2563 12218 2597
rect 12252 2563 12270 2597
rect 12200 2537 12270 2563
rect 12300 2597 12370 2623
rect 12300 2563 12318 2597
rect 12352 2563 12370 2597
rect 12300 2537 12370 2563
rect 12400 2597 12470 2623
rect 12400 2563 12418 2597
rect 12452 2563 12470 2597
rect 12400 2537 12470 2563
rect 12500 2537 12570 2623
rect 12600 2597 12670 2623
rect 12600 2563 12618 2597
rect 12652 2563 12670 2597
rect 12600 2537 12670 2563
rect 12700 2597 12770 2623
rect 12700 2563 12718 2597
rect 12752 2563 12770 2597
rect 12700 2537 12770 2563
rect 12800 2537 12854 2623
rect 12912 2612 12970 2623
rect 12912 2578 12924 2612
rect 12958 2578 12970 2612
rect 12912 2537 12970 2578
rect 13000 2597 13070 2623
rect 13000 2563 13018 2597
rect 13052 2563 13070 2597
rect 13000 2537 13070 2563
rect 13100 2582 13158 2623
rect 13100 2548 13112 2582
rect 13146 2548 13158 2582
rect 13100 2537 13158 2548
rect 13220 2597 13280 2623
rect 13220 2563 13228 2597
rect 13262 2563 13280 2597
rect 13220 2537 13280 2563
rect 13310 2597 13380 2623
rect 13310 2563 13328 2597
rect 13362 2563 13380 2597
rect 13310 2537 13380 2563
rect 13410 2597 13480 2623
rect 13410 2563 13428 2597
rect 13462 2563 13480 2597
rect 13410 2537 13480 2563
rect 13510 2597 13580 2623
rect 13510 2563 13528 2597
rect 13562 2563 13580 2597
rect 13510 2537 13580 2563
rect 13610 2597 13670 2623
rect 13610 2563 13628 2597
rect 13662 2563 13670 2597
rect 13610 2537 13670 2563
rect 9716 2367 9770 2393
rect 9716 2333 9724 2367
rect 9758 2333 9770 2367
rect 9716 2307 9770 2333
rect 9800 2367 9870 2393
rect 9800 2333 9818 2367
rect 9852 2333 9870 2367
rect 9800 2307 9870 2333
rect 9900 2307 9970 2393
rect 10000 2367 10070 2393
rect 10000 2333 10018 2367
rect 10052 2333 10070 2367
rect 10000 2307 10070 2333
rect 10100 2367 10170 2393
rect 10100 2333 10118 2367
rect 10152 2333 10170 2367
rect 10100 2307 10170 2333
rect 10200 2307 10270 2393
rect 10300 2367 10370 2393
rect 10300 2333 10318 2367
rect 10352 2333 10370 2367
rect 10300 2307 10370 2333
rect 10400 2367 10470 2393
rect 10400 2333 10418 2367
rect 10452 2333 10470 2367
rect 10400 2307 10470 2333
rect 10500 2367 10570 2393
rect 10500 2333 10518 2367
rect 10552 2333 10570 2367
rect 10500 2307 10570 2333
rect 10600 2367 10670 2393
rect 10600 2333 10618 2367
rect 10652 2333 10670 2367
rect 10600 2307 10670 2333
rect 10700 2367 10770 2393
rect 10700 2333 10718 2367
rect 10752 2333 10770 2367
rect 10700 2307 10770 2333
rect 10800 2367 10870 2393
rect 10800 2333 10818 2367
rect 10852 2333 10870 2367
rect 10800 2307 10870 2333
rect 10900 2367 10970 2393
rect 10900 2333 10918 2367
rect 10952 2333 10970 2367
rect 10900 2307 10970 2333
rect 11000 2307 11070 2393
rect 11100 2367 11170 2393
rect 11100 2333 11118 2367
rect 11152 2333 11170 2367
rect 11100 2307 11170 2333
rect 11200 2367 11270 2393
rect 11200 2333 11218 2367
rect 11252 2333 11270 2367
rect 11200 2307 11270 2333
rect 11300 2367 11370 2393
rect 11300 2333 11318 2367
rect 11352 2333 11370 2367
rect 11300 2307 11370 2333
rect 11400 2367 11470 2393
rect 11400 2333 11418 2367
rect 11452 2333 11470 2367
rect 11400 2307 11470 2333
rect 11500 2307 11570 2393
rect 11600 2367 11670 2393
rect 11600 2333 11618 2367
rect 11652 2333 11670 2367
rect 11600 2307 11670 2333
rect 11700 2367 11754 2393
rect 11700 2333 11712 2367
rect 11746 2333 11754 2367
rect 11700 2307 11754 2333
rect 9616 2227 9670 2253
rect 9616 2193 9624 2227
rect 9658 2193 9670 2227
rect 9616 2167 9670 2193
rect 9700 2227 9770 2253
rect 9700 2193 9718 2227
rect 9752 2193 9770 2227
rect 9700 2167 9770 2193
rect 9800 2227 9870 2253
rect 9800 2193 9818 2227
rect 9852 2193 9870 2227
rect 9800 2167 9870 2193
rect 9900 2167 9970 2253
rect 10000 2167 10070 2253
rect 10100 2167 10170 2253
rect 10200 2227 10270 2253
rect 10200 2193 10218 2227
rect 10252 2193 10270 2227
rect 10200 2167 10270 2193
rect 10300 2227 10370 2253
rect 10300 2193 10318 2227
rect 10352 2193 10370 2227
rect 10300 2167 10370 2193
rect 10400 2227 10470 2253
rect 10400 2193 10418 2227
rect 10452 2193 10470 2227
rect 10400 2167 10470 2193
rect 10500 2227 10554 2253
rect 10500 2193 10512 2227
rect 10546 2193 10554 2227
rect 10500 2167 10554 2193
rect 11816 2367 11870 2393
rect 11816 2333 11824 2367
rect 11858 2333 11870 2367
rect 11816 2307 11870 2333
rect 11900 2367 11954 2393
rect 11900 2333 11912 2367
rect 11946 2333 11954 2367
rect 11900 2307 11954 2333
rect 12016 2367 12070 2393
rect 12016 2333 12024 2367
rect 12058 2333 12070 2367
rect 12016 2307 12070 2333
rect 12100 2367 12170 2393
rect 12100 2333 12118 2367
rect 12152 2333 12170 2367
rect 12100 2307 12170 2333
rect 12200 2307 12270 2393
rect 12300 2367 12370 2393
rect 12300 2333 12318 2367
rect 12352 2333 12370 2367
rect 12300 2307 12370 2333
rect 12400 2367 12470 2393
rect 12400 2333 12418 2367
rect 12452 2333 12470 2367
rect 12400 2307 12470 2333
rect 12500 2367 12554 2393
rect 12500 2333 12512 2367
rect 12546 2333 12554 2367
rect 12500 2307 12554 2333
rect 10616 2227 10670 2253
rect 10616 2193 10624 2227
rect 10658 2193 10670 2227
rect 10616 2167 10670 2193
rect 10700 2227 10770 2253
rect 10700 2193 10718 2227
rect 10752 2193 10770 2227
rect 10700 2167 10770 2193
rect 10800 2227 10870 2253
rect 10800 2193 10818 2227
rect 10852 2193 10870 2227
rect 10800 2167 10870 2193
rect 10900 2227 10970 2253
rect 10900 2193 10918 2227
rect 10952 2193 10970 2227
rect 10900 2167 10970 2193
rect 11000 2167 11070 2253
rect 11100 2167 11170 2253
rect 11200 2167 11270 2253
rect 11300 2227 11370 2253
rect 11300 2193 11318 2227
rect 11352 2193 11370 2227
rect 11300 2167 11370 2193
rect 11400 2227 11470 2253
rect 11400 2193 11418 2227
rect 11452 2193 11470 2227
rect 11400 2167 11470 2193
rect 11500 2227 11570 2253
rect 11500 2193 11518 2227
rect 11552 2193 11570 2227
rect 11500 2167 11570 2193
rect 11600 2167 11670 2253
rect 11700 2167 11770 2253
rect 11800 2227 11870 2253
rect 11800 2193 11818 2227
rect 11852 2193 11870 2227
rect 11800 2167 11870 2193
rect 11900 2227 11970 2253
rect 11900 2193 11918 2227
rect 11952 2193 11970 2227
rect 11900 2167 11970 2193
rect 12000 2227 12054 2253
rect 12000 2193 12012 2227
rect 12046 2193 12054 2227
rect 12000 2167 12054 2193
rect 9316 2087 9370 2113
rect 9316 2053 9324 2087
rect 9358 2053 9370 2087
rect 9316 2027 9370 2053
rect 9400 2087 9470 2113
rect 9400 2053 9418 2087
rect 9452 2053 9470 2087
rect 9400 2027 9470 2053
rect 9500 2027 9570 2113
rect 9600 2027 9670 2113
rect 9700 2027 9770 2113
rect 9800 2027 9870 2113
rect 9900 2027 9970 2113
rect 10000 2027 10070 2113
rect 10100 2087 10170 2113
rect 10100 2053 10118 2087
rect 10152 2053 10170 2087
rect 10100 2027 10170 2053
rect 10200 2087 10270 2113
rect 10200 2053 10218 2087
rect 10252 2053 10270 2087
rect 10200 2027 10270 2053
rect 10300 2087 10370 2113
rect 10300 2053 10318 2087
rect 10352 2053 10370 2087
rect 10300 2027 10370 2053
rect 10400 2087 10470 2113
rect 10400 2053 10418 2087
rect 10452 2053 10470 2087
rect 10400 2027 10470 2053
rect 10500 2027 10570 2113
rect 10600 2087 10670 2113
rect 10600 2053 10618 2087
rect 10652 2053 10670 2087
rect 10600 2027 10670 2053
rect 10700 2087 10770 2113
rect 10700 2053 10718 2087
rect 10752 2053 10770 2087
rect 10700 2027 10770 2053
rect 10800 2027 10870 2113
rect 10900 2087 10970 2113
rect 10900 2053 10918 2087
rect 10952 2053 10970 2087
rect 10900 2027 10970 2053
rect 11000 2087 11070 2113
rect 11000 2053 11018 2087
rect 11052 2053 11070 2087
rect 11000 2027 11070 2053
rect 11100 2087 11170 2113
rect 11100 2053 11118 2087
rect 11152 2053 11170 2087
rect 11100 2027 11170 2053
rect 11200 2087 11254 2113
rect 11200 2053 11212 2087
rect 11246 2053 11254 2087
rect 11200 2027 11254 2053
rect 7016 1947 7070 1973
rect 7016 1913 7024 1947
rect 7058 1913 7070 1947
rect 7016 1887 7070 1913
rect 7100 1947 7170 1973
rect 7100 1913 7118 1947
rect 7152 1913 7170 1947
rect 7100 1887 7170 1913
rect 7200 1947 7270 1973
rect 7200 1913 7218 1947
rect 7252 1913 7270 1947
rect 7200 1887 7270 1913
rect 7300 1947 7370 1973
rect 7300 1913 7318 1947
rect 7352 1913 7370 1947
rect 7300 1887 7370 1913
rect 7400 1887 7470 1973
rect 7500 1887 7570 1973
rect 7600 1887 7670 1973
rect 7700 1887 7770 1973
rect 7800 1887 7870 1973
rect 7900 1887 7970 1973
rect 8000 1887 8070 1973
rect 8100 1887 8170 1973
rect 8200 1947 8270 1973
rect 8200 1913 8218 1947
rect 8252 1913 8270 1947
rect 8200 1887 8270 1913
rect 8300 1947 8370 1973
rect 8300 1913 8318 1947
rect 8352 1913 8370 1947
rect 8300 1887 8370 1913
rect 8400 1947 8470 1973
rect 8400 1913 8418 1947
rect 8452 1913 8470 1947
rect 8400 1887 8470 1913
rect 8500 1887 8570 1973
rect 8600 1887 8670 1973
rect 8700 1887 8770 1973
rect 8800 1887 8870 1973
rect 8900 1887 8970 1973
rect 9000 1887 9070 1973
rect 9100 1887 9170 1973
rect 9200 1887 9270 1973
rect 9300 1947 9370 1973
rect 9300 1913 9318 1947
rect 9352 1913 9370 1947
rect 9300 1887 9370 1913
rect 9400 1947 9470 1973
rect 9400 1913 9418 1947
rect 9452 1913 9470 1947
rect 9400 1887 9470 1913
rect 9500 1887 9570 1973
rect 9600 1947 9670 1973
rect 9600 1913 9618 1947
rect 9652 1913 9670 1947
rect 9600 1887 9670 1913
rect 9700 1947 9770 1973
rect 9700 1913 9718 1947
rect 9752 1913 9770 1947
rect 9700 1887 9770 1913
rect 9800 1947 9870 1973
rect 9800 1913 9818 1947
rect 9852 1913 9870 1947
rect 9800 1887 9870 1913
rect 9900 1947 9970 1973
rect 9900 1913 9918 1947
rect 9952 1913 9970 1947
rect 9900 1887 9970 1913
rect 10000 1947 10070 1973
rect 10000 1913 10018 1947
rect 10052 1913 10070 1947
rect 10000 1887 10070 1913
rect 10100 1887 10170 1973
rect 10200 1887 10270 1973
rect 10300 1947 10370 1973
rect 10300 1913 10318 1947
rect 10352 1913 10370 1947
rect 10300 1887 10370 1913
rect 10400 1947 10470 1973
rect 10400 1913 10418 1947
rect 10452 1913 10470 1947
rect 10400 1887 10470 1913
rect 10500 1887 10570 1973
rect 10600 1947 10670 1973
rect 10600 1913 10618 1947
rect 10652 1913 10670 1947
rect 10600 1887 10670 1913
rect 10700 1947 10770 1973
rect 10700 1913 10718 1947
rect 10752 1913 10770 1947
rect 10700 1887 10770 1913
rect 10800 1947 10870 1973
rect 10800 1913 10818 1947
rect 10852 1913 10870 1947
rect 10800 1887 10870 1913
rect 10900 1947 10970 1973
rect 10900 1913 10918 1947
rect 10952 1913 10970 1947
rect 10900 1887 10970 1913
rect 11000 1947 11054 1973
rect 11000 1913 11012 1947
rect 11046 1913 11054 1947
rect 11000 1887 11054 1913
rect 6416 1807 6470 1833
rect 6416 1773 6424 1807
rect 6458 1773 6470 1807
rect 6416 1747 6470 1773
rect 6500 1807 6570 1833
rect 6500 1773 6518 1807
rect 6552 1773 6570 1807
rect 6500 1747 6570 1773
rect 6600 1747 6670 1833
rect 6700 1747 6770 1833
rect 6800 1807 6870 1833
rect 6800 1773 6818 1807
rect 6852 1773 6870 1807
rect 6800 1747 6870 1773
rect 6900 1807 6970 1833
rect 6900 1773 6918 1807
rect 6952 1773 6970 1807
rect 6900 1747 6970 1773
rect 7000 1807 7070 1833
rect 7000 1773 7018 1807
rect 7052 1773 7070 1807
rect 7000 1747 7070 1773
rect 7100 1807 7154 1833
rect 7100 1773 7112 1807
rect 7146 1773 7154 1807
rect 7100 1747 7154 1773
rect 6216 1667 6270 1693
rect 6216 1633 6224 1667
rect 6258 1633 6270 1667
rect 6216 1607 6270 1633
rect 6300 1667 6370 1693
rect 6300 1633 6318 1667
rect 6352 1633 6370 1667
rect 6300 1607 6370 1633
rect 6400 1667 6470 1693
rect 6400 1633 6418 1667
rect 6452 1633 6470 1667
rect 6400 1607 6470 1633
rect 6500 1667 6554 1693
rect 6500 1633 6512 1667
rect 6546 1633 6554 1667
rect 6500 1607 6554 1633
rect 6116 1527 6170 1553
rect 6116 1493 6124 1527
rect 6158 1493 6170 1527
rect 6116 1467 6170 1493
rect 6200 1527 6270 1553
rect 6200 1493 6218 1527
rect 6252 1493 6270 1527
rect 6200 1467 6270 1493
rect 6300 1527 6354 1553
rect 6300 1493 6312 1527
rect 6346 1493 6354 1527
rect 6300 1467 6354 1493
rect 5216 1387 5270 1413
rect 5216 1353 5224 1387
rect 5258 1353 5270 1387
rect 5216 1327 5270 1353
rect 5300 1387 5370 1413
rect 5300 1353 5318 1387
rect 5352 1353 5370 1387
rect 5300 1327 5370 1353
rect 5400 1327 5470 1413
rect 5500 1327 5570 1413
rect 5600 1387 5670 1413
rect 5600 1353 5618 1387
rect 5652 1353 5670 1387
rect 5600 1327 5670 1353
rect 5700 1387 5770 1413
rect 5700 1353 5718 1387
rect 5752 1353 5770 1387
rect 5700 1327 5770 1353
rect 5800 1387 5870 1413
rect 5800 1353 5818 1387
rect 5852 1353 5870 1387
rect 5800 1327 5870 1353
rect 5900 1327 5970 1413
rect 6000 1387 6070 1413
rect 6000 1353 6018 1387
rect 6052 1353 6070 1387
rect 6000 1327 6070 1353
rect 6100 1387 6170 1413
rect 6100 1353 6118 1387
rect 6152 1353 6170 1387
rect 6100 1327 6170 1353
rect 6200 1387 6254 1413
rect 6200 1353 6212 1387
rect 6246 1353 6254 1387
rect 6200 1327 6254 1353
rect 4716 1157 4770 1183
rect 4716 1123 4724 1157
rect 4758 1123 4770 1157
rect 4716 1097 4770 1123
rect 4800 1157 4870 1183
rect 4800 1123 4818 1157
rect 4852 1123 4870 1157
rect 4800 1097 4870 1123
rect 4900 1097 4970 1183
rect 5000 1097 5070 1183
rect 5100 1157 5170 1183
rect 5100 1123 5118 1157
rect 5152 1123 5170 1157
rect 5100 1097 5170 1123
rect 5200 1157 5270 1183
rect 5200 1123 5218 1157
rect 5252 1123 5270 1157
rect 5200 1097 5270 1123
rect 5300 1157 5370 1183
rect 5300 1123 5318 1157
rect 5352 1123 5370 1157
rect 5300 1097 5370 1123
rect 5400 1157 5454 1183
rect 5400 1123 5412 1157
rect 5446 1123 5454 1157
rect 5400 1097 5454 1123
rect 3916 1017 3970 1043
rect 3916 983 3924 1017
rect 3958 983 3970 1017
rect 3916 957 3970 983
rect 4000 1017 4070 1043
rect 4000 983 4018 1017
rect 4052 983 4070 1017
rect 4000 957 4070 983
rect 4100 1017 4170 1043
rect 4100 983 4118 1017
rect 4152 983 4170 1017
rect 4100 957 4170 983
rect 4200 1017 4270 1043
rect 4200 983 4218 1017
rect 4252 983 4270 1017
rect 4200 957 4270 983
rect 4300 1017 4370 1043
rect 4300 983 4318 1017
rect 4352 983 4370 1017
rect 4300 957 4370 983
rect 4400 1017 4470 1043
rect 4400 983 4418 1017
rect 4452 983 4470 1017
rect 4400 957 4470 983
rect 4500 957 4570 1043
rect 4600 957 4670 1043
rect 4700 1017 4770 1043
rect 4700 983 4718 1017
rect 4752 983 4770 1017
rect 4700 957 4770 983
rect 4800 1017 4854 1043
rect 4800 983 4812 1017
rect 4846 983 4854 1017
rect 4800 957 4854 983
rect 4916 1017 4970 1043
rect 4916 983 4924 1017
rect 4958 983 4970 1017
rect 4916 957 4970 983
rect 5000 1017 5070 1043
rect 5000 983 5018 1017
rect 5052 983 5070 1017
rect 5000 957 5070 983
rect 5100 957 5170 1043
rect 5200 1017 5270 1043
rect 5200 983 5218 1017
rect 5252 983 5270 1017
rect 5200 957 5270 983
rect 5300 1017 5354 1043
rect 5300 983 5312 1017
rect 5346 983 5354 1017
rect 5300 957 5354 983
rect 7216 1807 7270 1833
rect 7216 1773 7224 1807
rect 7258 1773 7270 1807
rect 7216 1747 7270 1773
rect 7300 1807 7370 1833
rect 7300 1773 7318 1807
rect 7352 1773 7370 1807
rect 7300 1747 7370 1773
rect 7400 1807 7454 1833
rect 7400 1773 7412 1807
rect 7446 1773 7454 1807
rect 7400 1747 7454 1773
rect 7516 1807 7570 1833
rect 7516 1773 7524 1807
rect 7558 1773 7570 1807
rect 7516 1747 7570 1773
rect 7600 1807 7670 1833
rect 7600 1773 7618 1807
rect 7652 1773 7670 1807
rect 7600 1747 7670 1773
rect 7700 1807 7754 1833
rect 7700 1773 7712 1807
rect 7746 1773 7754 1807
rect 7700 1747 7754 1773
rect 7816 1807 7870 1833
rect 7816 1773 7824 1807
rect 7858 1773 7870 1807
rect 7816 1747 7870 1773
rect 7900 1807 7970 1833
rect 7900 1773 7918 1807
rect 7952 1773 7970 1807
rect 7900 1747 7970 1773
rect 8000 1807 8054 1833
rect 8000 1773 8012 1807
rect 8046 1773 8054 1807
rect 8000 1747 8054 1773
rect 8116 1807 8170 1833
rect 8116 1773 8124 1807
rect 8158 1773 8170 1807
rect 8116 1747 8170 1773
rect 8200 1807 8270 1833
rect 8200 1773 8218 1807
rect 8252 1773 8270 1807
rect 8200 1747 8270 1773
rect 8300 1807 8370 1833
rect 8300 1773 8318 1807
rect 8352 1773 8370 1807
rect 8300 1747 8370 1773
rect 8400 1807 8470 1833
rect 8400 1773 8418 1807
rect 8452 1773 8470 1807
rect 8400 1747 8470 1773
rect 8500 1807 8570 1833
rect 8500 1773 8518 1807
rect 8552 1773 8570 1807
rect 8500 1747 8570 1773
rect 8600 1807 8654 1833
rect 8600 1773 8612 1807
rect 8646 1773 8654 1807
rect 8600 1747 8654 1773
rect 8716 1807 8770 1833
rect 8716 1773 8724 1807
rect 8758 1773 8770 1807
rect 8716 1747 8770 1773
rect 8800 1807 8870 1833
rect 8800 1773 8818 1807
rect 8852 1773 8870 1807
rect 8800 1747 8870 1773
rect 8900 1807 8970 1833
rect 8900 1773 8918 1807
rect 8952 1773 8970 1807
rect 8900 1747 8970 1773
rect 9000 1747 9070 1833
rect 9100 1747 9170 1833
rect 9200 1747 9270 1833
rect 9300 1807 9370 1833
rect 9300 1773 9318 1807
rect 9352 1773 9370 1807
rect 9300 1747 9370 1773
rect 9400 1807 9470 1833
rect 9400 1773 9418 1807
rect 9452 1773 9470 1807
rect 9400 1747 9470 1773
rect 9500 1807 9570 1833
rect 9500 1773 9518 1807
rect 9552 1773 9570 1807
rect 9500 1747 9570 1773
rect 9600 1747 9670 1833
rect 9700 1807 9770 1833
rect 9700 1773 9718 1807
rect 9752 1773 9770 1807
rect 9700 1747 9770 1773
rect 9800 1807 9854 1833
rect 9800 1773 9812 1807
rect 9846 1773 9854 1807
rect 9800 1747 9854 1773
rect 6616 1667 6670 1693
rect 6616 1633 6624 1667
rect 6658 1633 6670 1667
rect 6616 1607 6670 1633
rect 6700 1667 6770 1693
rect 6700 1633 6718 1667
rect 6752 1633 6770 1667
rect 6700 1607 6770 1633
rect 6800 1667 6870 1693
rect 6800 1633 6818 1667
rect 6852 1633 6870 1667
rect 6800 1607 6870 1633
rect 6900 1607 6970 1693
rect 7000 1667 7070 1693
rect 7000 1633 7018 1667
rect 7052 1633 7070 1667
rect 7000 1607 7070 1633
rect 7100 1667 7170 1693
rect 7100 1633 7118 1667
rect 7152 1633 7170 1667
rect 7100 1607 7170 1633
rect 7200 1607 7270 1693
rect 7300 1607 7370 1693
rect 7400 1607 7470 1693
rect 7500 1607 7570 1693
rect 7600 1667 7670 1693
rect 7600 1633 7618 1667
rect 7652 1633 7670 1667
rect 7600 1607 7670 1633
rect 7700 1667 7770 1693
rect 7700 1633 7718 1667
rect 7752 1633 7770 1667
rect 7700 1607 7770 1633
rect 7800 1607 7870 1693
rect 7900 1667 7970 1693
rect 7900 1633 7918 1667
rect 7952 1633 7970 1667
rect 7900 1607 7970 1633
rect 8000 1667 8070 1693
rect 8000 1633 8018 1667
rect 8052 1633 8070 1667
rect 8000 1607 8070 1633
rect 8100 1607 8170 1693
rect 8200 1667 8270 1693
rect 8200 1633 8218 1667
rect 8252 1633 8270 1667
rect 8200 1607 8270 1633
rect 8300 1667 8370 1693
rect 8300 1633 8318 1667
rect 8352 1633 8370 1667
rect 8300 1607 8370 1633
rect 8400 1667 8470 1693
rect 8400 1633 8418 1667
rect 8452 1633 8470 1667
rect 8400 1607 8470 1633
rect 8500 1607 8570 1693
rect 8600 1607 8670 1693
rect 8700 1607 8770 1693
rect 8800 1667 8870 1693
rect 8800 1633 8818 1667
rect 8852 1633 8870 1667
rect 8800 1607 8870 1633
rect 8900 1667 8970 1693
rect 8900 1633 8918 1667
rect 8952 1633 8970 1667
rect 8900 1607 8970 1633
rect 9000 1667 9070 1693
rect 9000 1633 9018 1667
rect 9052 1633 9070 1667
rect 9000 1607 9070 1633
rect 9100 1607 9170 1693
rect 9200 1607 9270 1693
rect 9300 1607 9370 1693
rect 9400 1667 9470 1693
rect 9400 1633 9418 1667
rect 9452 1633 9470 1667
rect 9400 1607 9470 1633
rect 9500 1667 9554 1693
rect 9500 1633 9512 1667
rect 9546 1633 9554 1667
rect 9500 1607 9554 1633
rect 6416 1527 6470 1553
rect 6416 1493 6424 1527
rect 6458 1493 6470 1527
rect 6416 1467 6470 1493
rect 6500 1527 6570 1553
rect 6500 1493 6518 1527
rect 6552 1493 6570 1527
rect 6500 1467 6570 1493
rect 6600 1527 6670 1553
rect 6600 1493 6618 1527
rect 6652 1493 6670 1527
rect 6600 1467 6670 1493
rect 6700 1467 6770 1553
rect 6800 1467 6870 1553
rect 6900 1467 6970 1553
rect 7000 1467 7070 1553
rect 7100 1467 7170 1553
rect 7200 1467 7270 1553
rect 7300 1467 7370 1553
rect 7400 1527 7470 1553
rect 7400 1493 7418 1527
rect 7452 1493 7470 1527
rect 7400 1467 7470 1493
rect 7500 1527 7570 1553
rect 7500 1493 7518 1527
rect 7552 1493 7570 1527
rect 7500 1467 7570 1493
rect 7600 1527 7670 1553
rect 7600 1493 7618 1527
rect 7652 1493 7670 1527
rect 7600 1467 7670 1493
rect 7700 1527 7754 1553
rect 7700 1493 7712 1527
rect 7746 1493 7754 1527
rect 7700 1467 7754 1493
rect 6316 1387 6370 1413
rect 6316 1353 6324 1387
rect 6358 1353 6370 1387
rect 6316 1327 6370 1353
rect 6400 1387 6454 1413
rect 6400 1353 6412 1387
rect 6446 1353 6454 1387
rect 6400 1327 6454 1353
rect 6516 1387 6570 1413
rect 6516 1353 6524 1387
rect 6558 1353 6570 1387
rect 6516 1327 6570 1353
rect 6600 1387 6670 1413
rect 6600 1353 6618 1387
rect 6652 1353 6670 1387
rect 6600 1327 6670 1353
rect 6700 1387 6754 1413
rect 6700 1353 6712 1387
rect 6746 1353 6754 1387
rect 6700 1327 6754 1353
rect 6816 1387 6870 1413
rect 6816 1353 6824 1387
rect 6858 1353 6870 1387
rect 6816 1327 6870 1353
rect 6900 1387 6954 1413
rect 6900 1353 6912 1387
rect 6946 1353 6954 1387
rect 6900 1327 6954 1353
rect 5516 1157 5570 1183
rect 5516 1123 5524 1157
rect 5558 1123 5570 1157
rect 5516 1097 5570 1123
rect 5600 1157 5670 1183
rect 5600 1123 5618 1157
rect 5652 1123 5670 1157
rect 5600 1097 5670 1123
rect 5700 1157 5770 1183
rect 5700 1123 5718 1157
rect 5752 1123 5770 1157
rect 5700 1097 5770 1123
rect 5800 1157 5870 1183
rect 5800 1123 5818 1157
rect 5852 1123 5870 1157
rect 5800 1097 5870 1123
rect 5900 1097 5970 1183
rect 6000 1097 6070 1183
rect 6100 1097 6170 1183
rect 6200 1097 6270 1183
rect 6300 1097 6370 1183
rect 6400 1097 6470 1183
rect 6500 1157 6570 1183
rect 6500 1123 6518 1157
rect 6552 1123 6570 1157
rect 6500 1097 6570 1123
rect 6600 1157 6670 1183
rect 6600 1123 6618 1157
rect 6652 1123 6670 1157
rect 6600 1097 6670 1123
rect 6700 1157 6754 1183
rect 6700 1123 6712 1157
rect 6746 1123 6754 1157
rect 6700 1097 6754 1123
rect 5416 1017 5470 1043
rect 5416 983 5424 1017
rect 5458 983 5470 1017
rect 5416 957 5470 983
rect 5500 1017 5570 1043
rect 5500 983 5518 1017
rect 5552 983 5570 1017
rect 5500 957 5570 983
rect 5600 1017 5670 1043
rect 5600 983 5618 1017
rect 5652 983 5670 1017
rect 5600 957 5670 983
rect 5700 1017 5770 1043
rect 5700 983 5718 1017
rect 5752 983 5770 1017
rect 5700 957 5770 983
rect 5800 1017 5870 1043
rect 5800 983 5818 1017
rect 5852 983 5870 1017
rect 5800 957 5870 983
rect 5900 1017 5970 1043
rect 5900 983 5918 1017
rect 5952 983 5970 1017
rect 5900 957 5970 983
rect 6000 957 6070 1043
rect 6100 1017 6170 1043
rect 6100 983 6118 1017
rect 6152 983 6170 1017
rect 6100 957 6170 983
rect 6200 1017 6270 1043
rect 6200 983 6218 1017
rect 6252 983 6270 1017
rect 6200 957 6270 983
rect 6300 1017 6370 1043
rect 6300 983 6318 1017
rect 6352 983 6370 1017
rect 6300 957 6370 983
rect 6400 1017 6454 1043
rect 6400 983 6412 1017
rect 6446 983 6454 1017
rect 6400 957 6454 983
rect 7816 1527 7870 1553
rect 7816 1493 7824 1527
rect 7858 1493 7870 1527
rect 7816 1467 7870 1493
rect 7900 1527 7954 1553
rect 7900 1493 7912 1527
rect 7946 1493 7954 1527
rect 7900 1467 7954 1493
rect 7016 1387 7070 1413
rect 7016 1353 7024 1387
rect 7058 1353 7070 1387
rect 7016 1327 7070 1353
rect 7100 1387 7170 1413
rect 7100 1353 7118 1387
rect 7152 1353 7170 1387
rect 7100 1327 7170 1353
rect 7200 1387 7270 1413
rect 7200 1353 7218 1387
rect 7252 1353 7270 1387
rect 7200 1327 7270 1353
rect 7300 1387 7370 1413
rect 7300 1353 7318 1387
rect 7352 1353 7370 1387
rect 7300 1327 7370 1353
rect 7400 1387 7470 1413
rect 7400 1353 7418 1387
rect 7452 1353 7470 1387
rect 7400 1327 7470 1353
rect 7500 1387 7570 1413
rect 7500 1353 7518 1387
rect 7552 1353 7570 1387
rect 7500 1327 7570 1353
rect 7600 1327 7670 1413
rect 7700 1327 7770 1413
rect 7800 1387 7870 1413
rect 7800 1353 7818 1387
rect 7852 1353 7870 1387
rect 7800 1327 7870 1353
rect 7900 1387 7954 1413
rect 7900 1353 7912 1387
rect 7946 1353 7954 1387
rect 7900 1327 7954 1353
rect 8016 1527 8070 1553
rect 8016 1493 8024 1527
rect 8058 1493 8070 1527
rect 8016 1467 8070 1493
rect 8100 1527 8170 1553
rect 8100 1493 8118 1527
rect 8152 1493 8170 1527
rect 8100 1467 8170 1493
rect 8200 1467 8270 1553
rect 8300 1467 8370 1553
rect 8400 1527 8470 1553
rect 8400 1493 8418 1527
rect 8452 1493 8470 1527
rect 8400 1467 8470 1493
rect 8500 1527 8554 1553
rect 8500 1493 8512 1527
rect 8546 1493 8554 1527
rect 8500 1467 8554 1493
rect 8616 1527 8670 1553
rect 8616 1493 8624 1527
rect 8658 1493 8670 1527
rect 8616 1467 8670 1493
rect 8700 1527 8770 1553
rect 8700 1493 8718 1527
rect 8752 1493 8770 1527
rect 8700 1467 8770 1493
rect 8800 1467 8870 1553
rect 8900 1527 8970 1553
rect 8900 1493 8918 1527
rect 8952 1493 8970 1527
rect 8900 1467 8970 1493
rect 9000 1527 9070 1553
rect 9000 1493 9018 1527
rect 9052 1493 9070 1527
rect 9000 1467 9070 1493
rect 9100 1527 9170 1553
rect 9100 1493 9118 1527
rect 9152 1493 9170 1527
rect 9100 1467 9170 1493
rect 9200 1527 9270 1553
rect 9200 1493 9218 1527
rect 9252 1493 9270 1527
rect 9200 1467 9270 1493
rect 9300 1527 9354 1553
rect 9300 1493 9312 1527
rect 9346 1493 9354 1527
rect 9300 1467 9354 1493
rect 8016 1387 8070 1413
rect 8016 1353 8024 1387
rect 8058 1353 8070 1387
rect 8016 1327 8070 1353
rect 8100 1387 8170 1413
rect 8100 1353 8118 1387
rect 8152 1353 8170 1387
rect 8100 1327 8170 1353
rect 8200 1387 8270 1413
rect 8200 1353 8218 1387
rect 8252 1353 8270 1387
rect 8200 1327 8270 1353
rect 8300 1387 8370 1413
rect 8300 1353 8318 1387
rect 8352 1353 8370 1387
rect 8300 1327 8370 1353
rect 8400 1327 8470 1413
rect 8500 1327 8570 1413
rect 8600 1327 8670 1413
rect 8700 1387 8770 1413
rect 8700 1353 8718 1387
rect 8752 1353 8770 1387
rect 8700 1327 8770 1353
rect 8800 1387 8870 1413
rect 8800 1353 8818 1387
rect 8852 1353 8870 1387
rect 8800 1327 8870 1353
rect 8900 1387 8970 1413
rect 8900 1353 8918 1387
rect 8952 1353 8970 1387
rect 8900 1327 8970 1353
rect 9000 1327 9070 1413
rect 9100 1387 9170 1413
rect 9100 1353 9118 1387
rect 9152 1353 9170 1387
rect 9100 1327 9170 1353
rect 9200 1387 9270 1413
rect 9200 1353 9218 1387
rect 9252 1353 9270 1387
rect 9200 1327 9270 1353
rect 9300 1387 9354 1413
rect 9300 1353 9312 1387
rect 9346 1353 9354 1387
rect 9300 1327 9354 1353
rect 9916 1807 9970 1833
rect 9916 1773 9924 1807
rect 9958 1773 9970 1807
rect 9916 1747 9970 1773
rect 10000 1807 10054 1833
rect 10000 1773 10012 1807
rect 10046 1773 10054 1807
rect 10000 1747 10054 1773
rect 10116 1807 10170 1833
rect 10116 1773 10124 1807
rect 10158 1773 10170 1807
rect 10116 1747 10170 1773
rect 10200 1807 10254 1833
rect 10200 1773 10212 1807
rect 10246 1773 10254 1807
rect 10200 1747 10254 1773
rect 10316 1807 10370 1833
rect 10316 1773 10324 1807
rect 10358 1773 10370 1807
rect 10316 1747 10370 1773
rect 10400 1807 10454 1833
rect 10400 1773 10412 1807
rect 10446 1773 10454 1807
rect 10400 1747 10454 1773
rect 10516 1807 10570 1833
rect 10516 1773 10524 1807
rect 10558 1773 10570 1807
rect 10516 1747 10570 1773
rect 10600 1807 10670 1833
rect 10600 1773 10618 1807
rect 10652 1773 10670 1807
rect 10600 1747 10670 1773
rect 10700 1807 10754 1833
rect 10700 1773 10712 1807
rect 10746 1773 10754 1807
rect 10700 1747 10754 1773
rect 11116 1947 11170 1973
rect 11116 1913 11124 1947
rect 11158 1913 11170 1947
rect 11116 1887 11170 1913
rect 11200 1947 11254 1973
rect 11200 1913 11212 1947
rect 11246 1913 11254 1947
rect 11200 1887 11254 1913
rect 11316 2087 11370 2113
rect 11316 2053 11324 2087
rect 11358 2053 11370 2087
rect 11316 2027 11370 2053
rect 11400 2087 11454 2113
rect 11400 2053 11412 2087
rect 11446 2053 11454 2087
rect 11400 2027 11454 2053
rect 12116 2227 12170 2253
rect 12116 2193 12124 2227
rect 12158 2193 12170 2227
rect 12116 2167 12170 2193
rect 12200 2227 12270 2253
rect 12200 2193 12218 2227
rect 12252 2193 12270 2227
rect 12200 2167 12270 2193
rect 12300 2227 12354 2253
rect 12300 2193 12312 2227
rect 12346 2193 12354 2227
rect 12300 2167 12354 2193
rect 12616 2367 12670 2393
rect 12616 2333 12624 2367
rect 12658 2333 12670 2367
rect 12616 2307 12670 2333
rect 12700 2367 12770 2393
rect 12700 2333 12718 2367
rect 12752 2333 12770 2367
rect 12700 2307 12770 2333
rect 12800 2307 12854 2393
rect 12912 2382 12970 2393
rect 12912 2348 12924 2382
rect 12958 2348 12970 2382
rect 12912 2307 12970 2348
rect 13000 2367 13070 2393
rect 13000 2333 13018 2367
rect 13052 2333 13070 2367
rect 13000 2307 13070 2333
rect 13100 2352 13158 2393
rect 13100 2318 13112 2352
rect 13146 2318 13158 2352
rect 13100 2307 13158 2318
rect 13220 2367 13280 2393
rect 13220 2333 13228 2367
rect 13262 2333 13280 2367
rect 13220 2307 13280 2333
rect 13310 2367 13380 2393
rect 13310 2333 13328 2367
rect 13362 2333 13380 2367
rect 13310 2307 13380 2333
rect 13410 2367 13480 2393
rect 13410 2333 13428 2367
rect 13462 2333 13480 2367
rect 13410 2307 13480 2333
rect 13510 2367 13580 2393
rect 13510 2333 13528 2367
rect 13562 2333 13580 2367
rect 13510 2307 13580 2333
rect 13610 2367 13670 2393
rect 13610 2333 13628 2367
rect 13662 2333 13670 2367
rect 13610 2307 13670 2333
rect 12416 2227 12470 2253
rect 12416 2193 12424 2227
rect 12458 2193 12470 2227
rect 12416 2167 12470 2193
rect 12500 2227 12570 2253
rect 12500 2193 12518 2227
rect 12552 2193 12570 2227
rect 12500 2167 12570 2193
rect 12600 2227 12654 2253
rect 12600 2193 12612 2227
rect 12646 2193 12654 2227
rect 12600 2167 12654 2193
rect 11516 2087 11570 2113
rect 11516 2053 11524 2087
rect 11558 2053 11570 2087
rect 11516 2027 11570 2053
rect 11600 2087 11670 2113
rect 11600 2053 11618 2087
rect 11652 2053 11670 2087
rect 11600 2027 11670 2053
rect 11700 2087 11770 2113
rect 11700 2053 11718 2087
rect 11752 2053 11770 2087
rect 11700 2027 11770 2053
rect 11800 2087 11870 2113
rect 11800 2053 11818 2087
rect 11852 2053 11870 2087
rect 11800 2027 11870 2053
rect 11900 2087 11970 2113
rect 11900 2053 11918 2087
rect 11952 2053 11970 2087
rect 11900 2027 11970 2053
rect 12000 2027 12070 2113
rect 12100 2087 12170 2113
rect 12100 2053 12118 2087
rect 12152 2053 12170 2087
rect 12100 2027 12170 2053
rect 12200 2087 12270 2113
rect 12200 2053 12218 2087
rect 12252 2053 12270 2087
rect 12200 2027 12270 2053
rect 12300 2087 12370 2113
rect 12300 2053 12318 2087
rect 12352 2053 12370 2087
rect 12300 2027 12370 2053
rect 12400 2027 12470 2113
rect 12500 2087 12570 2113
rect 12500 2053 12518 2087
rect 12552 2053 12570 2087
rect 12500 2027 12570 2053
rect 12600 2087 12654 2113
rect 12600 2053 12612 2087
rect 12646 2053 12654 2087
rect 12600 2027 12654 2053
rect 11316 1947 11370 1973
rect 11316 1913 11324 1947
rect 11358 1913 11370 1947
rect 11316 1887 11370 1913
rect 11400 1947 11470 1973
rect 11400 1913 11418 1947
rect 11452 1913 11470 1947
rect 11400 1887 11470 1913
rect 11500 1887 11570 1973
rect 11600 1887 11670 1973
rect 11700 1887 11770 1973
rect 11800 1887 11870 1973
rect 11900 1947 11970 1973
rect 11900 1913 11918 1947
rect 11952 1913 11970 1947
rect 11900 1887 11970 1913
rect 12000 1947 12070 1973
rect 12000 1913 12018 1947
rect 12052 1913 12070 1947
rect 12000 1887 12070 1913
rect 12100 1947 12170 1973
rect 12100 1913 12118 1947
rect 12152 1913 12170 1947
rect 12100 1887 12170 1913
rect 12200 1947 12270 1973
rect 12200 1913 12218 1947
rect 12252 1913 12270 1947
rect 12200 1887 12270 1913
rect 12300 1947 12370 1973
rect 12300 1913 12318 1947
rect 12352 1913 12370 1947
rect 12300 1887 12370 1913
rect 12400 1887 12470 1973
rect 12500 1947 12570 1973
rect 12500 1913 12518 1947
rect 12552 1913 12570 1947
rect 12500 1887 12570 1913
rect 12600 1947 12654 1973
rect 12600 1913 12612 1947
rect 12646 1913 12654 1947
rect 12600 1887 12654 1913
rect 10816 1807 10870 1833
rect 10816 1773 10824 1807
rect 10858 1773 10870 1807
rect 10816 1747 10870 1773
rect 10900 1807 10970 1833
rect 10900 1773 10918 1807
rect 10952 1773 10970 1807
rect 10900 1747 10970 1773
rect 11000 1807 11070 1833
rect 11000 1773 11018 1807
rect 11052 1773 11070 1807
rect 11000 1747 11070 1773
rect 11100 1807 11170 1833
rect 11100 1773 11118 1807
rect 11152 1773 11170 1807
rect 11100 1747 11170 1773
rect 11200 1807 11270 1833
rect 11200 1773 11218 1807
rect 11252 1773 11270 1807
rect 11200 1747 11270 1773
rect 11300 1747 11370 1833
rect 11400 1807 11470 1833
rect 11400 1773 11418 1807
rect 11452 1773 11470 1807
rect 11400 1747 11470 1773
rect 11500 1807 11570 1833
rect 11500 1773 11518 1807
rect 11552 1773 11570 1807
rect 11500 1747 11570 1773
rect 11600 1807 11654 1833
rect 11600 1773 11612 1807
rect 11646 1773 11654 1807
rect 11600 1747 11654 1773
rect 9616 1667 9670 1693
rect 9616 1633 9624 1667
rect 9658 1633 9670 1667
rect 9616 1607 9670 1633
rect 9700 1667 9770 1693
rect 9700 1633 9718 1667
rect 9752 1633 9770 1667
rect 9700 1607 9770 1633
rect 9800 1667 9870 1693
rect 9800 1633 9818 1667
rect 9852 1633 9870 1667
rect 9800 1607 9870 1633
rect 9900 1607 9970 1693
rect 10000 1667 10070 1693
rect 10000 1633 10018 1667
rect 10052 1633 10070 1667
rect 10000 1607 10070 1633
rect 10100 1667 10170 1693
rect 10100 1633 10118 1667
rect 10152 1633 10170 1667
rect 10100 1607 10170 1633
rect 10200 1667 10270 1693
rect 10200 1633 10218 1667
rect 10252 1633 10270 1667
rect 10200 1607 10270 1633
rect 10300 1667 10370 1693
rect 10300 1633 10318 1667
rect 10352 1633 10370 1667
rect 10300 1607 10370 1633
rect 10400 1667 10470 1693
rect 10400 1633 10418 1667
rect 10452 1633 10470 1667
rect 10400 1607 10470 1633
rect 10500 1607 10570 1693
rect 10600 1667 10670 1693
rect 10600 1633 10618 1667
rect 10652 1633 10670 1667
rect 10600 1607 10670 1633
rect 10700 1667 10770 1693
rect 10700 1633 10718 1667
rect 10752 1633 10770 1667
rect 10700 1607 10770 1633
rect 10800 1667 10870 1693
rect 10800 1633 10818 1667
rect 10852 1633 10870 1667
rect 10800 1607 10870 1633
rect 10900 1667 10954 1693
rect 10900 1633 10912 1667
rect 10946 1633 10954 1667
rect 10900 1607 10954 1633
rect 9416 1527 9470 1553
rect 9416 1493 9424 1527
rect 9458 1493 9470 1527
rect 9416 1467 9470 1493
rect 9500 1527 9570 1553
rect 9500 1493 9518 1527
rect 9552 1493 9570 1527
rect 9500 1467 9570 1493
rect 9600 1527 9670 1553
rect 9600 1493 9618 1527
rect 9652 1493 9670 1527
rect 9600 1467 9670 1493
rect 9700 1467 9770 1553
rect 9800 1527 9870 1553
rect 9800 1493 9818 1527
rect 9852 1493 9870 1527
rect 9800 1467 9870 1493
rect 9900 1527 9970 1553
rect 9900 1493 9918 1527
rect 9952 1493 9970 1527
rect 9900 1467 9970 1493
rect 10000 1467 10070 1553
rect 10100 1527 10170 1553
rect 10100 1493 10118 1527
rect 10152 1493 10170 1527
rect 10100 1467 10170 1493
rect 10200 1527 10270 1553
rect 10200 1493 10218 1527
rect 10252 1493 10270 1527
rect 10200 1467 10270 1493
rect 10300 1467 10370 1553
rect 10400 1467 10470 1553
rect 10500 1527 10570 1553
rect 10500 1493 10518 1527
rect 10552 1493 10570 1527
rect 10500 1467 10570 1493
rect 10600 1527 10670 1553
rect 10600 1493 10618 1527
rect 10652 1493 10670 1527
rect 10600 1467 10670 1493
rect 10700 1527 10770 1553
rect 10700 1493 10718 1527
rect 10752 1493 10770 1527
rect 10700 1467 10770 1493
rect 10800 1527 10870 1553
rect 10800 1493 10818 1527
rect 10852 1493 10870 1527
rect 10800 1467 10870 1493
rect 10900 1527 10954 1553
rect 10900 1493 10912 1527
rect 10946 1493 10954 1527
rect 10900 1467 10954 1493
rect 9416 1387 9470 1413
rect 9416 1353 9424 1387
rect 9458 1353 9470 1387
rect 9416 1327 9470 1353
rect 9500 1387 9570 1413
rect 9500 1353 9518 1387
rect 9552 1353 9570 1387
rect 9500 1327 9570 1353
rect 9600 1327 9670 1413
rect 9700 1327 9770 1413
rect 9800 1387 9870 1413
rect 9800 1353 9818 1387
rect 9852 1353 9870 1387
rect 9800 1327 9870 1353
rect 9900 1387 9970 1413
rect 9900 1353 9918 1387
rect 9952 1353 9970 1387
rect 9900 1327 9970 1353
rect 10000 1387 10070 1413
rect 10000 1353 10018 1387
rect 10052 1353 10070 1387
rect 10000 1327 10070 1353
rect 10100 1387 10170 1413
rect 10100 1353 10118 1387
rect 10152 1353 10170 1387
rect 10100 1327 10170 1353
rect 10200 1387 10254 1413
rect 10200 1353 10212 1387
rect 10246 1353 10254 1387
rect 10200 1327 10254 1353
rect 6816 1157 6870 1183
rect 6816 1123 6824 1157
rect 6858 1123 6870 1157
rect 6816 1097 6870 1123
rect 6900 1157 6970 1183
rect 6900 1123 6918 1157
rect 6952 1123 6970 1157
rect 6900 1097 6970 1123
rect 7000 1097 7070 1183
rect 7100 1097 7170 1183
rect 7200 1097 7270 1183
rect 7300 1157 7370 1183
rect 7300 1123 7318 1157
rect 7352 1123 7370 1157
rect 7300 1097 7370 1123
rect 7400 1157 7470 1183
rect 7400 1123 7418 1157
rect 7452 1123 7470 1157
rect 7400 1097 7470 1123
rect 7500 1097 7570 1183
rect 7600 1097 7670 1183
rect 7700 1157 7770 1183
rect 7700 1123 7718 1157
rect 7752 1123 7770 1157
rect 7700 1097 7770 1123
rect 7800 1157 7870 1183
rect 7800 1123 7818 1157
rect 7852 1123 7870 1157
rect 7800 1097 7870 1123
rect 7900 1097 7970 1183
rect 8000 1157 8070 1183
rect 8000 1123 8018 1157
rect 8052 1123 8070 1157
rect 8000 1097 8070 1123
rect 8100 1157 8170 1183
rect 8100 1123 8118 1157
rect 8152 1123 8170 1157
rect 8100 1097 8170 1123
rect 8200 1097 8270 1183
rect 8300 1157 8370 1183
rect 8300 1123 8318 1157
rect 8352 1123 8370 1157
rect 8300 1097 8370 1123
rect 8400 1157 8470 1183
rect 8400 1123 8418 1157
rect 8452 1123 8470 1157
rect 8400 1097 8470 1123
rect 8500 1157 8570 1183
rect 8500 1123 8518 1157
rect 8552 1123 8570 1157
rect 8500 1097 8570 1123
rect 8600 1097 8670 1183
rect 8700 1157 8770 1183
rect 8700 1123 8718 1157
rect 8752 1123 8770 1157
rect 8700 1097 8770 1123
rect 8800 1157 8870 1183
rect 8800 1123 8818 1157
rect 8852 1123 8870 1157
rect 8800 1097 8870 1123
rect 8900 1157 8970 1183
rect 8900 1123 8918 1157
rect 8952 1123 8970 1157
rect 8900 1097 8970 1123
rect 9000 1097 9070 1183
rect 9100 1097 9170 1183
rect 9200 1157 9270 1183
rect 9200 1123 9218 1157
rect 9252 1123 9270 1157
rect 9200 1097 9270 1123
rect 9300 1157 9370 1183
rect 9300 1123 9318 1157
rect 9352 1123 9370 1157
rect 9300 1097 9370 1123
rect 9400 1097 9470 1183
rect 9500 1157 9570 1183
rect 9500 1123 9518 1157
rect 9552 1123 9570 1157
rect 9500 1097 9570 1123
rect 9600 1157 9654 1183
rect 9600 1123 9612 1157
rect 9646 1123 9654 1157
rect 9600 1097 9654 1123
rect 6516 1017 6570 1043
rect 6516 983 6524 1017
rect 6558 983 6570 1017
rect 6516 957 6570 983
rect 6600 1017 6670 1043
rect 6600 983 6618 1017
rect 6652 983 6670 1017
rect 6600 957 6670 983
rect 6700 1017 6770 1043
rect 6700 983 6718 1017
rect 6752 983 6770 1017
rect 6700 957 6770 983
rect 6800 1017 6870 1043
rect 6800 983 6818 1017
rect 6852 983 6870 1017
rect 6800 957 6870 983
rect 6900 1017 6954 1043
rect 6900 983 6912 1017
rect 6946 983 6954 1017
rect 6900 957 6954 983
rect 3916 877 3970 903
rect 3916 843 3924 877
rect 3958 843 3970 877
rect 3916 817 3970 843
rect 4000 877 4070 903
rect 4000 843 4018 877
rect 4052 843 4070 877
rect 4000 817 4070 843
rect 4100 877 4170 903
rect 4100 843 4118 877
rect 4152 843 4170 877
rect 4100 817 4170 843
rect 4200 877 4270 903
rect 4200 843 4218 877
rect 4252 843 4270 877
rect 4200 817 4270 843
rect 4300 877 4370 903
rect 4300 843 4318 877
rect 4352 843 4370 877
rect 4300 817 4370 843
rect 4400 877 4470 903
rect 4400 843 4418 877
rect 4452 843 4470 877
rect 4400 817 4470 843
rect 4500 817 4570 903
rect 4600 817 4670 903
rect 4700 877 4770 903
rect 4700 843 4718 877
rect 4752 843 4770 877
rect 4700 817 4770 843
rect 4800 877 4870 903
rect 4800 843 4818 877
rect 4852 843 4870 877
rect 4800 817 4870 843
rect 4900 877 4970 903
rect 4900 843 4918 877
rect 4952 843 4970 877
rect 4900 817 4970 843
rect 5000 877 5070 903
rect 5000 843 5018 877
rect 5052 843 5070 877
rect 5000 817 5070 843
rect 5100 877 5170 903
rect 5100 843 5118 877
rect 5152 843 5170 877
rect 5100 817 5170 843
rect 5200 817 5270 903
rect 5300 877 5370 903
rect 5300 843 5318 877
rect 5352 843 5370 877
rect 5300 817 5370 843
rect 5400 877 5470 903
rect 5400 843 5418 877
rect 5452 843 5470 877
rect 5400 817 5470 843
rect 5500 877 5570 903
rect 5500 843 5518 877
rect 5552 843 5570 877
rect 5500 817 5570 843
rect 5600 877 5670 903
rect 5600 843 5618 877
rect 5652 843 5670 877
rect 5600 817 5670 843
rect 5700 817 5770 903
rect 5800 817 5870 903
rect 5900 877 5970 903
rect 5900 843 5918 877
rect 5952 843 5970 877
rect 5900 817 5970 843
rect 6000 877 6070 903
rect 6000 843 6018 877
rect 6052 843 6070 877
rect 6000 817 6070 843
rect 6100 877 6170 903
rect 6100 843 6118 877
rect 6152 843 6170 877
rect 6100 817 6170 843
rect 6200 877 6270 903
rect 6200 843 6218 877
rect 6252 843 6270 877
rect 6200 817 6270 843
rect 6300 817 6370 903
rect 6400 877 6470 903
rect 6400 843 6418 877
rect 6452 843 6470 877
rect 6400 817 6470 843
rect 6500 877 6570 903
rect 6500 843 6518 877
rect 6552 843 6570 877
rect 6500 817 6570 843
rect 6600 877 6654 903
rect 6600 843 6612 877
rect 6646 843 6654 877
rect 6600 817 6654 843
rect 3716 737 3770 763
rect 3716 703 3724 737
rect 3758 703 3770 737
rect 3716 677 3770 703
rect 3800 737 3870 763
rect 3800 703 3818 737
rect 3852 703 3870 737
rect 3800 677 3870 703
rect 3900 737 3970 763
rect 3900 703 3918 737
rect 3952 703 3970 737
rect 3900 677 3970 703
rect 4000 737 4070 763
rect 4000 703 4018 737
rect 4052 703 4070 737
rect 4000 677 4070 703
rect 4100 677 4170 763
rect 4200 677 4270 763
rect 4300 677 4370 763
rect 4400 737 4470 763
rect 4400 703 4418 737
rect 4452 703 4470 737
rect 4400 677 4470 703
rect 4500 737 4570 763
rect 4500 703 4518 737
rect 4552 703 4570 737
rect 4500 677 4570 703
rect 4600 737 4654 763
rect 4600 703 4612 737
rect 4646 703 4654 737
rect 4600 677 4654 703
rect 2816 597 2870 623
rect 2816 563 2824 597
rect 2858 563 2870 597
rect 2816 537 2870 563
rect 2900 597 2970 623
rect 2900 563 2918 597
rect 2952 563 2970 597
rect 2900 537 2970 563
rect 3000 537 3070 623
rect 3100 537 3170 623
rect 3200 537 3270 623
rect 3300 537 3370 623
rect 3400 597 3470 623
rect 3400 563 3418 597
rect 3452 563 3470 597
rect 3400 537 3470 563
rect 3500 597 3570 623
rect 3500 563 3518 597
rect 3552 563 3570 597
rect 3500 537 3570 563
rect 3600 597 3670 623
rect 3600 563 3618 597
rect 3652 563 3670 597
rect 3600 537 3670 563
rect 3700 597 3770 623
rect 3700 563 3718 597
rect 3752 563 3770 597
rect 3700 537 3770 563
rect 3800 597 3870 623
rect 3800 563 3818 597
rect 3852 563 3870 597
rect 3800 537 3870 563
rect 3900 597 3954 623
rect 3900 563 3912 597
rect 3946 563 3954 597
rect 3900 537 3954 563
rect 4016 597 4070 623
rect 4016 563 4024 597
rect 4058 563 4070 597
rect 4016 537 4070 563
rect 4100 597 4154 623
rect 4100 563 4112 597
rect 4146 563 4154 597
rect 4100 537 4154 563
rect 4716 737 4770 763
rect 4716 703 4724 737
rect 4758 703 4770 737
rect 4716 677 4770 703
rect 4800 737 4870 763
rect 4800 703 4818 737
rect 4852 703 4870 737
rect 4800 677 4870 703
rect 4900 677 4970 763
rect 5000 737 5070 763
rect 5000 703 5018 737
rect 5052 703 5070 737
rect 5000 677 5070 703
rect 5100 737 5154 763
rect 5100 703 5112 737
rect 5146 703 5154 737
rect 5100 677 5154 703
rect 4216 597 4270 623
rect 4216 563 4224 597
rect 4258 563 4270 597
rect 4216 537 4270 563
rect 4300 597 4370 623
rect 4300 563 4318 597
rect 4352 563 4370 597
rect 4300 537 4370 563
rect 4400 537 4470 623
rect 4500 537 4570 623
rect 4600 597 4670 623
rect 4600 563 4618 597
rect 4652 563 4670 597
rect 4600 537 4670 563
rect 4700 597 4770 623
rect 4700 563 4718 597
rect 4752 563 4770 597
rect 4700 537 4770 563
rect 4800 597 4854 623
rect 4800 563 4812 597
rect 4846 563 4854 597
rect 4800 537 4854 563
rect 2716 457 2770 483
rect 2716 423 2724 457
rect 2758 423 2770 457
rect 2716 397 2770 423
rect 2800 457 2870 483
rect 2800 423 2818 457
rect 2852 423 2870 457
rect 2800 397 2870 423
rect 2900 457 2970 483
rect 2900 423 2918 457
rect 2952 423 2970 457
rect 2900 397 2970 423
rect 3000 397 3070 483
rect 3100 457 3170 483
rect 3100 423 3118 457
rect 3152 423 3170 457
rect 3100 397 3170 423
rect 3200 457 3270 483
rect 3200 423 3218 457
rect 3252 423 3270 457
rect 3200 397 3270 423
rect 3300 397 3370 483
rect 3400 397 3470 483
rect 3500 397 3570 483
rect 3600 457 3670 483
rect 3600 423 3618 457
rect 3652 423 3670 457
rect 3600 397 3670 423
rect 3700 457 3770 483
rect 3700 423 3718 457
rect 3752 423 3770 457
rect 3700 397 3770 423
rect 3800 457 3870 483
rect 3800 423 3818 457
rect 3852 423 3870 457
rect 3800 397 3870 423
rect 3900 457 3970 483
rect 3900 423 3918 457
rect 3952 423 3970 457
rect 3900 397 3970 423
rect 4000 457 4070 483
rect 4000 423 4018 457
rect 4052 423 4070 457
rect 4000 397 4070 423
rect 4100 397 4170 483
rect 4200 397 4270 483
rect 4300 457 4370 483
rect 4300 423 4318 457
rect 4352 423 4370 457
rect 4300 397 4370 423
rect 4400 457 4454 483
rect 4400 423 4412 457
rect 4446 423 4454 457
rect 4400 397 4454 423
rect 1816 317 1870 343
rect 1816 283 1824 317
rect 1858 283 1870 317
rect 1816 257 1870 283
rect 1900 317 1970 343
rect 1900 283 1918 317
rect 1952 283 1970 317
rect 1900 257 1970 283
rect 2000 257 2070 343
rect 2100 257 2170 343
rect 2200 257 2270 343
rect 2300 317 2370 343
rect 2300 283 2318 317
rect 2352 283 2370 317
rect 2300 257 2370 283
rect 2400 317 2470 343
rect 2400 283 2418 317
rect 2452 283 2470 317
rect 2400 257 2470 283
rect 2500 257 2570 343
rect 2600 257 2670 343
rect 2700 317 2770 343
rect 2700 283 2718 317
rect 2752 283 2770 317
rect 2700 257 2770 283
rect 2800 317 2854 343
rect 2800 283 2812 317
rect 2846 283 2854 317
rect 2800 257 2854 283
rect 1716 177 1770 203
rect 1716 143 1724 177
rect 1758 143 1770 177
rect 1716 117 1770 143
rect 1800 177 1854 203
rect 1800 143 1812 177
rect 1846 143 1854 177
rect 1800 117 1854 143
rect 2916 317 2970 343
rect 2916 283 2924 317
rect 2958 283 2970 317
rect 2916 257 2970 283
rect 3000 317 3054 343
rect 3000 283 3012 317
rect 3046 283 3054 317
rect 3000 257 3054 283
rect 4916 597 4970 623
rect 4916 563 4924 597
rect 4958 563 4970 597
rect 4916 537 4970 563
rect 5000 597 5054 623
rect 5000 563 5012 597
rect 5046 563 5054 597
rect 5000 537 5054 563
rect 5216 737 5270 763
rect 5216 703 5224 737
rect 5258 703 5270 737
rect 5216 677 5270 703
rect 5300 737 5370 763
rect 5300 703 5318 737
rect 5352 703 5370 737
rect 5300 677 5370 703
rect 5400 677 5470 763
rect 5500 677 5570 763
rect 5600 737 5670 763
rect 5600 703 5618 737
rect 5652 703 5670 737
rect 5600 677 5670 703
rect 5700 737 5754 763
rect 5700 703 5712 737
rect 5746 703 5754 737
rect 5700 677 5754 703
rect 5116 597 5170 623
rect 5116 563 5124 597
rect 5158 563 5170 597
rect 5116 537 5170 563
rect 5200 597 5254 623
rect 5200 563 5212 597
rect 5246 563 5254 597
rect 5200 537 5254 563
rect 4516 457 4570 483
rect 4516 423 4524 457
rect 4558 423 4570 457
rect 4516 397 4570 423
rect 4600 457 4670 483
rect 4600 423 4618 457
rect 4652 423 4670 457
rect 4600 397 4670 423
rect 4700 457 4770 483
rect 4700 423 4718 457
rect 4752 423 4770 457
rect 4700 397 4770 423
rect 4800 457 4870 483
rect 4800 423 4818 457
rect 4852 423 4870 457
rect 4800 397 4870 423
rect 4900 397 4970 483
rect 5000 457 5070 483
rect 5000 423 5018 457
rect 5052 423 5070 457
rect 5000 397 5070 423
rect 5100 457 5154 483
rect 5100 423 5112 457
rect 5146 423 5154 457
rect 5100 397 5154 423
rect 3116 317 3170 343
rect 3116 283 3124 317
rect 3158 283 3170 317
rect 3116 257 3170 283
rect 3200 317 3270 343
rect 3200 283 3218 317
rect 3252 283 3270 317
rect 3200 257 3270 283
rect 3300 317 3370 343
rect 3300 283 3318 317
rect 3352 283 3370 317
rect 3300 257 3370 283
rect 3400 257 3470 343
rect 3500 317 3570 343
rect 3500 283 3518 317
rect 3552 283 3570 317
rect 3500 257 3570 283
rect 3600 317 3670 343
rect 3600 283 3618 317
rect 3652 283 3670 317
rect 3600 257 3670 283
rect 3700 257 3770 343
rect 3800 317 3870 343
rect 3800 283 3818 317
rect 3852 283 3870 317
rect 3800 257 3870 283
rect 3900 317 3970 343
rect 3900 283 3918 317
rect 3952 283 3970 317
rect 3900 257 3970 283
rect 4000 317 4070 343
rect 4000 283 4018 317
rect 4052 283 4070 317
rect 4000 257 4070 283
rect 4100 317 4170 343
rect 4100 283 4118 317
rect 4152 283 4170 317
rect 4100 257 4170 283
rect 4200 317 4270 343
rect 4200 283 4218 317
rect 4252 283 4270 317
rect 4200 257 4270 283
rect 4300 317 4370 343
rect 4300 283 4318 317
rect 4352 283 4370 317
rect 4300 257 4370 283
rect 4400 317 4470 343
rect 4400 283 4418 317
rect 4452 283 4470 317
rect 4400 257 4470 283
rect 4500 317 4554 343
rect 4500 283 4512 317
rect 4546 283 4554 317
rect 4500 257 4554 283
rect 4616 317 4670 343
rect 4616 283 4624 317
rect 4658 283 4670 317
rect 4616 257 4670 283
rect 4700 317 4770 343
rect 4700 283 4718 317
rect 4752 283 4770 317
rect 4700 257 4770 283
rect 4800 317 4854 343
rect 4800 283 4812 317
rect 4846 283 4854 317
rect 4800 257 4854 283
rect 4916 317 4970 343
rect 4916 283 4924 317
rect 4958 283 4970 317
rect 4916 257 4970 283
rect 5000 317 5054 343
rect 5000 283 5012 317
rect 5046 283 5054 317
rect 5000 257 5054 283
rect 5816 737 5870 763
rect 5816 703 5824 737
rect 5858 703 5870 737
rect 5816 677 5870 703
rect 5900 737 5970 763
rect 5900 703 5918 737
rect 5952 703 5970 737
rect 5900 677 5970 703
rect 6000 677 6070 763
rect 6100 737 6170 763
rect 6100 703 6118 737
rect 6152 703 6170 737
rect 6100 677 6170 703
rect 6200 737 6254 763
rect 6200 703 6212 737
rect 6246 703 6254 737
rect 6200 677 6254 703
rect 6316 737 6370 763
rect 6316 703 6324 737
rect 6358 703 6370 737
rect 6316 677 6370 703
rect 6400 737 6454 763
rect 6400 703 6412 737
rect 6446 703 6454 737
rect 6400 677 6454 703
rect 7016 1017 7070 1043
rect 7016 983 7024 1017
rect 7058 983 7070 1017
rect 7016 957 7070 983
rect 7100 1017 7154 1043
rect 7100 983 7112 1017
rect 7146 983 7154 1017
rect 7100 957 7154 983
rect 7216 1017 7270 1043
rect 7216 983 7224 1017
rect 7258 983 7270 1017
rect 7216 957 7270 983
rect 7300 1017 7354 1043
rect 7300 983 7312 1017
rect 7346 983 7354 1017
rect 7300 957 7354 983
rect 6716 877 6770 903
rect 6716 843 6724 877
rect 6758 843 6770 877
rect 6716 817 6770 843
rect 6800 877 6870 903
rect 6800 843 6818 877
rect 6852 843 6870 877
rect 6800 817 6870 843
rect 6900 817 6970 903
rect 7000 877 7070 903
rect 7000 843 7018 877
rect 7052 843 7070 877
rect 7000 817 7070 843
rect 7100 877 7170 903
rect 7100 843 7118 877
rect 7152 843 7170 877
rect 7100 817 7170 843
rect 7200 877 7270 903
rect 7200 843 7218 877
rect 7252 843 7270 877
rect 7200 817 7270 843
rect 7300 877 7354 903
rect 7300 843 7312 877
rect 7346 843 7354 877
rect 7300 817 7354 843
rect 6516 737 6570 763
rect 6516 703 6524 737
rect 6558 703 6570 737
rect 6516 677 6570 703
rect 6600 737 6670 763
rect 6600 703 6618 737
rect 6652 703 6670 737
rect 6600 677 6670 703
rect 6700 677 6770 763
rect 6800 677 6870 763
rect 6900 737 6970 763
rect 6900 703 6918 737
rect 6952 703 6970 737
rect 6900 677 6970 703
rect 7000 737 7054 763
rect 7000 703 7012 737
rect 7046 703 7054 737
rect 7000 677 7054 703
rect 7416 1017 7470 1043
rect 7416 983 7424 1017
rect 7458 983 7470 1017
rect 7416 957 7470 983
rect 7500 1017 7570 1043
rect 7500 983 7518 1017
rect 7552 983 7570 1017
rect 7500 957 7570 983
rect 7600 1017 7670 1043
rect 7600 983 7618 1017
rect 7652 983 7670 1017
rect 7600 957 7670 983
rect 7700 1017 7770 1043
rect 7700 983 7718 1017
rect 7752 983 7770 1017
rect 7700 957 7770 983
rect 7800 1017 7870 1043
rect 7800 983 7818 1017
rect 7852 983 7870 1017
rect 7800 957 7870 983
rect 7900 957 7970 1043
rect 8000 957 8070 1043
rect 8100 957 8170 1043
rect 8200 1017 8270 1043
rect 8200 983 8218 1017
rect 8252 983 8270 1017
rect 8200 957 8270 983
rect 8300 1017 8370 1043
rect 8300 983 8318 1017
rect 8352 983 8370 1017
rect 8300 957 8370 983
rect 8400 1017 8470 1043
rect 8400 983 8418 1017
rect 8452 983 8470 1017
rect 8400 957 8470 983
rect 8500 1017 8570 1043
rect 8500 983 8518 1017
rect 8552 983 8570 1017
rect 8500 957 8570 983
rect 8600 1017 8654 1043
rect 8600 983 8612 1017
rect 8646 983 8654 1017
rect 8600 957 8654 983
rect 7416 877 7470 903
rect 7416 843 7424 877
rect 7458 843 7470 877
rect 7416 817 7470 843
rect 7500 877 7554 903
rect 7500 843 7512 877
rect 7546 843 7554 877
rect 7500 817 7554 843
rect 7616 877 7670 903
rect 7616 843 7624 877
rect 7658 843 7670 877
rect 7616 817 7670 843
rect 7700 877 7754 903
rect 7700 843 7712 877
rect 7746 843 7754 877
rect 7700 817 7754 843
rect 7816 877 7870 903
rect 7816 843 7824 877
rect 7858 843 7870 877
rect 7816 817 7870 843
rect 7900 877 7954 903
rect 7900 843 7912 877
rect 7946 843 7954 877
rect 7900 817 7954 843
rect 8016 877 8070 903
rect 8016 843 8024 877
rect 8058 843 8070 877
rect 8016 817 8070 843
rect 8100 877 8170 903
rect 8100 843 8118 877
rect 8152 843 8170 877
rect 8100 817 8170 843
rect 8200 817 8270 903
rect 8300 877 8370 903
rect 8300 843 8318 877
rect 8352 843 8370 877
rect 8300 817 8370 843
rect 8400 877 8470 903
rect 8400 843 8418 877
rect 8452 843 8470 877
rect 8400 817 8470 843
rect 8500 877 8570 903
rect 8500 843 8518 877
rect 8552 843 8570 877
rect 8500 817 8570 843
rect 8600 877 8654 903
rect 8600 843 8612 877
rect 8646 843 8654 877
rect 8600 817 8654 843
rect 8716 1017 8770 1043
rect 8716 983 8724 1017
rect 8758 983 8770 1017
rect 8716 957 8770 983
rect 8800 1017 8854 1043
rect 8800 983 8812 1017
rect 8846 983 8854 1017
rect 8800 957 8854 983
rect 8716 877 8770 903
rect 8716 843 8724 877
rect 8758 843 8770 877
rect 8716 817 8770 843
rect 8800 877 8854 903
rect 8800 843 8812 877
rect 8846 843 8854 877
rect 8800 817 8854 843
rect 8916 1017 8970 1043
rect 8916 983 8924 1017
rect 8958 983 8970 1017
rect 8916 957 8970 983
rect 9000 1017 9070 1043
rect 9000 983 9018 1017
rect 9052 983 9070 1017
rect 9000 957 9070 983
rect 9100 1017 9170 1043
rect 9100 983 9118 1017
rect 9152 983 9170 1017
rect 9100 957 9170 983
rect 9200 957 9270 1043
rect 9300 957 9370 1043
rect 9400 1017 9470 1043
rect 9400 983 9418 1017
rect 9452 983 9470 1017
rect 9400 957 9470 983
rect 9500 1017 9554 1043
rect 9500 983 9512 1017
rect 9546 983 9554 1017
rect 9500 957 9554 983
rect 11716 1807 11770 1833
rect 11716 1773 11724 1807
rect 11758 1773 11770 1807
rect 11716 1747 11770 1773
rect 11800 1807 11870 1833
rect 11800 1773 11818 1807
rect 11852 1773 11870 1807
rect 11800 1747 11870 1773
rect 11900 1807 11954 1833
rect 11900 1773 11912 1807
rect 11946 1773 11954 1807
rect 11900 1747 11954 1773
rect 11016 1667 11070 1693
rect 11016 1633 11024 1667
rect 11058 1633 11070 1667
rect 11016 1607 11070 1633
rect 11100 1667 11170 1693
rect 11100 1633 11118 1667
rect 11152 1633 11170 1667
rect 11100 1607 11170 1633
rect 11200 1667 11270 1693
rect 11200 1633 11218 1667
rect 11252 1633 11270 1667
rect 11200 1607 11270 1633
rect 11300 1607 11370 1693
rect 11400 1607 11470 1693
rect 11500 1607 11570 1693
rect 11600 1667 11670 1693
rect 11600 1633 11618 1667
rect 11652 1633 11670 1667
rect 11600 1607 11670 1633
rect 11700 1667 11754 1693
rect 11700 1633 11712 1667
rect 11746 1633 11754 1667
rect 11700 1607 11754 1633
rect 11016 1527 11070 1553
rect 11016 1493 11024 1527
rect 11058 1493 11070 1527
rect 11016 1467 11070 1493
rect 11100 1527 11154 1553
rect 11100 1493 11112 1527
rect 11146 1493 11154 1527
rect 11100 1467 11154 1493
rect 10316 1387 10370 1413
rect 10316 1353 10324 1387
rect 10358 1353 10370 1387
rect 10316 1327 10370 1353
rect 10400 1387 10470 1413
rect 10400 1353 10418 1387
rect 10452 1353 10470 1387
rect 10400 1327 10470 1353
rect 10500 1327 10570 1413
rect 10600 1327 10670 1413
rect 10700 1327 10770 1413
rect 10800 1327 10870 1413
rect 10900 1387 10970 1413
rect 10900 1353 10918 1387
rect 10952 1353 10970 1387
rect 10900 1327 10970 1353
rect 11000 1387 11070 1413
rect 11000 1353 11018 1387
rect 11052 1353 11070 1387
rect 11000 1327 11070 1353
rect 11100 1387 11154 1413
rect 11100 1353 11112 1387
rect 11146 1353 11154 1387
rect 11100 1327 11154 1353
rect 12716 2227 12770 2253
rect 12716 2193 12724 2227
rect 12758 2193 12770 2227
rect 12716 2167 12770 2193
rect 12800 2227 12854 2253
rect 12800 2193 12812 2227
rect 12846 2193 12854 2227
rect 12800 2167 12854 2193
rect 12912 2242 12970 2253
rect 12912 2208 12924 2242
rect 12958 2208 12970 2242
rect 12912 2167 12970 2208
rect 13000 2227 13070 2253
rect 13000 2193 13018 2227
rect 13052 2193 13070 2227
rect 13000 2167 13070 2193
rect 13100 2212 13158 2253
rect 13100 2178 13112 2212
rect 13146 2178 13158 2212
rect 13100 2167 13158 2178
rect 13220 2227 13280 2253
rect 13220 2193 13228 2227
rect 13262 2193 13280 2227
rect 13220 2167 13280 2193
rect 13310 2227 13380 2253
rect 13310 2193 13328 2227
rect 13362 2193 13380 2227
rect 13310 2167 13380 2193
rect 13410 2227 13480 2253
rect 13410 2193 13428 2227
rect 13462 2193 13480 2227
rect 13410 2167 13480 2193
rect 13510 2227 13580 2253
rect 13510 2193 13528 2227
rect 13562 2193 13580 2227
rect 13510 2167 13580 2193
rect 13610 2227 13670 2253
rect 13610 2193 13628 2227
rect 13662 2193 13670 2227
rect 13610 2167 13670 2193
rect 12716 2087 12770 2113
rect 12716 2053 12724 2087
rect 12758 2053 12770 2087
rect 12716 2027 12770 2053
rect 12800 2087 12854 2113
rect 12800 2053 12812 2087
rect 12846 2053 12854 2087
rect 12800 2027 12854 2053
rect 12912 2102 12970 2113
rect 12912 2068 12924 2102
rect 12958 2068 12970 2102
rect 12912 2027 12970 2068
rect 13000 2087 13070 2113
rect 13000 2053 13018 2087
rect 13052 2053 13070 2087
rect 13000 2027 13070 2053
rect 13100 2072 13158 2113
rect 13100 2038 13112 2072
rect 13146 2038 13158 2072
rect 13100 2027 13158 2038
rect 13220 2087 13280 2113
rect 13220 2053 13228 2087
rect 13262 2053 13280 2087
rect 13220 2027 13280 2053
rect 13310 2087 13380 2113
rect 13310 2053 13328 2087
rect 13362 2053 13380 2087
rect 13310 2027 13380 2053
rect 13410 2087 13480 2113
rect 13410 2053 13428 2087
rect 13462 2053 13480 2087
rect 13410 2027 13480 2053
rect 13510 2087 13580 2113
rect 13510 2053 13528 2087
rect 13562 2053 13580 2087
rect 13510 2027 13580 2053
rect 13610 2087 13670 2113
rect 13610 2053 13628 2087
rect 13662 2053 13670 2087
rect 13610 2027 13670 2053
rect 12716 1947 12770 1973
rect 12716 1913 12724 1947
rect 12758 1913 12770 1947
rect 12716 1887 12770 1913
rect 12800 1947 12854 1973
rect 12800 1913 12812 1947
rect 12846 1913 12854 1947
rect 12800 1887 12854 1913
rect 12912 1962 12970 1973
rect 12912 1928 12924 1962
rect 12958 1928 12970 1962
rect 12912 1887 12970 1928
rect 13000 1947 13070 1973
rect 13000 1913 13018 1947
rect 13052 1913 13070 1947
rect 13000 1887 13070 1913
rect 13100 1932 13158 1973
rect 13100 1898 13112 1932
rect 13146 1898 13158 1932
rect 13100 1887 13158 1898
rect 13220 1947 13280 1973
rect 13220 1913 13228 1947
rect 13262 1913 13280 1947
rect 13220 1887 13280 1913
rect 13310 1947 13380 1973
rect 13310 1913 13328 1947
rect 13362 1913 13380 1947
rect 13310 1887 13380 1913
rect 13410 1947 13480 1973
rect 13410 1913 13428 1947
rect 13462 1913 13480 1947
rect 13410 1887 13480 1913
rect 13510 1947 13580 1973
rect 13510 1913 13528 1947
rect 13562 1913 13580 1947
rect 13510 1887 13580 1913
rect 13610 1947 13670 1973
rect 13610 1913 13628 1947
rect 13662 1913 13670 1947
rect 13610 1887 13670 1913
rect 12016 1807 12070 1833
rect 12016 1773 12024 1807
rect 12058 1773 12070 1807
rect 12016 1747 12070 1773
rect 12100 1807 12170 1833
rect 12100 1773 12118 1807
rect 12152 1773 12170 1807
rect 12100 1747 12170 1773
rect 12200 1807 12270 1833
rect 12200 1773 12218 1807
rect 12252 1773 12270 1807
rect 12200 1747 12270 1773
rect 12300 1747 12370 1833
rect 12400 1747 12470 1833
rect 12500 1747 12570 1833
rect 12600 1807 12670 1833
rect 12600 1773 12618 1807
rect 12652 1773 12670 1807
rect 12600 1747 12670 1773
rect 12700 1807 12770 1833
rect 12700 1773 12718 1807
rect 12752 1773 12770 1807
rect 12700 1747 12770 1773
rect 12800 1807 12854 1833
rect 12800 1773 12812 1807
rect 12846 1773 12854 1807
rect 12800 1747 12854 1773
rect 12912 1822 12970 1833
rect 12912 1788 12924 1822
rect 12958 1788 12970 1822
rect 12912 1747 12970 1788
rect 13000 1807 13070 1833
rect 13000 1773 13018 1807
rect 13052 1773 13070 1807
rect 13000 1747 13070 1773
rect 13100 1792 13158 1833
rect 13100 1758 13112 1792
rect 13146 1758 13158 1792
rect 13100 1747 13158 1758
rect 13220 1807 13280 1833
rect 13220 1773 13228 1807
rect 13262 1773 13280 1807
rect 13220 1747 13280 1773
rect 13310 1807 13380 1833
rect 13310 1773 13328 1807
rect 13362 1773 13380 1807
rect 13310 1747 13380 1773
rect 13410 1807 13480 1833
rect 13410 1773 13428 1807
rect 13462 1773 13480 1807
rect 13410 1747 13480 1773
rect 13510 1807 13580 1833
rect 13510 1773 13528 1807
rect 13562 1773 13580 1807
rect 13510 1747 13580 1773
rect 13610 1807 13670 1833
rect 13610 1773 13628 1807
rect 13662 1773 13670 1807
rect 13610 1747 13670 1773
rect 11816 1667 11870 1693
rect 11816 1633 11824 1667
rect 11858 1633 11870 1667
rect 11816 1607 11870 1633
rect 11900 1667 11970 1693
rect 11900 1633 11918 1667
rect 11952 1633 11970 1667
rect 11900 1607 11970 1633
rect 12000 1607 12070 1693
rect 12100 1667 12170 1693
rect 12100 1633 12118 1667
rect 12152 1633 12170 1667
rect 12100 1607 12170 1633
rect 12200 1667 12270 1693
rect 12200 1633 12218 1667
rect 12252 1633 12270 1667
rect 12200 1607 12270 1633
rect 12300 1667 12370 1693
rect 12300 1633 12318 1667
rect 12352 1633 12370 1667
rect 12300 1607 12370 1633
rect 12400 1667 12470 1693
rect 12400 1633 12418 1667
rect 12452 1633 12470 1667
rect 12400 1607 12470 1633
rect 12500 1667 12570 1693
rect 12500 1633 12518 1667
rect 12552 1633 12570 1667
rect 12500 1607 12570 1633
rect 12600 1667 12670 1693
rect 12600 1633 12618 1667
rect 12652 1633 12670 1667
rect 12600 1607 12670 1633
rect 12700 1667 12770 1693
rect 12700 1633 12718 1667
rect 12752 1633 12770 1667
rect 12700 1607 12770 1633
rect 12800 1607 12854 1693
rect 12912 1682 12970 1693
rect 12912 1648 12924 1682
rect 12958 1648 12970 1682
rect 12912 1607 12970 1648
rect 13000 1667 13070 1693
rect 13000 1633 13018 1667
rect 13052 1633 13070 1667
rect 13000 1607 13070 1633
rect 13100 1652 13158 1693
rect 13100 1618 13112 1652
rect 13146 1618 13158 1652
rect 13100 1607 13158 1618
rect 13220 1667 13280 1693
rect 13220 1633 13228 1667
rect 13262 1633 13280 1667
rect 13220 1607 13280 1633
rect 13310 1667 13380 1693
rect 13310 1633 13328 1667
rect 13362 1633 13380 1667
rect 13310 1607 13380 1633
rect 13410 1667 13480 1693
rect 13410 1633 13428 1667
rect 13462 1633 13480 1667
rect 13410 1607 13480 1633
rect 13510 1667 13580 1693
rect 13510 1633 13528 1667
rect 13562 1633 13580 1667
rect 13510 1607 13580 1633
rect 13610 1667 13670 1693
rect 13610 1633 13628 1667
rect 13662 1633 13670 1667
rect 13610 1607 13670 1633
rect 11216 1527 11270 1553
rect 11216 1493 11224 1527
rect 11258 1493 11270 1527
rect 11216 1467 11270 1493
rect 11300 1527 11370 1553
rect 11300 1493 11318 1527
rect 11352 1493 11370 1527
rect 11300 1467 11370 1493
rect 11400 1467 11470 1553
rect 11500 1527 11570 1553
rect 11500 1493 11518 1527
rect 11552 1493 11570 1527
rect 11500 1467 11570 1493
rect 11600 1527 11670 1553
rect 11600 1493 11618 1527
rect 11652 1493 11670 1527
rect 11600 1467 11670 1493
rect 11700 1467 11770 1553
rect 11800 1467 11870 1553
rect 11900 1527 11970 1553
rect 11900 1493 11918 1527
rect 11952 1493 11970 1527
rect 11900 1467 11970 1493
rect 12000 1527 12054 1553
rect 12000 1493 12012 1527
rect 12046 1493 12054 1527
rect 12000 1467 12054 1493
rect 11216 1387 11270 1413
rect 11216 1353 11224 1387
rect 11258 1353 11270 1387
rect 11216 1327 11270 1353
rect 11300 1387 11370 1413
rect 11300 1353 11318 1387
rect 11352 1353 11370 1387
rect 11300 1327 11370 1353
rect 11400 1327 11470 1413
rect 11500 1387 11570 1413
rect 11500 1353 11518 1387
rect 11552 1353 11570 1387
rect 11500 1327 11570 1353
rect 11600 1387 11670 1413
rect 11600 1353 11618 1387
rect 11652 1353 11670 1387
rect 11600 1327 11670 1353
rect 11700 1387 11754 1413
rect 11700 1353 11712 1387
rect 11746 1353 11754 1387
rect 11700 1327 11754 1353
rect 9716 1157 9770 1183
rect 9716 1123 9724 1157
rect 9758 1123 9770 1157
rect 9716 1097 9770 1123
rect 9800 1157 9870 1183
rect 9800 1123 9818 1157
rect 9852 1123 9870 1157
rect 9800 1097 9870 1123
rect 9900 1157 9970 1183
rect 9900 1123 9918 1157
rect 9952 1123 9970 1157
rect 9900 1097 9970 1123
rect 10000 1157 10070 1183
rect 10000 1123 10018 1157
rect 10052 1123 10070 1157
rect 10000 1097 10070 1123
rect 10100 1097 10170 1183
rect 10200 1097 10270 1183
rect 10300 1097 10370 1183
rect 10400 1097 10470 1183
rect 10500 1157 10570 1183
rect 10500 1123 10518 1157
rect 10552 1123 10570 1157
rect 10500 1097 10570 1123
rect 10600 1157 10670 1183
rect 10600 1123 10618 1157
rect 10652 1123 10670 1157
rect 10600 1097 10670 1123
rect 10700 1157 10770 1183
rect 10700 1123 10718 1157
rect 10752 1123 10770 1157
rect 10700 1097 10770 1123
rect 10800 1097 10870 1183
rect 10900 1157 10970 1183
rect 10900 1123 10918 1157
rect 10952 1123 10970 1157
rect 10900 1097 10970 1123
rect 11000 1157 11054 1183
rect 11000 1123 11012 1157
rect 11046 1123 11054 1157
rect 11000 1097 11054 1123
rect 9616 1017 9670 1043
rect 9616 983 9624 1017
rect 9658 983 9670 1017
rect 9616 957 9670 983
rect 9700 1017 9770 1043
rect 9700 983 9718 1017
rect 9752 983 9770 1017
rect 9700 957 9770 983
rect 9800 1017 9870 1043
rect 9800 983 9818 1017
rect 9852 983 9870 1017
rect 9800 957 9870 983
rect 9900 1017 9954 1043
rect 9900 983 9912 1017
rect 9946 983 9954 1017
rect 9900 957 9954 983
rect 8916 877 8970 903
rect 8916 843 8924 877
rect 8958 843 8970 877
rect 8916 817 8970 843
rect 9000 877 9070 903
rect 9000 843 9018 877
rect 9052 843 9070 877
rect 9000 817 9070 843
rect 9100 877 9170 903
rect 9100 843 9118 877
rect 9152 843 9170 877
rect 9100 817 9170 843
rect 9200 817 9270 903
rect 9300 817 9370 903
rect 9400 877 9470 903
rect 9400 843 9418 877
rect 9452 843 9470 877
rect 9400 817 9470 843
rect 9500 877 9570 903
rect 9500 843 9518 877
rect 9552 843 9570 877
rect 9500 817 9570 843
rect 9600 817 9670 903
rect 9700 877 9770 903
rect 9700 843 9718 877
rect 9752 843 9770 877
rect 9700 817 9770 843
rect 9800 877 9870 903
rect 9800 843 9818 877
rect 9852 843 9870 877
rect 9800 817 9870 843
rect 9900 877 9954 903
rect 9900 843 9912 877
rect 9946 843 9954 877
rect 9900 817 9954 843
rect 7116 737 7170 763
rect 7116 703 7124 737
rect 7158 703 7170 737
rect 7116 677 7170 703
rect 7200 737 7270 763
rect 7200 703 7218 737
rect 7252 703 7270 737
rect 7200 677 7270 703
rect 7300 737 7370 763
rect 7300 703 7318 737
rect 7352 703 7370 737
rect 7300 677 7370 703
rect 7400 737 7470 763
rect 7400 703 7418 737
rect 7452 703 7470 737
rect 7400 677 7470 703
rect 7500 737 7570 763
rect 7500 703 7518 737
rect 7552 703 7570 737
rect 7500 677 7570 703
rect 7600 737 7670 763
rect 7600 703 7618 737
rect 7652 703 7670 737
rect 7600 677 7670 703
rect 7700 737 7770 763
rect 7700 703 7718 737
rect 7752 703 7770 737
rect 7700 677 7770 703
rect 7800 677 7870 763
rect 7900 737 7970 763
rect 7900 703 7918 737
rect 7952 703 7970 737
rect 7900 677 7970 703
rect 8000 737 8070 763
rect 8000 703 8018 737
rect 8052 703 8070 737
rect 8000 677 8070 703
rect 8100 737 8170 763
rect 8100 703 8118 737
rect 8152 703 8170 737
rect 8100 677 8170 703
rect 8200 737 8270 763
rect 8200 703 8218 737
rect 8252 703 8270 737
rect 8200 677 8270 703
rect 8300 737 8370 763
rect 8300 703 8318 737
rect 8352 703 8370 737
rect 8300 677 8370 703
rect 8400 737 8470 763
rect 8400 703 8418 737
rect 8452 703 8470 737
rect 8400 677 8470 703
rect 8500 677 8570 763
rect 8600 737 8670 763
rect 8600 703 8618 737
rect 8652 703 8670 737
rect 8600 677 8670 703
rect 8700 737 8770 763
rect 8700 703 8718 737
rect 8752 703 8770 737
rect 8700 677 8770 703
rect 8800 737 8870 763
rect 8800 703 8818 737
rect 8852 703 8870 737
rect 8800 677 8870 703
rect 8900 677 8970 763
rect 9000 737 9070 763
rect 9000 703 9018 737
rect 9052 703 9070 737
rect 9000 677 9070 703
rect 9100 737 9154 763
rect 9100 703 9112 737
rect 9146 703 9154 737
rect 9100 677 9154 703
rect 5316 597 5370 623
rect 5316 563 5324 597
rect 5358 563 5370 597
rect 5316 537 5370 563
rect 5400 597 5470 623
rect 5400 563 5418 597
rect 5452 563 5470 597
rect 5400 537 5470 563
rect 5500 597 5570 623
rect 5500 563 5518 597
rect 5552 563 5570 597
rect 5500 537 5570 563
rect 5600 537 5670 623
rect 5700 537 5770 623
rect 5800 537 5870 623
rect 5900 597 5970 623
rect 5900 563 5918 597
rect 5952 563 5970 597
rect 5900 537 5970 563
rect 6000 597 6070 623
rect 6000 563 6018 597
rect 6052 563 6070 597
rect 6000 537 6070 563
rect 6100 597 6170 623
rect 6100 563 6118 597
rect 6152 563 6170 597
rect 6100 537 6170 563
rect 6200 537 6270 623
rect 6300 597 6370 623
rect 6300 563 6318 597
rect 6352 563 6370 597
rect 6300 537 6370 563
rect 6400 597 6470 623
rect 6400 563 6418 597
rect 6452 563 6470 597
rect 6400 537 6470 563
rect 6500 537 6570 623
rect 6600 537 6670 623
rect 6700 597 6770 623
rect 6700 563 6718 597
rect 6752 563 6770 597
rect 6700 537 6770 563
rect 6800 597 6870 623
rect 6800 563 6818 597
rect 6852 563 6870 597
rect 6800 537 6870 563
rect 6900 597 6970 623
rect 6900 563 6918 597
rect 6952 563 6970 597
rect 6900 537 6970 563
rect 7000 537 7070 623
rect 7100 537 7170 623
rect 7200 597 7270 623
rect 7200 563 7218 597
rect 7252 563 7270 597
rect 7200 537 7270 563
rect 7300 597 7370 623
rect 7300 563 7318 597
rect 7352 563 7370 597
rect 7300 537 7370 563
rect 7400 537 7470 623
rect 7500 597 7570 623
rect 7500 563 7518 597
rect 7552 563 7570 597
rect 7500 537 7570 563
rect 7600 597 7670 623
rect 7600 563 7618 597
rect 7652 563 7670 597
rect 7600 537 7670 563
rect 7700 597 7770 623
rect 7700 563 7718 597
rect 7752 563 7770 597
rect 7700 537 7770 563
rect 7800 597 7870 623
rect 7800 563 7818 597
rect 7852 563 7870 597
rect 7800 537 7870 563
rect 7900 537 7970 623
rect 8000 537 8070 623
rect 8100 597 8170 623
rect 8100 563 8118 597
rect 8152 563 8170 597
rect 8100 537 8170 563
rect 8200 597 8270 623
rect 8200 563 8218 597
rect 8252 563 8270 597
rect 8200 537 8270 563
rect 8300 597 8354 623
rect 8300 563 8312 597
rect 8346 563 8354 597
rect 8300 537 8354 563
rect 5216 457 5270 483
rect 5216 423 5224 457
rect 5258 423 5270 457
rect 5216 397 5270 423
rect 5300 457 5354 483
rect 5300 423 5312 457
rect 5346 423 5354 457
rect 5300 397 5354 423
rect 5416 457 5470 483
rect 5416 423 5424 457
rect 5458 423 5470 457
rect 5416 397 5470 423
rect 5500 457 5570 483
rect 5500 423 5518 457
rect 5552 423 5570 457
rect 5500 397 5570 423
rect 5600 457 5670 483
rect 5600 423 5618 457
rect 5652 423 5670 457
rect 5600 397 5670 423
rect 5700 457 5770 483
rect 5700 423 5718 457
rect 5752 423 5770 457
rect 5700 397 5770 423
rect 5800 457 5870 483
rect 5800 423 5818 457
rect 5852 423 5870 457
rect 5800 397 5870 423
rect 5900 397 5970 483
rect 6000 457 6070 483
rect 6000 423 6018 457
rect 6052 423 6070 457
rect 6000 397 6070 423
rect 6100 457 6154 483
rect 6100 423 6112 457
rect 6146 423 6154 457
rect 6100 397 6154 423
rect 5116 317 5170 343
rect 5116 283 5124 317
rect 5158 283 5170 317
rect 5116 257 5170 283
rect 5200 317 5270 343
rect 5200 283 5218 317
rect 5252 283 5270 317
rect 5200 257 5270 283
rect 5300 317 5370 343
rect 5300 283 5318 317
rect 5352 283 5370 317
rect 5300 257 5370 283
rect 5400 257 5470 343
rect 5500 257 5570 343
rect 5600 257 5670 343
rect 5700 317 5770 343
rect 5700 283 5718 317
rect 5752 283 5770 317
rect 5700 257 5770 283
rect 5800 317 5854 343
rect 5800 283 5812 317
rect 5846 283 5854 317
rect 5800 257 5854 283
rect 5916 317 5970 343
rect 5916 283 5924 317
rect 5958 283 5970 317
rect 5916 257 5970 283
rect 6000 317 6054 343
rect 6000 283 6012 317
rect 6046 283 6054 317
rect 6000 257 6054 283
rect 6216 457 6270 483
rect 6216 423 6224 457
rect 6258 423 6270 457
rect 6216 397 6270 423
rect 6300 457 6370 483
rect 6300 423 6318 457
rect 6352 423 6370 457
rect 6300 397 6370 423
rect 6400 457 6454 483
rect 6400 423 6412 457
rect 6446 423 6454 457
rect 6400 397 6454 423
rect 6116 317 6170 343
rect 6116 283 6124 317
rect 6158 283 6170 317
rect 6116 257 6170 283
rect 6200 317 6254 343
rect 6200 283 6212 317
rect 6246 283 6254 317
rect 6200 257 6254 283
rect 6316 317 6370 343
rect 6316 283 6324 317
rect 6358 283 6370 317
rect 6316 257 6370 283
rect 6400 317 6454 343
rect 6400 283 6412 317
rect 6446 283 6454 317
rect 6400 257 6454 283
rect 6516 457 6570 483
rect 6516 423 6524 457
rect 6558 423 6570 457
rect 6516 397 6570 423
rect 6600 457 6670 483
rect 6600 423 6618 457
rect 6652 423 6670 457
rect 6600 397 6670 423
rect 6700 397 6770 483
rect 6800 397 6870 483
rect 6900 457 6970 483
rect 6900 423 6918 457
rect 6952 423 6970 457
rect 6900 397 6970 423
rect 7000 457 7070 483
rect 7000 423 7018 457
rect 7052 423 7070 457
rect 7000 397 7070 423
rect 7100 457 7154 483
rect 7100 423 7112 457
rect 7146 423 7154 457
rect 7100 397 7154 423
rect 6516 317 6570 343
rect 6516 283 6524 317
rect 6558 283 6570 317
rect 6516 257 6570 283
rect 6600 317 6654 343
rect 6600 283 6612 317
rect 6646 283 6654 317
rect 6600 257 6654 283
rect 6716 317 6770 343
rect 6716 283 6724 317
rect 6758 283 6770 317
rect 6716 257 6770 283
rect 6800 317 6854 343
rect 6800 283 6812 317
rect 6846 283 6854 317
rect 6800 257 6854 283
rect 7216 457 7270 483
rect 7216 423 7224 457
rect 7258 423 7270 457
rect 7216 397 7270 423
rect 7300 457 7354 483
rect 7300 423 7312 457
rect 7346 423 7354 457
rect 7300 397 7354 423
rect 7416 457 7470 483
rect 7416 423 7424 457
rect 7458 423 7470 457
rect 7416 397 7470 423
rect 7500 457 7554 483
rect 7500 423 7512 457
rect 7546 423 7554 457
rect 7500 397 7554 423
rect 7616 457 7670 483
rect 7616 423 7624 457
rect 7658 423 7670 457
rect 7616 397 7670 423
rect 7700 457 7770 483
rect 7700 423 7718 457
rect 7752 423 7770 457
rect 7700 397 7770 423
rect 7800 457 7870 483
rect 7800 423 7818 457
rect 7852 423 7870 457
rect 7800 397 7870 423
rect 7900 397 7970 483
rect 8000 397 8070 483
rect 8100 397 8170 483
rect 8200 457 8270 483
rect 8200 423 8218 457
rect 8252 423 8270 457
rect 8200 397 8270 423
rect 8300 457 8354 483
rect 8300 423 8312 457
rect 8346 423 8354 457
rect 8300 397 8354 423
rect 6916 317 6970 343
rect 6916 283 6924 317
rect 6958 283 6970 317
rect 6916 257 6970 283
rect 7000 317 7070 343
rect 7000 283 7018 317
rect 7052 283 7070 317
rect 7000 257 7070 283
rect 7100 257 7170 343
rect 7200 317 7270 343
rect 7200 283 7218 317
rect 7252 283 7270 317
rect 7200 257 7270 283
rect 7300 317 7370 343
rect 7300 283 7318 317
rect 7352 283 7370 317
rect 7300 257 7370 283
rect 7400 317 7470 343
rect 7400 283 7418 317
rect 7452 283 7470 317
rect 7400 257 7470 283
rect 7500 257 7570 343
rect 7600 257 7670 343
rect 7700 317 7770 343
rect 7700 283 7718 317
rect 7752 283 7770 317
rect 7700 257 7770 283
rect 7800 317 7854 343
rect 7800 283 7812 317
rect 7846 283 7854 317
rect 7800 257 7854 283
rect 1916 177 1970 203
rect 1916 143 1924 177
rect 1958 143 1970 177
rect 1916 117 1970 143
rect 2000 177 2070 203
rect 2000 143 2018 177
rect 2052 143 2070 177
rect 2000 117 2070 143
rect 2100 117 2170 203
rect 2200 177 2270 203
rect 2200 143 2218 177
rect 2252 143 2270 177
rect 2200 117 2270 143
rect 2300 177 2370 203
rect 2300 143 2318 177
rect 2352 143 2370 177
rect 2300 117 2370 143
rect 2400 117 2470 203
rect 2500 177 2570 203
rect 2500 143 2518 177
rect 2552 143 2570 177
rect 2500 117 2570 143
rect 2600 177 2670 203
rect 2600 143 2618 177
rect 2652 143 2670 177
rect 2600 117 2670 143
rect 2700 117 2770 203
rect 2800 117 2870 203
rect 2900 177 2970 203
rect 2900 143 2918 177
rect 2952 143 2970 177
rect 2900 117 2970 143
rect 3000 177 3070 203
rect 3000 143 3018 177
rect 3052 143 3070 177
rect 3000 117 3070 143
rect 3100 117 3170 203
rect 3200 117 3270 203
rect 3300 177 3370 203
rect 3300 143 3318 177
rect 3352 143 3370 177
rect 3300 117 3370 143
rect 3400 177 3470 203
rect 3400 143 3418 177
rect 3452 143 3470 177
rect 3400 117 3470 143
rect 3500 117 3570 203
rect 3600 117 3670 203
rect 3700 177 3770 203
rect 3700 143 3718 177
rect 3752 143 3770 177
rect 3700 117 3770 143
rect 3800 177 3870 203
rect 3800 143 3818 177
rect 3852 143 3870 177
rect 3800 117 3870 143
rect 3900 177 3970 203
rect 3900 143 3918 177
rect 3952 143 3970 177
rect 3900 117 3970 143
rect 4000 177 4070 203
rect 4000 143 4018 177
rect 4052 143 4070 177
rect 4000 117 4070 143
rect 4100 177 4170 203
rect 4100 143 4118 177
rect 4152 143 4170 177
rect 4100 117 4170 143
rect 4200 177 4270 203
rect 4200 143 4218 177
rect 4252 143 4270 177
rect 4200 117 4270 143
rect 4300 177 4370 203
rect 4300 143 4318 177
rect 4352 143 4370 177
rect 4300 117 4370 143
rect 4400 117 4470 203
rect 4500 117 4570 203
rect 4600 117 4670 203
rect 4700 177 4770 203
rect 4700 143 4718 177
rect 4752 143 4770 177
rect 4700 117 4770 143
rect 4800 177 4870 203
rect 4800 143 4818 177
rect 4852 143 4870 177
rect 4800 117 4870 143
rect 4900 177 4970 203
rect 4900 143 4918 177
rect 4952 143 4970 177
rect 4900 117 4970 143
rect 5000 177 5070 203
rect 5000 143 5018 177
rect 5052 143 5070 177
rect 5000 117 5070 143
rect 5100 117 5170 203
rect 5200 117 5270 203
rect 5300 117 5370 203
rect 5400 117 5470 203
rect 5500 177 5570 203
rect 5500 143 5518 177
rect 5552 143 5570 177
rect 5500 117 5570 143
rect 5600 177 5670 203
rect 5600 143 5618 177
rect 5652 143 5670 177
rect 5600 117 5670 143
rect 5700 117 5770 203
rect 5800 177 5870 203
rect 5800 143 5818 177
rect 5852 143 5870 177
rect 5800 117 5870 143
rect 5900 177 5970 203
rect 5900 143 5918 177
rect 5952 143 5970 177
rect 5900 117 5970 143
rect 6000 177 6070 203
rect 6000 143 6018 177
rect 6052 143 6070 177
rect 6000 117 6070 143
rect 6100 177 6170 203
rect 6100 143 6118 177
rect 6152 143 6170 177
rect 6100 117 6170 143
rect 6200 177 6270 203
rect 6200 143 6218 177
rect 6252 143 6270 177
rect 6200 117 6270 143
rect 6300 177 6370 203
rect 6300 143 6318 177
rect 6352 143 6370 177
rect 6300 117 6370 143
rect 6400 177 6470 203
rect 6400 143 6418 177
rect 6452 143 6470 177
rect 6400 117 6470 143
rect 6500 117 6570 203
rect 6600 117 6670 203
rect 6700 117 6770 203
rect 6800 117 6870 203
rect 6900 177 6970 203
rect 6900 143 6918 177
rect 6952 143 6970 177
rect 6900 117 6970 143
rect 7000 177 7054 203
rect 7000 143 7012 177
rect 7046 143 7054 177
rect 7000 117 7054 143
rect 7916 317 7970 343
rect 7916 283 7924 317
rect 7958 283 7970 317
rect 7916 257 7970 283
rect 8000 317 8054 343
rect 8000 283 8012 317
rect 8046 283 8054 317
rect 8000 257 8054 283
rect 9216 737 9270 763
rect 9216 703 9224 737
rect 9258 703 9270 737
rect 9216 677 9270 703
rect 9300 737 9354 763
rect 9300 703 9312 737
rect 9346 703 9354 737
rect 9300 677 9354 703
rect 9416 737 9470 763
rect 9416 703 9424 737
rect 9458 703 9470 737
rect 9416 677 9470 703
rect 9500 737 9570 763
rect 9500 703 9518 737
rect 9552 703 9570 737
rect 9500 677 9570 703
rect 9600 737 9654 763
rect 9600 703 9612 737
rect 9646 703 9654 737
rect 9600 677 9654 703
rect 9716 737 9770 763
rect 9716 703 9724 737
rect 9758 703 9770 737
rect 9716 677 9770 703
rect 9800 737 9854 763
rect 9800 703 9812 737
rect 9846 703 9854 737
rect 9800 677 9854 703
rect 10016 1017 10070 1043
rect 10016 983 10024 1017
rect 10058 983 10070 1017
rect 10016 957 10070 983
rect 10100 1017 10170 1043
rect 10100 983 10118 1017
rect 10152 983 10170 1017
rect 10100 957 10170 983
rect 10200 1017 10270 1043
rect 10200 983 10218 1017
rect 10252 983 10270 1017
rect 10200 957 10270 983
rect 10300 1017 10354 1043
rect 10300 983 10312 1017
rect 10346 983 10354 1017
rect 10300 957 10354 983
rect 11116 1157 11170 1183
rect 11116 1123 11124 1157
rect 11158 1123 11170 1157
rect 11116 1097 11170 1123
rect 11200 1157 11254 1183
rect 11200 1123 11212 1157
rect 11246 1123 11254 1157
rect 11200 1097 11254 1123
rect 11316 1157 11370 1183
rect 11316 1123 11324 1157
rect 11358 1123 11370 1157
rect 11316 1097 11370 1123
rect 11400 1157 11454 1183
rect 11400 1123 11412 1157
rect 11446 1123 11454 1157
rect 11400 1097 11454 1123
rect 10416 1017 10470 1043
rect 10416 983 10424 1017
rect 10458 983 10470 1017
rect 10416 957 10470 983
rect 10500 1017 10570 1043
rect 10500 983 10518 1017
rect 10552 983 10570 1017
rect 10500 957 10570 983
rect 10600 957 10670 1043
rect 10700 957 10770 1043
rect 10800 1017 10870 1043
rect 10800 983 10818 1017
rect 10852 983 10870 1017
rect 10800 957 10870 983
rect 10900 1017 10970 1043
rect 10900 983 10918 1017
rect 10952 983 10970 1017
rect 10900 957 10970 983
rect 11000 1017 11070 1043
rect 11000 983 11018 1017
rect 11052 983 11070 1017
rect 11000 957 11070 983
rect 11100 1017 11170 1043
rect 11100 983 11118 1017
rect 11152 983 11170 1017
rect 11100 957 11170 983
rect 11200 1017 11270 1043
rect 11200 983 11218 1017
rect 11252 983 11270 1017
rect 11200 957 11270 983
rect 11300 1017 11354 1043
rect 11300 983 11312 1017
rect 11346 983 11354 1017
rect 11300 957 11354 983
rect 10016 877 10070 903
rect 10016 843 10024 877
rect 10058 843 10070 877
rect 10016 817 10070 843
rect 10100 877 10170 903
rect 10100 843 10118 877
rect 10152 843 10170 877
rect 10100 817 10170 843
rect 10200 817 10270 903
rect 10300 817 10370 903
rect 10400 817 10470 903
rect 10500 877 10570 903
rect 10500 843 10518 877
rect 10552 843 10570 877
rect 10500 817 10570 843
rect 10600 877 10670 903
rect 10600 843 10618 877
rect 10652 843 10670 877
rect 10600 817 10670 843
rect 10700 877 10754 903
rect 10700 843 10712 877
rect 10746 843 10754 877
rect 10700 817 10754 843
rect 9916 737 9970 763
rect 9916 703 9924 737
rect 9958 703 9970 737
rect 9916 677 9970 703
rect 10000 737 10070 763
rect 10000 703 10018 737
rect 10052 703 10070 737
rect 10000 677 10070 703
rect 10100 737 10154 763
rect 10100 703 10112 737
rect 10146 703 10154 737
rect 10100 677 10154 703
rect 10816 877 10870 903
rect 10816 843 10824 877
rect 10858 843 10870 877
rect 10816 817 10870 843
rect 10900 877 10954 903
rect 10900 843 10912 877
rect 10946 843 10954 877
rect 10900 817 10954 843
rect 10216 737 10270 763
rect 10216 703 10224 737
rect 10258 703 10270 737
rect 10216 677 10270 703
rect 10300 737 10370 763
rect 10300 703 10318 737
rect 10352 703 10370 737
rect 10300 677 10370 703
rect 10400 677 10470 763
rect 10500 677 10570 763
rect 10600 677 10670 763
rect 10700 737 10770 763
rect 10700 703 10718 737
rect 10752 703 10770 737
rect 10700 677 10770 703
rect 10800 737 10870 763
rect 10800 703 10818 737
rect 10852 703 10870 737
rect 10800 677 10870 703
rect 10900 737 10954 763
rect 10900 703 10912 737
rect 10946 703 10954 737
rect 10900 677 10954 703
rect 8416 597 8470 623
rect 8416 563 8424 597
rect 8458 563 8470 597
rect 8416 537 8470 563
rect 8500 597 8570 623
rect 8500 563 8518 597
rect 8552 563 8570 597
rect 8500 537 8570 563
rect 8600 537 8670 623
rect 8700 597 8770 623
rect 8700 563 8718 597
rect 8752 563 8770 597
rect 8700 537 8770 563
rect 8800 597 8870 623
rect 8800 563 8818 597
rect 8852 563 8870 597
rect 8800 537 8870 563
rect 8900 597 8970 623
rect 8900 563 8918 597
rect 8952 563 8970 597
rect 8900 537 8970 563
rect 9000 597 9070 623
rect 9000 563 9018 597
rect 9052 563 9070 597
rect 9000 537 9070 563
rect 9100 537 9170 623
rect 9200 597 9270 623
rect 9200 563 9218 597
rect 9252 563 9270 597
rect 9200 537 9270 563
rect 9300 597 9370 623
rect 9300 563 9318 597
rect 9352 563 9370 597
rect 9300 537 9370 563
rect 9400 537 9470 623
rect 9500 597 9570 623
rect 9500 563 9518 597
rect 9552 563 9570 597
rect 9500 537 9570 563
rect 9600 597 9670 623
rect 9600 563 9618 597
rect 9652 563 9670 597
rect 9600 537 9670 563
rect 9700 537 9770 623
rect 9800 537 9870 623
rect 9900 597 9970 623
rect 9900 563 9918 597
rect 9952 563 9970 597
rect 9900 537 9970 563
rect 10000 597 10070 623
rect 10000 563 10018 597
rect 10052 563 10070 597
rect 10000 537 10070 563
rect 10100 597 10170 623
rect 10100 563 10118 597
rect 10152 563 10170 597
rect 10100 537 10170 563
rect 10200 597 10254 623
rect 10200 563 10212 597
rect 10246 563 10254 597
rect 10200 537 10254 563
rect 8416 457 8470 483
rect 8416 423 8424 457
rect 8458 423 8470 457
rect 8416 397 8470 423
rect 8500 457 8570 483
rect 8500 423 8518 457
rect 8552 423 8570 457
rect 8500 397 8570 423
rect 8600 397 8670 483
rect 8700 457 8770 483
rect 8700 423 8718 457
rect 8752 423 8770 457
rect 8700 397 8770 423
rect 8800 457 8870 483
rect 8800 423 8818 457
rect 8852 423 8870 457
rect 8800 397 8870 423
rect 8900 457 8970 483
rect 8900 423 8918 457
rect 8952 423 8970 457
rect 8900 397 8970 423
rect 9000 457 9070 483
rect 9000 423 9018 457
rect 9052 423 9070 457
rect 9000 397 9070 423
rect 9100 457 9170 483
rect 9100 423 9118 457
rect 9152 423 9170 457
rect 9100 397 9170 423
rect 9200 457 9270 483
rect 9200 423 9218 457
rect 9252 423 9270 457
rect 9200 397 9270 423
rect 9300 397 9370 483
rect 9400 457 9470 483
rect 9400 423 9418 457
rect 9452 423 9470 457
rect 9400 397 9470 423
rect 9500 457 9570 483
rect 9500 423 9518 457
rect 9552 423 9570 457
rect 9500 397 9570 423
rect 9600 457 9670 483
rect 9600 423 9618 457
rect 9652 423 9670 457
rect 9600 397 9670 423
rect 9700 457 9770 483
rect 9700 423 9718 457
rect 9752 423 9770 457
rect 9700 397 9770 423
rect 9800 457 9870 483
rect 9800 423 9818 457
rect 9852 423 9870 457
rect 9800 397 9870 423
rect 9900 457 9954 483
rect 9900 423 9912 457
rect 9946 423 9954 457
rect 9900 397 9954 423
rect 8116 317 8170 343
rect 8116 283 8124 317
rect 8158 283 8170 317
rect 8116 257 8170 283
rect 8200 317 8270 343
rect 8200 283 8218 317
rect 8252 283 8270 317
rect 8200 257 8270 283
rect 8300 317 8370 343
rect 8300 283 8318 317
rect 8352 283 8370 317
rect 8300 257 8370 283
rect 8400 317 8470 343
rect 8400 283 8418 317
rect 8452 283 8470 317
rect 8400 257 8470 283
rect 8500 317 8570 343
rect 8500 283 8518 317
rect 8552 283 8570 317
rect 8500 257 8570 283
rect 8600 317 8670 343
rect 8600 283 8618 317
rect 8652 283 8670 317
rect 8600 257 8670 283
rect 8700 317 8754 343
rect 8700 283 8712 317
rect 8746 283 8754 317
rect 8700 257 8754 283
rect 8816 317 8870 343
rect 8816 283 8824 317
rect 8858 283 8870 317
rect 8816 257 8870 283
rect 8900 317 8970 343
rect 8900 283 8918 317
rect 8952 283 8970 317
rect 8900 257 8970 283
rect 9000 317 9054 343
rect 9000 283 9012 317
rect 9046 283 9054 317
rect 9000 257 9054 283
rect 9116 317 9170 343
rect 9116 283 9124 317
rect 9158 283 9170 317
rect 9116 257 9170 283
rect 9200 317 9254 343
rect 9200 283 9212 317
rect 9246 283 9254 317
rect 9200 257 9254 283
rect 10016 457 10070 483
rect 10016 423 10024 457
rect 10058 423 10070 457
rect 10016 397 10070 423
rect 10100 457 10170 483
rect 10100 423 10118 457
rect 10152 423 10170 457
rect 10100 397 10170 423
rect 10200 457 10254 483
rect 10200 423 10212 457
rect 10246 423 10254 457
rect 10200 397 10254 423
rect 9316 317 9370 343
rect 9316 283 9324 317
rect 9358 283 9370 317
rect 9316 257 9370 283
rect 9400 317 9470 343
rect 9400 283 9418 317
rect 9452 283 9470 317
rect 9400 257 9470 283
rect 9500 317 9570 343
rect 9500 283 9518 317
rect 9552 283 9570 317
rect 9500 257 9570 283
rect 9600 317 9670 343
rect 9600 283 9618 317
rect 9652 283 9670 317
rect 9600 257 9670 283
rect 9700 257 9770 343
rect 9800 257 9870 343
rect 9900 257 9970 343
rect 10000 317 10070 343
rect 10000 283 10018 317
rect 10052 283 10070 317
rect 10000 257 10070 283
rect 10100 317 10154 343
rect 10100 283 10112 317
rect 10146 283 10154 317
rect 10100 257 10154 283
rect 10316 597 10370 623
rect 10316 563 10324 597
rect 10358 563 10370 597
rect 10316 537 10370 563
rect 10400 597 10454 623
rect 10400 563 10412 597
rect 10446 563 10454 597
rect 10400 537 10454 563
rect 12116 1527 12170 1553
rect 12116 1493 12124 1527
rect 12158 1493 12170 1527
rect 12116 1467 12170 1493
rect 12200 1527 12270 1553
rect 12200 1493 12218 1527
rect 12252 1493 12270 1527
rect 12200 1467 12270 1493
rect 12300 1527 12370 1553
rect 12300 1493 12318 1527
rect 12352 1493 12370 1527
rect 12300 1467 12370 1493
rect 12400 1527 12454 1553
rect 12400 1493 12412 1527
rect 12446 1493 12454 1527
rect 12400 1467 12454 1493
rect 11816 1387 11870 1413
rect 11816 1353 11824 1387
rect 11858 1353 11870 1387
rect 11816 1327 11870 1353
rect 11900 1387 11970 1413
rect 11900 1353 11918 1387
rect 11952 1353 11970 1387
rect 11900 1327 11970 1353
rect 12000 1387 12070 1413
rect 12000 1353 12018 1387
rect 12052 1353 12070 1387
rect 12000 1327 12070 1353
rect 12100 1327 12170 1413
rect 12200 1327 12270 1413
rect 12300 1387 12370 1413
rect 12300 1353 12318 1387
rect 12352 1353 12370 1387
rect 12300 1327 12370 1353
rect 12400 1387 12454 1413
rect 12400 1353 12412 1387
rect 12446 1353 12454 1387
rect 12400 1327 12454 1353
rect 11516 1157 11570 1183
rect 11516 1123 11524 1157
rect 11558 1123 11570 1157
rect 11516 1097 11570 1123
rect 11600 1157 11670 1183
rect 11600 1123 11618 1157
rect 11652 1123 11670 1157
rect 11600 1097 11670 1123
rect 11700 1097 11770 1183
rect 11800 1097 11870 1183
rect 11900 1157 11970 1183
rect 11900 1123 11918 1157
rect 11952 1123 11970 1157
rect 11900 1097 11970 1123
rect 12000 1157 12054 1183
rect 12000 1123 12012 1157
rect 12046 1123 12054 1157
rect 12000 1097 12054 1123
rect 11416 1017 11470 1043
rect 11416 983 11424 1017
rect 11458 983 11470 1017
rect 11416 957 11470 983
rect 11500 1017 11570 1043
rect 11500 983 11518 1017
rect 11552 983 11570 1017
rect 11500 957 11570 983
rect 11600 1017 11654 1043
rect 11600 983 11612 1017
rect 11646 983 11654 1017
rect 11600 957 11654 983
rect 11716 1017 11770 1043
rect 11716 983 11724 1017
rect 11758 983 11770 1017
rect 11716 957 11770 983
rect 11800 1017 11870 1043
rect 11800 983 11818 1017
rect 11852 983 11870 1017
rect 11800 957 11870 983
rect 11900 1017 11954 1043
rect 11900 983 11912 1017
rect 11946 983 11954 1017
rect 11900 957 11954 983
rect 11016 877 11070 903
rect 11016 843 11024 877
rect 11058 843 11070 877
rect 11016 817 11070 843
rect 11100 877 11170 903
rect 11100 843 11118 877
rect 11152 843 11170 877
rect 11100 817 11170 843
rect 11200 877 11270 903
rect 11200 843 11218 877
rect 11252 843 11270 877
rect 11200 817 11270 843
rect 11300 877 11370 903
rect 11300 843 11318 877
rect 11352 843 11370 877
rect 11300 817 11370 843
rect 11400 817 11470 903
rect 11500 817 11570 903
rect 11600 817 11670 903
rect 11700 877 11770 903
rect 11700 843 11718 877
rect 11752 843 11770 877
rect 11700 817 11770 843
rect 11800 877 11870 903
rect 11800 843 11818 877
rect 11852 843 11870 877
rect 11800 817 11870 843
rect 11900 877 11954 903
rect 11900 843 11912 877
rect 11946 843 11954 877
rect 11900 817 11954 843
rect 11016 737 11070 763
rect 11016 703 11024 737
rect 11058 703 11070 737
rect 11016 677 11070 703
rect 11100 737 11170 763
rect 11100 703 11118 737
rect 11152 703 11170 737
rect 11100 677 11170 703
rect 11200 737 11270 763
rect 11200 703 11218 737
rect 11252 703 11270 737
rect 11200 677 11270 703
rect 11300 737 11370 763
rect 11300 703 11318 737
rect 11352 703 11370 737
rect 11300 677 11370 703
rect 11400 677 11470 763
rect 11500 737 11570 763
rect 11500 703 11518 737
rect 11552 703 11570 737
rect 11500 677 11570 703
rect 11600 737 11670 763
rect 11600 703 11618 737
rect 11652 703 11670 737
rect 11600 677 11670 703
rect 11700 737 11754 763
rect 11700 703 11712 737
rect 11746 703 11754 737
rect 11700 677 11754 703
rect 10516 597 10570 623
rect 10516 563 10524 597
rect 10558 563 10570 597
rect 10516 537 10570 563
rect 10600 597 10670 623
rect 10600 563 10618 597
rect 10652 563 10670 597
rect 10600 537 10670 563
rect 10700 597 10770 623
rect 10700 563 10718 597
rect 10752 563 10770 597
rect 10700 537 10770 563
rect 10800 597 10870 623
rect 10800 563 10818 597
rect 10852 563 10870 597
rect 10800 537 10870 563
rect 10900 537 10970 623
rect 11000 537 11070 623
rect 11100 597 11170 623
rect 11100 563 11118 597
rect 11152 563 11170 597
rect 11100 537 11170 563
rect 11200 597 11254 623
rect 11200 563 11212 597
rect 11246 563 11254 597
rect 11200 537 11254 563
rect 10316 457 10370 483
rect 10316 423 10324 457
rect 10358 423 10370 457
rect 10316 397 10370 423
rect 10400 457 10470 483
rect 10400 423 10418 457
rect 10452 423 10470 457
rect 10400 397 10470 423
rect 10500 457 10570 483
rect 10500 423 10518 457
rect 10552 423 10570 457
rect 10500 397 10570 423
rect 10600 457 10670 483
rect 10600 423 10618 457
rect 10652 423 10670 457
rect 10600 397 10670 423
rect 10700 457 10770 483
rect 10700 423 10718 457
rect 10752 423 10770 457
rect 10700 397 10770 423
rect 10800 457 10854 483
rect 10800 423 10812 457
rect 10846 423 10854 457
rect 10800 397 10854 423
rect 10916 457 10970 483
rect 10916 423 10924 457
rect 10958 423 10970 457
rect 10916 397 10970 423
rect 11000 457 11070 483
rect 11000 423 11018 457
rect 11052 423 11070 457
rect 11000 397 11070 423
rect 11100 457 11154 483
rect 11100 423 11112 457
rect 11146 423 11154 457
rect 11100 397 11154 423
rect 12516 1527 12570 1553
rect 12516 1493 12524 1527
rect 12558 1493 12570 1527
rect 12516 1467 12570 1493
rect 12600 1527 12670 1553
rect 12600 1493 12618 1527
rect 12652 1493 12670 1527
rect 12600 1467 12670 1493
rect 12700 1527 12770 1553
rect 12700 1493 12718 1527
rect 12752 1493 12770 1527
rect 12700 1467 12770 1493
rect 12800 1467 12854 1553
rect 12912 1542 12970 1553
rect 12912 1508 12924 1542
rect 12958 1508 12970 1542
rect 12912 1467 12970 1508
rect 13000 1527 13070 1553
rect 13000 1493 13018 1527
rect 13052 1493 13070 1527
rect 13000 1467 13070 1493
rect 13100 1512 13158 1553
rect 13100 1478 13112 1512
rect 13146 1478 13158 1512
rect 13100 1467 13158 1478
rect 13220 1527 13280 1553
rect 13220 1493 13228 1527
rect 13262 1493 13280 1527
rect 13220 1467 13280 1493
rect 13310 1527 13380 1553
rect 13310 1493 13328 1527
rect 13362 1493 13380 1527
rect 13310 1467 13380 1493
rect 13410 1527 13480 1553
rect 13410 1493 13428 1527
rect 13462 1493 13480 1527
rect 13410 1467 13480 1493
rect 13510 1527 13580 1553
rect 13510 1493 13528 1527
rect 13562 1493 13580 1527
rect 13510 1467 13580 1493
rect 13610 1527 13670 1553
rect 13610 1493 13628 1527
rect 13662 1493 13670 1527
rect 13610 1467 13670 1493
rect 12516 1387 12570 1413
rect 12516 1353 12524 1387
rect 12558 1353 12570 1387
rect 12516 1327 12570 1353
rect 12600 1387 12670 1413
rect 12600 1353 12618 1387
rect 12652 1353 12670 1387
rect 12600 1327 12670 1353
rect 12700 1327 12770 1413
rect 12800 1327 12854 1413
rect 12912 1402 12970 1413
rect 12912 1368 12924 1402
rect 12958 1368 12970 1402
rect 12912 1327 12970 1368
rect 13000 1387 13070 1413
rect 13000 1353 13018 1387
rect 13052 1353 13070 1387
rect 13000 1327 13070 1353
rect 13100 1372 13158 1413
rect 13100 1338 13112 1372
rect 13146 1338 13158 1372
rect 13100 1327 13158 1338
rect 13220 1387 13280 1413
rect 13220 1353 13228 1387
rect 13262 1353 13280 1387
rect 13220 1327 13280 1353
rect 13310 1387 13380 1413
rect 13310 1353 13328 1387
rect 13362 1353 13380 1387
rect 13310 1327 13380 1353
rect 13410 1387 13480 1413
rect 13410 1353 13428 1387
rect 13462 1353 13480 1387
rect 13410 1327 13480 1353
rect 13510 1387 13580 1413
rect 13510 1353 13528 1387
rect 13562 1353 13580 1387
rect 13510 1327 13580 1353
rect 13610 1387 13670 1413
rect 13610 1353 13628 1387
rect 13662 1353 13670 1387
rect 13610 1327 13670 1353
rect 12116 1157 12170 1183
rect 12116 1123 12124 1157
rect 12158 1123 12170 1157
rect 12116 1097 12170 1123
rect 12200 1157 12270 1183
rect 12200 1123 12218 1157
rect 12252 1123 12270 1157
rect 12200 1097 12270 1123
rect 12300 1097 12370 1183
rect 12400 1097 12470 1183
rect 12500 1157 12570 1183
rect 12500 1123 12518 1157
rect 12552 1123 12570 1157
rect 12500 1097 12570 1123
rect 12600 1157 12654 1183
rect 12600 1123 12612 1157
rect 12646 1123 12654 1157
rect 12600 1097 12654 1123
rect 12716 1157 12770 1183
rect 12716 1123 12724 1157
rect 12758 1123 12770 1157
rect 12716 1097 12770 1123
rect 12800 1157 12854 1183
rect 12800 1123 12812 1157
rect 12846 1123 12854 1157
rect 12800 1097 12854 1123
rect 12912 1172 12970 1183
rect 12912 1138 12924 1172
rect 12958 1138 12970 1172
rect 12912 1097 12970 1138
rect 13000 1157 13070 1183
rect 13000 1123 13018 1157
rect 13052 1123 13070 1157
rect 13000 1097 13070 1123
rect 13100 1142 13158 1183
rect 13100 1108 13112 1142
rect 13146 1108 13158 1142
rect 13100 1097 13158 1108
rect 13220 1157 13280 1183
rect 13220 1123 13228 1157
rect 13262 1123 13280 1157
rect 13220 1097 13280 1123
rect 13310 1157 13380 1183
rect 13310 1123 13328 1157
rect 13362 1123 13380 1157
rect 13310 1097 13380 1123
rect 13410 1157 13480 1183
rect 13410 1123 13428 1157
rect 13462 1123 13480 1157
rect 13410 1097 13480 1123
rect 13510 1157 13580 1183
rect 13510 1123 13528 1157
rect 13562 1123 13580 1157
rect 13510 1097 13580 1123
rect 13610 1157 13670 1183
rect 13610 1123 13628 1157
rect 13662 1123 13670 1157
rect 13610 1097 13670 1123
rect 12016 1017 12070 1043
rect 12016 983 12024 1017
rect 12058 983 12070 1017
rect 12016 957 12070 983
rect 12100 1017 12170 1043
rect 12100 983 12118 1017
rect 12152 983 12170 1017
rect 12100 957 12170 983
rect 12200 1017 12270 1043
rect 12200 983 12218 1017
rect 12252 983 12270 1017
rect 12200 957 12270 983
rect 12300 957 12370 1043
rect 12400 957 12470 1043
rect 12500 957 12570 1043
rect 12600 1017 12670 1043
rect 12600 983 12618 1017
rect 12652 983 12670 1017
rect 12600 957 12670 983
rect 12700 1017 12770 1043
rect 12700 983 12718 1017
rect 12752 983 12770 1017
rect 12700 957 12770 983
rect 12800 1017 12854 1043
rect 12800 983 12812 1017
rect 12846 983 12854 1017
rect 12800 957 12854 983
rect 12912 1032 12970 1043
rect 12912 998 12924 1032
rect 12958 998 12970 1032
rect 12912 957 12970 998
rect 13000 1017 13070 1043
rect 13000 983 13018 1017
rect 13052 983 13070 1017
rect 13000 957 13070 983
rect 13100 1002 13158 1043
rect 13100 968 13112 1002
rect 13146 968 13158 1002
rect 13100 957 13158 968
rect 13220 1017 13280 1043
rect 13220 983 13228 1017
rect 13262 983 13280 1017
rect 13220 957 13280 983
rect 13310 1017 13380 1043
rect 13310 983 13328 1017
rect 13362 983 13380 1017
rect 13310 957 13380 983
rect 13410 1017 13480 1043
rect 13410 983 13428 1017
rect 13462 983 13480 1017
rect 13410 957 13480 983
rect 13510 1017 13580 1043
rect 13510 983 13528 1017
rect 13562 983 13580 1017
rect 13510 957 13580 983
rect 13610 1017 13670 1043
rect 13610 983 13628 1017
rect 13662 983 13670 1017
rect 13610 957 13670 983
rect 12016 877 12070 903
rect 12016 843 12024 877
rect 12058 843 12070 877
rect 12016 817 12070 843
rect 12100 877 12170 903
rect 12100 843 12118 877
rect 12152 843 12170 877
rect 12100 817 12170 843
rect 12200 877 12270 903
rect 12200 843 12218 877
rect 12252 843 12270 877
rect 12200 817 12270 843
rect 12300 877 12354 903
rect 12300 843 12312 877
rect 12346 843 12354 877
rect 12300 817 12354 843
rect 11816 737 11870 763
rect 11816 703 11824 737
rect 11858 703 11870 737
rect 11816 677 11870 703
rect 11900 737 11970 763
rect 11900 703 11918 737
rect 11952 703 11970 737
rect 11900 677 11970 703
rect 12000 737 12070 763
rect 12000 703 12018 737
rect 12052 703 12070 737
rect 12000 677 12070 703
rect 12100 737 12154 763
rect 12100 703 12112 737
rect 12146 703 12154 737
rect 12100 677 12154 703
rect 12416 877 12470 903
rect 12416 843 12424 877
rect 12458 843 12470 877
rect 12416 817 12470 843
rect 12500 877 12554 903
rect 12500 843 12512 877
rect 12546 843 12554 877
rect 12500 817 12554 843
rect 12616 877 12670 903
rect 12616 843 12624 877
rect 12658 843 12670 877
rect 12616 817 12670 843
rect 12700 877 12770 903
rect 12700 843 12718 877
rect 12752 843 12770 877
rect 12700 817 12770 843
rect 12800 817 12854 903
rect 12912 892 12970 903
rect 12912 858 12924 892
rect 12958 858 12970 892
rect 12912 817 12970 858
rect 13000 877 13070 903
rect 13000 843 13018 877
rect 13052 843 13070 877
rect 13000 817 13070 843
rect 13100 862 13158 903
rect 13100 828 13112 862
rect 13146 828 13158 862
rect 13100 817 13158 828
rect 13220 877 13280 903
rect 13220 843 13228 877
rect 13262 843 13280 877
rect 13220 817 13280 843
rect 13310 877 13380 903
rect 13310 843 13328 877
rect 13362 843 13380 877
rect 13310 817 13380 843
rect 13410 877 13480 903
rect 13410 843 13428 877
rect 13462 843 13480 877
rect 13410 817 13480 843
rect 13510 877 13580 903
rect 13510 843 13528 877
rect 13562 843 13580 877
rect 13510 817 13580 843
rect 13610 877 13670 903
rect 13610 843 13628 877
rect 13662 843 13670 877
rect 13610 817 13670 843
rect 12216 737 12270 763
rect 12216 703 12224 737
rect 12258 703 12270 737
rect 12216 677 12270 703
rect 12300 737 12370 763
rect 12300 703 12318 737
rect 12352 703 12370 737
rect 12300 677 12370 703
rect 12400 677 12470 763
rect 12500 737 12570 763
rect 12500 703 12518 737
rect 12552 703 12570 737
rect 12500 677 12570 703
rect 12600 737 12670 763
rect 12600 703 12618 737
rect 12652 703 12670 737
rect 12600 677 12670 703
rect 12700 677 12770 763
rect 12800 677 12854 763
rect 12912 752 12970 763
rect 12912 718 12924 752
rect 12958 718 12970 752
rect 12912 677 12970 718
rect 13000 737 13070 763
rect 13000 703 13018 737
rect 13052 703 13070 737
rect 13000 677 13070 703
rect 13100 722 13158 763
rect 13100 688 13112 722
rect 13146 688 13158 722
rect 13100 677 13158 688
rect 13220 737 13280 763
rect 13220 703 13228 737
rect 13262 703 13280 737
rect 13220 677 13280 703
rect 13310 737 13380 763
rect 13310 703 13328 737
rect 13362 703 13380 737
rect 13310 677 13380 703
rect 13410 737 13480 763
rect 13410 703 13428 737
rect 13462 703 13480 737
rect 13410 677 13480 703
rect 13510 737 13580 763
rect 13510 703 13528 737
rect 13562 703 13580 737
rect 13510 677 13580 703
rect 13610 737 13670 763
rect 13610 703 13628 737
rect 13662 703 13670 737
rect 13610 677 13670 703
rect 11316 597 11370 623
rect 11316 563 11324 597
rect 11358 563 11370 597
rect 11316 537 11370 563
rect 11400 597 11470 623
rect 11400 563 11418 597
rect 11452 563 11470 597
rect 11400 537 11470 563
rect 11500 597 11570 623
rect 11500 563 11518 597
rect 11552 563 11570 597
rect 11500 537 11570 563
rect 11600 597 11670 623
rect 11600 563 11618 597
rect 11652 563 11670 597
rect 11600 537 11670 563
rect 11700 597 11770 623
rect 11700 563 11718 597
rect 11752 563 11770 597
rect 11700 537 11770 563
rect 11800 597 11870 623
rect 11800 563 11818 597
rect 11852 563 11870 597
rect 11800 537 11870 563
rect 11900 597 11970 623
rect 11900 563 11918 597
rect 11952 563 11970 597
rect 11900 537 11970 563
rect 12000 537 12070 623
rect 12100 597 12170 623
rect 12100 563 12118 597
rect 12152 563 12170 597
rect 12100 537 12170 563
rect 12200 597 12270 623
rect 12200 563 12218 597
rect 12252 563 12270 597
rect 12200 537 12270 563
rect 12300 597 12370 623
rect 12300 563 12318 597
rect 12352 563 12370 597
rect 12300 537 12370 563
rect 12400 597 12470 623
rect 12400 563 12418 597
rect 12452 563 12470 597
rect 12400 537 12470 563
rect 12500 597 12570 623
rect 12500 563 12518 597
rect 12552 563 12570 597
rect 12500 537 12570 563
rect 12600 597 12670 623
rect 12600 563 12618 597
rect 12652 563 12670 597
rect 12600 537 12670 563
rect 12700 597 12770 623
rect 12700 563 12718 597
rect 12752 563 12770 597
rect 12700 537 12770 563
rect 12800 597 12854 623
rect 12800 563 12812 597
rect 12846 563 12854 597
rect 12800 537 12854 563
rect 12912 612 12970 623
rect 12912 578 12924 612
rect 12958 578 12970 612
rect 12912 537 12970 578
rect 13000 597 13070 623
rect 13000 563 13018 597
rect 13052 563 13070 597
rect 13000 537 13070 563
rect 13100 582 13158 623
rect 13100 548 13112 582
rect 13146 548 13158 582
rect 13100 537 13158 548
rect 13220 597 13280 623
rect 13220 563 13228 597
rect 13262 563 13280 597
rect 13220 537 13280 563
rect 13310 597 13380 623
rect 13310 563 13328 597
rect 13362 563 13380 597
rect 13310 537 13380 563
rect 13410 597 13480 623
rect 13410 563 13428 597
rect 13462 563 13480 597
rect 13410 537 13480 563
rect 13510 597 13580 623
rect 13510 563 13528 597
rect 13562 563 13580 597
rect 13510 537 13580 563
rect 13610 597 13670 623
rect 13610 563 13628 597
rect 13662 563 13670 597
rect 13610 537 13670 563
rect 11216 457 11270 483
rect 11216 423 11224 457
rect 11258 423 11270 457
rect 11216 397 11270 423
rect 11300 457 11354 483
rect 11300 423 11312 457
rect 11346 423 11354 457
rect 11300 397 11354 423
rect 11416 457 11470 483
rect 11416 423 11424 457
rect 11458 423 11470 457
rect 11416 397 11470 423
rect 11500 457 11570 483
rect 11500 423 11518 457
rect 11552 423 11570 457
rect 11500 397 11570 423
rect 11600 397 11670 483
rect 11700 397 11770 483
rect 11800 397 11870 483
rect 11900 397 11970 483
rect 12000 457 12070 483
rect 12000 423 12018 457
rect 12052 423 12070 457
rect 12000 397 12070 423
rect 12100 457 12170 483
rect 12100 423 12118 457
rect 12152 423 12170 457
rect 12100 397 12170 423
rect 12200 457 12270 483
rect 12200 423 12218 457
rect 12252 423 12270 457
rect 12200 397 12270 423
rect 12300 457 12354 483
rect 12300 423 12312 457
rect 12346 423 12354 457
rect 12300 397 12354 423
rect 10216 317 10270 343
rect 10216 283 10224 317
rect 10258 283 10270 317
rect 10216 257 10270 283
rect 10300 317 10370 343
rect 10300 283 10318 317
rect 10352 283 10370 317
rect 10300 257 10370 283
rect 10400 317 10470 343
rect 10400 283 10418 317
rect 10452 283 10470 317
rect 10400 257 10470 283
rect 10500 257 10570 343
rect 10600 257 10670 343
rect 10700 317 10770 343
rect 10700 283 10718 317
rect 10752 283 10770 317
rect 10700 257 10770 283
rect 10800 317 10870 343
rect 10800 283 10818 317
rect 10852 283 10870 317
rect 10800 257 10870 283
rect 10900 317 10970 343
rect 10900 283 10918 317
rect 10952 283 10970 317
rect 10900 257 10970 283
rect 11000 257 11070 343
rect 11100 257 11170 343
rect 11200 257 11270 343
rect 11300 317 11370 343
rect 11300 283 11318 317
rect 11352 283 11370 317
rect 11300 257 11370 283
rect 11400 317 11454 343
rect 11400 283 11412 317
rect 11446 283 11454 317
rect 11400 257 11454 283
rect 7116 177 7170 203
rect 7116 143 7124 177
rect 7158 143 7170 177
rect 7116 117 7170 143
rect 7200 177 7270 203
rect 7200 143 7218 177
rect 7252 143 7270 177
rect 7200 117 7270 143
rect 7300 177 7370 203
rect 7300 143 7318 177
rect 7352 143 7370 177
rect 7300 117 7370 143
rect 7400 117 7470 203
rect 7500 117 7570 203
rect 7600 177 7670 203
rect 7600 143 7618 177
rect 7652 143 7670 177
rect 7600 117 7670 143
rect 7700 177 7770 203
rect 7700 143 7718 177
rect 7752 143 7770 177
rect 7700 117 7770 143
rect 7800 117 7870 203
rect 7900 177 7970 203
rect 7900 143 7918 177
rect 7952 143 7970 177
rect 7900 117 7970 143
rect 8000 177 8070 203
rect 8000 143 8018 177
rect 8052 143 8070 177
rect 8000 117 8070 143
rect 8100 117 8170 203
rect 8200 117 8270 203
rect 8300 177 8370 203
rect 8300 143 8318 177
rect 8352 143 8370 177
rect 8300 117 8370 143
rect 8400 177 8470 203
rect 8400 143 8418 177
rect 8452 143 8470 177
rect 8400 117 8470 143
rect 8500 117 8570 203
rect 8600 117 8670 203
rect 8700 177 8770 203
rect 8700 143 8718 177
rect 8752 143 8770 177
rect 8700 117 8770 143
rect 8800 177 8870 203
rect 8800 143 8818 177
rect 8852 143 8870 177
rect 8800 117 8870 143
rect 8900 177 8970 203
rect 8900 143 8918 177
rect 8952 143 8970 177
rect 8900 117 8970 143
rect 9000 177 9070 203
rect 9000 143 9018 177
rect 9052 143 9070 177
rect 9000 117 9070 143
rect 9100 177 9170 203
rect 9100 143 9118 177
rect 9152 143 9170 177
rect 9100 117 9170 143
rect 9200 117 9270 203
rect 9300 177 9370 203
rect 9300 143 9318 177
rect 9352 143 9370 177
rect 9300 117 9370 143
rect 9400 177 9470 203
rect 9400 143 9418 177
rect 9452 143 9470 177
rect 9400 117 9470 143
rect 9500 117 9570 203
rect 9600 177 9670 203
rect 9600 143 9618 177
rect 9652 143 9670 177
rect 9600 117 9670 143
rect 9700 177 9770 203
rect 9700 143 9718 177
rect 9752 143 9770 177
rect 9700 117 9770 143
rect 9800 177 9870 203
rect 9800 143 9818 177
rect 9852 143 9870 177
rect 9800 117 9870 143
rect 9900 177 9970 203
rect 9900 143 9918 177
rect 9952 143 9970 177
rect 9900 117 9970 143
rect 10000 177 10070 203
rect 10000 143 10018 177
rect 10052 143 10070 177
rect 10000 117 10070 143
rect 10100 177 10170 203
rect 10100 143 10118 177
rect 10152 143 10170 177
rect 10100 117 10170 143
rect 10200 177 10270 203
rect 10200 143 10218 177
rect 10252 143 10270 177
rect 10200 117 10270 143
rect 10300 117 10370 203
rect 10400 117 10470 203
rect 10500 117 10570 203
rect 10600 177 10670 203
rect 10600 143 10618 177
rect 10652 143 10670 177
rect 10600 117 10670 143
rect 10700 177 10770 203
rect 10700 143 10718 177
rect 10752 143 10770 177
rect 10700 117 10770 143
rect 10800 117 10870 203
rect 10900 177 10970 203
rect 10900 143 10918 177
rect 10952 143 10970 177
rect 10900 117 10970 143
rect 11000 177 11070 203
rect 11000 143 11018 177
rect 11052 143 11070 177
rect 11000 117 11070 143
rect 11100 177 11170 203
rect 11100 143 11118 177
rect 11152 143 11170 177
rect 11100 117 11170 143
rect 11200 117 11270 203
rect 11300 177 11370 203
rect 11300 143 11318 177
rect 11352 143 11370 177
rect 11300 117 11370 143
rect 11400 177 11454 203
rect 11400 143 11412 177
rect 11446 143 11454 177
rect 11400 117 11454 143
rect 11516 317 11570 343
rect 11516 283 11524 317
rect 11558 283 11570 317
rect 11516 257 11570 283
rect 11600 317 11670 343
rect 11600 283 11618 317
rect 11652 283 11670 317
rect 11600 257 11670 283
rect 11700 317 11770 343
rect 11700 283 11718 317
rect 11752 283 11770 317
rect 11700 257 11770 283
rect 11800 317 11870 343
rect 11800 283 11818 317
rect 11852 283 11870 317
rect 11800 257 11870 283
rect 11900 257 11970 343
rect 12000 317 12070 343
rect 12000 283 12018 317
rect 12052 283 12070 317
rect 12000 257 12070 283
rect 12100 317 12170 343
rect 12100 283 12118 317
rect 12152 283 12170 317
rect 12100 257 12170 283
rect 12200 317 12254 343
rect 12200 283 12212 317
rect 12246 283 12254 317
rect 12200 257 12254 283
rect 12416 457 12470 483
rect 12416 423 12424 457
rect 12458 423 12470 457
rect 12416 397 12470 423
rect 12500 457 12570 483
rect 12500 423 12518 457
rect 12552 423 12570 457
rect 12500 397 12570 423
rect 12600 397 12670 483
rect 12700 457 12770 483
rect 12700 423 12718 457
rect 12752 423 12770 457
rect 12700 397 12770 423
rect 12800 457 12854 483
rect 12800 423 12812 457
rect 12846 423 12854 457
rect 12800 397 12854 423
rect 12912 472 12970 483
rect 12912 438 12924 472
rect 12958 438 12970 472
rect 12912 397 12970 438
rect 13000 457 13070 483
rect 13000 423 13018 457
rect 13052 423 13070 457
rect 13000 397 13070 423
rect 13100 442 13158 483
rect 13100 408 13112 442
rect 13146 408 13158 442
rect 13100 397 13158 408
rect 13220 457 13280 483
rect 13220 423 13228 457
rect 13262 423 13280 457
rect 13220 397 13280 423
rect 13310 457 13380 483
rect 13310 423 13328 457
rect 13362 423 13380 457
rect 13310 397 13380 423
rect 13410 457 13480 483
rect 13410 423 13428 457
rect 13462 423 13480 457
rect 13410 397 13480 423
rect 13510 457 13580 483
rect 13510 423 13528 457
rect 13562 423 13580 457
rect 13510 397 13580 423
rect 13610 457 13670 483
rect 13610 423 13628 457
rect 13662 423 13670 457
rect 13610 397 13670 423
rect 12316 317 12370 343
rect 12316 283 12324 317
rect 12358 283 12370 317
rect 12316 257 12370 283
rect 12400 317 12470 343
rect 12400 283 12418 317
rect 12452 283 12470 317
rect 12400 257 12470 283
rect 12500 317 12570 343
rect 12500 283 12518 317
rect 12552 283 12570 317
rect 12500 257 12570 283
rect 12600 317 12670 343
rect 12600 283 12618 317
rect 12652 283 12670 317
rect 12600 257 12670 283
rect 12700 257 12770 343
rect 12800 257 12854 343
rect 12912 332 12970 343
rect 12912 298 12924 332
rect 12958 298 12970 332
rect 12912 257 12970 298
rect 13000 317 13070 343
rect 13000 283 13018 317
rect 13052 283 13070 317
rect 13000 257 13070 283
rect 13100 302 13158 343
rect 13100 268 13112 302
rect 13146 268 13158 302
rect 13100 257 13158 268
rect 13220 317 13280 343
rect 13220 283 13228 317
rect 13262 283 13280 317
rect 13220 257 13280 283
rect 13310 317 13380 343
rect 13310 283 13328 317
rect 13362 283 13380 317
rect 13310 257 13380 283
rect 13410 317 13480 343
rect 13410 283 13428 317
rect 13462 283 13480 317
rect 13410 257 13480 283
rect 13510 317 13580 343
rect 13510 283 13528 317
rect 13562 283 13580 317
rect 13510 257 13580 283
rect 13610 317 13670 343
rect 13610 283 13628 317
rect 13662 283 13670 317
rect 13610 257 13670 283
rect 11516 177 11570 203
rect 11516 143 11524 177
rect 11558 143 11570 177
rect 11516 117 11570 143
rect 11600 177 11670 203
rect 11600 143 11618 177
rect 11652 143 11670 177
rect 11600 117 11670 143
rect 11700 117 11770 203
rect 11800 177 11870 203
rect 11800 143 11818 177
rect 11852 143 11870 177
rect 11800 117 11870 143
rect 11900 177 11970 203
rect 11900 143 11918 177
rect 11952 143 11970 177
rect 11900 117 11970 143
rect 12000 177 12070 203
rect 12000 143 12018 177
rect 12052 143 12070 177
rect 12000 117 12070 143
rect 12100 177 12170 203
rect 12100 143 12118 177
rect 12152 143 12170 177
rect 12100 117 12170 143
rect 12200 117 12270 203
rect 12300 117 12370 203
rect 12400 177 12470 203
rect 12400 143 12418 177
rect 12452 143 12470 177
rect 12400 117 12470 143
rect 12500 177 12570 203
rect 12500 143 12518 177
rect 12552 143 12570 177
rect 12500 117 12570 143
rect 12600 177 12670 203
rect 12600 143 12618 177
rect 12652 143 12670 177
rect 12600 117 12670 143
rect 12700 177 12770 203
rect 12700 143 12718 177
rect 12752 143 12770 177
rect 12700 117 12770 143
rect 12800 117 12854 203
rect 12912 192 12970 203
rect 12912 158 12924 192
rect 12958 158 12970 192
rect 12912 117 12970 158
rect 13000 177 13070 203
rect 13000 143 13018 177
rect 13052 143 13070 177
rect 13000 117 13070 143
rect 13100 162 13158 203
rect 13100 128 13112 162
rect 13146 128 13158 162
rect 13100 117 13158 128
rect 13220 177 13280 203
rect 13220 143 13228 177
rect 13262 143 13280 177
rect 13220 117 13280 143
rect 13310 177 13380 203
rect 13310 143 13328 177
rect 13362 143 13380 177
rect 13310 117 13380 143
rect 13410 177 13480 203
rect 13410 143 13428 177
rect 13462 143 13480 177
rect 13410 117 13480 143
rect 13510 177 13580 203
rect 13510 143 13528 177
rect 13562 143 13580 177
rect 13510 117 13580 143
rect 13610 177 13670 203
rect 13610 143 13628 177
rect 13662 143 13670 177
rect 13610 117 13670 143
rect -94 -149 -30 -126
rect -94 -183 -82 -149
rect -48 -183 -30 -149
rect -94 -210 -30 -183
rect 0 -149 70 -126
rect 0 -183 18 -149
rect 52 -183 70 -149
rect 0 -210 70 -183
rect 100 -149 170 -126
rect 100 -183 118 -149
rect 152 -183 170 -149
rect 100 -210 170 -183
rect 200 -149 270 -126
rect 200 -183 218 -149
rect 252 -183 270 -149
rect 200 -210 270 -183
rect 300 -149 370 -126
rect 300 -183 318 -149
rect 352 -183 370 -149
rect 300 -210 370 -183
rect 400 -149 470 -126
rect 400 -183 418 -149
rect 452 -183 470 -149
rect 400 -210 470 -183
rect 500 -149 570 -126
rect 500 -183 518 -149
rect 552 -183 570 -149
rect 500 -210 570 -183
rect 600 -149 670 -126
rect 600 -183 618 -149
rect 652 -183 670 -149
rect 600 -210 670 -183
rect 700 -149 770 -126
rect 700 -183 718 -149
rect 752 -183 770 -149
rect 700 -210 770 -183
rect 800 -149 870 -126
rect 800 -183 818 -149
rect 852 -183 870 -149
rect 800 -210 870 -183
rect 900 -149 970 -126
rect 900 -183 918 -149
rect 952 -183 970 -149
rect 900 -210 970 -183
rect 1000 -149 1070 -126
rect 1000 -183 1018 -149
rect 1052 -183 1070 -149
rect 1000 -210 1070 -183
rect 1100 -149 1170 -126
rect 1100 -183 1118 -149
rect 1152 -183 1170 -149
rect 1100 -210 1170 -183
rect 1200 -149 1270 -126
rect 1200 -183 1218 -149
rect 1252 -183 1270 -149
rect 1200 -210 1270 -183
rect 1300 -149 1370 -126
rect 1300 -183 1318 -149
rect 1352 -183 1370 -149
rect 1300 -210 1370 -183
rect 1400 -149 1470 -126
rect 1400 -183 1418 -149
rect 1452 -183 1470 -149
rect 1400 -210 1470 -183
rect 1500 -149 1570 -126
rect 1500 -183 1518 -149
rect 1552 -183 1570 -149
rect 1500 -210 1570 -183
rect 1600 -149 1670 -126
rect 1600 -183 1618 -149
rect 1652 -183 1670 -149
rect 1600 -210 1670 -183
rect 1700 -149 1770 -126
rect 1700 -183 1718 -149
rect 1752 -183 1770 -149
rect 1700 -210 1770 -183
rect 1800 -149 1870 -126
rect 1800 -183 1818 -149
rect 1852 -183 1870 -149
rect 1800 -210 1870 -183
rect 1900 -149 1970 -126
rect 1900 -183 1918 -149
rect 1952 -183 1970 -149
rect 1900 -210 1970 -183
rect 2000 -149 2070 -126
rect 2000 -183 2018 -149
rect 2052 -183 2070 -149
rect 2000 -210 2070 -183
rect 2100 -149 2170 -126
rect 2100 -183 2118 -149
rect 2152 -183 2170 -149
rect 2100 -210 2170 -183
rect 2200 -149 2270 -126
rect 2200 -183 2218 -149
rect 2252 -183 2270 -149
rect 2200 -210 2270 -183
rect 2300 -149 2370 -126
rect 2300 -183 2318 -149
rect 2352 -183 2370 -149
rect 2300 -210 2370 -183
rect 2400 -149 2470 -126
rect 2400 -183 2418 -149
rect 2452 -183 2470 -149
rect 2400 -210 2470 -183
rect 2500 -149 2570 -126
rect 2500 -183 2518 -149
rect 2552 -183 2570 -149
rect 2500 -210 2570 -183
rect 2600 -149 2670 -126
rect 2600 -183 2618 -149
rect 2652 -183 2670 -149
rect 2600 -210 2670 -183
rect 2700 -149 2770 -126
rect 2700 -183 2718 -149
rect 2752 -183 2770 -149
rect 2700 -210 2770 -183
rect 2800 -149 2870 -126
rect 2800 -183 2818 -149
rect 2852 -183 2870 -149
rect 2800 -210 2870 -183
rect 2900 -149 2970 -126
rect 2900 -183 2918 -149
rect 2952 -183 2970 -149
rect 2900 -210 2970 -183
rect 3000 -149 3070 -126
rect 3000 -183 3018 -149
rect 3052 -183 3070 -149
rect 3000 -210 3070 -183
rect 3100 -149 3170 -126
rect 3100 -183 3118 -149
rect 3152 -183 3170 -149
rect 3100 -210 3170 -183
rect 3200 -149 3270 -126
rect 3200 -183 3218 -149
rect 3252 -183 3270 -149
rect 3200 -210 3270 -183
rect 3300 -149 3370 -126
rect 3300 -183 3318 -149
rect 3352 -183 3370 -149
rect 3300 -210 3370 -183
rect 3400 -149 3470 -126
rect 3400 -183 3418 -149
rect 3452 -183 3470 -149
rect 3400 -210 3470 -183
rect 3500 -149 3570 -126
rect 3500 -183 3518 -149
rect 3552 -183 3570 -149
rect 3500 -210 3570 -183
rect 3600 -149 3670 -126
rect 3600 -183 3618 -149
rect 3652 -183 3670 -149
rect 3600 -210 3670 -183
rect 3700 -149 3770 -126
rect 3700 -183 3718 -149
rect 3752 -183 3770 -149
rect 3700 -210 3770 -183
rect 3800 -149 3870 -126
rect 3800 -183 3818 -149
rect 3852 -183 3870 -149
rect 3800 -210 3870 -183
rect 3900 -149 3970 -126
rect 3900 -183 3918 -149
rect 3952 -183 3970 -149
rect 3900 -210 3970 -183
rect 4000 -149 4070 -126
rect 4000 -183 4018 -149
rect 4052 -183 4070 -149
rect 4000 -210 4070 -183
rect 4100 -149 4170 -126
rect 4100 -183 4118 -149
rect 4152 -183 4170 -149
rect 4100 -210 4170 -183
rect 4200 -149 4270 -126
rect 4200 -183 4218 -149
rect 4252 -183 4270 -149
rect 4200 -210 4270 -183
rect 4300 -149 4370 -126
rect 4300 -183 4318 -149
rect 4352 -183 4370 -149
rect 4300 -210 4370 -183
rect 4400 -149 4470 -126
rect 4400 -183 4418 -149
rect 4452 -183 4470 -149
rect 4400 -210 4470 -183
rect 4500 -149 4570 -126
rect 4500 -183 4518 -149
rect 4552 -183 4570 -149
rect 4500 -210 4570 -183
rect 4600 -149 4670 -126
rect 4600 -183 4618 -149
rect 4652 -183 4670 -149
rect 4600 -210 4670 -183
rect 4700 -149 4770 -126
rect 4700 -183 4718 -149
rect 4752 -183 4770 -149
rect 4700 -210 4770 -183
rect 4800 -149 4870 -126
rect 4800 -183 4818 -149
rect 4852 -183 4870 -149
rect 4800 -210 4870 -183
rect 4900 -149 4970 -126
rect 4900 -183 4918 -149
rect 4952 -183 4970 -149
rect 4900 -210 4970 -183
rect 5000 -149 5070 -126
rect 5000 -183 5018 -149
rect 5052 -183 5070 -149
rect 5000 -210 5070 -183
rect 5100 -149 5170 -126
rect 5100 -183 5118 -149
rect 5152 -183 5170 -149
rect 5100 -210 5170 -183
rect 5200 -149 5270 -126
rect 5200 -183 5218 -149
rect 5252 -183 5270 -149
rect 5200 -210 5270 -183
rect 5300 -149 5370 -126
rect 5300 -183 5318 -149
rect 5352 -183 5370 -149
rect 5300 -210 5370 -183
rect 5400 -149 5470 -126
rect 5400 -183 5418 -149
rect 5452 -183 5470 -149
rect 5400 -210 5470 -183
rect 5500 -149 5570 -126
rect 5500 -183 5518 -149
rect 5552 -183 5570 -149
rect 5500 -210 5570 -183
rect 5600 -149 5670 -126
rect 5600 -183 5618 -149
rect 5652 -183 5670 -149
rect 5600 -210 5670 -183
rect 5700 -149 5770 -126
rect 5700 -183 5718 -149
rect 5752 -183 5770 -149
rect 5700 -210 5770 -183
rect 5800 -149 5870 -126
rect 5800 -183 5818 -149
rect 5852 -183 5870 -149
rect 5800 -210 5870 -183
rect 5900 -149 5970 -126
rect 5900 -183 5918 -149
rect 5952 -183 5970 -149
rect 5900 -210 5970 -183
rect 6000 -149 6070 -126
rect 6000 -183 6018 -149
rect 6052 -183 6070 -149
rect 6000 -210 6070 -183
rect 6100 -149 6170 -126
rect 6100 -183 6118 -149
rect 6152 -183 6170 -149
rect 6100 -210 6170 -183
rect 6200 -149 6270 -126
rect 6200 -183 6218 -149
rect 6252 -183 6270 -149
rect 6200 -210 6270 -183
rect 6300 -149 6370 -126
rect 6300 -183 6318 -149
rect 6352 -183 6370 -149
rect 6300 -210 6370 -183
rect 6400 -149 6470 -126
rect 6400 -183 6418 -149
rect 6452 -183 6470 -149
rect 6400 -210 6470 -183
rect 6500 -149 6570 -126
rect 6500 -183 6518 -149
rect 6552 -183 6570 -149
rect 6500 -210 6570 -183
rect 6600 -149 6670 -126
rect 6600 -183 6618 -149
rect 6652 -183 6670 -149
rect 6600 -210 6670 -183
rect 6700 -149 6770 -126
rect 6700 -183 6718 -149
rect 6752 -183 6770 -149
rect 6700 -210 6770 -183
rect 6800 -149 6870 -126
rect 6800 -183 6818 -149
rect 6852 -183 6870 -149
rect 6800 -210 6870 -183
rect 6900 -149 6970 -126
rect 6900 -183 6918 -149
rect 6952 -183 6970 -149
rect 6900 -210 6970 -183
rect 7000 -149 7070 -126
rect 7000 -183 7018 -149
rect 7052 -183 7070 -149
rect 7000 -210 7070 -183
rect 7100 -149 7170 -126
rect 7100 -183 7118 -149
rect 7152 -183 7170 -149
rect 7100 -210 7170 -183
rect 7200 -149 7270 -126
rect 7200 -183 7218 -149
rect 7252 -183 7270 -149
rect 7200 -210 7270 -183
rect 7300 -149 7370 -126
rect 7300 -183 7318 -149
rect 7352 -183 7370 -149
rect 7300 -210 7370 -183
rect 7400 -149 7470 -126
rect 7400 -183 7418 -149
rect 7452 -183 7470 -149
rect 7400 -210 7470 -183
rect 7500 -149 7570 -126
rect 7500 -183 7518 -149
rect 7552 -183 7570 -149
rect 7500 -210 7570 -183
rect 7600 -149 7670 -126
rect 7600 -183 7618 -149
rect 7652 -183 7670 -149
rect 7600 -210 7670 -183
rect 7700 -149 7770 -126
rect 7700 -183 7718 -149
rect 7752 -183 7770 -149
rect 7700 -210 7770 -183
rect 7800 -149 7870 -126
rect 7800 -183 7818 -149
rect 7852 -183 7870 -149
rect 7800 -210 7870 -183
rect 7900 -149 7970 -126
rect 7900 -183 7918 -149
rect 7952 -183 7970 -149
rect 7900 -210 7970 -183
rect 8000 -149 8070 -126
rect 8000 -183 8018 -149
rect 8052 -183 8070 -149
rect 8000 -210 8070 -183
rect 8100 -149 8170 -126
rect 8100 -183 8118 -149
rect 8152 -183 8170 -149
rect 8100 -210 8170 -183
rect 8200 -149 8270 -126
rect 8200 -183 8218 -149
rect 8252 -183 8270 -149
rect 8200 -210 8270 -183
rect 8300 -149 8370 -126
rect 8300 -183 8318 -149
rect 8352 -183 8370 -149
rect 8300 -210 8370 -183
rect 8400 -149 8470 -126
rect 8400 -183 8418 -149
rect 8452 -183 8470 -149
rect 8400 -210 8470 -183
rect 8500 -149 8570 -126
rect 8500 -183 8518 -149
rect 8552 -183 8570 -149
rect 8500 -210 8570 -183
rect 8600 -149 8670 -126
rect 8600 -183 8618 -149
rect 8652 -183 8670 -149
rect 8600 -210 8670 -183
rect 8700 -149 8770 -126
rect 8700 -183 8718 -149
rect 8752 -183 8770 -149
rect 8700 -210 8770 -183
rect 8800 -149 8870 -126
rect 8800 -183 8818 -149
rect 8852 -183 8870 -149
rect 8800 -210 8870 -183
rect 8900 -149 8970 -126
rect 8900 -183 8918 -149
rect 8952 -183 8970 -149
rect 8900 -210 8970 -183
rect 9000 -149 9070 -126
rect 9000 -183 9018 -149
rect 9052 -183 9070 -149
rect 9000 -210 9070 -183
rect 9100 -149 9170 -126
rect 9100 -183 9118 -149
rect 9152 -183 9170 -149
rect 9100 -210 9170 -183
rect 9200 -149 9270 -126
rect 9200 -183 9218 -149
rect 9252 -183 9270 -149
rect 9200 -210 9270 -183
rect 9300 -149 9370 -126
rect 9300 -183 9318 -149
rect 9352 -183 9370 -149
rect 9300 -210 9370 -183
rect 9400 -149 9470 -126
rect 9400 -183 9418 -149
rect 9452 -183 9470 -149
rect 9400 -210 9470 -183
rect 9500 -149 9570 -126
rect 9500 -183 9518 -149
rect 9552 -183 9570 -149
rect 9500 -210 9570 -183
rect 9600 -149 9670 -126
rect 9600 -183 9618 -149
rect 9652 -183 9670 -149
rect 9600 -210 9670 -183
rect 9700 -149 9770 -126
rect 9700 -183 9718 -149
rect 9752 -183 9770 -149
rect 9700 -210 9770 -183
rect 9800 -149 9870 -126
rect 9800 -183 9818 -149
rect 9852 -183 9870 -149
rect 9800 -210 9870 -183
rect 9900 -149 9970 -126
rect 9900 -183 9918 -149
rect 9952 -183 9970 -149
rect 9900 -210 9970 -183
rect 10000 -149 10070 -126
rect 10000 -183 10018 -149
rect 10052 -183 10070 -149
rect 10000 -210 10070 -183
rect 10100 -149 10170 -126
rect 10100 -183 10118 -149
rect 10152 -183 10170 -149
rect 10100 -210 10170 -183
rect 10200 -149 10270 -126
rect 10200 -183 10218 -149
rect 10252 -183 10270 -149
rect 10200 -210 10270 -183
rect 10300 -149 10370 -126
rect 10300 -183 10318 -149
rect 10352 -183 10370 -149
rect 10300 -210 10370 -183
rect 10400 -149 10470 -126
rect 10400 -183 10418 -149
rect 10452 -183 10470 -149
rect 10400 -210 10470 -183
rect 10500 -149 10570 -126
rect 10500 -183 10518 -149
rect 10552 -183 10570 -149
rect 10500 -210 10570 -183
rect 10600 -149 10670 -126
rect 10600 -183 10618 -149
rect 10652 -183 10670 -149
rect 10600 -210 10670 -183
rect 10700 -149 10770 -126
rect 10700 -183 10718 -149
rect 10752 -183 10770 -149
rect 10700 -210 10770 -183
rect 10800 -149 10870 -126
rect 10800 -183 10818 -149
rect 10852 -183 10870 -149
rect 10800 -210 10870 -183
rect 10900 -149 10970 -126
rect 10900 -183 10918 -149
rect 10952 -183 10970 -149
rect 10900 -210 10970 -183
rect 11000 -149 11070 -126
rect 11000 -183 11018 -149
rect 11052 -183 11070 -149
rect 11000 -210 11070 -183
rect 11100 -149 11170 -126
rect 11100 -183 11118 -149
rect 11152 -183 11170 -149
rect 11100 -210 11170 -183
rect 11200 -149 11270 -126
rect 11200 -183 11218 -149
rect 11252 -183 11270 -149
rect 11200 -210 11270 -183
rect 11300 -149 11370 -126
rect 11300 -183 11318 -149
rect 11352 -183 11370 -149
rect 11300 -210 11370 -183
rect 11400 -149 11470 -126
rect 11400 -183 11418 -149
rect 11452 -183 11470 -149
rect 11400 -210 11470 -183
rect 11500 -149 11570 -126
rect 11500 -183 11518 -149
rect 11552 -183 11570 -149
rect 11500 -210 11570 -183
rect 11600 -149 11670 -126
rect 11600 -183 11618 -149
rect 11652 -183 11670 -149
rect 11600 -210 11670 -183
rect 11700 -149 11770 -126
rect 11700 -183 11718 -149
rect 11752 -183 11770 -149
rect 11700 -210 11770 -183
rect 11800 -149 11870 -126
rect 11800 -183 11818 -149
rect 11852 -183 11870 -149
rect 11800 -210 11870 -183
rect 11900 -149 11970 -126
rect 11900 -183 11918 -149
rect 11952 -183 11970 -149
rect 11900 -210 11970 -183
rect 12000 -149 12070 -126
rect 12000 -183 12018 -149
rect 12052 -183 12070 -149
rect 12000 -210 12070 -183
rect 12100 -149 12170 -126
rect 12100 -183 12118 -149
rect 12152 -183 12170 -149
rect 12100 -210 12170 -183
rect 12200 -149 12270 -126
rect 12200 -183 12218 -149
rect 12252 -183 12270 -149
rect 12200 -210 12270 -183
rect 12300 -149 12370 -126
rect 12300 -183 12318 -149
rect 12352 -183 12370 -149
rect 12300 -210 12370 -183
rect 12400 -149 12470 -126
rect 12400 -183 12418 -149
rect 12452 -183 12470 -149
rect 12400 -210 12470 -183
rect 12500 -149 12570 -126
rect 12500 -183 12518 -149
rect 12552 -183 12570 -149
rect 12500 -210 12570 -183
rect 12600 -149 12670 -126
rect 12600 -183 12618 -149
rect 12652 -183 12670 -149
rect 12600 -210 12670 -183
rect 12700 -149 12764 -126
rect 12700 -183 12718 -149
rect 12752 -183 12764 -149
rect 12700 -210 12764 -183
rect 14540 -208 14690 -171
rect 14540 -242 14562 -208
rect 14596 -242 14630 -208
rect 14664 -242 14690 -208
rect 14540 -260 14690 -242
rect 15652 -208 15802 -171
rect 15652 -242 15678 -208
rect 15712 -242 15746 -208
rect 15780 -242 15802 -208
rect 15652 -260 15802 -242
rect 14540 -308 14690 -290
rect 14540 -342 14562 -308
rect 14596 -342 14630 -308
rect 14664 -342 14690 -308
rect 14540 -360 14690 -342
rect 15652 -308 15802 -290
rect 15652 -342 15678 -308
rect 15712 -342 15746 -308
rect 15780 -342 15802 -308
rect 15652 -360 15802 -342
rect 14540 -408 14690 -390
rect 14540 -442 14562 -408
rect 14596 -442 14630 -408
rect 14664 -442 14690 -408
rect 14540 -460 14690 -442
rect 15652 -408 15802 -390
rect 15652 -442 15678 -408
rect 15712 -442 15746 -408
rect 15780 -442 15802 -408
rect 15652 -460 15802 -442
rect 14540 -508 14690 -490
rect 14540 -542 14562 -508
rect 14596 -542 14630 -508
rect 14664 -542 14690 -508
rect 14540 -560 14690 -542
rect 15652 -508 15802 -490
rect 15652 -542 15678 -508
rect 15712 -542 15746 -508
rect 15780 -542 15802 -508
rect 15652 -560 15802 -542
rect 14540 -608 14690 -590
rect 14540 -642 14562 -608
rect 14596 -642 14630 -608
rect 14664 -642 14690 -608
rect 14540 -660 14690 -642
rect 15652 -608 15802 -590
rect 15652 -642 15678 -608
rect 15712 -642 15746 -608
rect 15780 -642 15802 -608
rect 15652 -660 15802 -642
rect 14540 -708 14690 -690
rect 14540 -742 14562 -708
rect 14596 -742 14630 -708
rect 14664 -742 14690 -708
rect 14540 -760 14690 -742
rect 15652 -708 15802 -690
rect 15652 -742 15678 -708
rect 15712 -742 15746 -708
rect 15780 -742 15802 -708
rect 15652 -760 15802 -742
rect 14540 -808 14690 -790
rect 14540 -842 14562 -808
rect 14596 -842 14630 -808
rect 14664 -842 14690 -808
rect -10 -858 108 -846
rect -10 -892 -2 -858
rect 32 -892 66 -858
rect 100 -892 108 -858
rect -10 -910 108 -892
rect 162 -858 280 -846
rect 162 -892 170 -858
rect 204 -892 238 -858
rect 272 -892 280 -858
rect 162 -910 280 -892
rect 390 -858 508 -846
rect 390 -892 398 -858
rect 432 -892 466 -858
rect 500 -892 508 -858
rect 390 -910 508 -892
rect 562 -858 680 -846
rect 562 -892 570 -858
rect 604 -892 638 -858
rect 672 -892 680 -858
rect 562 -910 680 -892
rect 790 -858 908 -846
rect 790 -892 798 -858
rect 832 -892 866 -858
rect 900 -892 908 -858
rect -10 -958 108 -940
rect -10 -992 -2 -958
rect 32 -992 66 -958
rect 100 -992 108 -958
rect -10 -1010 108 -992
rect 162 -958 280 -940
rect 162 -992 170 -958
rect 204 -992 238 -958
rect 272 -992 280 -958
rect 162 -1010 280 -992
rect 390 -958 508 -940
rect 390 -992 398 -958
rect 432 -992 466 -958
rect 500 -992 508 -958
rect 390 -1010 508 -992
rect 562 -958 680 -940
rect 790 -910 908 -892
rect 962 -858 1080 -846
rect 962 -892 970 -858
rect 1004 -892 1038 -858
rect 1072 -892 1080 -858
rect 962 -910 1080 -892
rect 1190 -858 1308 -846
rect 1190 -892 1198 -858
rect 1232 -892 1266 -858
rect 1300 -892 1308 -858
rect 1190 -910 1308 -892
rect 1362 -858 1480 -846
rect 1362 -892 1370 -858
rect 1404 -892 1438 -858
rect 1472 -892 1480 -858
rect 1362 -910 1480 -892
rect 1590 -858 1708 -846
rect 1590 -892 1598 -858
rect 1632 -892 1666 -858
rect 1700 -892 1708 -858
rect 562 -992 570 -958
rect 604 -992 638 -958
rect 672 -992 680 -958
rect 562 -1010 680 -992
rect 790 -958 908 -940
rect 790 -992 798 -958
rect 832 -992 866 -958
rect 900 -992 908 -958
rect -10 -1058 108 -1040
rect -10 -1092 -2 -1058
rect 32 -1092 66 -1058
rect 100 -1092 108 -1058
rect -10 -1110 108 -1092
rect 162 -1058 280 -1040
rect 162 -1092 170 -1058
rect 204 -1092 238 -1058
rect 272 -1092 280 -1058
rect 162 -1110 280 -1092
rect 390 -1058 508 -1040
rect 390 -1092 398 -1058
rect 432 -1092 466 -1058
rect 500 -1092 508 -1058
rect 390 -1110 508 -1092
rect 562 -1058 680 -1040
rect 790 -1010 908 -992
rect 962 -958 1080 -940
rect 962 -992 970 -958
rect 1004 -992 1038 -958
rect 1072 -992 1080 -958
rect 962 -1010 1080 -992
rect 1190 -958 1308 -940
rect 1190 -992 1198 -958
rect 1232 -992 1266 -958
rect 1300 -992 1308 -958
rect 1190 -1010 1308 -992
rect 1362 -958 1480 -940
rect 1590 -910 1708 -892
rect 1762 -858 1880 -846
rect 1762 -892 1770 -858
rect 1804 -892 1838 -858
rect 1872 -892 1880 -858
rect 1762 -910 1880 -892
rect 1990 -858 2108 -846
rect 1990 -892 1998 -858
rect 2032 -892 2066 -858
rect 2100 -892 2108 -858
rect 1990 -910 2108 -892
rect 2162 -858 2280 -846
rect 2162 -892 2170 -858
rect 2204 -892 2238 -858
rect 2272 -892 2280 -858
rect 2162 -910 2280 -892
rect 2390 -858 2508 -846
rect 2390 -892 2398 -858
rect 2432 -892 2466 -858
rect 2500 -892 2508 -858
rect 1362 -992 1370 -958
rect 1404 -992 1438 -958
rect 1472 -992 1480 -958
rect 1362 -1010 1480 -992
rect 1590 -958 1708 -940
rect 1590 -992 1598 -958
rect 1632 -992 1666 -958
rect 1700 -992 1708 -958
rect 562 -1092 570 -1058
rect 604 -1092 638 -1058
rect 672 -1092 680 -1058
rect 562 -1110 680 -1092
rect 790 -1058 908 -1040
rect 790 -1092 798 -1058
rect 832 -1092 866 -1058
rect 900 -1092 908 -1058
rect -10 -1158 108 -1140
rect -10 -1192 -2 -1158
rect 32 -1192 66 -1158
rect 100 -1192 108 -1158
rect -10 -1210 108 -1192
rect 162 -1158 280 -1140
rect 162 -1192 170 -1158
rect 204 -1192 238 -1158
rect 272 -1192 280 -1158
rect 162 -1210 280 -1192
rect 390 -1158 508 -1140
rect 390 -1192 398 -1158
rect 432 -1192 466 -1158
rect 500 -1192 508 -1158
rect 390 -1210 508 -1192
rect 562 -1158 680 -1140
rect 790 -1110 908 -1092
rect 962 -1058 1080 -1040
rect 962 -1092 970 -1058
rect 1004 -1092 1038 -1058
rect 1072 -1092 1080 -1058
rect 962 -1110 1080 -1092
rect 1190 -1058 1308 -1040
rect 1190 -1092 1198 -1058
rect 1232 -1092 1266 -1058
rect 1300 -1092 1308 -1058
rect 1190 -1110 1308 -1092
rect 1362 -1058 1480 -1040
rect 1590 -1010 1708 -992
rect 1762 -958 1880 -940
rect 1762 -992 1770 -958
rect 1804 -992 1838 -958
rect 1872 -992 1880 -958
rect 1762 -1010 1880 -992
rect 1990 -958 2108 -940
rect 1990 -992 1998 -958
rect 2032 -992 2066 -958
rect 2100 -992 2108 -958
rect 1990 -1010 2108 -992
rect 2162 -958 2280 -940
rect 2390 -910 2508 -892
rect 2562 -858 2680 -846
rect 2562 -892 2570 -858
rect 2604 -892 2638 -858
rect 2672 -892 2680 -858
rect 2562 -910 2680 -892
rect 2790 -858 2908 -846
rect 2790 -892 2798 -858
rect 2832 -892 2866 -858
rect 2900 -892 2908 -858
rect 2790 -910 2908 -892
rect 2962 -858 3080 -846
rect 2962 -892 2970 -858
rect 3004 -892 3038 -858
rect 3072 -892 3080 -858
rect 2962 -910 3080 -892
rect 3190 -858 3308 -846
rect 3190 -892 3198 -858
rect 3232 -892 3266 -858
rect 3300 -892 3308 -858
rect 2162 -992 2170 -958
rect 2204 -992 2238 -958
rect 2272 -992 2280 -958
rect 2162 -1010 2280 -992
rect 2390 -958 2508 -940
rect 2390 -992 2398 -958
rect 2432 -992 2466 -958
rect 2500 -992 2508 -958
rect 1362 -1092 1370 -1058
rect 1404 -1092 1438 -1058
rect 1472 -1092 1480 -1058
rect 1362 -1110 1480 -1092
rect 1590 -1058 1708 -1040
rect 1590 -1092 1598 -1058
rect 1632 -1092 1666 -1058
rect 1700 -1092 1708 -1058
rect 562 -1192 570 -1158
rect 604 -1192 638 -1158
rect 672 -1192 680 -1158
rect 562 -1210 680 -1192
rect 790 -1158 908 -1140
rect 790 -1192 798 -1158
rect 832 -1192 866 -1158
rect 900 -1192 908 -1158
rect -10 -1258 108 -1240
rect -10 -1292 -2 -1258
rect 32 -1292 66 -1258
rect 100 -1292 108 -1258
rect -10 -1310 108 -1292
rect 162 -1258 280 -1240
rect 162 -1292 170 -1258
rect 204 -1292 238 -1258
rect 272 -1292 280 -1258
rect 162 -1310 280 -1292
rect 390 -1258 508 -1240
rect 390 -1292 398 -1258
rect 432 -1292 466 -1258
rect 500 -1292 508 -1258
rect 390 -1310 508 -1292
rect 562 -1258 680 -1240
rect 790 -1210 908 -1192
rect 962 -1158 1080 -1140
rect 962 -1192 970 -1158
rect 1004 -1192 1038 -1158
rect 1072 -1192 1080 -1158
rect 962 -1210 1080 -1192
rect 1190 -1158 1308 -1140
rect 1190 -1192 1198 -1158
rect 1232 -1192 1266 -1158
rect 1300 -1192 1308 -1158
rect 1190 -1210 1308 -1192
rect 1362 -1158 1480 -1140
rect 1590 -1110 1708 -1092
rect 1762 -1058 1880 -1040
rect 1762 -1092 1770 -1058
rect 1804 -1092 1838 -1058
rect 1872 -1092 1880 -1058
rect 1762 -1110 1880 -1092
rect 1990 -1058 2108 -1040
rect 1990 -1092 1998 -1058
rect 2032 -1092 2066 -1058
rect 2100 -1092 2108 -1058
rect 1990 -1110 2108 -1092
rect 2162 -1058 2280 -1040
rect 2390 -1010 2508 -992
rect 2562 -958 2680 -940
rect 2562 -992 2570 -958
rect 2604 -992 2638 -958
rect 2672 -992 2680 -958
rect 2562 -1010 2680 -992
rect 2790 -958 2908 -940
rect 2790 -992 2798 -958
rect 2832 -992 2866 -958
rect 2900 -992 2908 -958
rect 2790 -1010 2908 -992
rect 2962 -958 3080 -940
rect 3190 -910 3308 -892
rect 3362 -858 3480 -846
rect 3362 -892 3370 -858
rect 3404 -892 3438 -858
rect 3472 -892 3480 -858
rect 3362 -910 3480 -892
rect 3590 -858 3708 -846
rect 3590 -892 3598 -858
rect 3632 -892 3666 -858
rect 3700 -892 3708 -858
rect 3590 -910 3708 -892
rect 3762 -858 3880 -846
rect 3762 -892 3770 -858
rect 3804 -892 3838 -858
rect 3872 -892 3880 -858
rect 3762 -910 3880 -892
rect 3990 -858 4108 -846
rect 3990 -892 3998 -858
rect 4032 -892 4066 -858
rect 4100 -892 4108 -858
rect 2962 -992 2970 -958
rect 3004 -992 3038 -958
rect 3072 -992 3080 -958
rect 2962 -1010 3080 -992
rect 3190 -958 3308 -940
rect 3190 -992 3198 -958
rect 3232 -992 3266 -958
rect 3300 -992 3308 -958
rect 2162 -1092 2170 -1058
rect 2204 -1092 2238 -1058
rect 2272 -1092 2280 -1058
rect 2162 -1110 2280 -1092
rect 2390 -1058 2508 -1040
rect 2390 -1092 2398 -1058
rect 2432 -1092 2466 -1058
rect 2500 -1092 2508 -1058
rect 1362 -1192 1370 -1158
rect 1404 -1192 1438 -1158
rect 1472 -1192 1480 -1158
rect 1362 -1210 1480 -1192
rect 1590 -1158 1708 -1140
rect 1590 -1192 1598 -1158
rect 1632 -1192 1666 -1158
rect 1700 -1192 1708 -1158
rect 562 -1292 570 -1258
rect 604 -1292 638 -1258
rect 672 -1292 680 -1258
rect 562 -1310 680 -1292
rect 790 -1258 908 -1240
rect 790 -1292 798 -1258
rect 832 -1292 866 -1258
rect 900 -1292 908 -1258
rect -10 -1358 108 -1340
rect -10 -1392 -2 -1358
rect 32 -1392 66 -1358
rect 100 -1392 108 -1358
rect -10 -1410 108 -1392
rect 162 -1358 280 -1340
rect 162 -1392 170 -1358
rect 204 -1392 238 -1358
rect 272 -1392 280 -1358
rect 162 -1410 280 -1392
rect 390 -1358 508 -1340
rect 390 -1392 398 -1358
rect 432 -1392 466 -1358
rect 500 -1392 508 -1358
rect 390 -1410 508 -1392
rect 562 -1358 680 -1340
rect 790 -1310 908 -1292
rect 962 -1258 1080 -1240
rect 962 -1292 970 -1258
rect 1004 -1292 1038 -1258
rect 1072 -1292 1080 -1258
rect 962 -1310 1080 -1292
rect 1190 -1258 1308 -1240
rect 1190 -1292 1198 -1258
rect 1232 -1292 1266 -1258
rect 1300 -1292 1308 -1258
rect 1190 -1310 1308 -1292
rect 1362 -1258 1480 -1240
rect 1590 -1210 1708 -1192
rect 1762 -1158 1880 -1140
rect 1762 -1192 1770 -1158
rect 1804 -1192 1838 -1158
rect 1872 -1192 1880 -1158
rect 1762 -1210 1880 -1192
rect 1990 -1158 2108 -1140
rect 1990 -1192 1998 -1158
rect 2032 -1192 2066 -1158
rect 2100 -1192 2108 -1158
rect 1990 -1210 2108 -1192
rect 2162 -1158 2280 -1140
rect 2390 -1110 2508 -1092
rect 2562 -1058 2680 -1040
rect 2562 -1092 2570 -1058
rect 2604 -1092 2638 -1058
rect 2672 -1092 2680 -1058
rect 2562 -1110 2680 -1092
rect 2790 -1058 2908 -1040
rect 2790 -1092 2798 -1058
rect 2832 -1092 2866 -1058
rect 2900 -1092 2908 -1058
rect 2790 -1110 2908 -1092
rect 2962 -1058 3080 -1040
rect 3190 -1010 3308 -992
rect 3362 -958 3480 -940
rect 3362 -992 3370 -958
rect 3404 -992 3438 -958
rect 3472 -992 3480 -958
rect 3362 -1010 3480 -992
rect 3590 -958 3708 -940
rect 3590 -992 3598 -958
rect 3632 -992 3666 -958
rect 3700 -992 3708 -958
rect 3590 -1010 3708 -992
rect 3762 -958 3880 -940
rect 3990 -910 4108 -892
rect 4162 -858 4280 -846
rect 4162 -892 4170 -858
rect 4204 -892 4238 -858
rect 4272 -892 4280 -858
rect 4162 -910 4280 -892
rect 4390 -858 4508 -846
rect 4390 -892 4398 -858
rect 4432 -892 4466 -858
rect 4500 -892 4508 -858
rect 4390 -910 4508 -892
rect 4562 -858 4680 -846
rect 4562 -892 4570 -858
rect 4604 -892 4638 -858
rect 4672 -892 4680 -858
rect 4562 -910 4680 -892
rect 4790 -858 4908 -846
rect 4790 -892 4798 -858
rect 4832 -892 4866 -858
rect 4900 -892 4908 -858
rect 3762 -992 3770 -958
rect 3804 -992 3838 -958
rect 3872 -992 3880 -958
rect 3762 -1010 3880 -992
rect 3990 -958 4108 -940
rect 3990 -992 3998 -958
rect 4032 -992 4066 -958
rect 4100 -992 4108 -958
rect 2962 -1092 2970 -1058
rect 3004 -1092 3038 -1058
rect 3072 -1092 3080 -1058
rect 2962 -1110 3080 -1092
rect 3190 -1058 3308 -1040
rect 3190 -1092 3198 -1058
rect 3232 -1092 3266 -1058
rect 3300 -1092 3308 -1058
rect 2162 -1192 2170 -1158
rect 2204 -1192 2238 -1158
rect 2272 -1192 2280 -1158
rect 2162 -1210 2280 -1192
rect 2390 -1158 2508 -1140
rect 2390 -1192 2398 -1158
rect 2432 -1192 2466 -1158
rect 2500 -1192 2508 -1158
rect 1362 -1292 1370 -1258
rect 1404 -1292 1438 -1258
rect 1472 -1292 1480 -1258
rect 1362 -1310 1480 -1292
rect 1590 -1258 1708 -1240
rect 1590 -1292 1598 -1258
rect 1632 -1292 1666 -1258
rect 1700 -1292 1708 -1258
rect 562 -1392 570 -1358
rect 604 -1392 638 -1358
rect 672 -1392 680 -1358
rect 562 -1410 680 -1392
rect 790 -1358 908 -1340
rect 790 -1392 798 -1358
rect 832 -1392 866 -1358
rect 900 -1392 908 -1358
rect -10 -1458 108 -1440
rect -10 -1492 -2 -1458
rect 32 -1492 66 -1458
rect 100 -1492 108 -1458
rect -10 -1510 108 -1492
rect 162 -1458 280 -1440
rect 162 -1492 170 -1458
rect 204 -1492 238 -1458
rect 272 -1492 280 -1458
rect 162 -1510 280 -1492
rect 390 -1458 508 -1440
rect 390 -1492 398 -1458
rect 432 -1492 466 -1458
rect 500 -1492 508 -1458
rect 390 -1510 508 -1492
rect 562 -1458 680 -1440
rect 790 -1410 908 -1392
rect 962 -1358 1080 -1340
rect 962 -1392 970 -1358
rect 1004 -1392 1038 -1358
rect 1072 -1392 1080 -1358
rect 962 -1410 1080 -1392
rect 1190 -1358 1308 -1340
rect 1190 -1392 1198 -1358
rect 1232 -1392 1266 -1358
rect 1300 -1392 1308 -1358
rect 1190 -1410 1308 -1392
rect 1362 -1358 1480 -1340
rect 1590 -1310 1708 -1292
rect 1762 -1258 1880 -1240
rect 1762 -1292 1770 -1258
rect 1804 -1292 1838 -1258
rect 1872 -1292 1880 -1258
rect 1762 -1310 1880 -1292
rect 1990 -1258 2108 -1240
rect 1990 -1292 1998 -1258
rect 2032 -1292 2066 -1258
rect 2100 -1292 2108 -1258
rect 1990 -1310 2108 -1292
rect 2162 -1258 2280 -1240
rect 2390 -1210 2508 -1192
rect 2562 -1158 2680 -1140
rect 2562 -1192 2570 -1158
rect 2604 -1192 2638 -1158
rect 2672 -1192 2680 -1158
rect 2562 -1210 2680 -1192
rect 2790 -1158 2908 -1140
rect 2790 -1192 2798 -1158
rect 2832 -1192 2866 -1158
rect 2900 -1192 2908 -1158
rect 2790 -1210 2908 -1192
rect 2962 -1158 3080 -1140
rect 3190 -1110 3308 -1092
rect 3362 -1058 3480 -1040
rect 3362 -1092 3370 -1058
rect 3404 -1092 3438 -1058
rect 3472 -1092 3480 -1058
rect 3362 -1110 3480 -1092
rect 3590 -1058 3708 -1040
rect 3590 -1092 3598 -1058
rect 3632 -1092 3666 -1058
rect 3700 -1092 3708 -1058
rect 3590 -1110 3708 -1092
rect 3762 -1058 3880 -1040
rect 3990 -1010 4108 -992
rect 4162 -958 4280 -940
rect 4162 -992 4170 -958
rect 4204 -992 4238 -958
rect 4272 -992 4280 -958
rect 4162 -1010 4280 -992
rect 4390 -958 4508 -940
rect 4390 -992 4398 -958
rect 4432 -992 4466 -958
rect 4500 -992 4508 -958
rect 4390 -1010 4508 -992
rect 4562 -958 4680 -940
rect 4790 -910 4908 -892
rect 4962 -858 5080 -846
rect 4962 -892 4970 -858
rect 5004 -892 5038 -858
rect 5072 -892 5080 -858
rect 4962 -910 5080 -892
rect 5190 -858 5308 -846
rect 5190 -892 5198 -858
rect 5232 -892 5266 -858
rect 5300 -892 5308 -858
rect 5190 -910 5308 -892
rect 5362 -858 5480 -846
rect 5362 -892 5370 -858
rect 5404 -892 5438 -858
rect 5472 -892 5480 -858
rect 5362 -910 5480 -892
rect 5590 -858 5708 -846
rect 5590 -892 5598 -858
rect 5632 -892 5666 -858
rect 5700 -892 5708 -858
rect 4562 -992 4570 -958
rect 4604 -992 4638 -958
rect 4672 -992 4680 -958
rect 4562 -1010 4680 -992
rect 4790 -958 4908 -940
rect 4790 -992 4798 -958
rect 4832 -992 4866 -958
rect 4900 -992 4908 -958
rect 3762 -1092 3770 -1058
rect 3804 -1092 3838 -1058
rect 3872 -1092 3880 -1058
rect 3762 -1110 3880 -1092
rect 3990 -1058 4108 -1040
rect 3990 -1092 3998 -1058
rect 4032 -1092 4066 -1058
rect 4100 -1092 4108 -1058
rect 2962 -1192 2970 -1158
rect 3004 -1192 3038 -1158
rect 3072 -1192 3080 -1158
rect 2962 -1210 3080 -1192
rect 3190 -1158 3308 -1140
rect 3190 -1192 3198 -1158
rect 3232 -1192 3266 -1158
rect 3300 -1192 3308 -1158
rect 2162 -1292 2170 -1258
rect 2204 -1292 2238 -1258
rect 2272 -1292 2280 -1258
rect 2162 -1310 2280 -1292
rect 2390 -1258 2508 -1240
rect 2390 -1292 2398 -1258
rect 2432 -1292 2466 -1258
rect 2500 -1292 2508 -1258
rect 1362 -1392 1370 -1358
rect 1404 -1392 1438 -1358
rect 1472 -1392 1480 -1358
rect 1362 -1410 1480 -1392
rect 1590 -1358 1708 -1340
rect 1590 -1392 1598 -1358
rect 1632 -1392 1666 -1358
rect 1700 -1392 1708 -1358
rect 562 -1492 570 -1458
rect 604 -1492 638 -1458
rect 672 -1492 680 -1458
rect 562 -1510 680 -1492
rect 790 -1458 908 -1440
rect 790 -1492 798 -1458
rect 832 -1492 866 -1458
rect 900 -1492 908 -1458
rect -10 -1558 108 -1540
rect -10 -1592 -2 -1558
rect 32 -1592 66 -1558
rect 100 -1592 108 -1558
rect -10 -1610 108 -1592
rect 162 -1558 280 -1540
rect 162 -1592 170 -1558
rect 204 -1592 238 -1558
rect 272 -1592 280 -1558
rect 162 -1610 280 -1592
rect 390 -1558 508 -1540
rect 390 -1592 398 -1558
rect 432 -1592 466 -1558
rect 500 -1592 508 -1558
rect 390 -1610 508 -1592
rect 562 -1558 680 -1540
rect 790 -1510 908 -1492
rect 962 -1458 1080 -1440
rect 962 -1492 970 -1458
rect 1004 -1492 1038 -1458
rect 1072 -1492 1080 -1458
rect 962 -1510 1080 -1492
rect 1190 -1458 1308 -1440
rect 1190 -1492 1198 -1458
rect 1232 -1492 1266 -1458
rect 1300 -1492 1308 -1458
rect 1190 -1510 1308 -1492
rect 1362 -1458 1480 -1440
rect 1590 -1410 1708 -1392
rect 1762 -1358 1880 -1340
rect 1762 -1392 1770 -1358
rect 1804 -1392 1838 -1358
rect 1872 -1392 1880 -1358
rect 1762 -1410 1880 -1392
rect 1990 -1358 2108 -1340
rect 1990 -1392 1998 -1358
rect 2032 -1392 2066 -1358
rect 2100 -1392 2108 -1358
rect 1990 -1410 2108 -1392
rect 2162 -1358 2280 -1340
rect 2390 -1310 2508 -1292
rect 2562 -1258 2680 -1240
rect 2562 -1292 2570 -1258
rect 2604 -1292 2638 -1258
rect 2672 -1292 2680 -1258
rect 2562 -1310 2680 -1292
rect 2790 -1258 2908 -1240
rect 2790 -1292 2798 -1258
rect 2832 -1292 2866 -1258
rect 2900 -1292 2908 -1258
rect 2790 -1310 2908 -1292
rect 2962 -1258 3080 -1240
rect 3190 -1210 3308 -1192
rect 3362 -1158 3480 -1140
rect 3362 -1192 3370 -1158
rect 3404 -1192 3438 -1158
rect 3472 -1192 3480 -1158
rect 3362 -1210 3480 -1192
rect 3590 -1158 3708 -1140
rect 3590 -1192 3598 -1158
rect 3632 -1192 3666 -1158
rect 3700 -1192 3708 -1158
rect 3590 -1210 3708 -1192
rect 3762 -1158 3880 -1140
rect 3990 -1110 4108 -1092
rect 4162 -1058 4280 -1040
rect 4162 -1092 4170 -1058
rect 4204 -1092 4238 -1058
rect 4272 -1092 4280 -1058
rect 4162 -1110 4280 -1092
rect 4390 -1058 4508 -1040
rect 4390 -1092 4398 -1058
rect 4432 -1092 4466 -1058
rect 4500 -1092 4508 -1058
rect 4390 -1110 4508 -1092
rect 4562 -1058 4680 -1040
rect 4790 -1010 4908 -992
rect 4962 -958 5080 -940
rect 4962 -992 4970 -958
rect 5004 -992 5038 -958
rect 5072 -992 5080 -958
rect 4962 -1010 5080 -992
rect 5190 -958 5308 -940
rect 5190 -992 5198 -958
rect 5232 -992 5266 -958
rect 5300 -992 5308 -958
rect 5190 -1010 5308 -992
rect 5362 -958 5480 -940
rect 5590 -910 5708 -892
rect 5762 -858 5880 -846
rect 5762 -892 5770 -858
rect 5804 -892 5838 -858
rect 5872 -892 5880 -858
rect 5762 -910 5880 -892
rect 5990 -858 6108 -846
rect 5990 -892 5998 -858
rect 6032 -892 6066 -858
rect 6100 -892 6108 -858
rect 5990 -910 6108 -892
rect 6162 -858 6280 -846
rect 6162 -892 6170 -858
rect 6204 -892 6238 -858
rect 6272 -892 6280 -858
rect 6162 -910 6280 -892
rect 6390 -858 6508 -846
rect 6390 -892 6398 -858
rect 6432 -892 6466 -858
rect 6500 -892 6508 -858
rect 5362 -992 5370 -958
rect 5404 -992 5438 -958
rect 5472 -992 5480 -958
rect 5362 -1010 5480 -992
rect 5590 -958 5708 -940
rect 5590 -992 5598 -958
rect 5632 -992 5666 -958
rect 5700 -992 5708 -958
rect 4562 -1092 4570 -1058
rect 4604 -1092 4638 -1058
rect 4672 -1092 4680 -1058
rect 4562 -1110 4680 -1092
rect 4790 -1058 4908 -1040
rect 4790 -1092 4798 -1058
rect 4832 -1092 4866 -1058
rect 4900 -1092 4908 -1058
rect 3762 -1192 3770 -1158
rect 3804 -1192 3838 -1158
rect 3872 -1192 3880 -1158
rect 3762 -1210 3880 -1192
rect 3990 -1158 4108 -1140
rect 3990 -1192 3998 -1158
rect 4032 -1192 4066 -1158
rect 4100 -1192 4108 -1158
rect 2962 -1292 2970 -1258
rect 3004 -1292 3038 -1258
rect 3072 -1292 3080 -1258
rect 2962 -1310 3080 -1292
rect 3190 -1258 3308 -1240
rect 3190 -1292 3198 -1258
rect 3232 -1292 3266 -1258
rect 3300 -1292 3308 -1258
rect 2162 -1392 2170 -1358
rect 2204 -1392 2238 -1358
rect 2272 -1392 2280 -1358
rect 2162 -1410 2280 -1392
rect 2390 -1358 2508 -1340
rect 2390 -1392 2398 -1358
rect 2432 -1392 2466 -1358
rect 2500 -1392 2508 -1358
rect 1362 -1492 1370 -1458
rect 1404 -1492 1438 -1458
rect 1472 -1492 1480 -1458
rect 1362 -1510 1480 -1492
rect 1590 -1458 1708 -1440
rect 1590 -1492 1598 -1458
rect 1632 -1492 1666 -1458
rect 1700 -1492 1708 -1458
rect 562 -1592 570 -1558
rect 604 -1592 638 -1558
rect 672 -1592 680 -1558
rect 562 -1610 680 -1592
rect 790 -1558 908 -1540
rect 790 -1592 798 -1558
rect 832 -1592 866 -1558
rect 900 -1592 908 -1558
rect -10 -1658 108 -1640
rect -10 -1692 -2 -1658
rect 32 -1692 66 -1658
rect 100 -1692 108 -1658
rect -10 -1710 108 -1692
rect 162 -1658 280 -1640
rect 162 -1692 170 -1658
rect 204 -1692 238 -1658
rect 272 -1692 280 -1658
rect 162 -1710 280 -1692
rect 390 -1658 508 -1640
rect 390 -1692 398 -1658
rect 432 -1692 466 -1658
rect 500 -1692 508 -1658
rect 390 -1710 508 -1692
rect 562 -1658 680 -1640
rect 790 -1610 908 -1592
rect 962 -1558 1080 -1540
rect 962 -1592 970 -1558
rect 1004 -1592 1038 -1558
rect 1072 -1592 1080 -1558
rect 962 -1610 1080 -1592
rect 1190 -1558 1308 -1540
rect 1190 -1592 1198 -1558
rect 1232 -1592 1266 -1558
rect 1300 -1592 1308 -1558
rect 1190 -1610 1308 -1592
rect 1362 -1558 1480 -1540
rect 1590 -1510 1708 -1492
rect 1762 -1458 1880 -1440
rect 1762 -1492 1770 -1458
rect 1804 -1492 1838 -1458
rect 1872 -1492 1880 -1458
rect 1762 -1510 1880 -1492
rect 1990 -1458 2108 -1440
rect 1990 -1492 1998 -1458
rect 2032 -1492 2066 -1458
rect 2100 -1492 2108 -1458
rect 1990 -1510 2108 -1492
rect 2162 -1458 2280 -1440
rect 2390 -1410 2508 -1392
rect 2562 -1358 2680 -1340
rect 2562 -1392 2570 -1358
rect 2604 -1392 2638 -1358
rect 2672 -1392 2680 -1358
rect 2562 -1410 2680 -1392
rect 2790 -1358 2908 -1340
rect 2790 -1392 2798 -1358
rect 2832 -1392 2866 -1358
rect 2900 -1392 2908 -1358
rect 2790 -1410 2908 -1392
rect 2962 -1358 3080 -1340
rect 3190 -1310 3308 -1292
rect 3362 -1258 3480 -1240
rect 3362 -1292 3370 -1258
rect 3404 -1292 3438 -1258
rect 3472 -1292 3480 -1258
rect 3362 -1310 3480 -1292
rect 3590 -1258 3708 -1240
rect 3590 -1292 3598 -1258
rect 3632 -1292 3666 -1258
rect 3700 -1292 3708 -1258
rect 3590 -1310 3708 -1292
rect 3762 -1258 3880 -1240
rect 3990 -1210 4108 -1192
rect 4162 -1158 4280 -1140
rect 4162 -1192 4170 -1158
rect 4204 -1192 4238 -1158
rect 4272 -1192 4280 -1158
rect 4162 -1210 4280 -1192
rect 4390 -1158 4508 -1140
rect 4390 -1192 4398 -1158
rect 4432 -1192 4466 -1158
rect 4500 -1192 4508 -1158
rect 4390 -1210 4508 -1192
rect 4562 -1158 4680 -1140
rect 4790 -1110 4908 -1092
rect 4962 -1058 5080 -1040
rect 4962 -1092 4970 -1058
rect 5004 -1092 5038 -1058
rect 5072 -1092 5080 -1058
rect 4962 -1110 5080 -1092
rect 5190 -1058 5308 -1040
rect 5190 -1092 5198 -1058
rect 5232 -1092 5266 -1058
rect 5300 -1092 5308 -1058
rect 5190 -1110 5308 -1092
rect 5362 -1058 5480 -1040
rect 5590 -1010 5708 -992
rect 5762 -958 5880 -940
rect 5762 -992 5770 -958
rect 5804 -992 5838 -958
rect 5872 -992 5880 -958
rect 5762 -1010 5880 -992
rect 5990 -958 6108 -940
rect 5990 -992 5998 -958
rect 6032 -992 6066 -958
rect 6100 -992 6108 -958
rect 5990 -1010 6108 -992
rect 6162 -958 6280 -940
rect 6390 -910 6508 -892
rect 6562 -858 6680 -846
rect 6562 -892 6570 -858
rect 6604 -892 6638 -858
rect 6672 -892 6680 -858
rect 6562 -910 6680 -892
rect 6790 -858 6908 -846
rect 6790 -892 6798 -858
rect 6832 -892 6866 -858
rect 6900 -892 6908 -858
rect 6790 -910 6908 -892
rect 6962 -858 7080 -846
rect 6962 -892 6970 -858
rect 7004 -892 7038 -858
rect 7072 -892 7080 -858
rect 6962 -910 7080 -892
rect 7190 -858 7308 -846
rect 7190 -892 7198 -858
rect 7232 -892 7266 -858
rect 7300 -892 7308 -858
rect 6162 -992 6170 -958
rect 6204 -992 6238 -958
rect 6272 -992 6280 -958
rect 6162 -1010 6280 -992
rect 6390 -958 6508 -940
rect 6390 -992 6398 -958
rect 6432 -992 6466 -958
rect 6500 -992 6508 -958
rect 5362 -1092 5370 -1058
rect 5404 -1092 5438 -1058
rect 5472 -1092 5480 -1058
rect 5362 -1110 5480 -1092
rect 5590 -1058 5708 -1040
rect 5590 -1092 5598 -1058
rect 5632 -1092 5666 -1058
rect 5700 -1092 5708 -1058
rect 4562 -1192 4570 -1158
rect 4604 -1192 4638 -1158
rect 4672 -1192 4680 -1158
rect 4562 -1210 4680 -1192
rect 4790 -1158 4908 -1140
rect 4790 -1192 4798 -1158
rect 4832 -1192 4866 -1158
rect 4900 -1192 4908 -1158
rect 3762 -1292 3770 -1258
rect 3804 -1292 3838 -1258
rect 3872 -1292 3880 -1258
rect 3762 -1310 3880 -1292
rect 3990 -1258 4108 -1240
rect 3990 -1292 3998 -1258
rect 4032 -1292 4066 -1258
rect 4100 -1292 4108 -1258
rect 2962 -1392 2970 -1358
rect 3004 -1392 3038 -1358
rect 3072 -1392 3080 -1358
rect 2962 -1410 3080 -1392
rect 3190 -1358 3308 -1340
rect 3190 -1392 3198 -1358
rect 3232 -1392 3266 -1358
rect 3300 -1392 3308 -1358
rect 2162 -1492 2170 -1458
rect 2204 -1492 2238 -1458
rect 2272 -1492 2280 -1458
rect 2162 -1510 2280 -1492
rect 2390 -1458 2508 -1440
rect 2390 -1492 2398 -1458
rect 2432 -1492 2466 -1458
rect 2500 -1492 2508 -1458
rect 1362 -1592 1370 -1558
rect 1404 -1592 1438 -1558
rect 1472 -1592 1480 -1558
rect 1362 -1610 1480 -1592
rect 1590 -1558 1708 -1540
rect 1590 -1592 1598 -1558
rect 1632 -1592 1666 -1558
rect 1700 -1592 1708 -1558
rect 562 -1692 570 -1658
rect 604 -1692 638 -1658
rect 672 -1692 680 -1658
rect 562 -1710 680 -1692
rect 790 -1658 908 -1640
rect 790 -1692 798 -1658
rect 832 -1692 866 -1658
rect 900 -1692 908 -1658
rect -10 -1758 108 -1740
rect -10 -1792 -2 -1758
rect 32 -1792 66 -1758
rect 100 -1792 108 -1758
rect -10 -1810 108 -1792
rect 162 -1758 280 -1740
rect 162 -1792 170 -1758
rect 204 -1792 238 -1758
rect 272 -1792 280 -1758
rect 162 -1810 280 -1792
rect 390 -1758 508 -1740
rect 390 -1792 398 -1758
rect 432 -1792 466 -1758
rect 500 -1792 508 -1758
rect 390 -1810 508 -1792
rect 562 -1758 680 -1740
rect 790 -1710 908 -1692
rect 962 -1658 1080 -1640
rect 962 -1692 970 -1658
rect 1004 -1692 1038 -1658
rect 1072 -1692 1080 -1658
rect 962 -1710 1080 -1692
rect 1190 -1658 1308 -1640
rect 1190 -1692 1198 -1658
rect 1232 -1692 1266 -1658
rect 1300 -1692 1308 -1658
rect 1190 -1710 1308 -1692
rect 1362 -1658 1480 -1640
rect 1590 -1610 1708 -1592
rect 1762 -1558 1880 -1540
rect 1762 -1592 1770 -1558
rect 1804 -1592 1838 -1558
rect 1872 -1592 1880 -1558
rect 1762 -1610 1880 -1592
rect 1990 -1558 2108 -1540
rect 1990 -1592 1998 -1558
rect 2032 -1592 2066 -1558
rect 2100 -1592 2108 -1558
rect 1990 -1610 2108 -1592
rect 2162 -1558 2280 -1540
rect 2390 -1510 2508 -1492
rect 2562 -1458 2680 -1440
rect 2562 -1492 2570 -1458
rect 2604 -1492 2638 -1458
rect 2672 -1492 2680 -1458
rect 2562 -1510 2680 -1492
rect 2790 -1458 2908 -1440
rect 2790 -1492 2798 -1458
rect 2832 -1492 2866 -1458
rect 2900 -1492 2908 -1458
rect 2790 -1510 2908 -1492
rect 2962 -1458 3080 -1440
rect 3190 -1410 3308 -1392
rect 3362 -1358 3480 -1340
rect 3362 -1392 3370 -1358
rect 3404 -1392 3438 -1358
rect 3472 -1392 3480 -1358
rect 3362 -1410 3480 -1392
rect 3590 -1358 3708 -1340
rect 3590 -1392 3598 -1358
rect 3632 -1392 3666 -1358
rect 3700 -1392 3708 -1358
rect 3590 -1410 3708 -1392
rect 3762 -1358 3880 -1340
rect 3990 -1310 4108 -1292
rect 4162 -1258 4280 -1240
rect 4162 -1292 4170 -1258
rect 4204 -1292 4238 -1258
rect 4272 -1292 4280 -1258
rect 4162 -1310 4280 -1292
rect 4390 -1258 4508 -1240
rect 4390 -1292 4398 -1258
rect 4432 -1292 4466 -1258
rect 4500 -1292 4508 -1258
rect 4390 -1310 4508 -1292
rect 4562 -1258 4680 -1240
rect 4790 -1210 4908 -1192
rect 4962 -1158 5080 -1140
rect 4962 -1192 4970 -1158
rect 5004 -1192 5038 -1158
rect 5072 -1192 5080 -1158
rect 4962 -1210 5080 -1192
rect 5190 -1158 5308 -1140
rect 5190 -1192 5198 -1158
rect 5232 -1192 5266 -1158
rect 5300 -1192 5308 -1158
rect 5190 -1210 5308 -1192
rect 5362 -1158 5480 -1140
rect 5590 -1110 5708 -1092
rect 5762 -1058 5880 -1040
rect 5762 -1092 5770 -1058
rect 5804 -1092 5838 -1058
rect 5872 -1092 5880 -1058
rect 5762 -1110 5880 -1092
rect 5990 -1058 6108 -1040
rect 5990 -1092 5998 -1058
rect 6032 -1092 6066 -1058
rect 6100 -1092 6108 -1058
rect 5990 -1110 6108 -1092
rect 6162 -1058 6280 -1040
rect 6390 -1010 6508 -992
rect 6562 -958 6680 -940
rect 6562 -992 6570 -958
rect 6604 -992 6638 -958
rect 6672 -992 6680 -958
rect 6562 -1010 6680 -992
rect 6790 -958 6908 -940
rect 6790 -992 6798 -958
rect 6832 -992 6866 -958
rect 6900 -992 6908 -958
rect 6790 -1010 6908 -992
rect 6962 -958 7080 -940
rect 7190 -910 7308 -892
rect 7362 -858 7480 -846
rect 7362 -892 7370 -858
rect 7404 -892 7438 -858
rect 7472 -892 7480 -858
rect 7362 -910 7480 -892
rect 7590 -858 7708 -846
rect 7590 -892 7598 -858
rect 7632 -892 7666 -858
rect 7700 -892 7708 -858
rect 7590 -910 7708 -892
rect 7762 -858 7880 -846
rect 7762 -892 7770 -858
rect 7804 -892 7838 -858
rect 7872 -892 7880 -858
rect 7762 -910 7880 -892
rect 7990 -858 8108 -846
rect 7990 -892 7998 -858
rect 8032 -892 8066 -858
rect 8100 -892 8108 -858
rect 6962 -992 6970 -958
rect 7004 -992 7038 -958
rect 7072 -992 7080 -958
rect 6962 -1010 7080 -992
rect 7190 -958 7308 -940
rect 7190 -992 7198 -958
rect 7232 -992 7266 -958
rect 7300 -992 7308 -958
rect 6162 -1092 6170 -1058
rect 6204 -1092 6238 -1058
rect 6272 -1092 6280 -1058
rect 6162 -1110 6280 -1092
rect 6390 -1058 6508 -1040
rect 6390 -1092 6398 -1058
rect 6432 -1092 6466 -1058
rect 6500 -1092 6508 -1058
rect 5362 -1192 5370 -1158
rect 5404 -1192 5438 -1158
rect 5472 -1192 5480 -1158
rect 5362 -1210 5480 -1192
rect 5590 -1158 5708 -1140
rect 5590 -1192 5598 -1158
rect 5632 -1192 5666 -1158
rect 5700 -1192 5708 -1158
rect 4562 -1292 4570 -1258
rect 4604 -1292 4638 -1258
rect 4672 -1292 4680 -1258
rect 4562 -1310 4680 -1292
rect 4790 -1258 4908 -1240
rect 4790 -1292 4798 -1258
rect 4832 -1292 4866 -1258
rect 4900 -1292 4908 -1258
rect 3762 -1392 3770 -1358
rect 3804 -1392 3838 -1358
rect 3872 -1392 3880 -1358
rect 3762 -1410 3880 -1392
rect 3990 -1358 4108 -1340
rect 3990 -1392 3998 -1358
rect 4032 -1392 4066 -1358
rect 4100 -1392 4108 -1358
rect 2962 -1492 2970 -1458
rect 3004 -1492 3038 -1458
rect 3072 -1492 3080 -1458
rect 2962 -1510 3080 -1492
rect 3190 -1458 3308 -1440
rect 3190 -1492 3198 -1458
rect 3232 -1492 3266 -1458
rect 3300 -1492 3308 -1458
rect 2162 -1592 2170 -1558
rect 2204 -1592 2238 -1558
rect 2272 -1592 2280 -1558
rect 2162 -1610 2280 -1592
rect 2390 -1558 2508 -1540
rect 2390 -1592 2398 -1558
rect 2432 -1592 2466 -1558
rect 2500 -1592 2508 -1558
rect 1362 -1692 1370 -1658
rect 1404 -1692 1438 -1658
rect 1472 -1692 1480 -1658
rect 1362 -1710 1480 -1692
rect 1590 -1658 1708 -1640
rect 1590 -1692 1598 -1658
rect 1632 -1692 1666 -1658
rect 1700 -1692 1708 -1658
rect 562 -1792 570 -1758
rect 604 -1792 638 -1758
rect 672 -1792 680 -1758
rect 562 -1810 680 -1792
rect 790 -1758 908 -1740
rect 790 -1792 798 -1758
rect 832 -1792 866 -1758
rect 900 -1792 908 -1758
rect -10 -1858 108 -1840
rect -10 -1892 -2 -1858
rect 32 -1892 66 -1858
rect 100 -1892 108 -1858
rect -10 -1910 108 -1892
rect 162 -1858 280 -1840
rect 162 -1892 170 -1858
rect 204 -1892 238 -1858
rect 272 -1892 280 -1858
rect 162 -1910 280 -1892
rect 390 -1858 508 -1840
rect 390 -1892 398 -1858
rect 432 -1892 466 -1858
rect 500 -1892 508 -1858
rect 390 -1910 508 -1892
rect 562 -1858 680 -1840
rect 790 -1810 908 -1792
rect 962 -1758 1080 -1740
rect 962 -1792 970 -1758
rect 1004 -1792 1038 -1758
rect 1072 -1792 1080 -1758
rect 962 -1810 1080 -1792
rect 1190 -1758 1308 -1740
rect 1190 -1792 1198 -1758
rect 1232 -1792 1266 -1758
rect 1300 -1792 1308 -1758
rect 1190 -1810 1308 -1792
rect 1362 -1758 1480 -1740
rect 1590 -1710 1708 -1692
rect 1762 -1658 1880 -1640
rect 1762 -1692 1770 -1658
rect 1804 -1692 1838 -1658
rect 1872 -1692 1880 -1658
rect 1762 -1710 1880 -1692
rect 1990 -1658 2108 -1640
rect 1990 -1692 1998 -1658
rect 2032 -1692 2066 -1658
rect 2100 -1692 2108 -1658
rect 1990 -1710 2108 -1692
rect 2162 -1658 2280 -1640
rect 2390 -1610 2508 -1592
rect 2562 -1558 2680 -1540
rect 2562 -1592 2570 -1558
rect 2604 -1592 2638 -1558
rect 2672 -1592 2680 -1558
rect 2562 -1610 2680 -1592
rect 2790 -1558 2908 -1540
rect 2790 -1592 2798 -1558
rect 2832 -1592 2866 -1558
rect 2900 -1592 2908 -1558
rect 2790 -1610 2908 -1592
rect 2962 -1558 3080 -1540
rect 3190 -1510 3308 -1492
rect 3362 -1458 3480 -1440
rect 3362 -1492 3370 -1458
rect 3404 -1492 3438 -1458
rect 3472 -1492 3480 -1458
rect 3362 -1510 3480 -1492
rect 3590 -1458 3708 -1440
rect 3590 -1492 3598 -1458
rect 3632 -1492 3666 -1458
rect 3700 -1492 3708 -1458
rect 3590 -1510 3708 -1492
rect 3762 -1458 3880 -1440
rect 3990 -1410 4108 -1392
rect 4162 -1358 4280 -1340
rect 4162 -1392 4170 -1358
rect 4204 -1392 4238 -1358
rect 4272 -1392 4280 -1358
rect 4162 -1410 4280 -1392
rect 4390 -1358 4508 -1340
rect 4390 -1392 4398 -1358
rect 4432 -1392 4466 -1358
rect 4500 -1392 4508 -1358
rect 4390 -1410 4508 -1392
rect 4562 -1358 4680 -1340
rect 4790 -1310 4908 -1292
rect 4962 -1258 5080 -1240
rect 4962 -1292 4970 -1258
rect 5004 -1292 5038 -1258
rect 5072 -1292 5080 -1258
rect 4962 -1310 5080 -1292
rect 5190 -1258 5308 -1240
rect 5190 -1292 5198 -1258
rect 5232 -1292 5266 -1258
rect 5300 -1292 5308 -1258
rect 5190 -1310 5308 -1292
rect 5362 -1258 5480 -1240
rect 5590 -1210 5708 -1192
rect 5762 -1158 5880 -1140
rect 5762 -1192 5770 -1158
rect 5804 -1192 5838 -1158
rect 5872 -1192 5880 -1158
rect 5762 -1210 5880 -1192
rect 5990 -1158 6108 -1140
rect 5990 -1192 5998 -1158
rect 6032 -1192 6066 -1158
rect 6100 -1192 6108 -1158
rect 5990 -1210 6108 -1192
rect 6162 -1158 6280 -1140
rect 6390 -1110 6508 -1092
rect 6562 -1058 6680 -1040
rect 6562 -1092 6570 -1058
rect 6604 -1092 6638 -1058
rect 6672 -1092 6680 -1058
rect 6562 -1110 6680 -1092
rect 6790 -1058 6908 -1040
rect 6790 -1092 6798 -1058
rect 6832 -1092 6866 -1058
rect 6900 -1092 6908 -1058
rect 6790 -1110 6908 -1092
rect 6962 -1058 7080 -1040
rect 7190 -1010 7308 -992
rect 7362 -958 7480 -940
rect 7362 -992 7370 -958
rect 7404 -992 7438 -958
rect 7472 -992 7480 -958
rect 7362 -1010 7480 -992
rect 7590 -958 7708 -940
rect 7590 -992 7598 -958
rect 7632 -992 7666 -958
rect 7700 -992 7708 -958
rect 7590 -1010 7708 -992
rect 7762 -958 7880 -940
rect 7990 -910 8108 -892
rect 8162 -858 8280 -846
rect 8162 -892 8170 -858
rect 8204 -892 8238 -858
rect 8272 -892 8280 -858
rect 8162 -910 8280 -892
rect 8390 -858 8508 -846
rect 8390 -892 8398 -858
rect 8432 -892 8466 -858
rect 8500 -892 8508 -858
rect 8390 -910 8508 -892
rect 8562 -858 8680 -846
rect 8562 -892 8570 -858
rect 8604 -892 8638 -858
rect 8672 -892 8680 -858
rect 8562 -910 8680 -892
rect 8790 -858 8908 -846
rect 8790 -892 8798 -858
rect 8832 -892 8866 -858
rect 8900 -892 8908 -858
rect 7762 -992 7770 -958
rect 7804 -992 7838 -958
rect 7872 -992 7880 -958
rect 7762 -1010 7880 -992
rect 7990 -958 8108 -940
rect 7990 -992 7998 -958
rect 8032 -992 8066 -958
rect 8100 -992 8108 -958
rect 6962 -1092 6970 -1058
rect 7004 -1092 7038 -1058
rect 7072 -1092 7080 -1058
rect 6962 -1110 7080 -1092
rect 7190 -1058 7308 -1040
rect 7190 -1092 7198 -1058
rect 7232 -1092 7266 -1058
rect 7300 -1092 7308 -1058
rect 6162 -1192 6170 -1158
rect 6204 -1192 6238 -1158
rect 6272 -1192 6280 -1158
rect 6162 -1210 6280 -1192
rect 6390 -1158 6508 -1140
rect 6390 -1192 6398 -1158
rect 6432 -1192 6466 -1158
rect 6500 -1192 6508 -1158
rect 5362 -1292 5370 -1258
rect 5404 -1292 5438 -1258
rect 5472 -1292 5480 -1258
rect 5362 -1310 5480 -1292
rect 5590 -1258 5708 -1240
rect 5590 -1292 5598 -1258
rect 5632 -1292 5666 -1258
rect 5700 -1292 5708 -1258
rect 4562 -1392 4570 -1358
rect 4604 -1392 4638 -1358
rect 4672 -1392 4680 -1358
rect 4562 -1410 4680 -1392
rect 4790 -1358 4908 -1340
rect 4790 -1392 4798 -1358
rect 4832 -1392 4866 -1358
rect 4900 -1392 4908 -1358
rect 3762 -1492 3770 -1458
rect 3804 -1492 3838 -1458
rect 3872 -1492 3880 -1458
rect 3762 -1510 3880 -1492
rect 3990 -1458 4108 -1440
rect 3990 -1492 3998 -1458
rect 4032 -1492 4066 -1458
rect 4100 -1492 4108 -1458
rect 2962 -1592 2970 -1558
rect 3004 -1592 3038 -1558
rect 3072 -1592 3080 -1558
rect 2962 -1610 3080 -1592
rect 3190 -1558 3308 -1540
rect 3190 -1592 3198 -1558
rect 3232 -1592 3266 -1558
rect 3300 -1592 3308 -1558
rect 2162 -1692 2170 -1658
rect 2204 -1692 2238 -1658
rect 2272 -1692 2280 -1658
rect 2162 -1710 2280 -1692
rect 2390 -1658 2508 -1640
rect 2390 -1692 2398 -1658
rect 2432 -1692 2466 -1658
rect 2500 -1692 2508 -1658
rect 1362 -1792 1370 -1758
rect 1404 -1792 1438 -1758
rect 1472 -1792 1480 -1758
rect 1362 -1810 1480 -1792
rect 1590 -1758 1708 -1740
rect 1590 -1792 1598 -1758
rect 1632 -1792 1666 -1758
rect 1700 -1792 1708 -1758
rect 562 -1892 570 -1858
rect 604 -1892 638 -1858
rect 672 -1892 680 -1858
rect 562 -1910 680 -1892
rect 790 -1858 908 -1840
rect 790 -1892 798 -1858
rect 832 -1892 866 -1858
rect 900 -1892 908 -1858
rect -10 -1958 108 -1940
rect -10 -1992 -2 -1958
rect 32 -1992 66 -1958
rect 100 -1992 108 -1958
rect -10 -2010 108 -1992
rect 162 -1958 280 -1940
rect 162 -1992 170 -1958
rect 204 -1992 238 -1958
rect 272 -1992 280 -1958
rect 162 -2010 280 -1992
rect 390 -1958 508 -1940
rect 390 -1992 398 -1958
rect 432 -1992 466 -1958
rect 500 -1992 508 -1958
rect 390 -2010 508 -1992
rect 562 -1958 680 -1940
rect 790 -1910 908 -1892
rect 962 -1858 1080 -1840
rect 962 -1892 970 -1858
rect 1004 -1892 1038 -1858
rect 1072 -1892 1080 -1858
rect 962 -1910 1080 -1892
rect 1190 -1858 1308 -1840
rect 1190 -1892 1198 -1858
rect 1232 -1892 1266 -1858
rect 1300 -1892 1308 -1858
rect 1190 -1910 1308 -1892
rect 1362 -1858 1480 -1840
rect 1590 -1810 1708 -1792
rect 1762 -1758 1880 -1740
rect 1762 -1792 1770 -1758
rect 1804 -1792 1838 -1758
rect 1872 -1792 1880 -1758
rect 1762 -1810 1880 -1792
rect 1990 -1758 2108 -1740
rect 1990 -1792 1998 -1758
rect 2032 -1792 2066 -1758
rect 2100 -1792 2108 -1758
rect 1990 -1810 2108 -1792
rect 2162 -1758 2280 -1740
rect 2390 -1710 2508 -1692
rect 2562 -1658 2680 -1640
rect 2562 -1692 2570 -1658
rect 2604 -1692 2638 -1658
rect 2672 -1692 2680 -1658
rect 2562 -1710 2680 -1692
rect 2790 -1658 2908 -1640
rect 2790 -1692 2798 -1658
rect 2832 -1692 2866 -1658
rect 2900 -1692 2908 -1658
rect 2790 -1710 2908 -1692
rect 2962 -1658 3080 -1640
rect 3190 -1610 3308 -1592
rect 3362 -1558 3480 -1540
rect 3362 -1592 3370 -1558
rect 3404 -1592 3438 -1558
rect 3472 -1592 3480 -1558
rect 3362 -1610 3480 -1592
rect 3590 -1558 3708 -1540
rect 3590 -1592 3598 -1558
rect 3632 -1592 3666 -1558
rect 3700 -1592 3708 -1558
rect 3590 -1610 3708 -1592
rect 3762 -1558 3880 -1540
rect 3990 -1510 4108 -1492
rect 4162 -1458 4280 -1440
rect 4162 -1492 4170 -1458
rect 4204 -1492 4238 -1458
rect 4272 -1492 4280 -1458
rect 4162 -1510 4280 -1492
rect 4390 -1458 4508 -1440
rect 4390 -1492 4398 -1458
rect 4432 -1492 4466 -1458
rect 4500 -1492 4508 -1458
rect 4390 -1510 4508 -1492
rect 4562 -1458 4680 -1440
rect 4790 -1410 4908 -1392
rect 4962 -1358 5080 -1340
rect 4962 -1392 4970 -1358
rect 5004 -1392 5038 -1358
rect 5072 -1392 5080 -1358
rect 4962 -1410 5080 -1392
rect 5190 -1358 5308 -1340
rect 5190 -1392 5198 -1358
rect 5232 -1392 5266 -1358
rect 5300 -1392 5308 -1358
rect 5190 -1410 5308 -1392
rect 5362 -1358 5480 -1340
rect 5590 -1310 5708 -1292
rect 5762 -1258 5880 -1240
rect 5762 -1292 5770 -1258
rect 5804 -1292 5838 -1258
rect 5872 -1292 5880 -1258
rect 5762 -1310 5880 -1292
rect 5990 -1258 6108 -1240
rect 5990 -1292 5998 -1258
rect 6032 -1292 6066 -1258
rect 6100 -1292 6108 -1258
rect 5990 -1310 6108 -1292
rect 6162 -1258 6280 -1240
rect 6390 -1210 6508 -1192
rect 6562 -1158 6680 -1140
rect 6562 -1192 6570 -1158
rect 6604 -1192 6638 -1158
rect 6672 -1192 6680 -1158
rect 6562 -1210 6680 -1192
rect 6790 -1158 6908 -1140
rect 6790 -1192 6798 -1158
rect 6832 -1192 6866 -1158
rect 6900 -1192 6908 -1158
rect 6790 -1210 6908 -1192
rect 6962 -1158 7080 -1140
rect 7190 -1110 7308 -1092
rect 7362 -1058 7480 -1040
rect 7362 -1092 7370 -1058
rect 7404 -1092 7438 -1058
rect 7472 -1092 7480 -1058
rect 7362 -1110 7480 -1092
rect 7590 -1058 7708 -1040
rect 7590 -1092 7598 -1058
rect 7632 -1092 7666 -1058
rect 7700 -1092 7708 -1058
rect 7590 -1110 7708 -1092
rect 7762 -1058 7880 -1040
rect 7990 -1010 8108 -992
rect 8162 -958 8280 -940
rect 8162 -992 8170 -958
rect 8204 -992 8238 -958
rect 8272 -992 8280 -958
rect 8162 -1010 8280 -992
rect 8390 -958 8508 -940
rect 8390 -992 8398 -958
rect 8432 -992 8466 -958
rect 8500 -992 8508 -958
rect 8390 -1010 8508 -992
rect 8562 -958 8680 -940
rect 8790 -910 8908 -892
rect 8962 -858 9080 -846
rect 8962 -892 8970 -858
rect 9004 -892 9038 -858
rect 9072 -892 9080 -858
rect 8962 -910 9080 -892
rect 9190 -858 9308 -846
rect 9190 -892 9198 -858
rect 9232 -892 9266 -858
rect 9300 -892 9308 -858
rect 9190 -910 9308 -892
rect 9362 -858 9480 -846
rect 9362 -892 9370 -858
rect 9404 -892 9438 -858
rect 9472 -892 9480 -858
rect 9362 -910 9480 -892
rect 9590 -858 9708 -846
rect 9590 -892 9598 -858
rect 9632 -892 9666 -858
rect 9700 -892 9708 -858
rect 8562 -992 8570 -958
rect 8604 -992 8638 -958
rect 8672 -992 8680 -958
rect 8562 -1010 8680 -992
rect 8790 -958 8908 -940
rect 8790 -992 8798 -958
rect 8832 -992 8866 -958
rect 8900 -992 8908 -958
rect 7762 -1092 7770 -1058
rect 7804 -1092 7838 -1058
rect 7872 -1092 7880 -1058
rect 7762 -1110 7880 -1092
rect 7990 -1058 8108 -1040
rect 7990 -1092 7998 -1058
rect 8032 -1092 8066 -1058
rect 8100 -1092 8108 -1058
rect 6962 -1192 6970 -1158
rect 7004 -1192 7038 -1158
rect 7072 -1192 7080 -1158
rect 6962 -1210 7080 -1192
rect 7190 -1158 7308 -1140
rect 7190 -1192 7198 -1158
rect 7232 -1192 7266 -1158
rect 7300 -1192 7308 -1158
rect 6162 -1292 6170 -1258
rect 6204 -1292 6238 -1258
rect 6272 -1292 6280 -1258
rect 6162 -1310 6280 -1292
rect 6390 -1258 6508 -1240
rect 6390 -1292 6398 -1258
rect 6432 -1292 6466 -1258
rect 6500 -1292 6508 -1258
rect 5362 -1392 5370 -1358
rect 5404 -1392 5438 -1358
rect 5472 -1392 5480 -1358
rect 5362 -1410 5480 -1392
rect 5590 -1358 5708 -1340
rect 5590 -1392 5598 -1358
rect 5632 -1392 5666 -1358
rect 5700 -1392 5708 -1358
rect 4562 -1492 4570 -1458
rect 4604 -1492 4638 -1458
rect 4672 -1492 4680 -1458
rect 4562 -1510 4680 -1492
rect 4790 -1458 4908 -1440
rect 4790 -1492 4798 -1458
rect 4832 -1492 4866 -1458
rect 4900 -1492 4908 -1458
rect 3762 -1592 3770 -1558
rect 3804 -1592 3838 -1558
rect 3872 -1592 3880 -1558
rect 3762 -1610 3880 -1592
rect 3990 -1558 4108 -1540
rect 3990 -1592 3998 -1558
rect 4032 -1592 4066 -1558
rect 4100 -1592 4108 -1558
rect 2962 -1692 2970 -1658
rect 3004 -1692 3038 -1658
rect 3072 -1692 3080 -1658
rect 2962 -1710 3080 -1692
rect 3190 -1658 3308 -1640
rect 3190 -1692 3198 -1658
rect 3232 -1692 3266 -1658
rect 3300 -1692 3308 -1658
rect 2162 -1792 2170 -1758
rect 2204 -1792 2238 -1758
rect 2272 -1792 2280 -1758
rect 2162 -1810 2280 -1792
rect 2390 -1758 2508 -1740
rect 2390 -1792 2398 -1758
rect 2432 -1792 2466 -1758
rect 2500 -1792 2508 -1758
rect 1362 -1892 1370 -1858
rect 1404 -1892 1438 -1858
rect 1472 -1892 1480 -1858
rect 1362 -1910 1480 -1892
rect 1590 -1858 1708 -1840
rect 1590 -1892 1598 -1858
rect 1632 -1892 1666 -1858
rect 1700 -1892 1708 -1858
rect 562 -1992 570 -1958
rect 604 -1992 638 -1958
rect 672 -1992 680 -1958
rect 562 -2010 680 -1992
rect 790 -1958 908 -1940
rect 790 -1992 798 -1958
rect 832 -1992 866 -1958
rect 900 -1992 908 -1958
rect -10 -2058 108 -2040
rect -10 -2092 -2 -2058
rect 32 -2092 66 -2058
rect 100 -2092 108 -2058
rect -10 -2129 108 -2092
rect 162 -2058 280 -2040
rect 162 -2092 170 -2058
rect 204 -2092 238 -2058
rect 272 -2092 280 -2058
rect 162 -2129 280 -2092
rect 390 -2058 508 -2040
rect 390 -2092 398 -2058
rect 432 -2092 466 -2058
rect 500 -2092 508 -2058
rect 390 -2129 508 -2092
rect 562 -2058 680 -2040
rect 790 -2010 908 -1992
rect 962 -1958 1080 -1940
rect 962 -1992 970 -1958
rect 1004 -1992 1038 -1958
rect 1072 -1992 1080 -1958
rect 962 -2010 1080 -1992
rect 1190 -1958 1308 -1940
rect 1190 -1992 1198 -1958
rect 1232 -1992 1266 -1958
rect 1300 -1992 1308 -1958
rect 1190 -2010 1308 -1992
rect 1362 -1958 1480 -1940
rect 1590 -1910 1708 -1892
rect 1762 -1858 1880 -1840
rect 1762 -1892 1770 -1858
rect 1804 -1892 1838 -1858
rect 1872 -1892 1880 -1858
rect 1762 -1910 1880 -1892
rect 1990 -1858 2108 -1840
rect 1990 -1892 1998 -1858
rect 2032 -1892 2066 -1858
rect 2100 -1892 2108 -1858
rect 1990 -1910 2108 -1892
rect 2162 -1858 2280 -1840
rect 2390 -1810 2508 -1792
rect 2562 -1758 2680 -1740
rect 2562 -1792 2570 -1758
rect 2604 -1792 2638 -1758
rect 2672 -1792 2680 -1758
rect 2562 -1810 2680 -1792
rect 2790 -1758 2908 -1740
rect 2790 -1792 2798 -1758
rect 2832 -1792 2866 -1758
rect 2900 -1792 2908 -1758
rect 2790 -1810 2908 -1792
rect 2962 -1758 3080 -1740
rect 3190 -1710 3308 -1692
rect 3362 -1658 3480 -1640
rect 3362 -1692 3370 -1658
rect 3404 -1692 3438 -1658
rect 3472 -1692 3480 -1658
rect 3362 -1710 3480 -1692
rect 3590 -1658 3708 -1640
rect 3590 -1692 3598 -1658
rect 3632 -1692 3666 -1658
rect 3700 -1692 3708 -1658
rect 3590 -1710 3708 -1692
rect 3762 -1658 3880 -1640
rect 3990 -1610 4108 -1592
rect 4162 -1558 4280 -1540
rect 4162 -1592 4170 -1558
rect 4204 -1592 4238 -1558
rect 4272 -1592 4280 -1558
rect 4162 -1610 4280 -1592
rect 4390 -1558 4508 -1540
rect 4390 -1592 4398 -1558
rect 4432 -1592 4466 -1558
rect 4500 -1592 4508 -1558
rect 4390 -1610 4508 -1592
rect 4562 -1558 4680 -1540
rect 4790 -1510 4908 -1492
rect 4962 -1458 5080 -1440
rect 4962 -1492 4970 -1458
rect 5004 -1492 5038 -1458
rect 5072 -1492 5080 -1458
rect 4962 -1510 5080 -1492
rect 5190 -1458 5308 -1440
rect 5190 -1492 5198 -1458
rect 5232 -1492 5266 -1458
rect 5300 -1492 5308 -1458
rect 5190 -1510 5308 -1492
rect 5362 -1458 5480 -1440
rect 5590 -1410 5708 -1392
rect 5762 -1358 5880 -1340
rect 5762 -1392 5770 -1358
rect 5804 -1392 5838 -1358
rect 5872 -1392 5880 -1358
rect 5762 -1410 5880 -1392
rect 5990 -1358 6108 -1340
rect 5990 -1392 5998 -1358
rect 6032 -1392 6066 -1358
rect 6100 -1392 6108 -1358
rect 5990 -1410 6108 -1392
rect 6162 -1358 6280 -1340
rect 6390 -1310 6508 -1292
rect 6562 -1258 6680 -1240
rect 6562 -1292 6570 -1258
rect 6604 -1292 6638 -1258
rect 6672 -1292 6680 -1258
rect 6562 -1310 6680 -1292
rect 6790 -1258 6908 -1240
rect 6790 -1292 6798 -1258
rect 6832 -1292 6866 -1258
rect 6900 -1292 6908 -1258
rect 6790 -1310 6908 -1292
rect 6962 -1258 7080 -1240
rect 7190 -1210 7308 -1192
rect 7362 -1158 7480 -1140
rect 7362 -1192 7370 -1158
rect 7404 -1192 7438 -1158
rect 7472 -1192 7480 -1158
rect 7362 -1210 7480 -1192
rect 7590 -1158 7708 -1140
rect 7590 -1192 7598 -1158
rect 7632 -1192 7666 -1158
rect 7700 -1192 7708 -1158
rect 7590 -1210 7708 -1192
rect 7762 -1158 7880 -1140
rect 7990 -1110 8108 -1092
rect 8162 -1058 8280 -1040
rect 8162 -1092 8170 -1058
rect 8204 -1092 8238 -1058
rect 8272 -1092 8280 -1058
rect 8162 -1110 8280 -1092
rect 8390 -1058 8508 -1040
rect 8390 -1092 8398 -1058
rect 8432 -1092 8466 -1058
rect 8500 -1092 8508 -1058
rect 8390 -1110 8508 -1092
rect 8562 -1058 8680 -1040
rect 8790 -1010 8908 -992
rect 8962 -958 9080 -940
rect 8962 -992 8970 -958
rect 9004 -992 9038 -958
rect 9072 -992 9080 -958
rect 8962 -1010 9080 -992
rect 9190 -958 9308 -940
rect 9190 -992 9198 -958
rect 9232 -992 9266 -958
rect 9300 -992 9308 -958
rect 9190 -1010 9308 -992
rect 9362 -958 9480 -940
rect 9590 -910 9708 -892
rect 9762 -858 9880 -846
rect 9762 -892 9770 -858
rect 9804 -892 9838 -858
rect 9872 -892 9880 -858
rect 9762 -910 9880 -892
rect 9990 -858 10108 -846
rect 9990 -892 9998 -858
rect 10032 -892 10066 -858
rect 10100 -892 10108 -858
rect 9990 -910 10108 -892
rect 10162 -858 10280 -846
rect 10162 -892 10170 -858
rect 10204 -892 10238 -858
rect 10272 -892 10280 -858
rect 10162 -910 10280 -892
rect 10390 -858 10508 -846
rect 10390 -892 10398 -858
rect 10432 -892 10466 -858
rect 10500 -892 10508 -858
rect 9362 -992 9370 -958
rect 9404 -992 9438 -958
rect 9472 -992 9480 -958
rect 9362 -1010 9480 -992
rect 9590 -958 9708 -940
rect 9590 -992 9598 -958
rect 9632 -992 9666 -958
rect 9700 -992 9708 -958
rect 8562 -1092 8570 -1058
rect 8604 -1092 8638 -1058
rect 8672 -1092 8680 -1058
rect 8562 -1110 8680 -1092
rect 8790 -1058 8908 -1040
rect 8790 -1092 8798 -1058
rect 8832 -1092 8866 -1058
rect 8900 -1092 8908 -1058
rect 7762 -1192 7770 -1158
rect 7804 -1192 7838 -1158
rect 7872 -1192 7880 -1158
rect 7762 -1210 7880 -1192
rect 7990 -1158 8108 -1140
rect 7990 -1192 7998 -1158
rect 8032 -1192 8066 -1158
rect 8100 -1192 8108 -1158
rect 6962 -1292 6970 -1258
rect 7004 -1292 7038 -1258
rect 7072 -1292 7080 -1258
rect 6962 -1310 7080 -1292
rect 7190 -1258 7308 -1240
rect 7190 -1292 7198 -1258
rect 7232 -1292 7266 -1258
rect 7300 -1292 7308 -1258
rect 6162 -1392 6170 -1358
rect 6204 -1392 6238 -1358
rect 6272 -1392 6280 -1358
rect 6162 -1410 6280 -1392
rect 6390 -1358 6508 -1340
rect 6390 -1392 6398 -1358
rect 6432 -1392 6466 -1358
rect 6500 -1392 6508 -1358
rect 5362 -1492 5370 -1458
rect 5404 -1492 5438 -1458
rect 5472 -1492 5480 -1458
rect 5362 -1510 5480 -1492
rect 5590 -1458 5708 -1440
rect 5590 -1492 5598 -1458
rect 5632 -1492 5666 -1458
rect 5700 -1492 5708 -1458
rect 4562 -1592 4570 -1558
rect 4604 -1592 4638 -1558
rect 4672 -1592 4680 -1558
rect 4562 -1610 4680 -1592
rect 4790 -1558 4908 -1540
rect 4790 -1592 4798 -1558
rect 4832 -1592 4866 -1558
rect 4900 -1592 4908 -1558
rect 3762 -1692 3770 -1658
rect 3804 -1692 3838 -1658
rect 3872 -1692 3880 -1658
rect 3762 -1710 3880 -1692
rect 3990 -1658 4108 -1640
rect 3990 -1692 3998 -1658
rect 4032 -1692 4066 -1658
rect 4100 -1692 4108 -1658
rect 2962 -1792 2970 -1758
rect 3004 -1792 3038 -1758
rect 3072 -1792 3080 -1758
rect 2962 -1810 3080 -1792
rect 3190 -1758 3308 -1740
rect 3190 -1792 3198 -1758
rect 3232 -1792 3266 -1758
rect 3300 -1792 3308 -1758
rect 2162 -1892 2170 -1858
rect 2204 -1892 2238 -1858
rect 2272 -1892 2280 -1858
rect 2162 -1910 2280 -1892
rect 2390 -1858 2508 -1840
rect 2390 -1892 2398 -1858
rect 2432 -1892 2466 -1858
rect 2500 -1892 2508 -1858
rect 1362 -1992 1370 -1958
rect 1404 -1992 1438 -1958
rect 1472 -1992 1480 -1958
rect 1362 -2010 1480 -1992
rect 1590 -1958 1708 -1940
rect 1590 -1992 1598 -1958
rect 1632 -1992 1666 -1958
rect 1700 -1992 1708 -1958
rect 562 -2092 570 -2058
rect 604 -2092 638 -2058
rect 672 -2092 680 -2058
rect 562 -2129 680 -2092
rect 790 -2058 908 -2040
rect 790 -2092 798 -2058
rect 832 -2092 866 -2058
rect 900 -2092 908 -2058
rect 790 -2129 908 -2092
rect 962 -2058 1080 -2040
rect 962 -2092 970 -2058
rect 1004 -2092 1038 -2058
rect 1072 -2092 1080 -2058
rect 962 -2129 1080 -2092
rect 1190 -2058 1308 -2040
rect 1190 -2092 1198 -2058
rect 1232 -2092 1266 -2058
rect 1300 -2092 1308 -2058
rect 1190 -2129 1308 -2092
rect 1362 -2058 1480 -2040
rect 1590 -2010 1708 -1992
rect 1762 -1958 1880 -1940
rect 1762 -1992 1770 -1958
rect 1804 -1992 1838 -1958
rect 1872 -1992 1880 -1958
rect 1762 -2010 1880 -1992
rect 1990 -1958 2108 -1940
rect 1990 -1992 1998 -1958
rect 2032 -1992 2066 -1958
rect 2100 -1992 2108 -1958
rect 1990 -2010 2108 -1992
rect 2162 -1958 2280 -1940
rect 2390 -1910 2508 -1892
rect 2562 -1858 2680 -1840
rect 2562 -1892 2570 -1858
rect 2604 -1892 2638 -1858
rect 2672 -1892 2680 -1858
rect 2562 -1910 2680 -1892
rect 2790 -1858 2908 -1840
rect 2790 -1892 2798 -1858
rect 2832 -1892 2866 -1858
rect 2900 -1892 2908 -1858
rect 2790 -1910 2908 -1892
rect 2962 -1858 3080 -1840
rect 3190 -1810 3308 -1792
rect 3362 -1758 3480 -1740
rect 3362 -1792 3370 -1758
rect 3404 -1792 3438 -1758
rect 3472 -1792 3480 -1758
rect 3362 -1810 3480 -1792
rect 3590 -1758 3708 -1740
rect 3590 -1792 3598 -1758
rect 3632 -1792 3666 -1758
rect 3700 -1792 3708 -1758
rect 3590 -1810 3708 -1792
rect 3762 -1758 3880 -1740
rect 3990 -1710 4108 -1692
rect 4162 -1658 4280 -1640
rect 4162 -1692 4170 -1658
rect 4204 -1692 4238 -1658
rect 4272 -1692 4280 -1658
rect 4162 -1710 4280 -1692
rect 4390 -1658 4508 -1640
rect 4390 -1692 4398 -1658
rect 4432 -1692 4466 -1658
rect 4500 -1692 4508 -1658
rect 4390 -1710 4508 -1692
rect 4562 -1658 4680 -1640
rect 4790 -1610 4908 -1592
rect 4962 -1558 5080 -1540
rect 4962 -1592 4970 -1558
rect 5004 -1592 5038 -1558
rect 5072 -1592 5080 -1558
rect 4962 -1610 5080 -1592
rect 5190 -1558 5308 -1540
rect 5190 -1592 5198 -1558
rect 5232 -1592 5266 -1558
rect 5300 -1592 5308 -1558
rect 5190 -1610 5308 -1592
rect 5362 -1558 5480 -1540
rect 5590 -1510 5708 -1492
rect 5762 -1458 5880 -1440
rect 5762 -1492 5770 -1458
rect 5804 -1492 5838 -1458
rect 5872 -1492 5880 -1458
rect 5762 -1510 5880 -1492
rect 5990 -1458 6108 -1440
rect 5990 -1492 5998 -1458
rect 6032 -1492 6066 -1458
rect 6100 -1492 6108 -1458
rect 5990 -1510 6108 -1492
rect 6162 -1458 6280 -1440
rect 6390 -1410 6508 -1392
rect 6562 -1358 6680 -1340
rect 6562 -1392 6570 -1358
rect 6604 -1392 6638 -1358
rect 6672 -1392 6680 -1358
rect 6562 -1410 6680 -1392
rect 6790 -1358 6908 -1340
rect 6790 -1392 6798 -1358
rect 6832 -1392 6866 -1358
rect 6900 -1392 6908 -1358
rect 6790 -1410 6908 -1392
rect 6962 -1358 7080 -1340
rect 7190 -1310 7308 -1292
rect 7362 -1258 7480 -1240
rect 7362 -1292 7370 -1258
rect 7404 -1292 7438 -1258
rect 7472 -1292 7480 -1258
rect 7362 -1310 7480 -1292
rect 7590 -1258 7708 -1240
rect 7590 -1292 7598 -1258
rect 7632 -1292 7666 -1258
rect 7700 -1292 7708 -1258
rect 7590 -1310 7708 -1292
rect 7762 -1258 7880 -1240
rect 7990 -1210 8108 -1192
rect 8162 -1158 8280 -1140
rect 8162 -1192 8170 -1158
rect 8204 -1192 8238 -1158
rect 8272 -1192 8280 -1158
rect 8162 -1210 8280 -1192
rect 8390 -1158 8508 -1140
rect 8390 -1192 8398 -1158
rect 8432 -1192 8466 -1158
rect 8500 -1192 8508 -1158
rect 8390 -1210 8508 -1192
rect 8562 -1158 8680 -1140
rect 8790 -1110 8908 -1092
rect 8962 -1058 9080 -1040
rect 8962 -1092 8970 -1058
rect 9004 -1092 9038 -1058
rect 9072 -1092 9080 -1058
rect 8962 -1110 9080 -1092
rect 9190 -1058 9308 -1040
rect 9190 -1092 9198 -1058
rect 9232 -1092 9266 -1058
rect 9300 -1092 9308 -1058
rect 9190 -1110 9308 -1092
rect 9362 -1058 9480 -1040
rect 9590 -1010 9708 -992
rect 9762 -958 9880 -940
rect 9762 -992 9770 -958
rect 9804 -992 9838 -958
rect 9872 -992 9880 -958
rect 9762 -1010 9880 -992
rect 9990 -958 10108 -940
rect 9990 -992 9998 -958
rect 10032 -992 10066 -958
rect 10100 -992 10108 -958
rect 9990 -1010 10108 -992
rect 10162 -958 10280 -940
rect 10390 -910 10508 -892
rect 10562 -858 10680 -846
rect 10562 -892 10570 -858
rect 10604 -892 10638 -858
rect 10672 -892 10680 -858
rect 10562 -910 10680 -892
rect 10790 -858 10908 -846
rect 10790 -892 10798 -858
rect 10832 -892 10866 -858
rect 10900 -892 10908 -858
rect 10790 -910 10908 -892
rect 10962 -858 11080 -846
rect 10962 -892 10970 -858
rect 11004 -892 11038 -858
rect 11072 -892 11080 -858
rect 10962 -910 11080 -892
rect 11190 -858 11308 -846
rect 11190 -892 11198 -858
rect 11232 -892 11266 -858
rect 11300 -892 11308 -858
rect 10162 -992 10170 -958
rect 10204 -992 10238 -958
rect 10272 -992 10280 -958
rect 10162 -1010 10280 -992
rect 10390 -958 10508 -940
rect 10390 -992 10398 -958
rect 10432 -992 10466 -958
rect 10500 -992 10508 -958
rect 9362 -1092 9370 -1058
rect 9404 -1092 9438 -1058
rect 9472 -1092 9480 -1058
rect 9362 -1110 9480 -1092
rect 9590 -1058 9708 -1040
rect 9590 -1092 9598 -1058
rect 9632 -1092 9666 -1058
rect 9700 -1092 9708 -1058
rect 8562 -1192 8570 -1158
rect 8604 -1192 8638 -1158
rect 8672 -1192 8680 -1158
rect 8562 -1210 8680 -1192
rect 8790 -1158 8908 -1140
rect 8790 -1192 8798 -1158
rect 8832 -1192 8866 -1158
rect 8900 -1192 8908 -1158
rect 7762 -1292 7770 -1258
rect 7804 -1292 7838 -1258
rect 7872 -1292 7880 -1258
rect 7762 -1310 7880 -1292
rect 7990 -1258 8108 -1240
rect 7990 -1292 7998 -1258
rect 8032 -1292 8066 -1258
rect 8100 -1292 8108 -1258
rect 6962 -1392 6970 -1358
rect 7004 -1392 7038 -1358
rect 7072 -1392 7080 -1358
rect 6962 -1410 7080 -1392
rect 7190 -1358 7308 -1340
rect 7190 -1392 7198 -1358
rect 7232 -1392 7266 -1358
rect 7300 -1392 7308 -1358
rect 6162 -1492 6170 -1458
rect 6204 -1492 6238 -1458
rect 6272 -1492 6280 -1458
rect 6162 -1510 6280 -1492
rect 6390 -1458 6508 -1440
rect 6390 -1492 6398 -1458
rect 6432 -1492 6466 -1458
rect 6500 -1492 6508 -1458
rect 5362 -1592 5370 -1558
rect 5404 -1592 5438 -1558
rect 5472 -1592 5480 -1558
rect 5362 -1610 5480 -1592
rect 5590 -1558 5708 -1540
rect 5590 -1592 5598 -1558
rect 5632 -1592 5666 -1558
rect 5700 -1592 5708 -1558
rect 4562 -1692 4570 -1658
rect 4604 -1692 4638 -1658
rect 4672 -1692 4680 -1658
rect 4562 -1710 4680 -1692
rect 4790 -1658 4908 -1640
rect 4790 -1692 4798 -1658
rect 4832 -1692 4866 -1658
rect 4900 -1692 4908 -1658
rect 3762 -1792 3770 -1758
rect 3804 -1792 3838 -1758
rect 3872 -1792 3880 -1758
rect 3762 -1810 3880 -1792
rect 3990 -1758 4108 -1740
rect 3990 -1792 3998 -1758
rect 4032 -1792 4066 -1758
rect 4100 -1792 4108 -1758
rect 2962 -1892 2970 -1858
rect 3004 -1892 3038 -1858
rect 3072 -1892 3080 -1858
rect 2962 -1910 3080 -1892
rect 3190 -1858 3308 -1840
rect 3190 -1892 3198 -1858
rect 3232 -1892 3266 -1858
rect 3300 -1892 3308 -1858
rect 2162 -1992 2170 -1958
rect 2204 -1992 2238 -1958
rect 2272 -1992 2280 -1958
rect 2162 -2010 2280 -1992
rect 2390 -1958 2508 -1940
rect 2390 -1992 2398 -1958
rect 2432 -1992 2466 -1958
rect 2500 -1992 2508 -1958
rect 1362 -2092 1370 -2058
rect 1404 -2092 1438 -2058
rect 1472 -2092 1480 -2058
rect 1362 -2129 1480 -2092
rect 1590 -2058 1708 -2040
rect 1590 -2092 1598 -2058
rect 1632 -2092 1666 -2058
rect 1700 -2092 1708 -2058
rect 1590 -2129 1708 -2092
rect 1762 -2058 1880 -2040
rect 1762 -2092 1770 -2058
rect 1804 -2092 1838 -2058
rect 1872 -2092 1880 -2058
rect 1762 -2129 1880 -2092
rect 1990 -2058 2108 -2040
rect 1990 -2092 1998 -2058
rect 2032 -2092 2066 -2058
rect 2100 -2092 2108 -2058
rect 1990 -2129 2108 -2092
rect 2162 -2058 2280 -2040
rect 2390 -2010 2508 -1992
rect 2562 -1958 2680 -1940
rect 2562 -1992 2570 -1958
rect 2604 -1992 2638 -1958
rect 2672 -1992 2680 -1958
rect 2562 -2010 2680 -1992
rect 2790 -1958 2908 -1940
rect 2790 -1992 2798 -1958
rect 2832 -1992 2866 -1958
rect 2900 -1992 2908 -1958
rect 2790 -2010 2908 -1992
rect 2962 -1958 3080 -1940
rect 3190 -1910 3308 -1892
rect 3362 -1858 3480 -1840
rect 3362 -1892 3370 -1858
rect 3404 -1892 3438 -1858
rect 3472 -1892 3480 -1858
rect 3362 -1910 3480 -1892
rect 3590 -1858 3708 -1840
rect 3590 -1892 3598 -1858
rect 3632 -1892 3666 -1858
rect 3700 -1892 3708 -1858
rect 3590 -1910 3708 -1892
rect 3762 -1858 3880 -1840
rect 3990 -1810 4108 -1792
rect 4162 -1758 4280 -1740
rect 4162 -1792 4170 -1758
rect 4204 -1792 4238 -1758
rect 4272 -1792 4280 -1758
rect 4162 -1810 4280 -1792
rect 4390 -1758 4508 -1740
rect 4390 -1792 4398 -1758
rect 4432 -1792 4466 -1758
rect 4500 -1792 4508 -1758
rect 4390 -1810 4508 -1792
rect 4562 -1758 4680 -1740
rect 4790 -1710 4908 -1692
rect 4962 -1658 5080 -1640
rect 4962 -1692 4970 -1658
rect 5004 -1692 5038 -1658
rect 5072 -1692 5080 -1658
rect 4962 -1710 5080 -1692
rect 5190 -1658 5308 -1640
rect 5190 -1692 5198 -1658
rect 5232 -1692 5266 -1658
rect 5300 -1692 5308 -1658
rect 5190 -1710 5308 -1692
rect 5362 -1658 5480 -1640
rect 5590 -1610 5708 -1592
rect 5762 -1558 5880 -1540
rect 5762 -1592 5770 -1558
rect 5804 -1592 5838 -1558
rect 5872 -1592 5880 -1558
rect 5762 -1610 5880 -1592
rect 5990 -1558 6108 -1540
rect 5990 -1592 5998 -1558
rect 6032 -1592 6066 -1558
rect 6100 -1592 6108 -1558
rect 5990 -1610 6108 -1592
rect 6162 -1558 6280 -1540
rect 6390 -1510 6508 -1492
rect 6562 -1458 6680 -1440
rect 6562 -1492 6570 -1458
rect 6604 -1492 6638 -1458
rect 6672 -1492 6680 -1458
rect 6562 -1510 6680 -1492
rect 6790 -1458 6908 -1440
rect 6790 -1492 6798 -1458
rect 6832 -1492 6866 -1458
rect 6900 -1492 6908 -1458
rect 6790 -1510 6908 -1492
rect 6962 -1458 7080 -1440
rect 7190 -1410 7308 -1392
rect 7362 -1358 7480 -1340
rect 7362 -1392 7370 -1358
rect 7404 -1392 7438 -1358
rect 7472 -1392 7480 -1358
rect 7362 -1410 7480 -1392
rect 7590 -1358 7708 -1340
rect 7590 -1392 7598 -1358
rect 7632 -1392 7666 -1358
rect 7700 -1392 7708 -1358
rect 7590 -1410 7708 -1392
rect 7762 -1358 7880 -1340
rect 7990 -1310 8108 -1292
rect 8162 -1258 8280 -1240
rect 8162 -1292 8170 -1258
rect 8204 -1292 8238 -1258
rect 8272 -1292 8280 -1258
rect 8162 -1310 8280 -1292
rect 8390 -1258 8508 -1240
rect 8390 -1292 8398 -1258
rect 8432 -1292 8466 -1258
rect 8500 -1292 8508 -1258
rect 8390 -1310 8508 -1292
rect 8562 -1258 8680 -1240
rect 8790 -1210 8908 -1192
rect 8962 -1158 9080 -1140
rect 8962 -1192 8970 -1158
rect 9004 -1192 9038 -1158
rect 9072 -1192 9080 -1158
rect 8962 -1210 9080 -1192
rect 9190 -1158 9308 -1140
rect 9190 -1192 9198 -1158
rect 9232 -1192 9266 -1158
rect 9300 -1192 9308 -1158
rect 9190 -1210 9308 -1192
rect 9362 -1158 9480 -1140
rect 9590 -1110 9708 -1092
rect 9762 -1058 9880 -1040
rect 9762 -1092 9770 -1058
rect 9804 -1092 9838 -1058
rect 9872 -1092 9880 -1058
rect 9762 -1110 9880 -1092
rect 9990 -1058 10108 -1040
rect 9990 -1092 9998 -1058
rect 10032 -1092 10066 -1058
rect 10100 -1092 10108 -1058
rect 9990 -1110 10108 -1092
rect 10162 -1058 10280 -1040
rect 10390 -1010 10508 -992
rect 10562 -958 10680 -940
rect 10562 -992 10570 -958
rect 10604 -992 10638 -958
rect 10672 -992 10680 -958
rect 10562 -1010 10680 -992
rect 10790 -958 10908 -940
rect 10790 -992 10798 -958
rect 10832 -992 10866 -958
rect 10900 -992 10908 -958
rect 10790 -1010 10908 -992
rect 10962 -958 11080 -940
rect 11190 -910 11308 -892
rect 11362 -858 11480 -846
rect 11362 -892 11370 -858
rect 11404 -892 11438 -858
rect 11472 -892 11480 -858
rect 11362 -910 11480 -892
rect 11590 -858 11708 -846
rect 11590 -892 11598 -858
rect 11632 -892 11666 -858
rect 11700 -892 11708 -858
rect 11590 -910 11708 -892
rect 11762 -858 11880 -846
rect 11762 -892 11770 -858
rect 11804 -892 11838 -858
rect 11872 -892 11880 -858
rect 11762 -910 11880 -892
rect 11990 -858 12108 -846
rect 11990 -892 11998 -858
rect 12032 -892 12066 -858
rect 12100 -892 12108 -858
rect 10962 -992 10970 -958
rect 11004 -992 11038 -958
rect 11072 -992 11080 -958
rect 10962 -1010 11080 -992
rect 11190 -958 11308 -940
rect 11190 -992 11198 -958
rect 11232 -992 11266 -958
rect 11300 -992 11308 -958
rect 10162 -1092 10170 -1058
rect 10204 -1092 10238 -1058
rect 10272 -1092 10280 -1058
rect 10162 -1110 10280 -1092
rect 10390 -1058 10508 -1040
rect 10390 -1092 10398 -1058
rect 10432 -1092 10466 -1058
rect 10500 -1092 10508 -1058
rect 9362 -1192 9370 -1158
rect 9404 -1192 9438 -1158
rect 9472 -1192 9480 -1158
rect 9362 -1210 9480 -1192
rect 9590 -1158 9708 -1140
rect 9590 -1192 9598 -1158
rect 9632 -1192 9666 -1158
rect 9700 -1192 9708 -1158
rect 8562 -1292 8570 -1258
rect 8604 -1292 8638 -1258
rect 8672 -1292 8680 -1258
rect 8562 -1310 8680 -1292
rect 8790 -1258 8908 -1240
rect 8790 -1292 8798 -1258
rect 8832 -1292 8866 -1258
rect 8900 -1292 8908 -1258
rect 7762 -1392 7770 -1358
rect 7804 -1392 7838 -1358
rect 7872 -1392 7880 -1358
rect 7762 -1410 7880 -1392
rect 7990 -1358 8108 -1340
rect 7990 -1392 7998 -1358
rect 8032 -1392 8066 -1358
rect 8100 -1392 8108 -1358
rect 6962 -1492 6970 -1458
rect 7004 -1492 7038 -1458
rect 7072 -1492 7080 -1458
rect 6962 -1510 7080 -1492
rect 7190 -1458 7308 -1440
rect 7190 -1492 7198 -1458
rect 7232 -1492 7266 -1458
rect 7300 -1492 7308 -1458
rect 6162 -1592 6170 -1558
rect 6204 -1592 6238 -1558
rect 6272 -1592 6280 -1558
rect 6162 -1610 6280 -1592
rect 6390 -1558 6508 -1540
rect 6390 -1592 6398 -1558
rect 6432 -1592 6466 -1558
rect 6500 -1592 6508 -1558
rect 5362 -1692 5370 -1658
rect 5404 -1692 5438 -1658
rect 5472 -1692 5480 -1658
rect 5362 -1710 5480 -1692
rect 5590 -1658 5708 -1640
rect 5590 -1692 5598 -1658
rect 5632 -1692 5666 -1658
rect 5700 -1692 5708 -1658
rect 4562 -1792 4570 -1758
rect 4604 -1792 4638 -1758
rect 4672 -1792 4680 -1758
rect 4562 -1810 4680 -1792
rect 4790 -1758 4908 -1740
rect 4790 -1792 4798 -1758
rect 4832 -1792 4866 -1758
rect 4900 -1792 4908 -1758
rect 3762 -1892 3770 -1858
rect 3804 -1892 3838 -1858
rect 3872 -1892 3880 -1858
rect 3762 -1910 3880 -1892
rect 3990 -1858 4108 -1840
rect 3990 -1892 3998 -1858
rect 4032 -1892 4066 -1858
rect 4100 -1892 4108 -1858
rect 2962 -1992 2970 -1958
rect 3004 -1992 3038 -1958
rect 3072 -1992 3080 -1958
rect 2962 -2010 3080 -1992
rect 3190 -1958 3308 -1940
rect 3190 -1992 3198 -1958
rect 3232 -1992 3266 -1958
rect 3300 -1992 3308 -1958
rect 2162 -2092 2170 -2058
rect 2204 -2092 2238 -2058
rect 2272 -2092 2280 -2058
rect 2162 -2129 2280 -2092
rect 2390 -2058 2508 -2040
rect 2390 -2092 2398 -2058
rect 2432 -2092 2466 -2058
rect 2500 -2092 2508 -2058
rect 2390 -2129 2508 -2092
rect 2562 -2058 2680 -2040
rect 2562 -2092 2570 -2058
rect 2604 -2092 2638 -2058
rect 2672 -2092 2680 -2058
rect 2562 -2129 2680 -2092
rect 2790 -2058 2908 -2040
rect 2790 -2092 2798 -2058
rect 2832 -2092 2866 -2058
rect 2900 -2092 2908 -2058
rect 2790 -2129 2908 -2092
rect 2962 -2058 3080 -2040
rect 3190 -2010 3308 -1992
rect 3362 -1958 3480 -1940
rect 3362 -1992 3370 -1958
rect 3404 -1992 3438 -1958
rect 3472 -1992 3480 -1958
rect 3362 -2010 3480 -1992
rect 3590 -1958 3708 -1940
rect 3590 -1992 3598 -1958
rect 3632 -1992 3666 -1958
rect 3700 -1992 3708 -1958
rect 3590 -2010 3708 -1992
rect 3762 -1958 3880 -1940
rect 3990 -1910 4108 -1892
rect 4162 -1858 4280 -1840
rect 4162 -1892 4170 -1858
rect 4204 -1892 4238 -1858
rect 4272 -1892 4280 -1858
rect 4162 -1910 4280 -1892
rect 4390 -1858 4508 -1840
rect 4390 -1892 4398 -1858
rect 4432 -1892 4466 -1858
rect 4500 -1892 4508 -1858
rect 4390 -1910 4508 -1892
rect 4562 -1858 4680 -1840
rect 4790 -1810 4908 -1792
rect 4962 -1758 5080 -1740
rect 4962 -1792 4970 -1758
rect 5004 -1792 5038 -1758
rect 5072 -1792 5080 -1758
rect 4962 -1810 5080 -1792
rect 5190 -1758 5308 -1740
rect 5190 -1792 5198 -1758
rect 5232 -1792 5266 -1758
rect 5300 -1792 5308 -1758
rect 5190 -1810 5308 -1792
rect 5362 -1758 5480 -1740
rect 5590 -1710 5708 -1692
rect 5762 -1658 5880 -1640
rect 5762 -1692 5770 -1658
rect 5804 -1692 5838 -1658
rect 5872 -1692 5880 -1658
rect 5762 -1710 5880 -1692
rect 5990 -1658 6108 -1640
rect 5990 -1692 5998 -1658
rect 6032 -1692 6066 -1658
rect 6100 -1692 6108 -1658
rect 5990 -1710 6108 -1692
rect 6162 -1658 6280 -1640
rect 6390 -1610 6508 -1592
rect 6562 -1558 6680 -1540
rect 6562 -1592 6570 -1558
rect 6604 -1592 6638 -1558
rect 6672 -1592 6680 -1558
rect 6562 -1610 6680 -1592
rect 6790 -1558 6908 -1540
rect 6790 -1592 6798 -1558
rect 6832 -1592 6866 -1558
rect 6900 -1592 6908 -1558
rect 6790 -1610 6908 -1592
rect 6962 -1558 7080 -1540
rect 7190 -1510 7308 -1492
rect 7362 -1458 7480 -1440
rect 7362 -1492 7370 -1458
rect 7404 -1492 7438 -1458
rect 7472 -1492 7480 -1458
rect 7362 -1510 7480 -1492
rect 7590 -1458 7708 -1440
rect 7590 -1492 7598 -1458
rect 7632 -1492 7666 -1458
rect 7700 -1492 7708 -1458
rect 7590 -1510 7708 -1492
rect 7762 -1458 7880 -1440
rect 7990 -1410 8108 -1392
rect 8162 -1358 8280 -1340
rect 8162 -1392 8170 -1358
rect 8204 -1392 8238 -1358
rect 8272 -1392 8280 -1358
rect 8162 -1410 8280 -1392
rect 8390 -1358 8508 -1340
rect 8390 -1392 8398 -1358
rect 8432 -1392 8466 -1358
rect 8500 -1392 8508 -1358
rect 8390 -1410 8508 -1392
rect 8562 -1358 8680 -1340
rect 8790 -1310 8908 -1292
rect 8962 -1258 9080 -1240
rect 8962 -1292 8970 -1258
rect 9004 -1292 9038 -1258
rect 9072 -1292 9080 -1258
rect 8962 -1310 9080 -1292
rect 9190 -1258 9308 -1240
rect 9190 -1292 9198 -1258
rect 9232 -1292 9266 -1258
rect 9300 -1292 9308 -1258
rect 9190 -1310 9308 -1292
rect 9362 -1258 9480 -1240
rect 9590 -1210 9708 -1192
rect 9762 -1158 9880 -1140
rect 9762 -1192 9770 -1158
rect 9804 -1192 9838 -1158
rect 9872 -1192 9880 -1158
rect 9762 -1210 9880 -1192
rect 9990 -1158 10108 -1140
rect 9990 -1192 9998 -1158
rect 10032 -1192 10066 -1158
rect 10100 -1192 10108 -1158
rect 9990 -1210 10108 -1192
rect 10162 -1158 10280 -1140
rect 10390 -1110 10508 -1092
rect 10562 -1058 10680 -1040
rect 10562 -1092 10570 -1058
rect 10604 -1092 10638 -1058
rect 10672 -1092 10680 -1058
rect 10562 -1110 10680 -1092
rect 10790 -1058 10908 -1040
rect 10790 -1092 10798 -1058
rect 10832 -1092 10866 -1058
rect 10900 -1092 10908 -1058
rect 10790 -1110 10908 -1092
rect 10962 -1058 11080 -1040
rect 11190 -1010 11308 -992
rect 11362 -958 11480 -940
rect 11362 -992 11370 -958
rect 11404 -992 11438 -958
rect 11472 -992 11480 -958
rect 11362 -1010 11480 -992
rect 11590 -958 11708 -940
rect 11590 -992 11598 -958
rect 11632 -992 11666 -958
rect 11700 -992 11708 -958
rect 11590 -1010 11708 -992
rect 11762 -958 11880 -940
rect 11990 -910 12108 -892
rect 12162 -858 12280 -846
rect 12162 -892 12170 -858
rect 12204 -892 12238 -858
rect 12272 -892 12280 -858
rect 12162 -910 12280 -892
rect 12390 -858 12508 -846
rect 12390 -892 12398 -858
rect 12432 -892 12466 -858
rect 12500 -892 12508 -858
rect 12390 -910 12508 -892
rect 12562 -858 12680 -846
rect 12562 -892 12570 -858
rect 12604 -892 12638 -858
rect 12672 -892 12680 -858
rect 14540 -860 14690 -842
rect 15652 -808 15802 -790
rect 15652 -842 15678 -808
rect 15712 -842 15746 -808
rect 15780 -842 15802 -808
rect 15652 -860 15802 -842
rect 12562 -910 12680 -892
rect 11762 -992 11770 -958
rect 11804 -992 11838 -958
rect 11872 -992 11880 -958
rect 11762 -1010 11880 -992
rect 11990 -958 12108 -940
rect 11990 -992 11998 -958
rect 12032 -992 12066 -958
rect 12100 -992 12108 -958
rect 10962 -1092 10970 -1058
rect 11004 -1092 11038 -1058
rect 11072 -1092 11080 -1058
rect 10962 -1110 11080 -1092
rect 11190 -1058 11308 -1040
rect 11190 -1092 11198 -1058
rect 11232 -1092 11266 -1058
rect 11300 -1092 11308 -1058
rect 10162 -1192 10170 -1158
rect 10204 -1192 10238 -1158
rect 10272 -1192 10280 -1158
rect 10162 -1210 10280 -1192
rect 10390 -1158 10508 -1140
rect 10390 -1192 10398 -1158
rect 10432 -1192 10466 -1158
rect 10500 -1192 10508 -1158
rect 9362 -1292 9370 -1258
rect 9404 -1292 9438 -1258
rect 9472 -1292 9480 -1258
rect 9362 -1310 9480 -1292
rect 9590 -1258 9708 -1240
rect 9590 -1292 9598 -1258
rect 9632 -1292 9666 -1258
rect 9700 -1292 9708 -1258
rect 8562 -1392 8570 -1358
rect 8604 -1392 8638 -1358
rect 8672 -1392 8680 -1358
rect 8562 -1410 8680 -1392
rect 8790 -1358 8908 -1340
rect 8790 -1392 8798 -1358
rect 8832 -1392 8866 -1358
rect 8900 -1392 8908 -1358
rect 7762 -1492 7770 -1458
rect 7804 -1492 7838 -1458
rect 7872 -1492 7880 -1458
rect 7762 -1510 7880 -1492
rect 7990 -1458 8108 -1440
rect 7990 -1492 7998 -1458
rect 8032 -1492 8066 -1458
rect 8100 -1492 8108 -1458
rect 6962 -1592 6970 -1558
rect 7004 -1592 7038 -1558
rect 7072 -1592 7080 -1558
rect 6962 -1610 7080 -1592
rect 7190 -1558 7308 -1540
rect 7190 -1592 7198 -1558
rect 7232 -1592 7266 -1558
rect 7300 -1592 7308 -1558
rect 6162 -1692 6170 -1658
rect 6204 -1692 6238 -1658
rect 6272 -1692 6280 -1658
rect 6162 -1710 6280 -1692
rect 6390 -1658 6508 -1640
rect 6390 -1692 6398 -1658
rect 6432 -1692 6466 -1658
rect 6500 -1692 6508 -1658
rect 5362 -1792 5370 -1758
rect 5404 -1792 5438 -1758
rect 5472 -1792 5480 -1758
rect 5362 -1810 5480 -1792
rect 5590 -1758 5708 -1740
rect 5590 -1792 5598 -1758
rect 5632 -1792 5666 -1758
rect 5700 -1792 5708 -1758
rect 4562 -1892 4570 -1858
rect 4604 -1892 4638 -1858
rect 4672 -1892 4680 -1858
rect 4562 -1910 4680 -1892
rect 4790 -1858 4908 -1840
rect 4790 -1892 4798 -1858
rect 4832 -1892 4866 -1858
rect 4900 -1892 4908 -1858
rect 3762 -1992 3770 -1958
rect 3804 -1992 3838 -1958
rect 3872 -1992 3880 -1958
rect 3762 -2010 3880 -1992
rect 3990 -1958 4108 -1940
rect 3990 -1992 3998 -1958
rect 4032 -1992 4066 -1958
rect 4100 -1992 4108 -1958
rect 2962 -2092 2970 -2058
rect 3004 -2092 3038 -2058
rect 3072 -2092 3080 -2058
rect 2962 -2129 3080 -2092
rect 3190 -2058 3308 -2040
rect 3190 -2092 3198 -2058
rect 3232 -2092 3266 -2058
rect 3300 -2092 3308 -2058
rect 3190 -2129 3308 -2092
rect 3362 -2058 3480 -2040
rect 3362 -2092 3370 -2058
rect 3404 -2092 3438 -2058
rect 3472 -2092 3480 -2058
rect 3362 -2129 3480 -2092
rect 3590 -2058 3708 -2040
rect 3590 -2092 3598 -2058
rect 3632 -2092 3666 -2058
rect 3700 -2092 3708 -2058
rect 3590 -2129 3708 -2092
rect 3762 -2058 3880 -2040
rect 3990 -2010 4108 -1992
rect 4162 -1958 4280 -1940
rect 4162 -1992 4170 -1958
rect 4204 -1992 4238 -1958
rect 4272 -1992 4280 -1958
rect 4162 -2010 4280 -1992
rect 4390 -1958 4508 -1940
rect 4390 -1992 4398 -1958
rect 4432 -1992 4466 -1958
rect 4500 -1992 4508 -1958
rect 4390 -2010 4508 -1992
rect 4562 -1958 4680 -1940
rect 4790 -1910 4908 -1892
rect 4962 -1858 5080 -1840
rect 4962 -1892 4970 -1858
rect 5004 -1892 5038 -1858
rect 5072 -1892 5080 -1858
rect 4962 -1910 5080 -1892
rect 5190 -1858 5308 -1840
rect 5190 -1892 5198 -1858
rect 5232 -1892 5266 -1858
rect 5300 -1892 5308 -1858
rect 5190 -1910 5308 -1892
rect 5362 -1858 5480 -1840
rect 5590 -1810 5708 -1792
rect 5762 -1758 5880 -1740
rect 5762 -1792 5770 -1758
rect 5804 -1792 5838 -1758
rect 5872 -1792 5880 -1758
rect 5762 -1810 5880 -1792
rect 5990 -1758 6108 -1740
rect 5990 -1792 5998 -1758
rect 6032 -1792 6066 -1758
rect 6100 -1792 6108 -1758
rect 5990 -1810 6108 -1792
rect 6162 -1758 6280 -1740
rect 6390 -1710 6508 -1692
rect 6562 -1658 6680 -1640
rect 6562 -1692 6570 -1658
rect 6604 -1692 6638 -1658
rect 6672 -1692 6680 -1658
rect 6562 -1710 6680 -1692
rect 6790 -1658 6908 -1640
rect 6790 -1692 6798 -1658
rect 6832 -1692 6866 -1658
rect 6900 -1692 6908 -1658
rect 6790 -1710 6908 -1692
rect 6962 -1658 7080 -1640
rect 7190 -1610 7308 -1592
rect 7362 -1558 7480 -1540
rect 7362 -1592 7370 -1558
rect 7404 -1592 7438 -1558
rect 7472 -1592 7480 -1558
rect 7362 -1610 7480 -1592
rect 7590 -1558 7708 -1540
rect 7590 -1592 7598 -1558
rect 7632 -1592 7666 -1558
rect 7700 -1592 7708 -1558
rect 7590 -1610 7708 -1592
rect 7762 -1558 7880 -1540
rect 7990 -1510 8108 -1492
rect 8162 -1458 8280 -1440
rect 8162 -1492 8170 -1458
rect 8204 -1492 8238 -1458
rect 8272 -1492 8280 -1458
rect 8162 -1510 8280 -1492
rect 8390 -1458 8508 -1440
rect 8390 -1492 8398 -1458
rect 8432 -1492 8466 -1458
rect 8500 -1492 8508 -1458
rect 8390 -1510 8508 -1492
rect 8562 -1458 8680 -1440
rect 8790 -1410 8908 -1392
rect 8962 -1358 9080 -1340
rect 8962 -1392 8970 -1358
rect 9004 -1392 9038 -1358
rect 9072 -1392 9080 -1358
rect 8962 -1410 9080 -1392
rect 9190 -1358 9308 -1340
rect 9190 -1392 9198 -1358
rect 9232 -1392 9266 -1358
rect 9300 -1392 9308 -1358
rect 9190 -1410 9308 -1392
rect 9362 -1358 9480 -1340
rect 9590 -1310 9708 -1292
rect 9762 -1258 9880 -1240
rect 9762 -1292 9770 -1258
rect 9804 -1292 9838 -1258
rect 9872 -1292 9880 -1258
rect 9762 -1310 9880 -1292
rect 9990 -1258 10108 -1240
rect 9990 -1292 9998 -1258
rect 10032 -1292 10066 -1258
rect 10100 -1292 10108 -1258
rect 9990 -1310 10108 -1292
rect 10162 -1258 10280 -1240
rect 10390 -1210 10508 -1192
rect 10562 -1158 10680 -1140
rect 10562 -1192 10570 -1158
rect 10604 -1192 10638 -1158
rect 10672 -1192 10680 -1158
rect 10562 -1210 10680 -1192
rect 10790 -1158 10908 -1140
rect 10790 -1192 10798 -1158
rect 10832 -1192 10866 -1158
rect 10900 -1192 10908 -1158
rect 10790 -1210 10908 -1192
rect 10962 -1158 11080 -1140
rect 11190 -1110 11308 -1092
rect 11362 -1058 11480 -1040
rect 11362 -1092 11370 -1058
rect 11404 -1092 11438 -1058
rect 11472 -1092 11480 -1058
rect 11362 -1110 11480 -1092
rect 11590 -1058 11708 -1040
rect 11590 -1092 11598 -1058
rect 11632 -1092 11666 -1058
rect 11700 -1092 11708 -1058
rect 11590 -1110 11708 -1092
rect 11762 -1058 11880 -1040
rect 11990 -1010 12108 -992
rect 12162 -958 12280 -940
rect 12162 -992 12170 -958
rect 12204 -992 12238 -958
rect 12272 -992 12280 -958
rect 12162 -1010 12280 -992
rect 12390 -958 12508 -940
rect 12390 -992 12398 -958
rect 12432 -992 12466 -958
rect 12500 -992 12508 -958
rect 12390 -1010 12508 -992
rect 12562 -958 12680 -940
rect 14540 -908 14690 -890
rect 14540 -942 14562 -908
rect 14596 -942 14630 -908
rect 14664 -942 14690 -908
rect 12562 -992 12570 -958
rect 12604 -992 12638 -958
rect 12672 -992 12680 -958
rect 14540 -960 14690 -942
rect 15652 -908 15802 -890
rect 15652 -942 15678 -908
rect 15712 -942 15746 -908
rect 15780 -942 15802 -908
rect 15652 -960 15802 -942
rect 12562 -1010 12680 -992
rect 11762 -1092 11770 -1058
rect 11804 -1092 11838 -1058
rect 11872 -1092 11880 -1058
rect 11762 -1110 11880 -1092
rect 11990 -1058 12108 -1040
rect 11990 -1092 11998 -1058
rect 12032 -1092 12066 -1058
rect 12100 -1092 12108 -1058
rect 10962 -1192 10970 -1158
rect 11004 -1192 11038 -1158
rect 11072 -1192 11080 -1158
rect 10962 -1210 11080 -1192
rect 11190 -1158 11308 -1140
rect 11190 -1192 11198 -1158
rect 11232 -1192 11266 -1158
rect 11300 -1192 11308 -1158
rect 10162 -1292 10170 -1258
rect 10204 -1292 10238 -1258
rect 10272 -1292 10280 -1258
rect 10162 -1310 10280 -1292
rect 10390 -1258 10508 -1240
rect 10390 -1292 10398 -1258
rect 10432 -1292 10466 -1258
rect 10500 -1292 10508 -1258
rect 9362 -1392 9370 -1358
rect 9404 -1392 9438 -1358
rect 9472 -1392 9480 -1358
rect 9362 -1410 9480 -1392
rect 9590 -1358 9708 -1340
rect 9590 -1392 9598 -1358
rect 9632 -1392 9666 -1358
rect 9700 -1392 9708 -1358
rect 8562 -1492 8570 -1458
rect 8604 -1492 8638 -1458
rect 8672 -1492 8680 -1458
rect 8562 -1510 8680 -1492
rect 8790 -1458 8908 -1440
rect 8790 -1492 8798 -1458
rect 8832 -1492 8866 -1458
rect 8900 -1492 8908 -1458
rect 7762 -1592 7770 -1558
rect 7804 -1592 7838 -1558
rect 7872 -1592 7880 -1558
rect 7762 -1610 7880 -1592
rect 7990 -1558 8108 -1540
rect 7990 -1592 7998 -1558
rect 8032 -1592 8066 -1558
rect 8100 -1592 8108 -1558
rect 6962 -1692 6970 -1658
rect 7004 -1692 7038 -1658
rect 7072 -1692 7080 -1658
rect 6962 -1710 7080 -1692
rect 7190 -1658 7308 -1640
rect 7190 -1692 7198 -1658
rect 7232 -1692 7266 -1658
rect 7300 -1692 7308 -1658
rect 6162 -1792 6170 -1758
rect 6204 -1792 6238 -1758
rect 6272 -1792 6280 -1758
rect 6162 -1810 6280 -1792
rect 6390 -1758 6508 -1740
rect 6390 -1792 6398 -1758
rect 6432 -1792 6466 -1758
rect 6500 -1792 6508 -1758
rect 5362 -1892 5370 -1858
rect 5404 -1892 5438 -1858
rect 5472 -1892 5480 -1858
rect 5362 -1910 5480 -1892
rect 5590 -1858 5708 -1840
rect 5590 -1892 5598 -1858
rect 5632 -1892 5666 -1858
rect 5700 -1892 5708 -1858
rect 4562 -1992 4570 -1958
rect 4604 -1992 4638 -1958
rect 4672 -1992 4680 -1958
rect 4562 -2010 4680 -1992
rect 4790 -1958 4908 -1940
rect 4790 -1992 4798 -1958
rect 4832 -1992 4866 -1958
rect 4900 -1992 4908 -1958
rect 3762 -2092 3770 -2058
rect 3804 -2092 3838 -2058
rect 3872 -2092 3880 -2058
rect 3762 -2129 3880 -2092
rect 3990 -2058 4108 -2040
rect 3990 -2092 3998 -2058
rect 4032 -2092 4066 -2058
rect 4100 -2092 4108 -2058
rect 3990 -2129 4108 -2092
rect 4162 -2058 4280 -2040
rect 4162 -2092 4170 -2058
rect 4204 -2092 4238 -2058
rect 4272 -2092 4280 -2058
rect 4162 -2129 4280 -2092
rect 4390 -2058 4508 -2040
rect 4390 -2092 4398 -2058
rect 4432 -2092 4466 -2058
rect 4500 -2092 4508 -2058
rect 4390 -2129 4508 -2092
rect 4562 -2058 4680 -2040
rect 4790 -2010 4908 -1992
rect 4962 -1958 5080 -1940
rect 4962 -1992 4970 -1958
rect 5004 -1992 5038 -1958
rect 5072 -1992 5080 -1958
rect 4962 -2010 5080 -1992
rect 5190 -1958 5308 -1940
rect 5190 -1992 5198 -1958
rect 5232 -1992 5266 -1958
rect 5300 -1992 5308 -1958
rect 5190 -2010 5308 -1992
rect 5362 -1958 5480 -1940
rect 5590 -1910 5708 -1892
rect 5762 -1858 5880 -1840
rect 5762 -1892 5770 -1858
rect 5804 -1892 5838 -1858
rect 5872 -1892 5880 -1858
rect 5762 -1910 5880 -1892
rect 5990 -1858 6108 -1840
rect 5990 -1892 5998 -1858
rect 6032 -1892 6066 -1858
rect 6100 -1892 6108 -1858
rect 5990 -1910 6108 -1892
rect 6162 -1858 6280 -1840
rect 6390 -1810 6508 -1792
rect 6562 -1758 6680 -1740
rect 6562 -1792 6570 -1758
rect 6604 -1792 6638 -1758
rect 6672 -1792 6680 -1758
rect 6562 -1810 6680 -1792
rect 6790 -1758 6908 -1740
rect 6790 -1792 6798 -1758
rect 6832 -1792 6866 -1758
rect 6900 -1792 6908 -1758
rect 6790 -1810 6908 -1792
rect 6962 -1758 7080 -1740
rect 7190 -1710 7308 -1692
rect 7362 -1658 7480 -1640
rect 7362 -1692 7370 -1658
rect 7404 -1692 7438 -1658
rect 7472 -1692 7480 -1658
rect 7362 -1710 7480 -1692
rect 7590 -1658 7708 -1640
rect 7590 -1692 7598 -1658
rect 7632 -1692 7666 -1658
rect 7700 -1692 7708 -1658
rect 7590 -1710 7708 -1692
rect 7762 -1658 7880 -1640
rect 7990 -1610 8108 -1592
rect 8162 -1558 8280 -1540
rect 8162 -1592 8170 -1558
rect 8204 -1592 8238 -1558
rect 8272 -1592 8280 -1558
rect 8162 -1610 8280 -1592
rect 8390 -1558 8508 -1540
rect 8390 -1592 8398 -1558
rect 8432 -1592 8466 -1558
rect 8500 -1592 8508 -1558
rect 8390 -1610 8508 -1592
rect 8562 -1558 8680 -1540
rect 8790 -1510 8908 -1492
rect 8962 -1458 9080 -1440
rect 8962 -1492 8970 -1458
rect 9004 -1492 9038 -1458
rect 9072 -1492 9080 -1458
rect 8962 -1510 9080 -1492
rect 9190 -1458 9308 -1440
rect 9190 -1492 9198 -1458
rect 9232 -1492 9266 -1458
rect 9300 -1492 9308 -1458
rect 9190 -1510 9308 -1492
rect 9362 -1458 9480 -1440
rect 9590 -1410 9708 -1392
rect 9762 -1358 9880 -1340
rect 9762 -1392 9770 -1358
rect 9804 -1392 9838 -1358
rect 9872 -1392 9880 -1358
rect 9762 -1410 9880 -1392
rect 9990 -1358 10108 -1340
rect 9990 -1392 9998 -1358
rect 10032 -1392 10066 -1358
rect 10100 -1392 10108 -1358
rect 9990 -1410 10108 -1392
rect 10162 -1358 10280 -1340
rect 10390 -1310 10508 -1292
rect 10562 -1258 10680 -1240
rect 10562 -1292 10570 -1258
rect 10604 -1292 10638 -1258
rect 10672 -1292 10680 -1258
rect 10562 -1310 10680 -1292
rect 10790 -1258 10908 -1240
rect 10790 -1292 10798 -1258
rect 10832 -1292 10866 -1258
rect 10900 -1292 10908 -1258
rect 10790 -1310 10908 -1292
rect 10962 -1258 11080 -1240
rect 11190 -1210 11308 -1192
rect 11362 -1158 11480 -1140
rect 11362 -1192 11370 -1158
rect 11404 -1192 11438 -1158
rect 11472 -1192 11480 -1158
rect 11362 -1210 11480 -1192
rect 11590 -1158 11708 -1140
rect 11590 -1192 11598 -1158
rect 11632 -1192 11666 -1158
rect 11700 -1192 11708 -1158
rect 11590 -1210 11708 -1192
rect 11762 -1158 11880 -1140
rect 11990 -1110 12108 -1092
rect 12162 -1058 12280 -1040
rect 12162 -1092 12170 -1058
rect 12204 -1092 12238 -1058
rect 12272 -1092 12280 -1058
rect 12162 -1110 12280 -1092
rect 12390 -1058 12508 -1040
rect 12390 -1092 12398 -1058
rect 12432 -1092 12466 -1058
rect 12500 -1092 12508 -1058
rect 12390 -1110 12508 -1092
rect 12562 -1058 12680 -1040
rect 14540 -1008 14690 -990
rect 14540 -1042 14562 -1008
rect 14596 -1042 14630 -1008
rect 14664 -1042 14690 -1008
rect 12562 -1092 12570 -1058
rect 12604 -1092 12638 -1058
rect 12672 -1092 12680 -1058
rect 14540 -1060 14690 -1042
rect 15652 -1008 15802 -990
rect 15652 -1042 15678 -1008
rect 15712 -1042 15746 -1008
rect 15780 -1042 15802 -1008
rect 15652 -1060 15802 -1042
rect 12562 -1110 12680 -1092
rect 11762 -1192 11770 -1158
rect 11804 -1192 11838 -1158
rect 11872 -1192 11880 -1158
rect 11762 -1210 11880 -1192
rect 11990 -1158 12108 -1140
rect 11990 -1192 11998 -1158
rect 12032 -1192 12066 -1158
rect 12100 -1192 12108 -1158
rect 10962 -1292 10970 -1258
rect 11004 -1292 11038 -1258
rect 11072 -1292 11080 -1258
rect 10962 -1310 11080 -1292
rect 11190 -1258 11308 -1240
rect 11190 -1292 11198 -1258
rect 11232 -1292 11266 -1258
rect 11300 -1292 11308 -1258
rect 10162 -1392 10170 -1358
rect 10204 -1392 10238 -1358
rect 10272 -1392 10280 -1358
rect 10162 -1410 10280 -1392
rect 10390 -1358 10508 -1340
rect 10390 -1392 10398 -1358
rect 10432 -1392 10466 -1358
rect 10500 -1392 10508 -1358
rect 9362 -1492 9370 -1458
rect 9404 -1492 9438 -1458
rect 9472 -1492 9480 -1458
rect 9362 -1510 9480 -1492
rect 9590 -1458 9708 -1440
rect 9590 -1492 9598 -1458
rect 9632 -1492 9666 -1458
rect 9700 -1492 9708 -1458
rect 8562 -1592 8570 -1558
rect 8604 -1592 8638 -1558
rect 8672 -1592 8680 -1558
rect 8562 -1610 8680 -1592
rect 8790 -1558 8908 -1540
rect 8790 -1592 8798 -1558
rect 8832 -1592 8866 -1558
rect 8900 -1592 8908 -1558
rect 7762 -1692 7770 -1658
rect 7804 -1692 7838 -1658
rect 7872 -1692 7880 -1658
rect 7762 -1710 7880 -1692
rect 7990 -1658 8108 -1640
rect 7990 -1692 7998 -1658
rect 8032 -1692 8066 -1658
rect 8100 -1692 8108 -1658
rect 6962 -1792 6970 -1758
rect 7004 -1792 7038 -1758
rect 7072 -1792 7080 -1758
rect 6962 -1810 7080 -1792
rect 7190 -1758 7308 -1740
rect 7190 -1792 7198 -1758
rect 7232 -1792 7266 -1758
rect 7300 -1792 7308 -1758
rect 6162 -1892 6170 -1858
rect 6204 -1892 6238 -1858
rect 6272 -1892 6280 -1858
rect 6162 -1910 6280 -1892
rect 6390 -1858 6508 -1840
rect 6390 -1892 6398 -1858
rect 6432 -1892 6466 -1858
rect 6500 -1892 6508 -1858
rect 5362 -1992 5370 -1958
rect 5404 -1992 5438 -1958
rect 5472 -1992 5480 -1958
rect 5362 -2010 5480 -1992
rect 5590 -1958 5708 -1940
rect 5590 -1992 5598 -1958
rect 5632 -1992 5666 -1958
rect 5700 -1992 5708 -1958
rect 4562 -2092 4570 -2058
rect 4604 -2092 4638 -2058
rect 4672 -2092 4680 -2058
rect 4562 -2129 4680 -2092
rect 4790 -2058 4908 -2040
rect 4790 -2092 4798 -2058
rect 4832 -2092 4866 -2058
rect 4900 -2092 4908 -2058
rect 4790 -2129 4908 -2092
rect 4962 -2058 5080 -2040
rect 4962 -2092 4970 -2058
rect 5004 -2092 5038 -2058
rect 5072 -2092 5080 -2058
rect 4962 -2129 5080 -2092
rect 5190 -2058 5308 -2040
rect 5190 -2092 5198 -2058
rect 5232 -2092 5266 -2058
rect 5300 -2092 5308 -2058
rect 5190 -2129 5308 -2092
rect 5362 -2058 5480 -2040
rect 5590 -2010 5708 -1992
rect 5762 -1958 5880 -1940
rect 5762 -1992 5770 -1958
rect 5804 -1992 5838 -1958
rect 5872 -1992 5880 -1958
rect 5762 -2010 5880 -1992
rect 5990 -1958 6108 -1940
rect 5990 -1992 5998 -1958
rect 6032 -1992 6066 -1958
rect 6100 -1992 6108 -1958
rect 5990 -2010 6108 -1992
rect 6162 -1958 6280 -1940
rect 6390 -1910 6508 -1892
rect 6562 -1858 6680 -1840
rect 6562 -1892 6570 -1858
rect 6604 -1892 6638 -1858
rect 6672 -1892 6680 -1858
rect 6562 -1910 6680 -1892
rect 6790 -1858 6908 -1840
rect 6790 -1892 6798 -1858
rect 6832 -1892 6866 -1858
rect 6900 -1892 6908 -1858
rect 6790 -1910 6908 -1892
rect 6962 -1858 7080 -1840
rect 7190 -1810 7308 -1792
rect 7362 -1758 7480 -1740
rect 7362 -1792 7370 -1758
rect 7404 -1792 7438 -1758
rect 7472 -1792 7480 -1758
rect 7362 -1810 7480 -1792
rect 7590 -1758 7708 -1740
rect 7590 -1792 7598 -1758
rect 7632 -1792 7666 -1758
rect 7700 -1792 7708 -1758
rect 7590 -1810 7708 -1792
rect 7762 -1758 7880 -1740
rect 7990 -1710 8108 -1692
rect 8162 -1658 8280 -1640
rect 8162 -1692 8170 -1658
rect 8204 -1692 8238 -1658
rect 8272 -1692 8280 -1658
rect 8162 -1710 8280 -1692
rect 8390 -1658 8508 -1640
rect 8390 -1692 8398 -1658
rect 8432 -1692 8466 -1658
rect 8500 -1692 8508 -1658
rect 8390 -1710 8508 -1692
rect 8562 -1658 8680 -1640
rect 8790 -1610 8908 -1592
rect 8962 -1558 9080 -1540
rect 8962 -1592 8970 -1558
rect 9004 -1592 9038 -1558
rect 9072 -1592 9080 -1558
rect 8962 -1610 9080 -1592
rect 9190 -1558 9308 -1540
rect 9190 -1592 9198 -1558
rect 9232 -1592 9266 -1558
rect 9300 -1592 9308 -1558
rect 9190 -1610 9308 -1592
rect 9362 -1558 9480 -1540
rect 9590 -1510 9708 -1492
rect 9762 -1458 9880 -1440
rect 9762 -1492 9770 -1458
rect 9804 -1492 9838 -1458
rect 9872 -1492 9880 -1458
rect 9762 -1510 9880 -1492
rect 9990 -1458 10108 -1440
rect 9990 -1492 9998 -1458
rect 10032 -1492 10066 -1458
rect 10100 -1492 10108 -1458
rect 9990 -1510 10108 -1492
rect 10162 -1458 10280 -1440
rect 10390 -1410 10508 -1392
rect 10562 -1358 10680 -1340
rect 10562 -1392 10570 -1358
rect 10604 -1392 10638 -1358
rect 10672 -1392 10680 -1358
rect 10562 -1410 10680 -1392
rect 10790 -1358 10908 -1340
rect 10790 -1392 10798 -1358
rect 10832 -1392 10866 -1358
rect 10900 -1392 10908 -1358
rect 10790 -1410 10908 -1392
rect 10962 -1358 11080 -1340
rect 11190 -1310 11308 -1292
rect 11362 -1258 11480 -1240
rect 11362 -1292 11370 -1258
rect 11404 -1292 11438 -1258
rect 11472 -1292 11480 -1258
rect 11362 -1310 11480 -1292
rect 11590 -1258 11708 -1240
rect 11590 -1292 11598 -1258
rect 11632 -1292 11666 -1258
rect 11700 -1292 11708 -1258
rect 11590 -1310 11708 -1292
rect 11762 -1258 11880 -1240
rect 11990 -1210 12108 -1192
rect 12162 -1158 12280 -1140
rect 12162 -1192 12170 -1158
rect 12204 -1192 12238 -1158
rect 12272 -1192 12280 -1158
rect 12162 -1210 12280 -1192
rect 12390 -1158 12508 -1140
rect 12390 -1192 12398 -1158
rect 12432 -1192 12466 -1158
rect 12500 -1192 12508 -1158
rect 12390 -1210 12508 -1192
rect 12562 -1158 12680 -1140
rect 14540 -1108 14690 -1090
rect 14540 -1142 14562 -1108
rect 14596 -1142 14630 -1108
rect 14664 -1142 14690 -1108
rect 12562 -1192 12570 -1158
rect 12604 -1192 12638 -1158
rect 12672 -1192 12680 -1158
rect 14540 -1160 14690 -1142
rect 15652 -1108 15802 -1090
rect 15652 -1142 15678 -1108
rect 15712 -1142 15746 -1108
rect 15780 -1142 15802 -1108
rect 15652 -1160 15802 -1142
rect 12562 -1210 12680 -1192
rect 11762 -1292 11770 -1258
rect 11804 -1292 11838 -1258
rect 11872 -1292 11880 -1258
rect 11762 -1310 11880 -1292
rect 11990 -1258 12108 -1240
rect 11990 -1292 11998 -1258
rect 12032 -1292 12066 -1258
rect 12100 -1292 12108 -1258
rect 10962 -1392 10970 -1358
rect 11004 -1392 11038 -1358
rect 11072 -1392 11080 -1358
rect 10962 -1410 11080 -1392
rect 11190 -1358 11308 -1340
rect 11190 -1392 11198 -1358
rect 11232 -1392 11266 -1358
rect 11300 -1392 11308 -1358
rect 10162 -1492 10170 -1458
rect 10204 -1492 10238 -1458
rect 10272 -1492 10280 -1458
rect 10162 -1510 10280 -1492
rect 10390 -1458 10508 -1440
rect 10390 -1492 10398 -1458
rect 10432 -1492 10466 -1458
rect 10500 -1492 10508 -1458
rect 9362 -1592 9370 -1558
rect 9404 -1592 9438 -1558
rect 9472 -1592 9480 -1558
rect 9362 -1610 9480 -1592
rect 9590 -1558 9708 -1540
rect 9590 -1592 9598 -1558
rect 9632 -1592 9666 -1558
rect 9700 -1592 9708 -1558
rect 8562 -1692 8570 -1658
rect 8604 -1692 8638 -1658
rect 8672 -1692 8680 -1658
rect 8562 -1710 8680 -1692
rect 8790 -1658 8908 -1640
rect 8790 -1692 8798 -1658
rect 8832 -1692 8866 -1658
rect 8900 -1692 8908 -1658
rect 7762 -1792 7770 -1758
rect 7804 -1792 7838 -1758
rect 7872 -1792 7880 -1758
rect 7762 -1810 7880 -1792
rect 7990 -1758 8108 -1740
rect 7990 -1792 7998 -1758
rect 8032 -1792 8066 -1758
rect 8100 -1792 8108 -1758
rect 6962 -1892 6970 -1858
rect 7004 -1892 7038 -1858
rect 7072 -1892 7080 -1858
rect 6962 -1910 7080 -1892
rect 7190 -1858 7308 -1840
rect 7190 -1892 7198 -1858
rect 7232 -1892 7266 -1858
rect 7300 -1892 7308 -1858
rect 6162 -1992 6170 -1958
rect 6204 -1992 6238 -1958
rect 6272 -1992 6280 -1958
rect 6162 -2010 6280 -1992
rect 6390 -1958 6508 -1940
rect 6390 -1992 6398 -1958
rect 6432 -1992 6466 -1958
rect 6500 -1992 6508 -1958
rect 5362 -2092 5370 -2058
rect 5404 -2092 5438 -2058
rect 5472 -2092 5480 -2058
rect 5362 -2129 5480 -2092
rect 5590 -2058 5708 -2040
rect 5590 -2092 5598 -2058
rect 5632 -2092 5666 -2058
rect 5700 -2092 5708 -2058
rect 5590 -2129 5708 -2092
rect 5762 -2058 5880 -2040
rect 5762 -2092 5770 -2058
rect 5804 -2092 5838 -2058
rect 5872 -2092 5880 -2058
rect 5762 -2129 5880 -2092
rect 5990 -2058 6108 -2040
rect 5990 -2092 5998 -2058
rect 6032 -2092 6066 -2058
rect 6100 -2092 6108 -2058
rect 5990 -2129 6108 -2092
rect 6162 -2058 6280 -2040
rect 6390 -2010 6508 -1992
rect 6562 -1958 6680 -1940
rect 6562 -1992 6570 -1958
rect 6604 -1992 6638 -1958
rect 6672 -1992 6680 -1958
rect 6562 -2010 6680 -1992
rect 6790 -1958 6908 -1940
rect 6790 -1992 6798 -1958
rect 6832 -1992 6866 -1958
rect 6900 -1992 6908 -1958
rect 6790 -2010 6908 -1992
rect 6962 -1958 7080 -1940
rect 7190 -1910 7308 -1892
rect 7362 -1858 7480 -1840
rect 7362 -1892 7370 -1858
rect 7404 -1892 7438 -1858
rect 7472 -1892 7480 -1858
rect 7362 -1910 7480 -1892
rect 7590 -1858 7708 -1840
rect 7590 -1892 7598 -1858
rect 7632 -1892 7666 -1858
rect 7700 -1892 7708 -1858
rect 7590 -1910 7708 -1892
rect 7762 -1858 7880 -1840
rect 7990 -1810 8108 -1792
rect 8162 -1758 8280 -1740
rect 8162 -1792 8170 -1758
rect 8204 -1792 8238 -1758
rect 8272 -1792 8280 -1758
rect 8162 -1810 8280 -1792
rect 8390 -1758 8508 -1740
rect 8390 -1792 8398 -1758
rect 8432 -1792 8466 -1758
rect 8500 -1792 8508 -1758
rect 8390 -1810 8508 -1792
rect 8562 -1758 8680 -1740
rect 8790 -1710 8908 -1692
rect 8962 -1658 9080 -1640
rect 8962 -1692 8970 -1658
rect 9004 -1692 9038 -1658
rect 9072 -1692 9080 -1658
rect 8962 -1710 9080 -1692
rect 9190 -1658 9308 -1640
rect 9190 -1692 9198 -1658
rect 9232 -1692 9266 -1658
rect 9300 -1692 9308 -1658
rect 9190 -1710 9308 -1692
rect 9362 -1658 9480 -1640
rect 9590 -1610 9708 -1592
rect 9762 -1558 9880 -1540
rect 9762 -1592 9770 -1558
rect 9804 -1592 9838 -1558
rect 9872 -1592 9880 -1558
rect 9762 -1610 9880 -1592
rect 9990 -1558 10108 -1540
rect 9990 -1592 9998 -1558
rect 10032 -1592 10066 -1558
rect 10100 -1592 10108 -1558
rect 9990 -1610 10108 -1592
rect 10162 -1558 10280 -1540
rect 10390 -1510 10508 -1492
rect 10562 -1458 10680 -1440
rect 10562 -1492 10570 -1458
rect 10604 -1492 10638 -1458
rect 10672 -1492 10680 -1458
rect 10562 -1510 10680 -1492
rect 10790 -1458 10908 -1440
rect 10790 -1492 10798 -1458
rect 10832 -1492 10866 -1458
rect 10900 -1492 10908 -1458
rect 10790 -1510 10908 -1492
rect 10962 -1458 11080 -1440
rect 11190 -1410 11308 -1392
rect 11362 -1358 11480 -1340
rect 11362 -1392 11370 -1358
rect 11404 -1392 11438 -1358
rect 11472 -1392 11480 -1358
rect 11362 -1410 11480 -1392
rect 11590 -1358 11708 -1340
rect 11590 -1392 11598 -1358
rect 11632 -1392 11666 -1358
rect 11700 -1392 11708 -1358
rect 11590 -1410 11708 -1392
rect 11762 -1358 11880 -1340
rect 11990 -1310 12108 -1292
rect 12162 -1258 12280 -1240
rect 12162 -1292 12170 -1258
rect 12204 -1292 12238 -1258
rect 12272 -1292 12280 -1258
rect 12162 -1310 12280 -1292
rect 12390 -1258 12508 -1240
rect 12390 -1292 12398 -1258
rect 12432 -1292 12466 -1258
rect 12500 -1292 12508 -1258
rect 12390 -1310 12508 -1292
rect 12562 -1258 12680 -1240
rect 14540 -1208 14690 -1190
rect 14540 -1242 14562 -1208
rect 14596 -1242 14630 -1208
rect 14664 -1242 14690 -1208
rect 12562 -1292 12570 -1258
rect 12604 -1292 12638 -1258
rect 12672 -1292 12680 -1258
rect 14540 -1260 14690 -1242
rect 15652 -1208 15802 -1190
rect 15652 -1242 15678 -1208
rect 15712 -1242 15746 -1208
rect 15780 -1242 15802 -1208
rect 15652 -1260 15802 -1242
rect 12562 -1310 12680 -1292
rect 11762 -1392 11770 -1358
rect 11804 -1392 11838 -1358
rect 11872 -1392 11880 -1358
rect 11762 -1410 11880 -1392
rect 11990 -1358 12108 -1340
rect 11990 -1392 11998 -1358
rect 12032 -1392 12066 -1358
rect 12100 -1392 12108 -1358
rect 10962 -1492 10970 -1458
rect 11004 -1492 11038 -1458
rect 11072 -1492 11080 -1458
rect 10962 -1510 11080 -1492
rect 11190 -1458 11308 -1440
rect 11190 -1492 11198 -1458
rect 11232 -1492 11266 -1458
rect 11300 -1492 11308 -1458
rect 10162 -1592 10170 -1558
rect 10204 -1592 10238 -1558
rect 10272 -1592 10280 -1558
rect 10162 -1610 10280 -1592
rect 10390 -1558 10508 -1540
rect 10390 -1592 10398 -1558
rect 10432 -1592 10466 -1558
rect 10500 -1592 10508 -1558
rect 9362 -1692 9370 -1658
rect 9404 -1692 9438 -1658
rect 9472 -1692 9480 -1658
rect 9362 -1710 9480 -1692
rect 9590 -1658 9708 -1640
rect 9590 -1692 9598 -1658
rect 9632 -1692 9666 -1658
rect 9700 -1692 9708 -1658
rect 8562 -1792 8570 -1758
rect 8604 -1792 8638 -1758
rect 8672 -1792 8680 -1758
rect 8562 -1810 8680 -1792
rect 8790 -1758 8908 -1740
rect 8790 -1792 8798 -1758
rect 8832 -1792 8866 -1758
rect 8900 -1792 8908 -1758
rect 7762 -1892 7770 -1858
rect 7804 -1892 7838 -1858
rect 7872 -1892 7880 -1858
rect 7762 -1910 7880 -1892
rect 7990 -1858 8108 -1840
rect 7990 -1892 7998 -1858
rect 8032 -1892 8066 -1858
rect 8100 -1892 8108 -1858
rect 6962 -1992 6970 -1958
rect 7004 -1992 7038 -1958
rect 7072 -1992 7080 -1958
rect 6962 -2010 7080 -1992
rect 7190 -1958 7308 -1940
rect 7190 -1992 7198 -1958
rect 7232 -1992 7266 -1958
rect 7300 -1992 7308 -1958
rect 6162 -2092 6170 -2058
rect 6204 -2092 6238 -2058
rect 6272 -2092 6280 -2058
rect 6162 -2129 6280 -2092
rect 6390 -2058 6508 -2040
rect 6390 -2092 6398 -2058
rect 6432 -2092 6466 -2058
rect 6500 -2092 6508 -2058
rect 6390 -2129 6508 -2092
rect 6562 -2058 6680 -2040
rect 6562 -2092 6570 -2058
rect 6604 -2092 6638 -2058
rect 6672 -2092 6680 -2058
rect 6562 -2129 6680 -2092
rect 6790 -2058 6908 -2040
rect 6790 -2092 6798 -2058
rect 6832 -2092 6866 -2058
rect 6900 -2092 6908 -2058
rect 6790 -2129 6908 -2092
rect 6962 -2058 7080 -2040
rect 7190 -2010 7308 -1992
rect 7362 -1958 7480 -1940
rect 7362 -1992 7370 -1958
rect 7404 -1992 7438 -1958
rect 7472 -1992 7480 -1958
rect 7362 -2010 7480 -1992
rect 7590 -1958 7708 -1940
rect 7590 -1992 7598 -1958
rect 7632 -1992 7666 -1958
rect 7700 -1992 7708 -1958
rect 7590 -2010 7708 -1992
rect 7762 -1958 7880 -1940
rect 7990 -1910 8108 -1892
rect 8162 -1858 8280 -1840
rect 8162 -1892 8170 -1858
rect 8204 -1892 8238 -1858
rect 8272 -1892 8280 -1858
rect 8162 -1910 8280 -1892
rect 8390 -1858 8508 -1840
rect 8390 -1892 8398 -1858
rect 8432 -1892 8466 -1858
rect 8500 -1892 8508 -1858
rect 8390 -1910 8508 -1892
rect 8562 -1858 8680 -1840
rect 8790 -1810 8908 -1792
rect 8962 -1758 9080 -1740
rect 8962 -1792 8970 -1758
rect 9004 -1792 9038 -1758
rect 9072 -1792 9080 -1758
rect 8962 -1810 9080 -1792
rect 9190 -1758 9308 -1740
rect 9190 -1792 9198 -1758
rect 9232 -1792 9266 -1758
rect 9300 -1792 9308 -1758
rect 9190 -1810 9308 -1792
rect 9362 -1758 9480 -1740
rect 9590 -1710 9708 -1692
rect 9762 -1658 9880 -1640
rect 9762 -1692 9770 -1658
rect 9804 -1692 9838 -1658
rect 9872 -1692 9880 -1658
rect 9762 -1710 9880 -1692
rect 9990 -1658 10108 -1640
rect 9990 -1692 9998 -1658
rect 10032 -1692 10066 -1658
rect 10100 -1692 10108 -1658
rect 9990 -1710 10108 -1692
rect 10162 -1658 10280 -1640
rect 10390 -1610 10508 -1592
rect 10562 -1558 10680 -1540
rect 10562 -1592 10570 -1558
rect 10604 -1592 10638 -1558
rect 10672 -1592 10680 -1558
rect 10562 -1610 10680 -1592
rect 10790 -1558 10908 -1540
rect 10790 -1592 10798 -1558
rect 10832 -1592 10866 -1558
rect 10900 -1592 10908 -1558
rect 10790 -1610 10908 -1592
rect 10962 -1558 11080 -1540
rect 11190 -1510 11308 -1492
rect 11362 -1458 11480 -1440
rect 11362 -1492 11370 -1458
rect 11404 -1492 11438 -1458
rect 11472 -1492 11480 -1458
rect 11362 -1510 11480 -1492
rect 11590 -1458 11708 -1440
rect 11590 -1492 11598 -1458
rect 11632 -1492 11666 -1458
rect 11700 -1492 11708 -1458
rect 11590 -1510 11708 -1492
rect 11762 -1458 11880 -1440
rect 11990 -1410 12108 -1392
rect 12162 -1358 12280 -1340
rect 12162 -1392 12170 -1358
rect 12204 -1392 12238 -1358
rect 12272 -1392 12280 -1358
rect 12162 -1410 12280 -1392
rect 12390 -1358 12508 -1340
rect 12390 -1392 12398 -1358
rect 12432 -1392 12466 -1358
rect 12500 -1392 12508 -1358
rect 12390 -1410 12508 -1392
rect 12562 -1358 12680 -1340
rect 14540 -1308 14690 -1290
rect 14540 -1342 14562 -1308
rect 14596 -1342 14630 -1308
rect 14664 -1342 14690 -1308
rect 12562 -1392 12570 -1358
rect 12604 -1392 12638 -1358
rect 12672 -1392 12680 -1358
rect 14540 -1360 14690 -1342
rect 15652 -1308 15802 -1290
rect 15652 -1342 15678 -1308
rect 15712 -1342 15746 -1308
rect 15780 -1342 15802 -1308
rect 15652 -1360 15802 -1342
rect 12562 -1410 12680 -1392
rect 11762 -1492 11770 -1458
rect 11804 -1492 11838 -1458
rect 11872 -1492 11880 -1458
rect 11762 -1510 11880 -1492
rect 11990 -1458 12108 -1440
rect 11990 -1492 11998 -1458
rect 12032 -1492 12066 -1458
rect 12100 -1492 12108 -1458
rect 10962 -1592 10970 -1558
rect 11004 -1592 11038 -1558
rect 11072 -1592 11080 -1558
rect 10962 -1610 11080 -1592
rect 11190 -1558 11308 -1540
rect 11190 -1592 11198 -1558
rect 11232 -1592 11266 -1558
rect 11300 -1592 11308 -1558
rect 10162 -1692 10170 -1658
rect 10204 -1692 10238 -1658
rect 10272 -1692 10280 -1658
rect 10162 -1710 10280 -1692
rect 10390 -1658 10508 -1640
rect 10390 -1692 10398 -1658
rect 10432 -1692 10466 -1658
rect 10500 -1692 10508 -1658
rect 9362 -1792 9370 -1758
rect 9404 -1792 9438 -1758
rect 9472 -1792 9480 -1758
rect 9362 -1810 9480 -1792
rect 9590 -1758 9708 -1740
rect 9590 -1792 9598 -1758
rect 9632 -1792 9666 -1758
rect 9700 -1792 9708 -1758
rect 8562 -1892 8570 -1858
rect 8604 -1892 8638 -1858
rect 8672 -1892 8680 -1858
rect 8562 -1910 8680 -1892
rect 8790 -1858 8908 -1840
rect 8790 -1892 8798 -1858
rect 8832 -1892 8866 -1858
rect 8900 -1892 8908 -1858
rect 7762 -1992 7770 -1958
rect 7804 -1992 7838 -1958
rect 7872 -1992 7880 -1958
rect 7762 -2010 7880 -1992
rect 7990 -1958 8108 -1940
rect 7990 -1992 7998 -1958
rect 8032 -1992 8066 -1958
rect 8100 -1992 8108 -1958
rect 6962 -2092 6970 -2058
rect 7004 -2092 7038 -2058
rect 7072 -2092 7080 -2058
rect 6962 -2129 7080 -2092
rect 7190 -2058 7308 -2040
rect 7190 -2092 7198 -2058
rect 7232 -2092 7266 -2058
rect 7300 -2092 7308 -2058
rect 7190 -2129 7308 -2092
rect 7362 -2058 7480 -2040
rect 7362 -2092 7370 -2058
rect 7404 -2092 7438 -2058
rect 7472 -2092 7480 -2058
rect 7362 -2129 7480 -2092
rect 7590 -2058 7708 -2040
rect 7590 -2092 7598 -2058
rect 7632 -2092 7666 -2058
rect 7700 -2092 7708 -2058
rect 7590 -2129 7708 -2092
rect 7762 -2058 7880 -2040
rect 7990 -2010 8108 -1992
rect 8162 -1958 8280 -1940
rect 8162 -1992 8170 -1958
rect 8204 -1992 8238 -1958
rect 8272 -1992 8280 -1958
rect 8162 -2010 8280 -1992
rect 8390 -1958 8508 -1940
rect 8390 -1992 8398 -1958
rect 8432 -1992 8466 -1958
rect 8500 -1992 8508 -1958
rect 8390 -2010 8508 -1992
rect 8562 -1958 8680 -1940
rect 8790 -1910 8908 -1892
rect 8962 -1858 9080 -1840
rect 8962 -1892 8970 -1858
rect 9004 -1892 9038 -1858
rect 9072 -1892 9080 -1858
rect 8962 -1910 9080 -1892
rect 9190 -1858 9308 -1840
rect 9190 -1892 9198 -1858
rect 9232 -1892 9266 -1858
rect 9300 -1892 9308 -1858
rect 9190 -1910 9308 -1892
rect 9362 -1858 9480 -1840
rect 9590 -1810 9708 -1792
rect 9762 -1758 9880 -1740
rect 9762 -1792 9770 -1758
rect 9804 -1792 9838 -1758
rect 9872 -1792 9880 -1758
rect 9762 -1810 9880 -1792
rect 9990 -1758 10108 -1740
rect 9990 -1792 9998 -1758
rect 10032 -1792 10066 -1758
rect 10100 -1792 10108 -1758
rect 9990 -1810 10108 -1792
rect 10162 -1758 10280 -1740
rect 10390 -1710 10508 -1692
rect 10562 -1658 10680 -1640
rect 10562 -1692 10570 -1658
rect 10604 -1692 10638 -1658
rect 10672 -1692 10680 -1658
rect 10562 -1710 10680 -1692
rect 10790 -1658 10908 -1640
rect 10790 -1692 10798 -1658
rect 10832 -1692 10866 -1658
rect 10900 -1692 10908 -1658
rect 10790 -1710 10908 -1692
rect 10962 -1658 11080 -1640
rect 11190 -1610 11308 -1592
rect 11362 -1558 11480 -1540
rect 11362 -1592 11370 -1558
rect 11404 -1592 11438 -1558
rect 11472 -1592 11480 -1558
rect 11362 -1610 11480 -1592
rect 11590 -1558 11708 -1540
rect 11590 -1592 11598 -1558
rect 11632 -1592 11666 -1558
rect 11700 -1592 11708 -1558
rect 11590 -1610 11708 -1592
rect 11762 -1558 11880 -1540
rect 11990 -1510 12108 -1492
rect 12162 -1458 12280 -1440
rect 12162 -1492 12170 -1458
rect 12204 -1492 12238 -1458
rect 12272 -1492 12280 -1458
rect 12162 -1510 12280 -1492
rect 12390 -1458 12508 -1440
rect 12390 -1492 12398 -1458
rect 12432 -1492 12466 -1458
rect 12500 -1492 12508 -1458
rect 12390 -1510 12508 -1492
rect 12562 -1458 12680 -1440
rect 14540 -1408 14690 -1390
rect 14540 -1442 14562 -1408
rect 14596 -1442 14630 -1408
rect 14664 -1442 14690 -1408
rect 12562 -1492 12570 -1458
rect 12604 -1492 12638 -1458
rect 12672 -1492 12680 -1458
rect 14540 -1460 14690 -1442
rect 15652 -1408 15802 -1390
rect 15652 -1442 15678 -1408
rect 15712 -1442 15746 -1408
rect 15780 -1442 15802 -1408
rect 15652 -1460 15802 -1442
rect 12562 -1510 12680 -1492
rect 11762 -1592 11770 -1558
rect 11804 -1592 11838 -1558
rect 11872 -1592 11880 -1558
rect 11762 -1610 11880 -1592
rect 11990 -1558 12108 -1540
rect 11990 -1592 11998 -1558
rect 12032 -1592 12066 -1558
rect 12100 -1592 12108 -1558
rect 10962 -1692 10970 -1658
rect 11004 -1692 11038 -1658
rect 11072 -1692 11080 -1658
rect 10962 -1710 11080 -1692
rect 11190 -1658 11308 -1640
rect 11190 -1692 11198 -1658
rect 11232 -1692 11266 -1658
rect 11300 -1692 11308 -1658
rect 10162 -1792 10170 -1758
rect 10204 -1792 10238 -1758
rect 10272 -1792 10280 -1758
rect 10162 -1810 10280 -1792
rect 10390 -1758 10508 -1740
rect 10390 -1792 10398 -1758
rect 10432 -1792 10466 -1758
rect 10500 -1792 10508 -1758
rect 9362 -1892 9370 -1858
rect 9404 -1892 9438 -1858
rect 9472 -1892 9480 -1858
rect 9362 -1910 9480 -1892
rect 9590 -1858 9708 -1840
rect 9590 -1892 9598 -1858
rect 9632 -1892 9666 -1858
rect 9700 -1892 9708 -1858
rect 8562 -1992 8570 -1958
rect 8604 -1992 8638 -1958
rect 8672 -1992 8680 -1958
rect 8562 -2010 8680 -1992
rect 8790 -1958 8908 -1940
rect 8790 -1992 8798 -1958
rect 8832 -1992 8866 -1958
rect 8900 -1992 8908 -1958
rect 7762 -2092 7770 -2058
rect 7804 -2092 7838 -2058
rect 7872 -2092 7880 -2058
rect 7762 -2129 7880 -2092
rect 7990 -2058 8108 -2040
rect 7990 -2092 7998 -2058
rect 8032 -2092 8066 -2058
rect 8100 -2092 8108 -2058
rect 7990 -2129 8108 -2092
rect 8162 -2058 8280 -2040
rect 8162 -2092 8170 -2058
rect 8204 -2092 8238 -2058
rect 8272 -2092 8280 -2058
rect 8162 -2129 8280 -2092
rect 8390 -2058 8508 -2040
rect 8390 -2092 8398 -2058
rect 8432 -2092 8466 -2058
rect 8500 -2092 8508 -2058
rect 8390 -2129 8508 -2092
rect 8562 -2058 8680 -2040
rect 8790 -2010 8908 -1992
rect 8962 -1958 9080 -1940
rect 8962 -1992 8970 -1958
rect 9004 -1992 9038 -1958
rect 9072 -1992 9080 -1958
rect 8962 -2010 9080 -1992
rect 9190 -1958 9308 -1940
rect 9190 -1992 9198 -1958
rect 9232 -1992 9266 -1958
rect 9300 -1992 9308 -1958
rect 9190 -2010 9308 -1992
rect 9362 -1958 9480 -1940
rect 9590 -1910 9708 -1892
rect 9762 -1858 9880 -1840
rect 9762 -1892 9770 -1858
rect 9804 -1892 9838 -1858
rect 9872 -1892 9880 -1858
rect 9762 -1910 9880 -1892
rect 9990 -1858 10108 -1840
rect 9990 -1892 9998 -1858
rect 10032 -1892 10066 -1858
rect 10100 -1892 10108 -1858
rect 9990 -1910 10108 -1892
rect 10162 -1858 10280 -1840
rect 10390 -1810 10508 -1792
rect 10562 -1758 10680 -1740
rect 10562 -1792 10570 -1758
rect 10604 -1792 10638 -1758
rect 10672 -1792 10680 -1758
rect 10562 -1810 10680 -1792
rect 10790 -1758 10908 -1740
rect 10790 -1792 10798 -1758
rect 10832 -1792 10866 -1758
rect 10900 -1792 10908 -1758
rect 10790 -1810 10908 -1792
rect 10962 -1758 11080 -1740
rect 11190 -1710 11308 -1692
rect 11362 -1658 11480 -1640
rect 11362 -1692 11370 -1658
rect 11404 -1692 11438 -1658
rect 11472 -1692 11480 -1658
rect 11362 -1710 11480 -1692
rect 11590 -1658 11708 -1640
rect 11590 -1692 11598 -1658
rect 11632 -1692 11666 -1658
rect 11700 -1692 11708 -1658
rect 11590 -1710 11708 -1692
rect 11762 -1658 11880 -1640
rect 11990 -1610 12108 -1592
rect 12162 -1558 12280 -1540
rect 12162 -1592 12170 -1558
rect 12204 -1592 12238 -1558
rect 12272 -1592 12280 -1558
rect 12162 -1610 12280 -1592
rect 12390 -1558 12508 -1540
rect 12390 -1592 12398 -1558
rect 12432 -1592 12466 -1558
rect 12500 -1592 12508 -1558
rect 12390 -1610 12508 -1592
rect 12562 -1558 12680 -1540
rect 14540 -1508 14690 -1490
rect 14540 -1542 14562 -1508
rect 14596 -1542 14630 -1508
rect 14664 -1542 14690 -1508
rect 12562 -1592 12570 -1558
rect 12604 -1592 12638 -1558
rect 12672 -1592 12680 -1558
rect 14540 -1560 14690 -1542
rect 15652 -1508 15802 -1490
rect 15652 -1542 15678 -1508
rect 15712 -1542 15746 -1508
rect 15780 -1542 15802 -1508
rect 15652 -1560 15802 -1542
rect 12562 -1610 12680 -1592
rect 11762 -1692 11770 -1658
rect 11804 -1692 11838 -1658
rect 11872 -1692 11880 -1658
rect 11762 -1710 11880 -1692
rect 11990 -1658 12108 -1640
rect 11990 -1692 11998 -1658
rect 12032 -1692 12066 -1658
rect 12100 -1692 12108 -1658
rect 10962 -1792 10970 -1758
rect 11004 -1792 11038 -1758
rect 11072 -1792 11080 -1758
rect 10962 -1810 11080 -1792
rect 11190 -1758 11308 -1740
rect 11190 -1792 11198 -1758
rect 11232 -1792 11266 -1758
rect 11300 -1792 11308 -1758
rect 10162 -1892 10170 -1858
rect 10204 -1892 10238 -1858
rect 10272 -1892 10280 -1858
rect 10162 -1910 10280 -1892
rect 10390 -1858 10508 -1840
rect 10390 -1892 10398 -1858
rect 10432 -1892 10466 -1858
rect 10500 -1892 10508 -1858
rect 9362 -1992 9370 -1958
rect 9404 -1992 9438 -1958
rect 9472 -1992 9480 -1958
rect 9362 -2010 9480 -1992
rect 9590 -1958 9708 -1940
rect 9590 -1992 9598 -1958
rect 9632 -1992 9666 -1958
rect 9700 -1992 9708 -1958
rect 8562 -2092 8570 -2058
rect 8604 -2092 8638 -2058
rect 8672 -2092 8680 -2058
rect 8562 -2129 8680 -2092
rect 8790 -2058 8908 -2040
rect 8790 -2092 8798 -2058
rect 8832 -2092 8866 -2058
rect 8900 -2092 8908 -2058
rect 8790 -2129 8908 -2092
rect 8962 -2058 9080 -2040
rect 8962 -2092 8970 -2058
rect 9004 -2092 9038 -2058
rect 9072 -2092 9080 -2058
rect 8962 -2129 9080 -2092
rect 9190 -2058 9308 -2040
rect 9190 -2092 9198 -2058
rect 9232 -2092 9266 -2058
rect 9300 -2092 9308 -2058
rect 9190 -2129 9308 -2092
rect 9362 -2058 9480 -2040
rect 9590 -2010 9708 -1992
rect 9762 -1958 9880 -1940
rect 9762 -1992 9770 -1958
rect 9804 -1992 9838 -1958
rect 9872 -1992 9880 -1958
rect 9762 -2010 9880 -1992
rect 9990 -1958 10108 -1940
rect 9990 -1992 9998 -1958
rect 10032 -1992 10066 -1958
rect 10100 -1992 10108 -1958
rect 9990 -2010 10108 -1992
rect 10162 -1958 10280 -1940
rect 10390 -1910 10508 -1892
rect 10562 -1858 10680 -1840
rect 10562 -1892 10570 -1858
rect 10604 -1892 10638 -1858
rect 10672 -1892 10680 -1858
rect 10562 -1910 10680 -1892
rect 10790 -1858 10908 -1840
rect 10790 -1892 10798 -1858
rect 10832 -1892 10866 -1858
rect 10900 -1892 10908 -1858
rect 10790 -1910 10908 -1892
rect 10962 -1858 11080 -1840
rect 11190 -1810 11308 -1792
rect 11362 -1758 11480 -1740
rect 11362 -1792 11370 -1758
rect 11404 -1792 11438 -1758
rect 11472 -1792 11480 -1758
rect 11362 -1810 11480 -1792
rect 11590 -1758 11708 -1740
rect 11590 -1792 11598 -1758
rect 11632 -1792 11666 -1758
rect 11700 -1792 11708 -1758
rect 11590 -1810 11708 -1792
rect 11762 -1758 11880 -1740
rect 11990 -1710 12108 -1692
rect 12162 -1658 12280 -1640
rect 12162 -1692 12170 -1658
rect 12204 -1692 12238 -1658
rect 12272 -1692 12280 -1658
rect 12162 -1710 12280 -1692
rect 12390 -1658 12508 -1640
rect 12390 -1692 12398 -1658
rect 12432 -1692 12466 -1658
rect 12500 -1692 12508 -1658
rect 12390 -1710 12508 -1692
rect 12562 -1658 12680 -1640
rect 14540 -1608 14690 -1590
rect 14540 -1642 14562 -1608
rect 14596 -1642 14630 -1608
rect 14664 -1642 14690 -1608
rect 12562 -1692 12570 -1658
rect 12604 -1692 12638 -1658
rect 12672 -1692 12680 -1658
rect 14540 -1660 14690 -1642
rect 15652 -1608 15802 -1590
rect 15652 -1642 15678 -1608
rect 15712 -1642 15746 -1608
rect 15780 -1642 15802 -1608
rect 15652 -1660 15802 -1642
rect 12562 -1710 12680 -1692
rect 11762 -1792 11770 -1758
rect 11804 -1792 11838 -1758
rect 11872 -1792 11880 -1758
rect 11762 -1810 11880 -1792
rect 11990 -1758 12108 -1740
rect 11990 -1792 11998 -1758
rect 12032 -1792 12066 -1758
rect 12100 -1792 12108 -1758
rect 10962 -1892 10970 -1858
rect 11004 -1892 11038 -1858
rect 11072 -1892 11080 -1858
rect 10962 -1910 11080 -1892
rect 11190 -1858 11308 -1840
rect 11190 -1892 11198 -1858
rect 11232 -1892 11266 -1858
rect 11300 -1892 11308 -1858
rect 10162 -1992 10170 -1958
rect 10204 -1992 10238 -1958
rect 10272 -1992 10280 -1958
rect 10162 -2010 10280 -1992
rect 10390 -1958 10508 -1940
rect 10390 -1992 10398 -1958
rect 10432 -1992 10466 -1958
rect 10500 -1992 10508 -1958
rect 9362 -2092 9370 -2058
rect 9404 -2092 9438 -2058
rect 9472 -2092 9480 -2058
rect 9362 -2129 9480 -2092
rect 9590 -2058 9708 -2040
rect 9590 -2092 9598 -2058
rect 9632 -2092 9666 -2058
rect 9700 -2092 9708 -2058
rect 9590 -2129 9708 -2092
rect 9762 -2058 9880 -2040
rect 9762 -2092 9770 -2058
rect 9804 -2092 9838 -2058
rect 9872 -2092 9880 -2058
rect 9762 -2129 9880 -2092
rect 9990 -2058 10108 -2040
rect 9990 -2092 9998 -2058
rect 10032 -2092 10066 -2058
rect 10100 -2092 10108 -2058
rect 9990 -2129 10108 -2092
rect 10162 -2058 10280 -2040
rect 10390 -2010 10508 -1992
rect 10562 -1958 10680 -1940
rect 10562 -1992 10570 -1958
rect 10604 -1992 10638 -1958
rect 10672 -1992 10680 -1958
rect 10562 -2010 10680 -1992
rect 10790 -1958 10908 -1940
rect 10790 -1992 10798 -1958
rect 10832 -1992 10866 -1958
rect 10900 -1992 10908 -1958
rect 10790 -2010 10908 -1992
rect 10962 -1958 11080 -1940
rect 11190 -1910 11308 -1892
rect 11362 -1858 11480 -1840
rect 11362 -1892 11370 -1858
rect 11404 -1892 11438 -1858
rect 11472 -1892 11480 -1858
rect 11362 -1910 11480 -1892
rect 11590 -1858 11708 -1840
rect 11590 -1892 11598 -1858
rect 11632 -1892 11666 -1858
rect 11700 -1892 11708 -1858
rect 11590 -1910 11708 -1892
rect 11762 -1858 11880 -1840
rect 11990 -1810 12108 -1792
rect 12162 -1758 12280 -1740
rect 12162 -1792 12170 -1758
rect 12204 -1792 12238 -1758
rect 12272 -1792 12280 -1758
rect 12162 -1810 12280 -1792
rect 12390 -1758 12508 -1740
rect 12390 -1792 12398 -1758
rect 12432 -1792 12466 -1758
rect 12500 -1792 12508 -1758
rect 12390 -1810 12508 -1792
rect 12562 -1758 12680 -1740
rect 14540 -1708 14690 -1690
rect 14540 -1742 14562 -1708
rect 14596 -1742 14630 -1708
rect 14664 -1742 14690 -1708
rect 12562 -1792 12570 -1758
rect 12604 -1792 12638 -1758
rect 12672 -1792 12680 -1758
rect 14540 -1760 14690 -1742
rect 15652 -1708 15802 -1690
rect 15652 -1742 15678 -1708
rect 15712 -1742 15746 -1708
rect 15780 -1742 15802 -1708
rect 15652 -1760 15802 -1742
rect 12562 -1810 12680 -1792
rect 11762 -1892 11770 -1858
rect 11804 -1892 11838 -1858
rect 11872 -1892 11880 -1858
rect 11762 -1910 11880 -1892
rect 11990 -1858 12108 -1840
rect 11990 -1892 11998 -1858
rect 12032 -1892 12066 -1858
rect 12100 -1892 12108 -1858
rect 10962 -1992 10970 -1958
rect 11004 -1992 11038 -1958
rect 11072 -1992 11080 -1958
rect 10962 -2010 11080 -1992
rect 11190 -1958 11308 -1940
rect 11190 -1992 11198 -1958
rect 11232 -1992 11266 -1958
rect 11300 -1992 11308 -1958
rect 10162 -2092 10170 -2058
rect 10204 -2092 10238 -2058
rect 10272 -2092 10280 -2058
rect 10162 -2129 10280 -2092
rect 10390 -2058 10508 -2040
rect 10390 -2092 10398 -2058
rect 10432 -2092 10466 -2058
rect 10500 -2092 10508 -2058
rect 10390 -2129 10508 -2092
rect 10562 -2058 10680 -2040
rect 10562 -2092 10570 -2058
rect 10604 -2092 10638 -2058
rect 10672 -2092 10680 -2058
rect 10562 -2129 10680 -2092
rect 10790 -2058 10908 -2040
rect 10790 -2092 10798 -2058
rect 10832 -2092 10866 -2058
rect 10900 -2092 10908 -2058
rect 10790 -2129 10908 -2092
rect 10962 -2058 11080 -2040
rect 11190 -2010 11308 -1992
rect 11362 -1958 11480 -1940
rect 11362 -1992 11370 -1958
rect 11404 -1992 11438 -1958
rect 11472 -1992 11480 -1958
rect 11362 -2010 11480 -1992
rect 11590 -1958 11708 -1940
rect 11590 -1992 11598 -1958
rect 11632 -1992 11666 -1958
rect 11700 -1992 11708 -1958
rect 11590 -2010 11708 -1992
rect 11762 -1958 11880 -1940
rect 11990 -1910 12108 -1892
rect 12162 -1858 12280 -1840
rect 12162 -1892 12170 -1858
rect 12204 -1892 12238 -1858
rect 12272 -1892 12280 -1858
rect 12162 -1910 12280 -1892
rect 12390 -1858 12508 -1840
rect 12390 -1892 12398 -1858
rect 12432 -1892 12466 -1858
rect 12500 -1892 12508 -1858
rect 12390 -1910 12508 -1892
rect 12562 -1858 12680 -1840
rect 14540 -1808 14690 -1790
rect 14540 -1842 14562 -1808
rect 14596 -1842 14630 -1808
rect 14664 -1842 14690 -1808
rect 12562 -1892 12570 -1858
rect 12604 -1892 12638 -1858
rect 12672 -1892 12680 -1858
rect 14540 -1860 14690 -1842
rect 15652 -1808 15802 -1790
rect 15652 -1842 15678 -1808
rect 15712 -1842 15746 -1808
rect 15780 -1842 15802 -1808
rect 15652 -1860 15802 -1842
rect 12562 -1910 12680 -1892
rect 11762 -1992 11770 -1958
rect 11804 -1992 11838 -1958
rect 11872 -1992 11880 -1958
rect 11762 -2010 11880 -1992
rect 11990 -1958 12108 -1940
rect 11990 -1992 11998 -1958
rect 12032 -1992 12066 -1958
rect 12100 -1992 12108 -1958
rect 10962 -2092 10970 -2058
rect 11004 -2092 11038 -2058
rect 11072 -2092 11080 -2058
rect 10962 -2129 11080 -2092
rect 11190 -2058 11308 -2040
rect 11190 -2092 11198 -2058
rect 11232 -2092 11266 -2058
rect 11300 -2092 11308 -2058
rect 11190 -2129 11308 -2092
rect 11362 -2058 11480 -2040
rect 11362 -2092 11370 -2058
rect 11404 -2092 11438 -2058
rect 11472 -2092 11480 -2058
rect 11362 -2129 11480 -2092
rect 11590 -2058 11708 -2040
rect 11590 -2092 11598 -2058
rect 11632 -2092 11666 -2058
rect 11700 -2092 11708 -2058
rect 11590 -2129 11708 -2092
rect 11762 -2058 11880 -2040
rect 11990 -2010 12108 -1992
rect 12162 -1958 12280 -1940
rect 12162 -1992 12170 -1958
rect 12204 -1992 12238 -1958
rect 12272 -1992 12280 -1958
rect 12162 -2010 12280 -1992
rect 12390 -1958 12508 -1940
rect 12390 -1992 12398 -1958
rect 12432 -1992 12466 -1958
rect 12500 -1992 12508 -1958
rect 12390 -2010 12508 -1992
rect 12562 -1958 12680 -1940
rect 14540 -1908 14690 -1890
rect 14540 -1942 14562 -1908
rect 14596 -1942 14630 -1908
rect 14664 -1942 14690 -1908
rect 12562 -1992 12570 -1958
rect 12604 -1992 12638 -1958
rect 12672 -1992 12680 -1958
rect 14540 -1960 14690 -1942
rect 15652 -1908 15802 -1890
rect 15652 -1942 15678 -1908
rect 15712 -1942 15746 -1908
rect 15780 -1942 15802 -1908
rect 15652 -1960 15802 -1942
rect 12562 -2010 12680 -1992
rect 11762 -2092 11770 -2058
rect 11804 -2092 11838 -2058
rect 11872 -2092 11880 -2058
rect 11762 -2129 11880 -2092
rect 11990 -2058 12108 -2040
rect 11990 -2092 11998 -2058
rect 12032 -2092 12066 -2058
rect 12100 -2092 12108 -2058
rect 11990 -2129 12108 -2092
rect 12162 -2058 12280 -2040
rect 12162 -2092 12170 -2058
rect 12204 -2092 12238 -2058
rect 12272 -2092 12280 -2058
rect 12162 -2129 12280 -2092
rect 12390 -2058 12508 -2040
rect 12390 -2092 12398 -2058
rect 12432 -2092 12466 -2058
rect 12500 -2092 12508 -2058
rect 12390 -2129 12508 -2092
rect 12562 -2058 12680 -2040
rect 14540 -2008 14690 -1990
rect 14540 -2042 14562 -2008
rect 14596 -2042 14630 -2008
rect 14664 -2042 14690 -2008
rect 12562 -2092 12570 -2058
rect 12604 -2092 12638 -2058
rect 12672 -2092 12680 -2058
rect 12562 -2129 12680 -2092
rect 14540 -2079 14690 -2042
rect 15652 -2008 15802 -1990
rect 15652 -2042 15678 -2008
rect 15712 -2042 15746 -2008
rect 15780 -2042 15802 -2008
rect 15652 -2079 15802 -2042
<< pdiff >>
rect 14816 -208 15116 -171
rect 14816 -242 14847 -208
rect 14881 -242 14915 -208
rect 14949 -242 14983 -208
rect 15017 -242 15051 -208
rect 15085 -242 15116 -208
rect 14816 -260 15116 -242
rect 15226 -208 15526 -171
rect 15226 -242 15257 -208
rect 15291 -242 15325 -208
rect 15359 -242 15393 -208
rect 15427 -242 15461 -208
rect 15495 -242 15526 -208
rect 15226 -260 15526 -242
rect -94 -363 -30 -330
rect -94 -397 -82 -363
rect -48 -397 -30 -363
rect -94 -431 -30 -397
rect -94 -465 -82 -431
rect -48 -465 -30 -431
rect -94 -498 -30 -465
rect 0 -363 70 -330
rect 0 -397 18 -363
rect 52 -397 70 -363
rect 0 -431 70 -397
rect 0 -465 18 -431
rect 52 -465 70 -431
rect 0 -498 70 -465
rect 100 -363 170 -330
rect 100 -397 118 -363
rect 152 -397 170 -363
rect 100 -431 170 -397
rect 100 -465 118 -431
rect 152 -465 170 -431
rect 100 -498 170 -465
rect 200 -363 270 -330
rect 200 -397 218 -363
rect 252 -397 270 -363
rect 200 -431 270 -397
rect 200 -465 218 -431
rect 252 -465 270 -431
rect 200 -498 270 -465
rect 300 -363 370 -330
rect 300 -397 318 -363
rect 352 -397 370 -363
rect 300 -431 370 -397
rect 300 -465 318 -431
rect 352 -465 370 -431
rect 300 -498 370 -465
rect 400 -363 470 -330
rect 400 -397 418 -363
rect 452 -397 470 -363
rect 400 -431 470 -397
rect 400 -465 418 -431
rect 452 -465 470 -431
rect 400 -498 470 -465
rect 500 -363 570 -330
rect 500 -397 518 -363
rect 552 -397 570 -363
rect 500 -431 570 -397
rect 500 -465 518 -431
rect 552 -465 570 -431
rect 500 -498 570 -465
rect 600 -363 670 -330
rect 600 -397 618 -363
rect 652 -397 670 -363
rect 600 -431 670 -397
rect 600 -465 618 -431
rect 652 -465 670 -431
rect 600 -498 670 -465
rect 700 -363 770 -330
rect 700 -397 718 -363
rect 752 -397 770 -363
rect 700 -431 770 -397
rect 700 -465 718 -431
rect 752 -465 770 -431
rect 700 -498 770 -465
rect 800 -363 870 -330
rect 800 -397 818 -363
rect 852 -397 870 -363
rect 800 -431 870 -397
rect 800 -465 818 -431
rect 852 -465 870 -431
rect 800 -498 870 -465
rect 900 -363 970 -330
rect 900 -397 918 -363
rect 952 -397 970 -363
rect 900 -431 970 -397
rect 900 -465 918 -431
rect 952 -465 970 -431
rect 900 -498 970 -465
rect 1000 -363 1070 -330
rect 1000 -397 1018 -363
rect 1052 -397 1070 -363
rect 1000 -431 1070 -397
rect 1000 -465 1018 -431
rect 1052 -465 1070 -431
rect 1000 -498 1070 -465
rect 1100 -363 1170 -330
rect 1100 -397 1118 -363
rect 1152 -397 1170 -363
rect 1100 -431 1170 -397
rect 1100 -465 1118 -431
rect 1152 -465 1170 -431
rect 1100 -498 1170 -465
rect 1200 -363 1270 -330
rect 1200 -397 1218 -363
rect 1252 -397 1270 -363
rect 1200 -431 1270 -397
rect 1200 -465 1218 -431
rect 1252 -465 1270 -431
rect 1200 -498 1270 -465
rect 1300 -363 1370 -330
rect 1300 -397 1318 -363
rect 1352 -397 1370 -363
rect 1300 -431 1370 -397
rect 1300 -465 1318 -431
rect 1352 -465 1370 -431
rect 1300 -498 1370 -465
rect 1400 -363 1470 -330
rect 1400 -397 1418 -363
rect 1452 -397 1470 -363
rect 1400 -431 1470 -397
rect 1400 -465 1418 -431
rect 1452 -465 1470 -431
rect 1400 -498 1470 -465
rect 1500 -363 1570 -330
rect 1500 -397 1518 -363
rect 1552 -397 1570 -363
rect 1500 -431 1570 -397
rect 1500 -465 1518 -431
rect 1552 -465 1570 -431
rect 1500 -498 1570 -465
rect 1600 -363 1670 -330
rect 1600 -397 1618 -363
rect 1652 -397 1670 -363
rect 1600 -431 1670 -397
rect 1600 -465 1618 -431
rect 1652 -465 1670 -431
rect 1600 -498 1670 -465
rect 1700 -363 1770 -330
rect 1700 -397 1718 -363
rect 1752 -397 1770 -363
rect 1700 -431 1770 -397
rect 1700 -465 1718 -431
rect 1752 -465 1770 -431
rect 1700 -498 1770 -465
rect 1800 -363 1870 -330
rect 1800 -397 1818 -363
rect 1852 -397 1870 -363
rect 1800 -431 1870 -397
rect 1800 -465 1818 -431
rect 1852 -465 1870 -431
rect 1800 -498 1870 -465
rect 1900 -363 1970 -330
rect 1900 -397 1918 -363
rect 1952 -397 1970 -363
rect 1900 -431 1970 -397
rect 1900 -465 1918 -431
rect 1952 -465 1970 -431
rect 1900 -498 1970 -465
rect 2000 -363 2070 -330
rect 2000 -397 2018 -363
rect 2052 -397 2070 -363
rect 2000 -431 2070 -397
rect 2000 -465 2018 -431
rect 2052 -465 2070 -431
rect 2000 -498 2070 -465
rect 2100 -363 2170 -330
rect 2100 -397 2118 -363
rect 2152 -397 2170 -363
rect 2100 -431 2170 -397
rect 2100 -465 2118 -431
rect 2152 -465 2170 -431
rect 2100 -498 2170 -465
rect 2200 -363 2270 -330
rect 2200 -397 2218 -363
rect 2252 -397 2270 -363
rect 2200 -431 2270 -397
rect 2200 -465 2218 -431
rect 2252 -465 2270 -431
rect 2200 -498 2270 -465
rect 2300 -363 2370 -330
rect 2300 -397 2318 -363
rect 2352 -397 2370 -363
rect 2300 -431 2370 -397
rect 2300 -465 2318 -431
rect 2352 -465 2370 -431
rect 2300 -498 2370 -465
rect 2400 -363 2470 -330
rect 2400 -397 2418 -363
rect 2452 -397 2470 -363
rect 2400 -431 2470 -397
rect 2400 -465 2418 -431
rect 2452 -465 2470 -431
rect 2400 -498 2470 -465
rect 2500 -363 2570 -330
rect 2500 -397 2518 -363
rect 2552 -397 2570 -363
rect 2500 -431 2570 -397
rect 2500 -465 2518 -431
rect 2552 -465 2570 -431
rect 2500 -498 2570 -465
rect 2600 -363 2670 -330
rect 2600 -397 2618 -363
rect 2652 -397 2670 -363
rect 2600 -431 2670 -397
rect 2600 -465 2618 -431
rect 2652 -465 2670 -431
rect 2600 -498 2670 -465
rect 2700 -363 2770 -330
rect 2700 -397 2718 -363
rect 2752 -397 2770 -363
rect 2700 -431 2770 -397
rect 2700 -465 2718 -431
rect 2752 -465 2770 -431
rect 2700 -498 2770 -465
rect 2800 -363 2870 -330
rect 2800 -397 2818 -363
rect 2852 -397 2870 -363
rect 2800 -431 2870 -397
rect 2800 -465 2818 -431
rect 2852 -465 2870 -431
rect 2800 -498 2870 -465
rect 2900 -363 2970 -330
rect 2900 -397 2918 -363
rect 2952 -397 2970 -363
rect 2900 -431 2970 -397
rect 2900 -465 2918 -431
rect 2952 -465 2970 -431
rect 2900 -498 2970 -465
rect 3000 -363 3070 -330
rect 3000 -397 3018 -363
rect 3052 -397 3070 -363
rect 3000 -431 3070 -397
rect 3000 -465 3018 -431
rect 3052 -465 3070 -431
rect 3000 -498 3070 -465
rect 3100 -363 3170 -330
rect 3100 -397 3118 -363
rect 3152 -397 3170 -363
rect 3100 -431 3170 -397
rect 3100 -465 3118 -431
rect 3152 -465 3170 -431
rect 3100 -498 3170 -465
rect 3200 -363 3270 -330
rect 3200 -397 3218 -363
rect 3252 -397 3270 -363
rect 3200 -431 3270 -397
rect 3200 -465 3218 -431
rect 3252 -465 3270 -431
rect 3200 -498 3270 -465
rect 3300 -363 3370 -330
rect 3300 -397 3318 -363
rect 3352 -397 3370 -363
rect 3300 -431 3370 -397
rect 3300 -465 3318 -431
rect 3352 -465 3370 -431
rect 3300 -498 3370 -465
rect 3400 -363 3470 -330
rect 3400 -397 3418 -363
rect 3452 -397 3470 -363
rect 3400 -431 3470 -397
rect 3400 -465 3418 -431
rect 3452 -465 3470 -431
rect 3400 -498 3470 -465
rect 3500 -363 3570 -330
rect 3500 -397 3518 -363
rect 3552 -397 3570 -363
rect 3500 -431 3570 -397
rect 3500 -465 3518 -431
rect 3552 -465 3570 -431
rect 3500 -498 3570 -465
rect 3600 -363 3670 -330
rect 3600 -397 3618 -363
rect 3652 -397 3670 -363
rect 3600 -431 3670 -397
rect 3600 -465 3618 -431
rect 3652 -465 3670 -431
rect 3600 -498 3670 -465
rect 3700 -363 3770 -330
rect 3700 -397 3718 -363
rect 3752 -397 3770 -363
rect 3700 -431 3770 -397
rect 3700 -465 3718 -431
rect 3752 -465 3770 -431
rect 3700 -498 3770 -465
rect 3800 -363 3870 -330
rect 3800 -397 3818 -363
rect 3852 -397 3870 -363
rect 3800 -431 3870 -397
rect 3800 -465 3818 -431
rect 3852 -465 3870 -431
rect 3800 -498 3870 -465
rect 3900 -363 3970 -330
rect 3900 -397 3918 -363
rect 3952 -397 3970 -363
rect 3900 -431 3970 -397
rect 3900 -465 3918 -431
rect 3952 -465 3970 -431
rect 3900 -498 3970 -465
rect 4000 -363 4070 -330
rect 4000 -397 4018 -363
rect 4052 -397 4070 -363
rect 4000 -431 4070 -397
rect 4000 -465 4018 -431
rect 4052 -465 4070 -431
rect 4000 -498 4070 -465
rect 4100 -363 4170 -330
rect 4100 -397 4118 -363
rect 4152 -397 4170 -363
rect 4100 -431 4170 -397
rect 4100 -465 4118 -431
rect 4152 -465 4170 -431
rect 4100 -498 4170 -465
rect 4200 -363 4270 -330
rect 4200 -397 4218 -363
rect 4252 -397 4270 -363
rect 4200 -431 4270 -397
rect 4200 -465 4218 -431
rect 4252 -465 4270 -431
rect 4200 -498 4270 -465
rect 4300 -363 4370 -330
rect 4300 -397 4318 -363
rect 4352 -397 4370 -363
rect 4300 -431 4370 -397
rect 4300 -465 4318 -431
rect 4352 -465 4370 -431
rect 4300 -498 4370 -465
rect 4400 -363 4470 -330
rect 4400 -397 4418 -363
rect 4452 -397 4470 -363
rect 4400 -431 4470 -397
rect 4400 -465 4418 -431
rect 4452 -465 4470 -431
rect 4400 -498 4470 -465
rect 4500 -363 4570 -330
rect 4500 -397 4518 -363
rect 4552 -397 4570 -363
rect 4500 -431 4570 -397
rect 4500 -465 4518 -431
rect 4552 -465 4570 -431
rect 4500 -498 4570 -465
rect 4600 -363 4670 -330
rect 4600 -397 4618 -363
rect 4652 -397 4670 -363
rect 4600 -431 4670 -397
rect 4600 -465 4618 -431
rect 4652 -465 4670 -431
rect 4600 -498 4670 -465
rect 4700 -363 4770 -330
rect 4700 -397 4718 -363
rect 4752 -397 4770 -363
rect 4700 -431 4770 -397
rect 4700 -465 4718 -431
rect 4752 -465 4770 -431
rect 4700 -498 4770 -465
rect 4800 -363 4870 -330
rect 4800 -397 4818 -363
rect 4852 -397 4870 -363
rect 4800 -431 4870 -397
rect 4800 -465 4818 -431
rect 4852 -465 4870 -431
rect 4800 -498 4870 -465
rect 4900 -363 4970 -330
rect 4900 -397 4918 -363
rect 4952 -397 4970 -363
rect 4900 -431 4970 -397
rect 4900 -465 4918 -431
rect 4952 -465 4970 -431
rect 4900 -498 4970 -465
rect 5000 -363 5070 -330
rect 5000 -397 5018 -363
rect 5052 -397 5070 -363
rect 5000 -431 5070 -397
rect 5000 -465 5018 -431
rect 5052 -465 5070 -431
rect 5000 -498 5070 -465
rect 5100 -363 5170 -330
rect 5100 -397 5118 -363
rect 5152 -397 5170 -363
rect 5100 -431 5170 -397
rect 5100 -465 5118 -431
rect 5152 -465 5170 -431
rect 5100 -498 5170 -465
rect 5200 -363 5270 -330
rect 5200 -397 5218 -363
rect 5252 -397 5270 -363
rect 5200 -431 5270 -397
rect 5200 -465 5218 -431
rect 5252 -465 5270 -431
rect 5200 -498 5270 -465
rect 5300 -363 5370 -330
rect 5300 -397 5318 -363
rect 5352 -397 5370 -363
rect 5300 -431 5370 -397
rect 5300 -465 5318 -431
rect 5352 -465 5370 -431
rect 5300 -498 5370 -465
rect 5400 -363 5470 -330
rect 5400 -397 5418 -363
rect 5452 -397 5470 -363
rect 5400 -431 5470 -397
rect 5400 -465 5418 -431
rect 5452 -465 5470 -431
rect 5400 -498 5470 -465
rect 5500 -363 5570 -330
rect 5500 -397 5518 -363
rect 5552 -397 5570 -363
rect 5500 -431 5570 -397
rect 5500 -465 5518 -431
rect 5552 -465 5570 -431
rect 5500 -498 5570 -465
rect 5600 -363 5670 -330
rect 5600 -397 5618 -363
rect 5652 -397 5670 -363
rect 5600 -431 5670 -397
rect 5600 -465 5618 -431
rect 5652 -465 5670 -431
rect 5600 -498 5670 -465
rect 5700 -363 5770 -330
rect 5700 -397 5718 -363
rect 5752 -397 5770 -363
rect 5700 -431 5770 -397
rect 5700 -465 5718 -431
rect 5752 -465 5770 -431
rect 5700 -498 5770 -465
rect 5800 -363 5870 -330
rect 5800 -397 5818 -363
rect 5852 -397 5870 -363
rect 5800 -431 5870 -397
rect 5800 -465 5818 -431
rect 5852 -465 5870 -431
rect 5800 -498 5870 -465
rect 5900 -363 5970 -330
rect 5900 -397 5918 -363
rect 5952 -397 5970 -363
rect 5900 -431 5970 -397
rect 5900 -465 5918 -431
rect 5952 -465 5970 -431
rect 5900 -498 5970 -465
rect 6000 -363 6070 -330
rect 6000 -397 6018 -363
rect 6052 -397 6070 -363
rect 6000 -431 6070 -397
rect 6000 -465 6018 -431
rect 6052 -465 6070 -431
rect 6000 -498 6070 -465
rect 6100 -363 6170 -330
rect 6100 -397 6118 -363
rect 6152 -397 6170 -363
rect 6100 -431 6170 -397
rect 6100 -465 6118 -431
rect 6152 -465 6170 -431
rect 6100 -498 6170 -465
rect 6200 -363 6270 -330
rect 6200 -397 6218 -363
rect 6252 -397 6270 -363
rect 6200 -431 6270 -397
rect 6200 -465 6218 -431
rect 6252 -465 6270 -431
rect 6200 -498 6270 -465
rect 6300 -363 6370 -330
rect 6300 -397 6318 -363
rect 6352 -397 6370 -363
rect 6300 -431 6370 -397
rect 6300 -465 6318 -431
rect 6352 -465 6370 -431
rect 6300 -498 6370 -465
rect 6400 -363 6470 -330
rect 6400 -397 6418 -363
rect 6452 -397 6470 -363
rect 6400 -431 6470 -397
rect 6400 -465 6418 -431
rect 6452 -465 6470 -431
rect 6400 -498 6470 -465
rect 6500 -363 6570 -330
rect 6500 -397 6518 -363
rect 6552 -397 6570 -363
rect 6500 -431 6570 -397
rect 6500 -465 6518 -431
rect 6552 -465 6570 -431
rect 6500 -498 6570 -465
rect 6600 -363 6670 -330
rect 6600 -397 6618 -363
rect 6652 -397 6670 -363
rect 6600 -431 6670 -397
rect 6600 -465 6618 -431
rect 6652 -465 6670 -431
rect 6600 -498 6670 -465
rect 6700 -363 6770 -330
rect 6700 -397 6718 -363
rect 6752 -397 6770 -363
rect 6700 -431 6770 -397
rect 6700 -465 6718 -431
rect 6752 -465 6770 -431
rect 6700 -498 6770 -465
rect 6800 -363 6870 -330
rect 6800 -397 6818 -363
rect 6852 -397 6870 -363
rect 6800 -431 6870 -397
rect 6800 -465 6818 -431
rect 6852 -465 6870 -431
rect 6800 -498 6870 -465
rect 6900 -363 6970 -330
rect 6900 -397 6918 -363
rect 6952 -397 6970 -363
rect 6900 -431 6970 -397
rect 6900 -465 6918 -431
rect 6952 -465 6970 -431
rect 6900 -498 6970 -465
rect 7000 -363 7070 -330
rect 7000 -397 7018 -363
rect 7052 -397 7070 -363
rect 7000 -431 7070 -397
rect 7000 -465 7018 -431
rect 7052 -465 7070 -431
rect 7000 -498 7070 -465
rect 7100 -363 7170 -330
rect 7100 -397 7118 -363
rect 7152 -397 7170 -363
rect 7100 -431 7170 -397
rect 7100 -465 7118 -431
rect 7152 -465 7170 -431
rect 7100 -498 7170 -465
rect 7200 -363 7270 -330
rect 7200 -397 7218 -363
rect 7252 -397 7270 -363
rect 7200 -431 7270 -397
rect 7200 -465 7218 -431
rect 7252 -465 7270 -431
rect 7200 -498 7270 -465
rect 7300 -363 7370 -330
rect 7300 -397 7318 -363
rect 7352 -397 7370 -363
rect 7300 -431 7370 -397
rect 7300 -465 7318 -431
rect 7352 -465 7370 -431
rect 7300 -498 7370 -465
rect 7400 -363 7470 -330
rect 7400 -397 7418 -363
rect 7452 -397 7470 -363
rect 7400 -431 7470 -397
rect 7400 -465 7418 -431
rect 7452 -465 7470 -431
rect 7400 -498 7470 -465
rect 7500 -363 7570 -330
rect 7500 -397 7518 -363
rect 7552 -397 7570 -363
rect 7500 -431 7570 -397
rect 7500 -465 7518 -431
rect 7552 -465 7570 -431
rect 7500 -498 7570 -465
rect 7600 -363 7670 -330
rect 7600 -397 7618 -363
rect 7652 -397 7670 -363
rect 7600 -431 7670 -397
rect 7600 -465 7618 -431
rect 7652 -465 7670 -431
rect 7600 -498 7670 -465
rect 7700 -363 7770 -330
rect 7700 -397 7718 -363
rect 7752 -397 7770 -363
rect 7700 -431 7770 -397
rect 7700 -465 7718 -431
rect 7752 -465 7770 -431
rect 7700 -498 7770 -465
rect 7800 -363 7870 -330
rect 7800 -397 7818 -363
rect 7852 -397 7870 -363
rect 7800 -431 7870 -397
rect 7800 -465 7818 -431
rect 7852 -465 7870 -431
rect 7800 -498 7870 -465
rect 7900 -363 7970 -330
rect 7900 -397 7918 -363
rect 7952 -397 7970 -363
rect 7900 -431 7970 -397
rect 7900 -465 7918 -431
rect 7952 -465 7970 -431
rect 7900 -498 7970 -465
rect 8000 -363 8070 -330
rect 8000 -397 8018 -363
rect 8052 -397 8070 -363
rect 8000 -431 8070 -397
rect 8000 -465 8018 -431
rect 8052 -465 8070 -431
rect 8000 -498 8070 -465
rect 8100 -363 8170 -330
rect 8100 -397 8118 -363
rect 8152 -397 8170 -363
rect 8100 -431 8170 -397
rect 8100 -465 8118 -431
rect 8152 -465 8170 -431
rect 8100 -498 8170 -465
rect 8200 -363 8270 -330
rect 8200 -397 8218 -363
rect 8252 -397 8270 -363
rect 8200 -431 8270 -397
rect 8200 -465 8218 -431
rect 8252 -465 8270 -431
rect 8200 -498 8270 -465
rect 8300 -363 8370 -330
rect 8300 -397 8318 -363
rect 8352 -397 8370 -363
rect 8300 -431 8370 -397
rect 8300 -465 8318 -431
rect 8352 -465 8370 -431
rect 8300 -498 8370 -465
rect 8400 -363 8470 -330
rect 8400 -397 8418 -363
rect 8452 -397 8470 -363
rect 8400 -431 8470 -397
rect 8400 -465 8418 -431
rect 8452 -465 8470 -431
rect 8400 -498 8470 -465
rect 8500 -363 8570 -330
rect 8500 -397 8518 -363
rect 8552 -397 8570 -363
rect 8500 -431 8570 -397
rect 8500 -465 8518 -431
rect 8552 -465 8570 -431
rect 8500 -498 8570 -465
rect 8600 -363 8670 -330
rect 8600 -397 8618 -363
rect 8652 -397 8670 -363
rect 8600 -431 8670 -397
rect 8600 -465 8618 -431
rect 8652 -465 8670 -431
rect 8600 -498 8670 -465
rect 8700 -363 8770 -330
rect 8700 -397 8718 -363
rect 8752 -397 8770 -363
rect 8700 -431 8770 -397
rect 8700 -465 8718 -431
rect 8752 -465 8770 -431
rect 8700 -498 8770 -465
rect 8800 -363 8870 -330
rect 8800 -397 8818 -363
rect 8852 -397 8870 -363
rect 8800 -431 8870 -397
rect 8800 -465 8818 -431
rect 8852 -465 8870 -431
rect 8800 -498 8870 -465
rect 8900 -363 8970 -330
rect 8900 -397 8918 -363
rect 8952 -397 8970 -363
rect 8900 -431 8970 -397
rect 8900 -465 8918 -431
rect 8952 -465 8970 -431
rect 8900 -498 8970 -465
rect 9000 -363 9070 -330
rect 9000 -397 9018 -363
rect 9052 -397 9070 -363
rect 9000 -431 9070 -397
rect 9000 -465 9018 -431
rect 9052 -465 9070 -431
rect 9000 -498 9070 -465
rect 9100 -363 9170 -330
rect 9100 -397 9118 -363
rect 9152 -397 9170 -363
rect 9100 -431 9170 -397
rect 9100 -465 9118 -431
rect 9152 -465 9170 -431
rect 9100 -498 9170 -465
rect 9200 -363 9270 -330
rect 9200 -397 9218 -363
rect 9252 -397 9270 -363
rect 9200 -431 9270 -397
rect 9200 -465 9218 -431
rect 9252 -465 9270 -431
rect 9200 -498 9270 -465
rect 9300 -363 9370 -330
rect 9300 -397 9318 -363
rect 9352 -397 9370 -363
rect 9300 -431 9370 -397
rect 9300 -465 9318 -431
rect 9352 -465 9370 -431
rect 9300 -498 9370 -465
rect 9400 -363 9470 -330
rect 9400 -397 9418 -363
rect 9452 -397 9470 -363
rect 9400 -431 9470 -397
rect 9400 -465 9418 -431
rect 9452 -465 9470 -431
rect 9400 -498 9470 -465
rect 9500 -363 9570 -330
rect 9500 -397 9518 -363
rect 9552 -397 9570 -363
rect 9500 -431 9570 -397
rect 9500 -465 9518 -431
rect 9552 -465 9570 -431
rect 9500 -498 9570 -465
rect 9600 -363 9670 -330
rect 9600 -397 9618 -363
rect 9652 -397 9670 -363
rect 9600 -431 9670 -397
rect 9600 -465 9618 -431
rect 9652 -465 9670 -431
rect 9600 -498 9670 -465
rect 9700 -363 9770 -330
rect 9700 -397 9718 -363
rect 9752 -397 9770 -363
rect 9700 -431 9770 -397
rect 9700 -465 9718 -431
rect 9752 -465 9770 -431
rect 9700 -498 9770 -465
rect 9800 -363 9870 -330
rect 9800 -397 9818 -363
rect 9852 -397 9870 -363
rect 9800 -431 9870 -397
rect 9800 -465 9818 -431
rect 9852 -465 9870 -431
rect 9800 -498 9870 -465
rect 9900 -363 9970 -330
rect 9900 -397 9918 -363
rect 9952 -397 9970 -363
rect 9900 -431 9970 -397
rect 9900 -465 9918 -431
rect 9952 -465 9970 -431
rect 9900 -498 9970 -465
rect 10000 -363 10070 -330
rect 10000 -397 10018 -363
rect 10052 -397 10070 -363
rect 10000 -431 10070 -397
rect 10000 -465 10018 -431
rect 10052 -465 10070 -431
rect 10000 -498 10070 -465
rect 10100 -363 10170 -330
rect 10100 -397 10118 -363
rect 10152 -397 10170 -363
rect 10100 -431 10170 -397
rect 10100 -465 10118 -431
rect 10152 -465 10170 -431
rect 10100 -498 10170 -465
rect 10200 -363 10270 -330
rect 10200 -397 10218 -363
rect 10252 -397 10270 -363
rect 10200 -431 10270 -397
rect 10200 -465 10218 -431
rect 10252 -465 10270 -431
rect 10200 -498 10270 -465
rect 10300 -363 10370 -330
rect 10300 -397 10318 -363
rect 10352 -397 10370 -363
rect 10300 -431 10370 -397
rect 10300 -465 10318 -431
rect 10352 -465 10370 -431
rect 10300 -498 10370 -465
rect 10400 -363 10470 -330
rect 10400 -397 10418 -363
rect 10452 -397 10470 -363
rect 10400 -431 10470 -397
rect 10400 -465 10418 -431
rect 10452 -465 10470 -431
rect 10400 -498 10470 -465
rect 10500 -363 10570 -330
rect 10500 -397 10518 -363
rect 10552 -397 10570 -363
rect 10500 -431 10570 -397
rect 10500 -465 10518 -431
rect 10552 -465 10570 -431
rect 10500 -498 10570 -465
rect 10600 -363 10670 -330
rect 10600 -397 10618 -363
rect 10652 -397 10670 -363
rect 10600 -431 10670 -397
rect 10600 -465 10618 -431
rect 10652 -465 10670 -431
rect 10600 -498 10670 -465
rect 10700 -363 10770 -330
rect 10700 -397 10718 -363
rect 10752 -397 10770 -363
rect 10700 -431 10770 -397
rect 10700 -465 10718 -431
rect 10752 -465 10770 -431
rect 10700 -498 10770 -465
rect 10800 -363 10870 -330
rect 10800 -397 10818 -363
rect 10852 -397 10870 -363
rect 10800 -431 10870 -397
rect 10800 -465 10818 -431
rect 10852 -465 10870 -431
rect 10800 -498 10870 -465
rect 10900 -363 10970 -330
rect 10900 -397 10918 -363
rect 10952 -397 10970 -363
rect 10900 -431 10970 -397
rect 10900 -465 10918 -431
rect 10952 -465 10970 -431
rect 10900 -498 10970 -465
rect 11000 -363 11070 -330
rect 11000 -397 11018 -363
rect 11052 -397 11070 -363
rect 11000 -431 11070 -397
rect 11000 -465 11018 -431
rect 11052 -465 11070 -431
rect 11000 -498 11070 -465
rect 11100 -363 11170 -330
rect 11100 -397 11118 -363
rect 11152 -397 11170 -363
rect 11100 -431 11170 -397
rect 11100 -465 11118 -431
rect 11152 -465 11170 -431
rect 11100 -498 11170 -465
rect 11200 -363 11270 -330
rect 11200 -397 11218 -363
rect 11252 -397 11270 -363
rect 11200 -431 11270 -397
rect 11200 -465 11218 -431
rect 11252 -465 11270 -431
rect 11200 -498 11270 -465
rect 11300 -363 11370 -330
rect 11300 -397 11318 -363
rect 11352 -397 11370 -363
rect 11300 -431 11370 -397
rect 11300 -465 11318 -431
rect 11352 -465 11370 -431
rect 11300 -498 11370 -465
rect 11400 -363 11470 -330
rect 11400 -397 11418 -363
rect 11452 -397 11470 -363
rect 11400 -431 11470 -397
rect 11400 -465 11418 -431
rect 11452 -465 11470 -431
rect 11400 -498 11470 -465
rect 11500 -363 11570 -330
rect 11500 -397 11518 -363
rect 11552 -397 11570 -363
rect 11500 -431 11570 -397
rect 11500 -465 11518 -431
rect 11552 -465 11570 -431
rect 11500 -498 11570 -465
rect 11600 -363 11670 -330
rect 11600 -397 11618 -363
rect 11652 -397 11670 -363
rect 11600 -431 11670 -397
rect 11600 -465 11618 -431
rect 11652 -465 11670 -431
rect 11600 -498 11670 -465
rect 11700 -363 11770 -330
rect 11700 -397 11718 -363
rect 11752 -397 11770 -363
rect 11700 -431 11770 -397
rect 11700 -465 11718 -431
rect 11752 -465 11770 -431
rect 11700 -498 11770 -465
rect 11800 -363 11870 -330
rect 11800 -397 11818 -363
rect 11852 -397 11870 -363
rect 11800 -431 11870 -397
rect 11800 -465 11818 -431
rect 11852 -465 11870 -431
rect 11800 -498 11870 -465
rect 11900 -363 11970 -330
rect 11900 -397 11918 -363
rect 11952 -397 11970 -363
rect 11900 -431 11970 -397
rect 11900 -465 11918 -431
rect 11952 -465 11970 -431
rect 11900 -498 11970 -465
rect 12000 -363 12070 -330
rect 12000 -397 12018 -363
rect 12052 -397 12070 -363
rect 12000 -431 12070 -397
rect 12000 -465 12018 -431
rect 12052 -465 12070 -431
rect 12000 -498 12070 -465
rect 12100 -363 12170 -330
rect 12100 -397 12118 -363
rect 12152 -397 12170 -363
rect 12100 -431 12170 -397
rect 12100 -465 12118 -431
rect 12152 -465 12170 -431
rect 12100 -498 12170 -465
rect 12200 -363 12270 -330
rect 12200 -397 12218 -363
rect 12252 -397 12270 -363
rect 12200 -431 12270 -397
rect 12200 -465 12218 -431
rect 12252 -465 12270 -431
rect 12200 -498 12270 -465
rect 12300 -363 12370 -330
rect 12300 -397 12318 -363
rect 12352 -397 12370 -363
rect 12300 -431 12370 -397
rect 12300 -465 12318 -431
rect 12352 -465 12370 -431
rect 12300 -498 12370 -465
rect 12400 -363 12470 -330
rect 12400 -397 12418 -363
rect 12452 -397 12470 -363
rect 12400 -431 12470 -397
rect 12400 -465 12418 -431
rect 12452 -465 12470 -431
rect 12400 -498 12470 -465
rect 12500 -363 12570 -330
rect 12500 -397 12518 -363
rect 12552 -397 12570 -363
rect 12500 -431 12570 -397
rect 12500 -465 12518 -431
rect 12552 -465 12570 -431
rect 12500 -498 12570 -465
rect 12600 -363 12670 -330
rect 12600 -397 12618 -363
rect 12652 -397 12670 -363
rect 12600 -431 12670 -397
rect 12600 -465 12618 -431
rect 12652 -465 12670 -431
rect 12600 -498 12670 -465
rect 12700 -363 12764 -330
rect 14816 -308 15116 -290
rect 14816 -342 14847 -308
rect 14881 -342 14915 -308
rect 14949 -342 14983 -308
rect 15017 -342 15051 -308
rect 15085 -342 15116 -308
rect 14816 -360 15116 -342
rect 15226 -308 15526 -290
rect 15226 -342 15257 -308
rect 15291 -342 15325 -308
rect 15359 -342 15393 -308
rect 15427 -342 15461 -308
rect 15495 -342 15526 -308
rect 15226 -360 15526 -342
rect 12700 -397 12718 -363
rect 12752 -397 12764 -363
rect 12700 -431 12764 -397
rect 12700 -465 12718 -431
rect 12752 -465 12764 -431
rect 14816 -408 15116 -390
rect 14816 -442 14847 -408
rect 14881 -442 14915 -408
rect 14949 -442 14983 -408
rect 15017 -442 15051 -408
rect 15085 -442 15116 -408
rect 14816 -460 15116 -442
rect 15226 -408 15526 -390
rect 15226 -442 15257 -408
rect 15291 -442 15325 -408
rect 15359 -442 15393 -408
rect 15427 -442 15461 -408
rect 15495 -442 15526 -408
rect 15226 -460 15526 -442
rect 12700 -498 12764 -465
rect 14816 -508 15116 -490
rect 14816 -542 14847 -508
rect 14881 -542 14915 -508
rect 14949 -542 14983 -508
rect 15017 -542 15051 -508
rect 15085 -542 15116 -508
rect 14816 -560 15116 -542
rect 15226 -508 15526 -490
rect 15226 -542 15257 -508
rect 15291 -542 15325 -508
rect 15359 -542 15393 -508
rect 15427 -542 15461 -508
rect 15495 -542 15526 -508
rect 15226 -560 15526 -542
rect -38 -683 15 -658
rect -38 -717 -30 -683
rect 4 -717 15 -683
rect -38 -742 15 -717
rect 107 -683 163 -658
rect 107 -717 118 -683
rect 152 -717 163 -683
rect 107 -742 163 -717
rect 255 -683 308 -658
rect 255 -717 266 -683
rect 300 -717 308 -683
rect 255 -742 308 -717
rect 362 -683 415 -658
rect 362 -717 370 -683
rect 404 -717 415 -683
rect 362 -742 415 -717
rect 507 -683 563 -658
rect 507 -717 518 -683
rect 552 -717 563 -683
rect 507 -742 563 -717
rect 655 -683 708 -658
rect 655 -717 666 -683
rect 700 -717 708 -683
rect 655 -742 708 -717
rect 762 -683 815 -658
rect 762 -717 770 -683
rect 804 -717 815 -683
rect 762 -742 815 -717
rect 907 -683 963 -658
rect 907 -717 918 -683
rect 952 -717 963 -683
rect 907 -742 963 -717
rect 1055 -683 1108 -658
rect 1055 -717 1066 -683
rect 1100 -717 1108 -683
rect 1055 -742 1108 -717
rect 1162 -683 1215 -658
rect 1162 -717 1170 -683
rect 1204 -717 1215 -683
rect 1162 -742 1215 -717
rect 1307 -683 1363 -658
rect 1307 -717 1318 -683
rect 1352 -717 1363 -683
rect 1307 -742 1363 -717
rect 1455 -683 1508 -658
rect 1455 -717 1466 -683
rect 1500 -717 1508 -683
rect 1455 -742 1508 -717
rect 1562 -683 1615 -658
rect 1562 -717 1570 -683
rect 1604 -717 1615 -683
rect 1562 -742 1615 -717
rect 1707 -683 1763 -658
rect 1707 -717 1718 -683
rect 1752 -717 1763 -683
rect 1707 -742 1763 -717
rect 1855 -683 1908 -658
rect 1855 -717 1866 -683
rect 1900 -717 1908 -683
rect 1855 -742 1908 -717
rect 1962 -683 2015 -658
rect 1962 -717 1970 -683
rect 2004 -717 2015 -683
rect 1962 -742 2015 -717
rect 2107 -683 2163 -658
rect 2107 -717 2118 -683
rect 2152 -717 2163 -683
rect 2107 -742 2163 -717
rect 2255 -683 2308 -658
rect 2255 -717 2266 -683
rect 2300 -717 2308 -683
rect 2255 -742 2308 -717
rect 2362 -683 2415 -658
rect 2362 -717 2370 -683
rect 2404 -717 2415 -683
rect 2362 -742 2415 -717
rect 2507 -683 2563 -658
rect 2507 -717 2518 -683
rect 2552 -717 2563 -683
rect 2507 -742 2563 -717
rect 2655 -683 2708 -658
rect 2655 -717 2666 -683
rect 2700 -717 2708 -683
rect 2655 -742 2708 -717
rect 2762 -683 2815 -658
rect 2762 -717 2770 -683
rect 2804 -717 2815 -683
rect 2762 -742 2815 -717
rect 2907 -683 2963 -658
rect 2907 -717 2918 -683
rect 2952 -717 2963 -683
rect 2907 -742 2963 -717
rect 3055 -683 3108 -658
rect 3055 -717 3066 -683
rect 3100 -717 3108 -683
rect 3055 -742 3108 -717
rect 3162 -683 3215 -658
rect 3162 -717 3170 -683
rect 3204 -717 3215 -683
rect 3162 -742 3215 -717
rect 3307 -683 3363 -658
rect 3307 -717 3318 -683
rect 3352 -717 3363 -683
rect 3307 -742 3363 -717
rect 3455 -683 3508 -658
rect 3455 -717 3466 -683
rect 3500 -717 3508 -683
rect 3455 -742 3508 -717
rect 3562 -683 3615 -658
rect 3562 -717 3570 -683
rect 3604 -717 3615 -683
rect 3562 -742 3615 -717
rect 3707 -683 3763 -658
rect 3707 -717 3718 -683
rect 3752 -717 3763 -683
rect 3707 -742 3763 -717
rect 3855 -683 3908 -658
rect 3855 -717 3866 -683
rect 3900 -717 3908 -683
rect 3855 -742 3908 -717
rect 3962 -683 4015 -658
rect 3962 -717 3970 -683
rect 4004 -717 4015 -683
rect 3962 -742 4015 -717
rect 4107 -683 4163 -658
rect 4107 -717 4118 -683
rect 4152 -717 4163 -683
rect 4107 -742 4163 -717
rect 4255 -683 4308 -658
rect 4255 -717 4266 -683
rect 4300 -717 4308 -683
rect 4255 -742 4308 -717
rect 4362 -683 4415 -658
rect 4362 -717 4370 -683
rect 4404 -717 4415 -683
rect 4362 -742 4415 -717
rect 4507 -683 4563 -658
rect 4507 -717 4518 -683
rect 4552 -717 4563 -683
rect 4507 -742 4563 -717
rect 4655 -683 4708 -658
rect 4655 -717 4666 -683
rect 4700 -717 4708 -683
rect 4655 -742 4708 -717
rect 4762 -683 4815 -658
rect 4762 -717 4770 -683
rect 4804 -717 4815 -683
rect 4762 -742 4815 -717
rect 4907 -683 4963 -658
rect 4907 -717 4918 -683
rect 4952 -717 4963 -683
rect 4907 -742 4963 -717
rect 5055 -683 5108 -658
rect 5055 -717 5066 -683
rect 5100 -717 5108 -683
rect 5055 -742 5108 -717
rect 5162 -683 5215 -658
rect 5162 -717 5170 -683
rect 5204 -717 5215 -683
rect 5162 -742 5215 -717
rect 5307 -683 5363 -658
rect 5307 -717 5318 -683
rect 5352 -717 5363 -683
rect 5307 -742 5363 -717
rect 5455 -683 5508 -658
rect 5455 -717 5466 -683
rect 5500 -717 5508 -683
rect 5455 -742 5508 -717
rect 5562 -683 5615 -658
rect 5562 -717 5570 -683
rect 5604 -717 5615 -683
rect 5562 -742 5615 -717
rect 5707 -683 5763 -658
rect 5707 -717 5718 -683
rect 5752 -717 5763 -683
rect 5707 -742 5763 -717
rect 5855 -683 5908 -658
rect 5855 -717 5866 -683
rect 5900 -717 5908 -683
rect 5855 -742 5908 -717
rect 5962 -683 6015 -658
rect 5962 -717 5970 -683
rect 6004 -717 6015 -683
rect 5962 -742 6015 -717
rect 6107 -683 6163 -658
rect 6107 -717 6118 -683
rect 6152 -717 6163 -683
rect 6107 -742 6163 -717
rect 6255 -683 6308 -658
rect 6255 -717 6266 -683
rect 6300 -717 6308 -683
rect 6255 -742 6308 -717
rect 6362 -683 6415 -658
rect 6362 -717 6370 -683
rect 6404 -717 6415 -683
rect 6362 -742 6415 -717
rect 6507 -683 6563 -658
rect 6507 -717 6518 -683
rect 6552 -717 6563 -683
rect 6507 -742 6563 -717
rect 6655 -683 6708 -658
rect 6655 -717 6666 -683
rect 6700 -717 6708 -683
rect 6655 -742 6708 -717
rect 6762 -683 6815 -658
rect 6762 -717 6770 -683
rect 6804 -717 6815 -683
rect 6762 -742 6815 -717
rect 6907 -683 6963 -658
rect 6907 -717 6918 -683
rect 6952 -717 6963 -683
rect 6907 -742 6963 -717
rect 7055 -683 7108 -658
rect 7055 -717 7066 -683
rect 7100 -717 7108 -683
rect 7055 -742 7108 -717
rect 7162 -683 7215 -658
rect 7162 -717 7170 -683
rect 7204 -717 7215 -683
rect 7162 -742 7215 -717
rect 7307 -683 7363 -658
rect 7307 -717 7318 -683
rect 7352 -717 7363 -683
rect 7307 -742 7363 -717
rect 7455 -683 7508 -658
rect 7455 -717 7466 -683
rect 7500 -717 7508 -683
rect 7455 -742 7508 -717
rect 7562 -683 7615 -658
rect 7562 -717 7570 -683
rect 7604 -717 7615 -683
rect 7562 -742 7615 -717
rect 7707 -683 7763 -658
rect 7707 -717 7718 -683
rect 7752 -717 7763 -683
rect 7707 -742 7763 -717
rect 7855 -683 7908 -658
rect 7855 -717 7866 -683
rect 7900 -717 7908 -683
rect 7855 -742 7908 -717
rect 7962 -683 8015 -658
rect 7962 -717 7970 -683
rect 8004 -717 8015 -683
rect 7962 -742 8015 -717
rect 8107 -683 8163 -658
rect 8107 -717 8118 -683
rect 8152 -717 8163 -683
rect 8107 -742 8163 -717
rect 8255 -683 8308 -658
rect 8255 -717 8266 -683
rect 8300 -717 8308 -683
rect 8255 -742 8308 -717
rect 8362 -683 8415 -658
rect 8362 -717 8370 -683
rect 8404 -717 8415 -683
rect 8362 -742 8415 -717
rect 8507 -683 8563 -658
rect 8507 -717 8518 -683
rect 8552 -717 8563 -683
rect 8507 -742 8563 -717
rect 8655 -683 8708 -658
rect 8655 -717 8666 -683
rect 8700 -717 8708 -683
rect 8655 -742 8708 -717
rect 8762 -683 8815 -658
rect 8762 -717 8770 -683
rect 8804 -717 8815 -683
rect 8762 -742 8815 -717
rect 8907 -683 8963 -658
rect 8907 -717 8918 -683
rect 8952 -717 8963 -683
rect 8907 -742 8963 -717
rect 9055 -683 9108 -658
rect 9055 -717 9066 -683
rect 9100 -717 9108 -683
rect 9055 -742 9108 -717
rect 9162 -683 9215 -658
rect 9162 -717 9170 -683
rect 9204 -717 9215 -683
rect 9162 -742 9215 -717
rect 9307 -683 9363 -658
rect 9307 -717 9318 -683
rect 9352 -717 9363 -683
rect 9307 -742 9363 -717
rect 9455 -683 9508 -658
rect 9455 -717 9466 -683
rect 9500 -717 9508 -683
rect 9455 -742 9508 -717
rect 9562 -683 9615 -658
rect 9562 -717 9570 -683
rect 9604 -717 9615 -683
rect 9562 -742 9615 -717
rect 9707 -683 9763 -658
rect 9707 -717 9718 -683
rect 9752 -717 9763 -683
rect 9707 -742 9763 -717
rect 9855 -683 9908 -658
rect 9855 -717 9866 -683
rect 9900 -717 9908 -683
rect 9855 -742 9908 -717
rect 9962 -683 10015 -658
rect 9962 -717 9970 -683
rect 10004 -717 10015 -683
rect 9962 -742 10015 -717
rect 10107 -683 10163 -658
rect 10107 -717 10118 -683
rect 10152 -717 10163 -683
rect 10107 -742 10163 -717
rect 10255 -683 10308 -658
rect 10255 -717 10266 -683
rect 10300 -717 10308 -683
rect 10255 -742 10308 -717
rect 10362 -683 10415 -658
rect 10362 -717 10370 -683
rect 10404 -717 10415 -683
rect 10362 -742 10415 -717
rect 10507 -683 10563 -658
rect 10507 -717 10518 -683
rect 10552 -717 10563 -683
rect 10507 -742 10563 -717
rect 10655 -683 10708 -658
rect 10655 -717 10666 -683
rect 10700 -717 10708 -683
rect 10655 -742 10708 -717
rect 10762 -683 10815 -658
rect 10762 -717 10770 -683
rect 10804 -717 10815 -683
rect 10762 -742 10815 -717
rect 10907 -683 10963 -658
rect 10907 -717 10918 -683
rect 10952 -717 10963 -683
rect 10907 -742 10963 -717
rect 11055 -683 11108 -658
rect 11055 -717 11066 -683
rect 11100 -717 11108 -683
rect 11055 -742 11108 -717
rect 11162 -683 11215 -658
rect 11162 -717 11170 -683
rect 11204 -717 11215 -683
rect 11162 -742 11215 -717
rect 11307 -683 11363 -658
rect 11307 -717 11318 -683
rect 11352 -717 11363 -683
rect 11307 -742 11363 -717
rect 11455 -683 11508 -658
rect 11455 -717 11466 -683
rect 11500 -717 11508 -683
rect 11455 -742 11508 -717
rect 11562 -683 11615 -658
rect 11562 -717 11570 -683
rect 11604 -717 11615 -683
rect 11562 -742 11615 -717
rect 11707 -683 11763 -658
rect 11707 -717 11718 -683
rect 11752 -717 11763 -683
rect 11707 -742 11763 -717
rect 11855 -683 11908 -658
rect 11855 -717 11866 -683
rect 11900 -717 11908 -683
rect 11855 -742 11908 -717
rect 11962 -683 12015 -658
rect 11962 -717 11970 -683
rect 12004 -717 12015 -683
rect 11962 -742 12015 -717
rect 12107 -683 12163 -658
rect 12107 -717 12118 -683
rect 12152 -717 12163 -683
rect 12107 -742 12163 -717
rect 12255 -683 12308 -658
rect 12255 -717 12266 -683
rect 12300 -717 12308 -683
rect 12255 -742 12308 -717
rect 12362 -683 12415 -658
rect 12362 -717 12370 -683
rect 12404 -717 12415 -683
rect 12362 -742 12415 -717
rect 12507 -683 12563 -658
rect 12507 -717 12518 -683
rect 12552 -717 12563 -683
rect 12507 -742 12563 -717
rect 12655 -683 12708 -658
rect 14816 -608 15116 -590
rect 14816 -642 14847 -608
rect 14881 -642 14915 -608
rect 14949 -642 14983 -608
rect 15017 -642 15051 -608
rect 15085 -642 15116 -608
rect 14816 -660 15116 -642
rect 15226 -608 15526 -590
rect 15226 -642 15257 -608
rect 15291 -642 15325 -608
rect 15359 -642 15393 -608
rect 15427 -642 15461 -608
rect 15495 -642 15526 -608
rect 15226 -660 15526 -642
rect 12655 -717 12666 -683
rect 12700 -717 12708 -683
rect 12655 -742 12708 -717
rect 14816 -708 15116 -690
rect 14816 -742 14847 -708
rect 14881 -742 14915 -708
rect 14949 -742 14983 -708
rect 15017 -742 15051 -708
rect 15085 -742 15116 -708
rect 14816 -760 15116 -742
rect 15226 -708 15526 -690
rect 15226 -742 15257 -708
rect 15291 -742 15325 -708
rect 15359 -742 15393 -708
rect 15427 -742 15461 -708
rect 15495 -742 15526 -708
rect 15226 -760 15526 -742
rect 14816 -808 15116 -790
rect 14816 -842 14847 -808
rect 14881 -842 14915 -808
rect 14949 -842 14983 -808
rect 15017 -842 15051 -808
rect 15085 -842 15116 -808
rect 14816 -860 15116 -842
rect 15226 -808 15526 -790
rect 15226 -842 15257 -808
rect 15291 -842 15325 -808
rect 15359 -842 15393 -808
rect 15427 -842 15461 -808
rect 15495 -842 15526 -808
rect 15226 -860 15526 -842
rect 14816 -908 15116 -890
rect 14816 -942 14847 -908
rect 14881 -942 14915 -908
rect 14949 -942 14983 -908
rect 15017 -942 15051 -908
rect 15085 -942 15116 -908
rect 14816 -960 15116 -942
rect 15226 -908 15526 -890
rect 15226 -942 15257 -908
rect 15291 -942 15325 -908
rect 15359 -942 15393 -908
rect 15427 -942 15461 -908
rect 15495 -942 15526 -908
rect 15226 -960 15526 -942
rect 14816 -1008 15116 -990
rect 14816 -1042 14847 -1008
rect 14881 -1042 14915 -1008
rect 14949 -1042 14983 -1008
rect 15017 -1042 15051 -1008
rect 15085 -1042 15116 -1008
rect 14816 -1060 15116 -1042
rect 15226 -1008 15526 -990
rect 15226 -1042 15257 -1008
rect 15291 -1042 15325 -1008
rect 15359 -1042 15393 -1008
rect 15427 -1042 15461 -1008
rect 15495 -1042 15526 -1008
rect 15226 -1060 15526 -1042
rect 14816 -1108 15116 -1090
rect 14816 -1142 14847 -1108
rect 14881 -1142 14915 -1108
rect 14949 -1142 14983 -1108
rect 15017 -1142 15051 -1108
rect 15085 -1142 15116 -1108
rect 14816 -1160 15116 -1142
rect 15226 -1108 15526 -1090
rect 15226 -1142 15257 -1108
rect 15291 -1142 15325 -1108
rect 15359 -1142 15393 -1108
rect 15427 -1142 15461 -1108
rect 15495 -1142 15526 -1108
rect 15226 -1160 15526 -1142
rect 14816 -1208 15116 -1190
rect 14816 -1242 14847 -1208
rect 14881 -1242 14915 -1208
rect 14949 -1242 14983 -1208
rect 15017 -1242 15051 -1208
rect 15085 -1242 15116 -1208
rect 14816 -1260 15116 -1242
rect 15226 -1208 15526 -1190
rect 15226 -1242 15257 -1208
rect 15291 -1242 15325 -1208
rect 15359 -1242 15393 -1208
rect 15427 -1242 15461 -1208
rect 15495 -1242 15526 -1208
rect 15226 -1260 15526 -1242
rect 14816 -1308 15116 -1290
rect 14816 -1342 14847 -1308
rect 14881 -1342 14915 -1308
rect 14949 -1342 14983 -1308
rect 15017 -1342 15051 -1308
rect 15085 -1342 15116 -1308
rect 14816 -1360 15116 -1342
rect 15226 -1308 15526 -1290
rect 15226 -1342 15257 -1308
rect 15291 -1342 15325 -1308
rect 15359 -1342 15393 -1308
rect 15427 -1342 15461 -1308
rect 15495 -1342 15526 -1308
rect 15226 -1360 15526 -1342
rect 14816 -1408 15116 -1390
rect 14816 -1442 14847 -1408
rect 14881 -1442 14915 -1408
rect 14949 -1442 14983 -1408
rect 15017 -1442 15051 -1408
rect 15085 -1442 15116 -1408
rect 14816 -1460 15116 -1442
rect 15226 -1408 15526 -1390
rect 15226 -1442 15257 -1408
rect 15291 -1442 15325 -1408
rect 15359 -1442 15393 -1408
rect 15427 -1442 15461 -1408
rect 15495 -1442 15526 -1408
rect 15226 -1460 15526 -1442
rect 14816 -1508 15116 -1490
rect 14816 -1542 14847 -1508
rect 14881 -1542 14915 -1508
rect 14949 -1542 14983 -1508
rect 15017 -1542 15051 -1508
rect 15085 -1542 15116 -1508
rect 14816 -1560 15116 -1542
rect 15226 -1508 15526 -1490
rect 15226 -1542 15257 -1508
rect 15291 -1542 15325 -1508
rect 15359 -1542 15393 -1508
rect 15427 -1542 15461 -1508
rect 15495 -1542 15526 -1508
rect 15226 -1560 15526 -1542
rect 14816 -1608 15116 -1590
rect 14816 -1642 14847 -1608
rect 14881 -1642 14915 -1608
rect 14949 -1642 14983 -1608
rect 15017 -1642 15051 -1608
rect 15085 -1642 15116 -1608
rect 14816 -1660 15116 -1642
rect 15226 -1608 15526 -1590
rect 15226 -1642 15257 -1608
rect 15291 -1642 15325 -1608
rect 15359 -1642 15393 -1608
rect 15427 -1642 15461 -1608
rect 15495 -1642 15526 -1608
rect 15226 -1660 15526 -1642
rect 14816 -1708 15116 -1690
rect 14816 -1742 14847 -1708
rect 14881 -1742 14915 -1708
rect 14949 -1742 14983 -1708
rect 15017 -1742 15051 -1708
rect 15085 -1742 15116 -1708
rect 14816 -1760 15116 -1742
rect 15226 -1708 15526 -1690
rect 15226 -1742 15257 -1708
rect 15291 -1742 15325 -1708
rect 15359 -1742 15393 -1708
rect 15427 -1742 15461 -1708
rect 15495 -1742 15526 -1708
rect 15226 -1760 15526 -1742
rect 14816 -1808 15116 -1790
rect 14816 -1842 14847 -1808
rect 14881 -1842 14915 -1808
rect 14949 -1842 14983 -1808
rect 15017 -1842 15051 -1808
rect 15085 -1842 15116 -1808
rect 14816 -1860 15116 -1842
rect 15226 -1808 15526 -1790
rect 15226 -1842 15257 -1808
rect 15291 -1842 15325 -1808
rect 15359 -1842 15393 -1808
rect 15427 -1842 15461 -1808
rect 15495 -1842 15526 -1808
rect 15226 -1860 15526 -1842
rect 14816 -1908 15116 -1890
rect 14816 -1942 14847 -1908
rect 14881 -1942 14915 -1908
rect 14949 -1942 14983 -1908
rect 15017 -1942 15051 -1908
rect 15085 -1942 15116 -1908
rect 14816 -1960 15116 -1942
rect 15226 -1908 15526 -1890
rect 15226 -1942 15257 -1908
rect 15291 -1942 15325 -1908
rect 15359 -1942 15393 -1908
rect 15427 -1942 15461 -1908
rect 15495 -1942 15526 -1908
rect 15226 -1960 15526 -1942
rect 14816 -2008 15116 -1990
rect 14816 -2042 14847 -2008
rect 14881 -2042 14915 -2008
rect 14949 -2042 14983 -2008
rect 15017 -2042 15051 -2008
rect 15085 -2042 15116 -2008
rect 14816 -2079 15116 -2042
rect 15226 -2008 15526 -1990
rect 15226 -2042 15257 -2008
rect 15291 -2042 15325 -2008
rect 15359 -2042 15393 -2008
rect 15427 -2042 15461 -2008
rect 15495 -2042 15526 -2008
rect 15226 -2079 15526 -2042
<< ndiffc >>
rect 24 4753 58 4787
rect 118 4753 152 4787
rect 218 4753 252 4787
rect 312 4753 346 4787
rect 424 4753 458 4787
rect 518 4753 552 4787
rect 618 4753 652 4787
rect 1018 4753 1052 4787
rect 1112 4753 1146 4787
rect 118 4613 152 4647
rect 218 4613 252 4647
rect 618 4613 652 4647
rect 718 4613 752 4647
rect 918 4613 952 4647
rect 1018 4613 1052 4647
rect 1112 4613 1146 4647
rect 218 4473 252 4507
rect 312 4473 346 4507
rect 1224 4753 1258 4787
rect 1318 4753 1352 4787
rect 1418 4753 1452 4787
rect 1618 4753 1652 4787
rect 1718 4753 1752 4787
rect 1818 4753 1852 4787
rect 1918 4753 1952 4787
rect 2218 4753 2252 4787
rect 2312 4753 2346 4787
rect 2424 4753 2458 4787
rect 2518 4753 2552 4787
rect 2618 4753 2652 4787
rect 2918 4753 2952 4787
rect 3018 4753 3052 4787
rect 3112 4753 3146 4787
rect 1224 4613 1258 4647
rect 1318 4613 1352 4647
rect 1518 4613 1552 4647
rect 1618 4613 1652 4647
rect 1718 4613 1752 4647
rect 2018 4613 2052 4647
rect 2118 4613 2152 4647
rect 2618 4613 2652 4647
rect 2718 4613 2752 4647
rect 2818 4613 2852 4647
rect 2912 4613 2946 4647
rect 424 4473 458 4507
rect 518 4473 552 4507
rect 618 4473 652 4507
rect 718 4473 752 4507
rect 818 4473 852 4507
rect 1018 4473 1052 4507
rect 1118 4473 1152 4507
rect 1418 4473 1452 4507
rect 1518 4473 1552 4507
rect 1612 4473 1646 4507
rect 24 4333 58 4367
rect 118 4333 152 4367
rect 218 4333 252 4367
rect 418 4333 452 4367
rect 518 4333 552 4367
rect 1018 4333 1052 4367
rect 1118 4333 1152 4367
rect 1212 4333 1246 4367
rect 118 4193 152 4227
rect 218 4193 252 4227
rect 418 4193 452 4227
rect 512 4193 546 4227
rect 24 4053 58 4087
rect 118 4053 152 4087
rect 212 4053 246 4087
rect 324 4053 358 4087
rect 412 4053 446 4087
rect 624 4193 658 4227
rect 718 4193 752 4227
rect 1018 4193 1052 4227
rect 1112 4193 1146 4227
rect 1724 4473 1758 4507
rect 1812 4473 1846 4507
rect 1924 4473 1958 4507
rect 2018 4473 2052 4507
rect 2118 4473 2152 4507
rect 2218 4473 2252 4507
rect 2312 4473 2346 4507
rect 1324 4333 1358 4367
rect 1418 4333 1452 4367
rect 1518 4333 1552 4367
rect 1718 4333 1752 4367
rect 1818 4333 1852 4367
rect 1912 4333 1946 4367
rect 1224 4193 1258 4227
rect 1318 4193 1352 4227
rect 1418 4193 1452 4227
rect 1518 4193 1552 4227
rect 1618 4193 1652 4227
rect 1718 4193 1752 4227
rect 1818 4193 1852 4227
rect 1912 4193 1946 4227
rect 524 4053 558 4087
rect 618 4053 652 4087
rect 918 4053 952 4087
rect 1018 4053 1052 4087
rect 1118 4053 1152 4087
rect 1218 4053 1252 4087
rect 1312 4053 1346 4087
rect 1424 4053 1458 4087
rect 1518 4053 1552 4087
rect 1612 4053 1646 4087
rect 2424 4473 2458 4507
rect 2518 4473 2552 4507
rect 2612 4473 2646 4507
rect 2724 4473 2758 4507
rect 2812 4473 2846 4507
rect 3224 4753 3258 4787
rect 3318 4753 3352 4787
rect 3412 4753 3446 4787
rect 3524 4753 3558 4787
rect 3618 4753 3652 4787
rect 3918 4753 3952 4787
rect 4018 4753 4052 4787
rect 4118 4753 4152 4787
rect 4212 4753 4246 4787
rect 3024 4613 3058 4647
rect 3118 4613 3152 4647
rect 3218 4613 3252 4647
rect 3318 4613 3352 4647
rect 3518 4613 3552 4647
rect 3612 4613 3646 4647
rect 4324 4753 4358 4787
rect 4418 4753 4452 4787
rect 4518 4753 4552 4787
rect 4618 4753 4652 4787
rect 4718 4753 4752 4787
rect 4918 4753 4952 4787
rect 5018 4753 5052 4787
rect 5318 4753 5352 4787
rect 5418 4753 5452 4787
rect 5518 4753 5552 4787
rect 5918 4753 5952 4787
rect 6018 4753 6052 4787
rect 6318 4753 6352 4787
rect 6412 4753 6446 4787
rect 3724 4613 3758 4647
rect 3818 4613 3852 4647
rect 4018 4613 4052 4647
rect 4118 4613 4152 4647
rect 4318 4613 4352 4647
rect 4418 4613 4452 4647
rect 4618 4613 4652 4647
rect 4712 4613 4746 4647
rect 2924 4473 2958 4507
rect 3018 4473 3052 4507
rect 3518 4473 3552 4507
rect 3618 4473 3652 4507
rect 3712 4473 3746 4507
rect 2024 4333 2058 4367
rect 2118 4333 2152 4367
rect 2218 4333 2252 4367
rect 2318 4333 2352 4367
rect 2418 4333 2452 4367
rect 2518 4333 2552 4367
rect 2818 4333 2852 4367
rect 2918 4333 2952 4367
rect 3118 4333 3152 4367
rect 3218 4333 3252 4367
rect 3318 4333 3352 4367
rect 3518 4333 3552 4367
rect 3618 4333 3652 4367
rect 3712 4333 3746 4367
rect 4824 4613 4858 4647
rect 4918 4613 4952 4647
rect 5012 4613 5046 4647
rect 3824 4473 3858 4507
rect 3918 4473 3952 4507
rect 4018 4473 4052 4507
rect 4118 4473 4152 4507
rect 4218 4473 4252 4507
rect 4318 4473 4352 4507
rect 4618 4473 4652 4507
rect 4718 4473 4752 4507
rect 4918 4473 4952 4507
rect 5012 4473 5046 4507
rect 5124 4613 5158 4647
rect 5218 4613 5252 4647
rect 5318 4613 5352 4647
rect 5718 4613 5752 4647
rect 5812 4613 5846 4647
rect 5124 4473 5158 4507
rect 5218 4473 5252 4507
rect 5312 4473 5346 4507
rect 5924 4613 5958 4647
rect 6018 4613 6052 4647
rect 6118 4613 6152 4647
rect 6218 4613 6252 4647
rect 6318 4613 6352 4647
rect 6412 4613 6446 4647
rect 5424 4473 5458 4507
rect 5518 4473 5552 4507
rect 5918 4473 5952 4507
rect 6012 4473 6046 4507
rect 3824 4333 3858 4367
rect 3918 4333 3952 4367
rect 4018 4333 4052 4367
rect 4118 4333 4152 4367
rect 4218 4333 4252 4367
rect 4418 4333 4452 4367
rect 4518 4333 4552 4367
rect 4618 4333 4652 4367
rect 4818 4333 4852 4367
rect 4918 4333 4952 4367
rect 5018 4333 5052 4367
rect 5218 4333 5252 4367
rect 5318 4333 5352 4367
rect 5518 4333 5552 4367
rect 5618 4333 5652 4367
rect 5918 4333 5952 4367
rect 6012 4333 6046 4367
rect 2024 4193 2058 4227
rect 2118 4193 2152 4227
rect 2318 4193 2352 4227
rect 2418 4193 2452 4227
rect 2518 4193 2552 4227
rect 2818 4193 2852 4227
rect 2918 4193 2952 4227
rect 3018 4193 3052 4227
rect 3218 4193 3252 4227
rect 3318 4193 3352 4227
rect 3618 4193 3652 4227
rect 3718 4193 3752 4227
rect 3818 4193 3852 4227
rect 3918 4193 3952 4227
rect 4012 4193 4046 4227
rect 1724 4053 1758 4087
rect 1818 4053 1852 4087
rect 2018 4053 2052 4087
rect 2118 4053 2152 4087
rect 2212 4053 2246 4087
rect 24 3913 58 3947
rect 118 3913 152 3947
rect 218 3913 252 3947
rect 318 3913 352 3947
rect 618 3913 652 3947
rect 718 3913 752 3947
rect 918 3913 952 3947
rect 1018 3913 1052 3947
rect 1118 3913 1152 3947
rect 1518 3913 1552 3947
rect 1618 3913 1652 3947
rect 1818 3913 1852 3947
rect 1912 3913 1946 3947
rect 2324 4053 2358 4087
rect 2418 4053 2452 4087
rect 2518 4053 2552 4087
rect 2612 4053 2646 4087
rect 2724 4053 2758 4087
rect 2818 4053 2852 4087
rect 2912 4053 2946 4087
rect 3024 4053 3058 4087
rect 3118 4053 3152 4087
rect 3212 4053 3246 4087
rect 4124 4193 4158 4227
rect 4212 4193 4246 4227
rect 3324 4053 3358 4087
rect 3418 4053 3452 4087
rect 3518 4053 3552 4087
rect 3618 4053 3652 4087
rect 3918 4053 3952 4087
rect 4018 4053 4052 4087
rect 4112 4053 4146 4087
rect 2024 3913 2058 3947
rect 2118 3913 2152 3947
rect 2918 3913 2952 3947
rect 3018 3913 3052 3947
rect 3118 3913 3152 3947
rect 3218 3913 3252 3947
rect 3318 3913 3352 3947
rect 3618 3913 3652 3947
rect 3718 3913 3752 3947
rect 3818 3913 3852 3947
rect 3912 3913 3946 3947
rect 24 3773 58 3807
rect 118 3773 152 3807
rect 218 3773 252 3807
rect 618 3773 652 3807
rect 718 3773 752 3807
rect 1018 3773 1052 3807
rect 1118 3773 1152 3807
rect 1718 3773 1752 3807
rect 1818 3773 1852 3807
rect 2018 3773 2052 3807
rect 2112 3773 2146 3807
rect 518 3543 552 3577
rect 618 3543 652 3577
rect 718 3543 752 3577
rect 812 3543 846 3577
rect 24 3403 58 3437
rect 118 3403 152 3437
rect 218 3403 252 3437
rect 312 3403 346 3437
rect 424 3403 458 3437
rect 512 3403 546 3437
rect 624 3403 658 3437
rect 712 3403 746 3437
rect 118 3263 152 3297
rect 218 3263 252 3297
rect 318 3263 352 3297
rect 418 3263 452 3297
rect 518 3263 552 3297
rect 618 3263 652 3297
rect 712 3263 746 3297
rect 24 3123 58 3157
rect 112 3123 146 3157
rect 924 3543 958 3577
rect 1012 3543 1046 3577
rect 824 3403 858 3437
rect 912 3403 946 3437
rect 824 3263 858 3297
rect 912 3263 946 3297
rect 2224 3773 2258 3807
rect 2318 3773 2352 3807
rect 2418 3773 2452 3807
rect 2512 3773 2546 3807
rect 2624 3773 2658 3807
rect 2712 3773 2746 3807
rect 1124 3543 1158 3577
rect 1218 3543 1252 3577
rect 1318 3543 1352 3577
rect 1418 3543 1452 3577
rect 1618 3543 1652 3577
rect 1718 3543 1752 3577
rect 1818 3543 1852 3577
rect 1918 3543 1952 3577
rect 2018 3543 2052 3577
rect 2118 3543 2152 3577
rect 2218 3543 2252 3577
rect 2318 3543 2352 3577
rect 2418 3543 2452 3577
rect 2512 3543 2546 3577
rect 2824 3773 2858 3807
rect 2918 3773 2952 3807
rect 3018 3773 3052 3807
rect 3112 3773 3146 3807
rect 4024 3913 4058 3947
rect 4112 3913 4146 3947
rect 4324 4193 4358 4227
rect 4412 4193 4446 4227
rect 4224 4053 4258 4087
rect 4312 4053 4346 4087
rect 4524 4193 4558 4227
rect 4612 4193 4646 4227
rect 4424 4053 4458 4087
rect 4512 4053 4546 4087
rect 4724 4193 4758 4227
rect 4812 4193 4846 4227
rect 4624 4053 4658 4087
rect 4712 4053 4746 4087
rect 4924 4193 4958 4227
rect 5018 4193 5052 4227
rect 5318 4193 5352 4227
rect 5418 4193 5452 4227
rect 5512 4193 5546 4227
rect 4824 4053 4858 4087
rect 4912 4053 4946 4087
rect 5024 4053 5058 4087
rect 5118 4053 5152 4087
rect 5212 4053 5246 4087
rect 4224 3913 4258 3947
rect 4318 3913 4352 3947
rect 4418 3913 4452 3947
rect 4618 3913 4652 3947
rect 4718 3913 4752 3947
rect 4918 3913 4952 3947
rect 5012 3913 5046 3947
rect 3224 3773 3258 3807
rect 3318 3773 3352 3807
rect 3618 3773 3652 3807
rect 3718 3773 3752 3807
rect 3918 3773 3952 3807
rect 4018 3773 4052 3807
rect 4218 3773 4252 3807
rect 4318 3773 4352 3807
rect 4418 3773 4452 3807
rect 4512 3773 4546 3807
rect 2624 3543 2658 3577
rect 2718 3543 2752 3577
rect 2918 3543 2952 3577
rect 3018 3543 3052 3577
rect 3112 3543 3146 3577
rect 5124 3913 5158 3947
rect 5212 3913 5246 3947
rect 5624 4193 5658 4227
rect 5718 4193 5752 4227
rect 5918 4193 5952 4227
rect 6012 4193 6046 4227
rect 5324 4053 5358 4087
rect 5418 4053 5452 4087
rect 5518 4053 5552 4087
rect 5612 4053 5646 4087
rect 5324 3913 5358 3947
rect 5418 3913 5452 3947
rect 5512 3913 5546 3947
rect 4624 3773 4658 3807
rect 4718 3773 4752 3807
rect 5018 3773 5052 3807
rect 5118 3773 5152 3807
rect 5318 3773 5352 3807
rect 5412 3773 5446 3807
rect 3224 3543 3258 3577
rect 3318 3543 3352 3577
rect 3518 3543 3552 3577
rect 3618 3543 3652 3577
rect 3718 3543 3752 3577
rect 4018 3543 4052 3577
rect 4118 3543 4152 3577
rect 4318 3543 4352 3577
rect 4412 3543 4446 3577
rect 1024 3403 1058 3437
rect 1118 3403 1152 3437
rect 1218 3403 1252 3437
rect 1418 3403 1452 3437
rect 1518 3403 1552 3437
rect 1618 3403 1652 3437
rect 1718 3403 1752 3437
rect 1818 3403 1852 3437
rect 1918 3403 1952 3437
rect 2018 3403 2052 3437
rect 2118 3403 2152 3437
rect 2518 3403 2552 3437
rect 2618 3403 2652 3437
rect 2718 3403 2752 3437
rect 3018 3403 3052 3437
rect 3118 3403 3152 3437
rect 3618 3403 3652 3437
rect 3718 3403 3752 3437
rect 3812 3403 3846 3437
rect 1024 3263 1058 3297
rect 1118 3263 1152 3297
rect 1218 3263 1252 3297
rect 1318 3263 1352 3297
rect 1418 3263 1452 3297
rect 1518 3263 1552 3297
rect 1618 3263 1652 3297
rect 1718 3263 1752 3297
rect 1818 3263 1852 3297
rect 1918 3263 1952 3297
rect 2018 3263 2052 3297
rect 2118 3263 2152 3297
rect 2218 3263 2252 3297
rect 2318 3263 2352 3297
rect 2418 3263 2452 3297
rect 2618 3263 2652 3297
rect 2712 3263 2746 3297
rect 224 3123 258 3157
rect 318 3123 352 3157
rect 418 3123 452 3157
rect 518 3123 552 3157
rect 618 3123 652 3157
rect 818 3123 852 3157
rect 918 3123 952 3157
rect 1218 3123 1252 3157
rect 1312 3123 1346 3157
rect 118 2983 152 3017
rect 218 2983 252 3017
rect 418 2983 452 3017
rect 518 2983 552 3017
rect 612 2983 646 3017
rect 1424 3123 1458 3157
rect 1518 3123 1552 3157
rect 1718 3123 1752 3157
rect 1818 3123 1852 3157
rect 2018 3123 2052 3157
rect 2118 3123 2152 3157
rect 2318 3123 2352 3157
rect 2418 3123 2452 3157
rect 2512 3123 2546 3157
rect 724 2983 758 3017
rect 818 2983 852 3017
rect 918 2983 952 3017
rect 1218 2983 1252 3017
rect 1318 2983 1352 3017
rect 1818 2983 1852 3017
rect 1918 2983 1952 3017
rect 2012 2983 2046 3017
rect 24 2843 58 2877
rect 118 2843 152 2877
rect 218 2843 252 2877
rect 418 2843 452 2877
rect 518 2843 552 2877
rect 618 2843 652 2877
rect 718 2843 752 2877
rect 812 2843 846 2877
rect 2824 3263 2858 3297
rect 2918 3263 2952 3297
rect 3018 3263 3052 3297
rect 3118 3263 3152 3297
rect 3212 3263 3246 3297
rect 2624 3123 2658 3157
rect 2718 3123 2752 3157
rect 2818 3123 2852 3157
rect 2918 3123 2952 3157
rect 3118 3123 3152 3157
rect 3212 3123 3246 3157
rect 2124 2983 2158 3017
rect 2218 2983 2252 3017
rect 2418 2983 2452 3017
rect 2518 2983 2552 3017
rect 2718 2983 2752 3017
rect 2818 2983 2852 3017
rect 2918 2983 2952 3017
rect 3012 2983 3046 3017
rect 924 2843 958 2877
rect 1018 2843 1052 2877
rect 1118 2843 1152 2877
rect 1318 2843 1352 2877
rect 1418 2843 1452 2877
rect 1818 2843 1852 2877
rect 1918 2843 1952 2877
rect 2018 2843 2052 2877
rect 2518 2843 2552 2877
rect 2612 2843 2646 2877
rect 218 2703 252 2737
rect 318 2703 352 2737
rect 418 2703 452 2737
rect 518 2703 552 2737
rect 1018 2703 1052 2737
rect 1112 2703 1146 2737
rect 1224 2703 1258 2737
rect 1318 2703 1352 2737
rect 1818 2703 1852 2737
rect 1918 2703 1952 2737
rect 2218 2703 2252 2737
rect 2312 2703 2346 2737
rect 2724 2843 2758 2877
rect 2818 2843 2852 2877
rect 2912 2843 2946 2877
rect 3324 3263 3358 3297
rect 3412 3263 3446 3297
rect 3924 3403 3958 3437
rect 4018 3403 4052 3437
rect 4118 3403 4152 3437
rect 4218 3403 4252 3437
rect 4318 3403 4352 3437
rect 4412 3403 4446 3437
rect 6524 4753 6558 4787
rect 6618 4753 6652 4787
rect 6718 4753 6752 4787
rect 7018 4753 7052 4787
rect 7118 4753 7152 4787
rect 7318 4753 7352 4787
rect 7418 4753 7452 4787
rect 7518 4753 7552 4787
rect 7618 4753 7652 4787
rect 7718 4753 7752 4787
rect 7818 4753 7852 4787
rect 8118 4753 8152 4787
rect 8218 4753 8252 4787
rect 8318 4753 8352 4787
rect 8418 4753 8452 4787
rect 8818 4753 8852 4787
rect 8918 4753 8952 4787
rect 9718 4753 9752 4787
rect 9812 4753 9846 4787
rect 6524 4613 6558 4647
rect 6618 4613 6652 4647
rect 6718 4613 6752 4647
rect 6818 4613 6852 4647
rect 6918 4613 6952 4647
rect 7018 4613 7052 4647
rect 7118 4613 7152 4647
rect 7218 4613 7252 4647
rect 7918 4613 7952 4647
rect 8018 4613 8052 4647
rect 8118 4613 8152 4647
rect 8218 4613 8252 4647
rect 8318 4613 8352 4647
rect 8618 4613 8652 4647
rect 8712 4613 8746 4647
rect 6124 4473 6158 4507
rect 6218 4473 6252 4507
rect 7018 4473 7052 4507
rect 7118 4473 7152 4507
rect 7218 4473 7252 4507
rect 7718 4473 7752 4507
rect 7818 4473 7852 4507
rect 7918 4473 7952 4507
rect 8012 4473 8046 4507
rect 6124 4333 6158 4367
rect 6218 4333 6252 4367
rect 6418 4333 6452 4367
rect 6518 4333 6552 4367
rect 6612 4333 6646 4367
rect 6124 4193 6158 4227
rect 6212 4193 6246 4227
rect 6324 4193 6358 4227
rect 6412 4193 6446 4227
rect 6524 4193 6558 4227
rect 6612 4193 6646 4227
rect 6724 4333 6758 4367
rect 6818 4333 6852 4367
rect 7118 4333 7152 4367
rect 7218 4333 7252 4367
rect 7312 4333 7346 4367
rect 6724 4193 6758 4227
rect 6818 4193 6852 4227
rect 7018 4193 7052 4227
rect 7112 4193 7146 4227
rect 8124 4473 8158 4507
rect 8218 4473 8252 4507
rect 8312 4473 8346 4507
rect 9924 4753 9958 4787
rect 10018 4753 10052 4787
rect 10118 4753 10152 4787
rect 10418 4753 10452 4787
rect 10518 4753 10552 4787
rect 10618 4753 10652 4787
rect 10712 4753 10746 4787
rect 10824 4753 10858 4787
rect 10918 4753 10952 4787
rect 11118 4753 11152 4787
rect 11218 4753 11252 4787
rect 11318 4753 11352 4787
rect 11518 4753 11552 4787
rect 11612 4753 11646 4787
rect 11724 4753 11758 4787
rect 11818 4753 11852 4787
rect 11918 4753 11952 4787
rect 12118 4753 12152 4787
rect 12218 4753 12252 4787
rect 12318 4753 12352 4787
rect 12412 4753 12446 4787
rect 12524 4753 12558 4787
rect 12618 4753 12652 4787
rect 12718 4753 12752 4787
rect 12812 4753 12846 4787
rect 12924 4768 12958 4802
rect 13018 4753 13052 4787
rect 13112 4738 13146 4772
rect 13228 4753 13262 4787
rect 13328 4753 13362 4787
rect 13428 4753 13462 4787
rect 13528 4753 13562 4787
rect 13628 4753 13662 4787
rect 8824 4613 8858 4647
rect 8918 4613 8952 4647
rect 9318 4613 9352 4647
rect 9418 4613 9452 4647
rect 9518 4613 9552 4647
rect 9618 4613 9652 4647
rect 9718 4613 9752 4647
rect 9918 4613 9952 4647
rect 10018 4613 10052 4647
rect 10118 4613 10152 4647
rect 10518 4613 10552 4647
rect 10618 4613 10652 4647
rect 11118 4613 11152 4647
rect 11218 4613 11252 4647
rect 11418 4613 11452 4647
rect 11518 4613 11552 4647
rect 11618 4613 11652 4647
rect 11718 4613 11752 4647
rect 11818 4613 11852 4647
rect 11918 4613 11952 4647
rect 12318 4613 12352 4647
rect 12418 4613 12452 4647
rect 12518 4613 12552 4647
rect 12612 4613 12646 4647
rect 8424 4473 8458 4507
rect 8518 4473 8552 4507
rect 8618 4473 8652 4507
rect 8718 4473 8752 4507
rect 8812 4473 8846 4507
rect 8924 4473 8958 4507
rect 9012 4473 9046 4507
rect 9124 4473 9158 4507
rect 9218 4473 9252 4507
rect 9312 4473 9346 4507
rect 9424 4473 9458 4507
rect 9518 4473 9552 4507
rect 9612 4473 9646 4507
rect 9724 4473 9758 4507
rect 9818 4473 9852 4507
rect 9912 4473 9946 4507
rect 10024 4473 10058 4507
rect 10118 4473 10152 4507
rect 10212 4473 10246 4507
rect 10324 4473 10358 4507
rect 10418 4473 10452 4507
rect 10512 4473 10546 4507
rect 10624 4473 10658 4507
rect 10712 4473 10746 4507
rect 10824 4473 10858 4507
rect 10912 4473 10946 4507
rect 7424 4333 7458 4367
rect 7518 4333 7552 4367
rect 7618 4333 7652 4367
rect 7718 4333 7752 4367
rect 8018 4333 8052 4367
rect 8118 4333 8152 4367
rect 8318 4333 8352 4367
rect 8418 4333 8452 4367
rect 8618 4333 8652 4367
rect 8718 4333 8752 4367
rect 8918 4333 8952 4367
rect 9018 4333 9052 4367
rect 9118 4333 9152 4367
rect 9318 4333 9352 4367
rect 9418 4333 9452 4367
rect 9918 4333 9952 4367
rect 10018 4333 10052 4367
rect 10118 4333 10152 4367
rect 10318 4333 10352 4367
rect 10418 4333 10452 4367
rect 10618 4333 10652 4367
rect 10718 4333 10752 4367
rect 10812 4333 10846 4367
rect 7224 4193 7258 4227
rect 7318 4193 7352 4227
rect 7518 4193 7552 4227
rect 7618 4193 7652 4227
rect 7718 4193 7752 4227
rect 7918 4193 7952 4227
rect 8018 4193 8052 4227
rect 8112 4193 8146 4227
rect 5724 4053 5758 4087
rect 5818 4053 5852 4087
rect 6218 4053 6252 4087
rect 6318 4053 6352 4087
rect 6418 4053 6452 4087
rect 6518 4053 6552 4087
rect 6818 4053 6852 4087
rect 6918 4053 6952 4087
rect 7018 4053 7052 4087
rect 7118 4053 7152 4087
rect 7218 4053 7252 4087
rect 7312 4053 7346 4087
rect 5624 3913 5658 3947
rect 5718 3913 5752 3947
rect 5818 3913 5852 3947
rect 5912 3913 5946 3947
rect 5524 3773 5558 3807
rect 5618 3773 5652 3807
rect 5718 3773 5752 3807
rect 5818 3773 5852 3807
rect 5912 3773 5946 3807
rect 4524 3543 4558 3577
rect 4618 3543 4652 3577
rect 4718 3543 4752 3577
rect 5118 3543 5152 3577
rect 5218 3543 5252 3577
rect 5418 3543 5452 3577
rect 5518 3543 5552 3577
rect 5618 3543 5652 3577
rect 5712 3543 5746 3577
rect 4524 3403 4558 3437
rect 4618 3403 4652 3437
rect 4718 3403 4752 3437
rect 4812 3403 4846 3437
rect 4924 3403 4958 3437
rect 5012 3403 5046 3437
rect 6024 3913 6058 3947
rect 6118 3913 6152 3947
rect 6218 3913 6252 3947
rect 6318 3913 6352 3947
rect 6618 3913 6652 3947
rect 6718 3913 6752 3947
rect 6818 3913 6852 3947
rect 6912 3913 6946 3947
rect 7024 3913 7058 3947
rect 7112 3913 7146 3947
rect 7424 4053 7458 4087
rect 7518 4053 7552 4087
rect 7612 4053 7646 4087
rect 7724 4053 7758 4087
rect 7812 4053 7846 4087
rect 8224 4193 8258 4227
rect 8312 4193 8346 4227
rect 8424 4193 8458 4227
rect 8512 4193 8546 4227
rect 8624 4193 8658 4227
rect 8712 4193 8746 4227
rect 7924 4053 7958 4087
rect 8018 4053 8052 4087
rect 8118 4053 8152 4087
rect 8418 4053 8452 4087
rect 8518 4053 8552 4087
rect 8618 4053 8652 4087
rect 8712 4053 8746 4087
rect 7224 3913 7258 3947
rect 7318 3913 7352 3947
rect 7418 3913 7452 3947
rect 7518 3913 7552 3947
rect 7618 3913 7652 3947
rect 8018 3913 8052 3947
rect 8118 3913 8152 3947
rect 8518 3913 8552 3947
rect 8618 3913 8652 3947
rect 8712 3913 8746 3947
rect 6024 3773 6058 3807
rect 6118 3773 6152 3807
rect 6518 3773 6552 3807
rect 6618 3773 6652 3807
rect 7118 3773 7152 3807
rect 7218 3773 7252 3807
rect 7518 3773 7552 3807
rect 7612 3773 7646 3807
rect 8824 4193 8858 4227
rect 8912 4193 8946 4227
rect 8824 4053 8858 4087
rect 8912 4053 8946 4087
rect 9024 4193 9058 4227
rect 9118 4193 9152 4227
rect 9218 4193 9252 4227
rect 9312 4193 9346 4227
rect 9424 4193 9458 4227
rect 9512 4193 9546 4227
rect 9024 4053 9058 4087
rect 9118 4053 9152 4087
rect 9318 4053 9352 4087
rect 9418 4053 9452 4087
rect 9512 4053 9546 4087
rect 8824 3913 8858 3947
rect 8918 3913 8952 3947
rect 9418 3913 9452 3947
rect 9512 3913 9546 3947
rect 7724 3773 7758 3807
rect 7818 3773 7852 3807
rect 7918 3773 7952 3807
rect 8018 3773 8052 3807
rect 8118 3773 8152 3807
rect 8218 3773 8252 3807
rect 8318 3773 8352 3807
rect 8418 3773 8452 3807
rect 8618 3773 8652 3807
rect 8718 3773 8752 3807
rect 8818 3773 8852 3807
rect 9218 3773 9252 3807
rect 9318 3773 9352 3807
rect 9412 3773 9446 3807
rect 5824 3543 5858 3577
rect 5918 3543 5952 3577
rect 6018 3543 6052 3577
rect 6618 3543 6652 3577
rect 6718 3543 6752 3577
rect 6818 3543 6852 3577
rect 7418 3543 7452 3577
rect 7518 3543 7552 3577
rect 7618 3543 7652 3577
rect 8018 3543 8052 3577
rect 8118 3543 8152 3577
rect 8318 3543 8352 3577
rect 8418 3543 8452 3577
rect 8518 3543 8552 3577
rect 8818 3543 8852 3577
rect 8912 3543 8946 3577
rect 5124 3403 5158 3437
rect 5218 3403 5252 3437
rect 5418 3403 5452 3437
rect 5518 3403 5552 3437
rect 5618 3403 5652 3437
rect 5918 3403 5952 3437
rect 6012 3403 6046 3437
rect 6124 3403 6158 3437
rect 6218 3403 6252 3437
rect 6318 3403 6352 3437
rect 6412 3403 6446 3437
rect 6524 3403 6558 3437
rect 6618 3403 6652 3437
rect 6712 3403 6746 3437
rect 9024 3543 9058 3577
rect 9112 3543 9146 3577
rect 9224 3543 9258 3577
rect 9312 3543 9346 3577
rect 9624 4193 9658 4227
rect 9712 4193 9746 4227
rect 9824 4193 9858 4227
rect 9918 4193 9952 4227
rect 10012 4193 10046 4227
rect 11024 4473 11058 4507
rect 11118 4473 11152 4507
rect 11212 4473 11246 4507
rect 10924 4333 10958 4367
rect 11018 4333 11052 4367
rect 11112 4333 11146 4367
rect 10124 4193 10158 4227
rect 10218 4193 10252 4227
rect 10618 4193 10652 4227
rect 10718 4193 10752 4227
rect 10818 4193 10852 4227
rect 10912 4193 10946 4227
rect 9624 4053 9658 4087
rect 9718 4053 9752 4087
rect 9918 4053 9952 4087
rect 10018 4053 10052 4087
rect 10118 4053 10152 4087
rect 10218 4053 10252 4087
rect 10318 4053 10352 4087
rect 10418 4053 10452 4087
rect 10518 4053 10552 4087
rect 10612 4053 10646 4087
rect 10724 4053 10758 4087
rect 10812 4053 10846 4087
rect 11324 4473 11358 4507
rect 11418 4473 11452 4507
rect 11518 4473 11552 4507
rect 11918 4473 11952 4507
rect 12018 4473 12052 4507
rect 12118 4473 12152 4507
rect 12318 4473 12352 4507
rect 12412 4473 12446 4507
rect 11224 4333 11258 4367
rect 11318 4333 11352 4367
rect 11418 4333 11452 4367
rect 11718 4333 11752 4367
rect 11818 4333 11852 4367
rect 11912 4333 11946 4367
rect 11024 4193 11058 4227
rect 11118 4193 11152 4227
rect 11218 4193 11252 4227
rect 11312 4193 11346 4227
rect 10924 4053 10958 4087
rect 11018 4053 11052 4087
rect 11218 4053 11252 4087
rect 11312 4053 11346 4087
rect 9624 3913 9658 3947
rect 9718 3913 9752 3947
rect 9818 3913 9852 3947
rect 10118 3913 10152 3947
rect 10218 3913 10252 3947
rect 10318 3913 10352 3947
rect 10418 3913 10452 3947
rect 10918 3913 10952 3947
rect 11012 3913 11046 3947
rect 9524 3773 9558 3807
rect 9618 3773 9652 3807
rect 9718 3773 9752 3807
rect 9918 3773 9952 3807
rect 10012 3773 10046 3807
rect 11424 4193 11458 4227
rect 11512 4193 11546 4227
rect 11424 4053 11458 4087
rect 11512 4053 11546 4087
rect 12724 4613 12758 4647
rect 12812 4613 12846 4647
rect 12924 4628 12958 4662
rect 13018 4613 13052 4647
rect 13112 4598 13146 4632
rect 13228 4613 13262 4647
rect 13328 4613 13362 4647
rect 13428 4613 13462 4647
rect 13528 4613 13562 4647
rect 13628 4613 13662 4647
rect 12524 4473 12558 4507
rect 12618 4473 12652 4507
rect 12718 4473 12752 4507
rect 12812 4473 12846 4507
rect 12924 4488 12958 4522
rect 13018 4473 13052 4507
rect 13112 4458 13146 4492
rect 13228 4473 13262 4507
rect 13328 4473 13362 4507
rect 13428 4473 13462 4507
rect 13528 4473 13562 4507
rect 13628 4473 13662 4507
rect 12024 4333 12058 4367
rect 12118 4333 12152 4367
rect 12218 4333 12252 4367
rect 12318 4333 12352 4367
rect 12518 4333 12552 4367
rect 12618 4333 12652 4367
rect 12718 4333 12752 4367
rect 12812 4333 12846 4367
rect 12924 4348 12958 4382
rect 13018 4333 13052 4367
rect 13112 4318 13146 4352
rect 13228 4333 13262 4367
rect 13328 4333 13362 4367
rect 13428 4333 13462 4367
rect 13528 4333 13562 4367
rect 13628 4333 13662 4367
rect 11624 4193 11658 4227
rect 11718 4193 11752 4227
rect 12618 4193 12652 4227
rect 12718 4193 12752 4227
rect 12924 4208 12958 4242
rect 13018 4193 13052 4227
rect 13112 4178 13146 4212
rect 13228 4193 13262 4227
rect 13328 4193 13362 4227
rect 13428 4193 13462 4227
rect 13528 4193 13562 4227
rect 13628 4193 13662 4227
rect 11624 4053 11658 4087
rect 11718 4053 11752 4087
rect 11812 4053 11846 4087
rect 11924 4053 11958 4087
rect 12018 4053 12052 4087
rect 12318 4053 12352 4087
rect 12418 4053 12452 4087
rect 12518 4053 12552 4087
rect 12612 4053 12646 4087
rect 12724 4053 12758 4087
rect 12812 4053 12846 4087
rect 12924 4068 12958 4102
rect 13018 4053 13052 4087
rect 13112 4038 13146 4072
rect 13228 4053 13262 4087
rect 13328 4053 13362 4087
rect 13428 4053 13462 4087
rect 13528 4053 13562 4087
rect 13628 4053 13662 4087
rect 11124 3913 11158 3947
rect 11218 3913 11252 3947
rect 11318 3913 11352 3947
rect 11718 3913 11752 3947
rect 11818 3913 11852 3947
rect 12118 3913 12152 3947
rect 12218 3913 12252 3947
rect 12318 3913 12352 3947
rect 12518 3913 12552 3947
rect 12618 3913 12652 3947
rect 12718 3913 12752 3947
rect 12812 3913 12846 3947
rect 12924 3928 12958 3962
rect 13018 3913 13052 3947
rect 13112 3898 13146 3932
rect 13228 3913 13262 3947
rect 13328 3913 13362 3947
rect 13428 3913 13462 3947
rect 13528 3913 13562 3947
rect 13628 3913 13662 3947
rect 10124 3773 10158 3807
rect 10218 3773 10252 3807
rect 10418 3773 10452 3807
rect 10518 3773 10552 3807
rect 10618 3773 10652 3807
rect 10718 3773 10752 3807
rect 10818 3773 10852 3807
rect 10918 3773 10952 3807
rect 11018 3773 11052 3807
rect 11112 3773 11146 3807
rect 9424 3543 9458 3577
rect 9518 3543 9552 3577
rect 9618 3543 9652 3577
rect 9718 3543 9752 3577
rect 9818 3543 9852 3577
rect 9918 3543 9952 3577
rect 10012 3543 10046 3577
rect 6824 3403 6858 3437
rect 6918 3403 6952 3437
rect 7318 3403 7352 3437
rect 7418 3403 7452 3437
rect 7718 3403 7752 3437
rect 7818 3403 7852 3437
rect 7918 3403 7952 3437
rect 8018 3403 8052 3437
rect 8418 3403 8452 3437
rect 8518 3403 8552 3437
rect 8618 3403 8652 3437
rect 8718 3403 8752 3437
rect 8918 3403 8952 3437
rect 9018 3403 9052 3437
rect 9118 3403 9152 3437
rect 9218 3403 9252 3437
rect 9318 3403 9352 3437
rect 9412 3403 9446 3437
rect 3524 3263 3558 3297
rect 3618 3263 3652 3297
rect 4118 3263 4152 3297
rect 4218 3263 4252 3297
rect 4318 3263 4352 3297
rect 4418 3263 4452 3297
rect 4718 3263 4752 3297
rect 4818 3263 4852 3297
rect 5018 3263 5052 3297
rect 5118 3263 5152 3297
rect 5218 3263 5252 3297
rect 5418 3263 5452 3297
rect 5518 3263 5552 3297
rect 5618 3263 5652 3297
rect 5818 3263 5852 3297
rect 5918 3263 5952 3297
rect 6018 3263 6052 3297
rect 6318 3263 6352 3297
rect 6418 3263 6452 3297
rect 6518 3263 6552 3297
rect 6618 3263 6652 3297
rect 6718 3263 6752 3297
rect 6818 3263 6852 3297
rect 7118 3263 7152 3297
rect 7218 3263 7252 3297
rect 7312 3263 7346 3297
rect 3324 3123 3358 3157
rect 3418 3123 3452 3157
rect 3518 3123 3552 3157
rect 3612 3123 3646 3157
rect 3724 3123 3758 3157
rect 3818 3123 3852 3157
rect 3918 3123 3952 3157
rect 4018 3123 4052 3157
rect 4118 3123 4152 3157
rect 4218 3123 4252 3157
rect 4318 3123 4352 3157
rect 4518 3123 4552 3157
rect 4618 3123 4652 3157
rect 4718 3123 4752 3157
rect 5218 3123 5252 3157
rect 5318 3123 5352 3157
rect 5412 3123 5446 3157
rect 3124 2983 3158 3017
rect 3218 2983 3252 3017
rect 3318 2983 3352 3017
rect 3418 2983 3452 3017
rect 3718 2983 3752 3017
rect 3812 2983 3846 3017
rect 3024 2843 3058 2877
rect 3118 2843 3152 2877
rect 3218 2843 3252 2877
rect 3312 2843 3346 2877
rect 3924 2983 3958 3017
rect 4018 2983 4052 3017
rect 4118 2983 4152 3017
rect 4218 2983 4252 3017
rect 4418 2983 4452 3017
rect 4512 2983 4546 3017
rect 3424 2843 3458 2877
rect 3518 2843 3552 2877
rect 3618 2843 3652 2877
rect 3718 2843 3752 2877
rect 3818 2843 3852 2877
rect 3912 2843 3946 2877
rect 4624 2983 4658 3017
rect 4718 2983 4752 3017
rect 4818 2983 4852 3017
rect 4912 2983 4946 3017
rect 5524 3123 5558 3157
rect 5612 3123 5646 3157
rect 5724 3123 5758 3157
rect 5812 3123 5846 3157
rect 5924 3123 5958 3157
rect 6018 3123 6052 3157
rect 6218 3123 6252 3157
rect 6312 3123 6346 3157
rect 5024 2983 5058 3017
rect 5118 2983 5152 3017
rect 5418 2983 5452 3017
rect 5518 2983 5552 3017
rect 5818 2983 5852 3017
rect 5912 2983 5946 3017
rect 4024 2843 4058 2877
rect 4118 2843 4152 2877
rect 4218 2843 4252 2877
rect 4418 2843 4452 2877
rect 4518 2843 4552 2877
rect 5218 2843 5252 2877
rect 5312 2843 5346 2877
rect 2424 2703 2458 2737
rect 2518 2703 2552 2737
rect 2618 2703 2652 2737
rect 2718 2703 2752 2737
rect 3018 2703 3052 2737
rect 3118 2703 3152 2737
rect 3218 2703 3252 2737
rect 3318 2703 3352 2737
rect 3518 2703 3552 2737
rect 3618 2703 3652 2737
rect 3918 2703 3952 2737
rect 4018 2703 4052 2737
rect 4112 2703 4146 2737
rect 118 2563 152 2597
rect 218 2563 252 2597
rect 418 2563 452 2597
rect 518 2563 552 2597
rect 618 2563 652 2597
rect 718 2563 752 2597
rect 1018 2563 1052 2597
rect 1118 2563 1152 2597
rect 1218 2563 1252 2597
rect 1318 2563 1352 2597
rect 1418 2563 1452 2597
rect 1518 2563 1552 2597
rect 1618 2563 1652 2597
rect 1818 2563 1852 2597
rect 1918 2563 1952 2597
rect 2018 2563 2052 2597
rect 2318 2563 2352 2597
rect 2418 2563 2452 2597
rect 2512 2563 2546 2597
rect 24 2333 58 2367
rect 112 2333 146 2367
rect 224 2333 258 2367
rect 318 2333 352 2367
rect 412 2333 446 2367
rect 524 2333 558 2367
rect 612 2333 646 2367
rect 724 2333 758 2367
rect 818 2333 852 2367
rect 918 2333 952 2367
rect 1418 2333 1452 2367
rect 1518 2333 1552 2367
rect 1718 2333 1752 2367
rect 1818 2333 1852 2367
rect 2018 2333 2052 2367
rect 2118 2333 2152 2367
rect 2218 2333 2252 2367
rect 2312 2333 2346 2367
rect 24 2193 58 2227
rect 118 2193 152 2227
rect 318 2193 352 2227
rect 418 2193 452 2227
rect 518 2193 552 2227
rect 718 2193 752 2227
rect 812 2193 846 2227
rect 318 2053 352 2087
rect 418 2053 452 2087
rect 518 2053 552 2087
rect 618 2053 652 2087
rect 712 2053 746 2087
rect 924 2193 958 2227
rect 1012 2193 1046 2227
rect 2624 2563 2658 2597
rect 2718 2563 2752 2597
rect 2818 2563 2852 2597
rect 2918 2563 2952 2597
rect 3018 2563 3052 2597
rect 3118 2563 3152 2597
rect 3218 2563 3252 2597
rect 3312 2563 3346 2597
rect 2424 2333 2458 2367
rect 2518 2333 2552 2367
rect 2612 2333 2646 2367
rect 1124 2193 1158 2227
rect 1218 2193 1252 2227
rect 1318 2193 1352 2227
rect 1618 2193 1652 2227
rect 1718 2193 1752 2227
rect 1918 2193 1952 2227
rect 2018 2193 2052 2227
rect 2518 2193 2552 2227
rect 2612 2193 2646 2227
rect 824 2053 858 2087
rect 918 2053 952 2087
rect 1318 2053 1352 2087
rect 1412 2053 1446 2087
rect 118 1913 152 1947
rect 218 1913 252 1947
rect 318 1913 352 1947
rect 418 1913 452 1947
rect 518 1913 552 1947
rect 618 1913 652 1947
rect 718 1913 752 1947
rect 818 1913 852 1947
rect 912 1913 946 1947
rect 3424 2563 3458 2597
rect 3518 2563 3552 2597
rect 3618 2563 3652 2597
rect 3818 2563 3852 2597
rect 3912 2563 3946 2597
rect 4024 2563 4058 2597
rect 4112 2563 4146 2597
rect 4224 2703 4258 2737
rect 4318 2703 4352 2737
rect 4518 2703 4552 2737
rect 4618 2703 4652 2737
rect 4712 2703 4746 2737
rect 4224 2563 4258 2597
rect 4312 2563 4346 2597
rect 4424 2563 4458 2597
rect 4518 2563 4552 2597
rect 4618 2563 4652 2597
rect 4712 2563 4746 2597
rect 4824 2703 4858 2737
rect 4918 2703 4952 2737
rect 5018 2703 5052 2737
rect 5112 2703 5146 2737
rect 5224 2703 5258 2737
rect 5312 2703 5346 2737
rect 6424 3123 6458 3157
rect 6512 3123 6546 3157
rect 6624 3123 6658 3157
rect 6718 3123 6752 3157
rect 6818 3123 6852 3157
rect 6918 3123 6952 3157
rect 7012 3123 7046 3157
rect 9524 3403 9558 3437
rect 9618 3403 9652 3437
rect 9712 3403 9746 3437
rect 7424 3263 7458 3297
rect 7518 3263 7552 3297
rect 7618 3263 7652 3297
rect 7718 3263 7752 3297
rect 7818 3263 7852 3297
rect 7918 3263 7952 3297
rect 8018 3263 8052 3297
rect 8118 3263 8152 3297
rect 8218 3263 8252 3297
rect 8318 3263 8352 3297
rect 8618 3263 8652 3297
rect 8718 3263 8752 3297
rect 9218 3263 9252 3297
rect 9318 3263 9352 3297
rect 9418 3263 9452 3297
rect 9512 3263 9546 3297
rect 7124 3123 7158 3157
rect 7218 3123 7252 3157
rect 7618 3123 7652 3157
rect 7718 3123 7752 3157
rect 7918 3123 7952 3157
rect 8018 3123 8052 3157
rect 8112 3123 8146 3157
rect 6024 2983 6058 3017
rect 6118 2983 6152 3017
rect 6218 2983 6252 3017
rect 6418 2983 6452 3017
rect 6518 2983 6552 3017
rect 6618 2983 6652 3017
rect 6718 2983 6752 3017
rect 6818 2983 6852 3017
rect 6918 2983 6952 3017
rect 7018 2983 7052 3017
rect 7518 2983 7552 3017
rect 7618 2983 7652 3017
rect 7718 2983 7752 3017
rect 7818 2983 7852 3017
rect 7918 2983 7952 3017
rect 8012 2983 8046 3017
rect 5424 2843 5458 2877
rect 5518 2843 5552 2877
rect 5618 2843 5652 2877
rect 5918 2843 5952 2877
rect 6012 2843 6046 2877
rect 5424 2703 5458 2737
rect 5518 2703 5552 2737
rect 5618 2703 5652 2737
rect 5718 2703 5752 2737
rect 5918 2703 5952 2737
rect 6012 2703 6046 2737
rect 6124 2843 6158 2877
rect 6218 2843 6252 2877
rect 6718 2843 6752 2877
rect 6818 2843 6852 2877
rect 6912 2843 6946 2877
rect 6124 2703 6158 2737
rect 6212 2703 6246 2737
rect 4824 2563 4858 2597
rect 4918 2563 4952 2597
rect 5518 2563 5552 2597
rect 5618 2563 5652 2597
rect 5718 2563 5752 2597
rect 5818 2563 5852 2597
rect 5918 2563 5952 2597
rect 6118 2563 6152 2597
rect 6212 2563 6246 2597
rect 6324 2703 6358 2737
rect 6418 2703 6452 2737
rect 6512 2703 6546 2737
rect 7024 2843 7058 2877
rect 7118 2843 7152 2877
rect 7218 2843 7252 2877
rect 7312 2843 7346 2877
rect 7424 2843 7458 2877
rect 7518 2843 7552 2877
rect 7618 2843 7652 2877
rect 7718 2843 7752 2877
rect 7818 2843 7852 2877
rect 7912 2843 7946 2877
rect 8224 3123 8258 3157
rect 8318 3123 8352 3157
rect 8418 3123 8452 3157
rect 8718 3123 8752 3157
rect 8812 3123 8846 3157
rect 8124 2983 8158 3017
rect 8218 2983 8252 3017
rect 8318 2983 8352 3017
rect 8618 2983 8652 3017
rect 8718 2983 8752 3017
rect 8812 2983 8846 3017
rect 8024 2843 8058 2877
rect 8118 2843 8152 2877
rect 8218 2843 8252 2877
rect 8618 2843 8652 2877
rect 8712 2843 8746 2877
rect 6624 2703 6658 2737
rect 6718 2703 6752 2737
rect 6818 2703 6852 2737
rect 6918 2703 6952 2737
rect 7118 2703 7152 2737
rect 7218 2703 7252 2737
rect 7518 2703 7552 2737
rect 7618 2703 7652 2737
rect 8018 2703 8052 2737
rect 8118 2703 8152 2737
rect 8212 2703 8246 2737
rect 6324 2563 6358 2597
rect 6418 2563 6452 2597
rect 6618 2563 6652 2597
rect 6712 2563 6746 2597
rect 6824 2563 6858 2597
rect 6918 2563 6952 2597
rect 7118 2563 7152 2597
rect 7218 2563 7252 2597
rect 7418 2563 7452 2597
rect 7518 2563 7552 2597
rect 8018 2563 8052 2597
rect 8118 2563 8152 2597
rect 8212 2563 8246 2597
rect 2724 2333 2758 2367
rect 2818 2333 2852 2367
rect 2918 2333 2952 2367
rect 3118 2333 3152 2367
rect 3218 2333 3252 2367
rect 3618 2333 3652 2367
rect 3718 2333 3752 2367
rect 4018 2333 4052 2367
rect 4118 2333 4152 2367
rect 4218 2333 4252 2367
rect 4318 2333 4352 2367
rect 4418 2333 4452 2367
rect 4918 2333 4952 2367
rect 5018 2333 5052 2367
rect 5518 2333 5552 2367
rect 5618 2333 5652 2367
rect 5718 2333 5752 2367
rect 5818 2333 5852 2367
rect 5918 2333 5952 2367
rect 6418 2333 6452 2367
rect 6518 2333 6552 2367
rect 6618 2333 6652 2367
rect 6818 2333 6852 2367
rect 6912 2333 6946 2367
rect 2724 2193 2758 2227
rect 2812 2193 2846 2227
rect 1524 2053 1558 2087
rect 1618 2053 1652 2087
rect 1918 2053 1952 2087
rect 2018 2053 2052 2087
rect 2118 2053 2152 2087
rect 2618 2053 2652 2087
rect 2712 2053 2746 2087
rect 1024 1913 1058 1947
rect 1118 1913 1152 1947
rect 1418 1913 1452 1947
rect 1512 1913 1546 1947
rect 2924 2193 2958 2227
rect 3012 2193 3046 2227
rect 2824 2053 2858 2087
rect 2912 2053 2946 2087
rect 3124 2193 3158 2227
rect 3218 2193 3252 2227
rect 3312 2193 3346 2227
rect 3424 2193 3458 2227
rect 3518 2193 3552 2227
rect 3612 2193 3646 2227
rect 3024 2053 3058 2087
rect 3118 2053 3152 2087
rect 3218 2053 3252 2087
rect 3418 2053 3452 2087
rect 3512 2053 3546 2087
rect 3724 2193 3758 2227
rect 3812 2193 3846 2227
rect 3924 2193 3958 2227
rect 4018 2193 4052 2227
rect 4118 2193 4152 2227
rect 4218 2193 4252 2227
rect 4312 2193 4346 2227
rect 4424 2193 4458 2227
rect 4518 2193 4552 2227
rect 4918 2193 4952 2227
rect 5018 2193 5052 2227
rect 5118 2193 5152 2227
rect 5818 2193 5852 2227
rect 5918 2193 5952 2227
rect 6018 2193 6052 2227
rect 6112 2193 6146 2227
rect 3624 2053 3658 2087
rect 3718 2053 3752 2087
rect 4018 2053 4052 2087
rect 4118 2053 4152 2087
rect 4318 2053 4352 2087
rect 4418 2053 4452 2087
rect 4518 2053 4552 2087
rect 4612 2053 4646 2087
rect 1624 1913 1658 1947
rect 1718 1913 1752 1947
rect 1818 1913 1852 1947
rect 1918 1913 1952 1947
rect 2018 1913 2052 1947
rect 2118 1913 2152 1947
rect 2218 1913 2252 1947
rect 2518 1913 2552 1947
rect 2618 1913 2652 1947
rect 2818 1913 2852 1947
rect 2918 1913 2952 1947
rect 3218 1913 3252 1947
rect 3318 1913 3352 1947
rect 3518 1913 3552 1947
rect 3612 1913 3646 1947
rect 118 1773 152 1807
rect 218 1773 252 1807
rect 318 1773 352 1807
rect 718 1773 752 1807
rect 818 1773 852 1807
rect 918 1773 952 1807
rect 1018 1773 1052 1807
rect 1118 1773 1152 1807
rect 1218 1773 1252 1807
rect 1318 1773 1352 1807
rect 1418 1773 1452 1807
rect 1518 1773 1552 1807
rect 1618 1773 1652 1807
rect 2118 1773 2152 1807
rect 2218 1773 2252 1807
rect 2318 1773 2352 1807
rect 2418 1773 2452 1807
rect 2718 1773 2752 1807
rect 2818 1773 2852 1807
rect 3018 1773 3052 1807
rect 3112 1773 3146 1807
rect 118 1633 152 1667
rect 218 1633 252 1667
rect 518 1633 552 1667
rect 612 1633 646 1667
rect 118 1493 152 1527
rect 218 1493 252 1527
rect 318 1493 352 1527
rect 412 1493 446 1527
rect 724 1633 758 1667
rect 818 1633 852 1667
rect 918 1633 952 1667
rect 1012 1633 1046 1667
rect 1124 1633 1158 1667
rect 1212 1633 1246 1667
rect 1324 1633 1358 1667
rect 1418 1633 1452 1667
rect 1512 1633 1546 1667
rect 1624 1633 1658 1667
rect 1718 1633 1752 1667
rect 1818 1633 1852 1667
rect 1918 1633 1952 1667
rect 2018 1633 2052 1667
rect 2118 1633 2152 1667
rect 2218 1633 2252 1667
rect 2418 1633 2452 1667
rect 2518 1633 2552 1667
rect 2612 1633 2646 1667
rect 524 1493 558 1527
rect 618 1493 652 1527
rect 718 1493 752 1527
rect 918 1493 952 1527
rect 1018 1493 1052 1527
rect 1518 1493 1552 1527
rect 1618 1493 1652 1527
rect 1718 1493 1752 1527
rect 1918 1493 1952 1527
rect 2018 1493 2052 1527
rect 2118 1493 2152 1527
rect 2318 1493 2352 1527
rect 2418 1493 2452 1527
rect 2512 1493 2546 1527
rect 518 1353 552 1387
rect 618 1353 652 1387
rect 718 1353 752 1387
rect 812 1353 846 1387
rect 3224 1773 3258 1807
rect 3312 1773 3346 1807
rect 3724 1913 3758 1947
rect 3818 1913 3852 1947
rect 4118 1913 4152 1947
rect 4212 1913 4246 1947
rect 3424 1773 3458 1807
rect 3518 1773 3552 1807
rect 3618 1773 3652 1807
rect 3818 1773 3852 1807
rect 3912 1773 3946 1807
rect 2724 1633 2758 1667
rect 2818 1633 2852 1667
rect 2918 1633 2952 1667
rect 3118 1633 3152 1667
rect 3218 1633 3252 1667
rect 3418 1633 3452 1667
rect 3518 1633 3552 1667
rect 3618 1633 3652 1667
rect 3712 1633 3746 1667
rect 2624 1493 2658 1527
rect 2718 1493 2752 1527
rect 2918 1493 2952 1527
rect 3018 1493 3052 1527
rect 3112 1493 3146 1527
rect 924 1353 958 1387
rect 1018 1353 1052 1387
rect 1118 1353 1152 1387
rect 1318 1353 1352 1387
rect 1418 1353 1452 1387
rect 1518 1353 1552 1387
rect 1818 1353 1852 1387
rect 1918 1353 1952 1387
rect 2118 1353 2152 1387
rect 2218 1353 2252 1387
rect 2318 1353 2352 1387
rect 2718 1353 2752 1387
rect 2812 1353 2846 1387
rect 118 1123 152 1157
rect 218 1123 252 1157
rect 1118 1123 1152 1157
rect 1218 1123 1252 1157
rect 1318 1123 1352 1157
rect 1618 1123 1652 1157
rect 1712 1123 1746 1157
rect 24 983 58 1017
rect 112 983 146 1017
rect 24 843 58 877
rect 112 843 146 877
rect 224 983 258 1017
rect 318 983 352 1017
rect 418 983 452 1017
rect 518 983 552 1017
rect 612 983 646 1017
rect 724 983 758 1017
rect 818 983 852 1017
rect 1018 983 1052 1017
rect 1118 983 1152 1017
rect 1212 983 1246 1017
rect 1824 1123 1858 1157
rect 1918 1123 1952 1157
rect 2012 1123 2046 1157
rect 3224 1493 3258 1527
rect 3318 1493 3352 1527
rect 3418 1493 3452 1527
rect 3512 1493 3546 1527
rect 3824 1633 3858 1667
rect 3912 1633 3946 1667
rect 4024 1773 4058 1807
rect 4112 1773 4146 1807
rect 4024 1633 4058 1667
rect 4112 1633 4146 1667
rect 3624 1493 3658 1527
rect 3718 1493 3752 1527
rect 3818 1493 3852 1527
rect 3918 1493 3952 1527
rect 4012 1493 4046 1527
rect 4324 1913 4358 1947
rect 4412 1913 4446 1947
rect 4524 1913 4558 1947
rect 4612 1913 4646 1947
rect 4724 2053 4758 2087
rect 4818 2053 4852 2087
rect 4912 2053 4946 2087
rect 5024 2053 5058 2087
rect 5118 2053 5152 2087
rect 5618 2053 5652 2087
rect 5712 2053 5746 2087
rect 4724 1913 4758 1947
rect 4818 1913 4852 1947
rect 5018 1913 5052 1947
rect 5112 1913 5146 1947
rect 4224 1773 4258 1807
rect 4318 1773 4352 1807
rect 4718 1773 4752 1807
rect 4812 1773 4846 1807
rect 4224 1633 4258 1667
rect 4318 1633 4352 1667
rect 4412 1633 4446 1667
rect 5224 1913 5258 1947
rect 5318 1913 5352 1947
rect 5418 1913 5452 1947
rect 5518 1913 5552 1947
rect 5618 1913 5652 1947
rect 5712 1913 5746 1947
rect 6224 2193 6258 2227
rect 6318 2193 6352 2227
rect 6412 2193 6446 2227
rect 6524 2193 6558 2227
rect 6618 2193 6652 2227
rect 6712 2193 6746 2227
rect 5824 2053 5858 2087
rect 5918 2053 5952 2087
rect 6018 2053 6052 2087
rect 6118 2053 6152 2087
rect 6518 2053 6552 2087
rect 6612 2053 6646 2087
rect 6824 2193 6858 2227
rect 6912 2193 6946 2227
rect 6724 2053 6758 2087
rect 6812 2053 6846 2087
rect 5824 1913 5858 1947
rect 5918 1913 5952 1947
rect 6218 1913 6252 1947
rect 6318 1913 6352 1947
rect 6418 1913 6452 1947
rect 6518 1913 6552 1947
rect 6618 1913 6652 1947
rect 6712 1913 6746 1947
rect 4924 1773 4958 1807
rect 5018 1773 5052 1807
rect 5118 1773 5152 1807
rect 5218 1773 5252 1807
rect 5318 1773 5352 1807
rect 5418 1773 5452 1807
rect 5518 1773 5552 1807
rect 6218 1773 6252 1807
rect 6312 1773 6346 1807
rect 4524 1633 4558 1667
rect 4618 1633 4652 1667
rect 4718 1633 4752 1667
rect 4818 1633 4852 1667
rect 4912 1633 4946 1667
rect 4124 1493 4158 1527
rect 4218 1493 4252 1527
rect 4318 1493 4352 1527
rect 4418 1493 4452 1527
rect 4618 1493 4652 1527
rect 4718 1493 4752 1527
rect 4812 1493 4846 1527
rect 2924 1353 2958 1387
rect 3018 1353 3052 1387
rect 3218 1353 3252 1387
rect 3318 1353 3352 1387
rect 3418 1353 3452 1387
rect 3518 1353 3552 1387
rect 3818 1353 3852 1387
rect 3918 1353 3952 1387
rect 4018 1353 4052 1387
rect 4118 1353 4152 1387
rect 4318 1353 4352 1387
rect 4418 1353 4452 1387
rect 4518 1353 4552 1387
rect 4612 1353 4646 1387
rect 2124 1123 2158 1157
rect 2218 1123 2252 1157
rect 2918 1123 2952 1157
rect 3012 1123 3046 1157
rect 1324 983 1358 1017
rect 1418 983 1452 1017
rect 1618 983 1652 1017
rect 1718 983 1752 1017
rect 2018 983 2052 1017
rect 2118 983 2152 1017
rect 2218 983 2252 1017
rect 2318 983 2352 1017
rect 2418 983 2452 1017
rect 2518 983 2552 1017
rect 2612 983 2646 1017
rect 2724 983 2758 1017
rect 2812 983 2846 1017
rect 3124 1123 3158 1157
rect 3212 1123 3246 1157
rect 2924 983 2958 1017
rect 3018 983 3052 1017
rect 3112 983 3146 1017
rect 224 843 258 877
rect 318 843 352 877
rect 418 843 452 877
rect 518 843 552 877
rect 618 843 652 877
rect 718 843 752 877
rect 918 843 952 877
rect 1018 843 1052 877
rect 1118 843 1152 877
rect 1218 843 1252 877
rect 1618 843 1652 877
rect 1718 843 1752 877
rect 1918 843 1952 877
rect 2018 843 2052 877
rect 2118 843 2152 877
rect 2418 843 2452 877
rect 2518 843 2552 877
rect 2718 843 2752 877
rect 2818 843 2852 877
rect 2912 843 2946 877
rect 118 703 152 737
rect 218 703 252 737
rect 418 703 452 737
rect 512 703 546 737
rect 624 703 658 737
rect 712 703 746 737
rect 418 563 452 597
rect 518 563 552 597
rect 618 563 652 597
rect 712 563 746 597
rect 118 423 152 457
rect 218 423 252 457
rect 312 423 346 457
rect 824 703 858 737
rect 918 703 952 737
rect 1118 703 1152 737
rect 1212 703 1246 737
rect 824 563 858 597
rect 918 563 952 597
rect 1118 563 1152 597
rect 1212 563 1246 597
rect 424 423 458 457
rect 518 423 552 457
rect 918 423 952 457
rect 1018 423 1052 457
rect 1112 423 1146 457
rect 1324 703 1358 737
rect 1412 703 1446 737
rect 1524 703 1558 737
rect 1618 703 1652 737
rect 1818 703 1852 737
rect 1918 703 1952 737
rect 2012 703 2046 737
rect 2124 703 2158 737
rect 2218 703 2252 737
rect 2318 703 2352 737
rect 2412 703 2446 737
rect 1324 563 1358 597
rect 1418 563 1452 597
rect 1518 563 1552 597
rect 1718 563 1752 597
rect 1818 563 1852 597
rect 1918 563 1952 597
rect 2018 563 2052 597
rect 2112 563 2146 597
rect 1224 423 1258 457
rect 1318 423 1352 457
rect 1418 423 1452 457
rect 1618 423 1652 457
rect 1718 423 1752 457
rect 1812 423 1846 457
rect 118 283 152 317
rect 218 283 252 317
rect 818 283 852 317
rect 918 283 952 317
rect 1018 283 1052 317
rect 1218 283 1252 317
rect 1318 283 1352 317
rect 1618 283 1652 317
rect 1712 283 1746 317
rect 24 143 58 177
rect 118 143 152 177
rect 218 143 252 177
rect 318 143 352 177
rect 418 143 452 177
rect 518 143 552 177
rect 618 143 652 177
rect 718 143 752 177
rect 1218 143 1252 177
rect 1318 143 1352 177
rect 1418 143 1452 177
rect 1518 143 1552 177
rect 1612 143 1646 177
rect 2524 703 2558 737
rect 2618 703 2652 737
rect 2718 703 2752 737
rect 2812 703 2846 737
rect 2224 563 2258 597
rect 2318 563 2352 597
rect 2418 563 2452 597
rect 2618 563 2652 597
rect 2712 563 2746 597
rect 1924 423 1958 457
rect 2018 423 2052 457
rect 2218 423 2252 457
rect 2312 423 2346 457
rect 2424 423 2458 457
rect 2518 423 2552 457
rect 2612 423 2646 457
rect 3324 1123 3358 1157
rect 3418 1123 3452 1157
rect 3618 1123 3652 1157
rect 3712 1123 3746 1157
rect 3224 983 3258 1017
rect 3312 983 3346 1017
rect 3424 983 3458 1017
rect 3518 983 3552 1017
rect 3612 983 3646 1017
rect 3824 1123 3858 1157
rect 3918 1123 3952 1157
rect 4018 1123 4052 1157
rect 4318 1123 4352 1157
rect 4412 1123 4446 1157
rect 3724 983 3758 1017
rect 3812 983 3846 1017
rect 3024 843 3058 877
rect 3118 843 3152 877
rect 3318 843 3352 877
rect 3418 843 3452 877
rect 3518 843 3552 877
rect 3618 843 3652 877
rect 3718 843 3752 877
rect 3812 843 3846 877
rect 2924 703 2958 737
rect 3012 703 3046 737
rect 3124 703 3158 737
rect 3218 703 3252 737
rect 3312 703 3346 737
rect 3424 703 3458 737
rect 3518 703 3552 737
rect 3612 703 3646 737
rect 4724 1353 4758 1387
rect 4812 1353 4846 1387
rect 4524 1123 4558 1157
rect 4612 1123 4646 1157
rect 5024 1633 5058 1667
rect 5118 1633 5152 1667
rect 5212 1633 5246 1667
rect 5324 1633 5358 1667
rect 5418 1633 5452 1667
rect 5518 1633 5552 1667
rect 5612 1633 5646 1667
rect 5724 1633 5758 1667
rect 5818 1633 5852 1667
rect 5912 1633 5946 1667
rect 4924 1493 4958 1527
rect 5018 1493 5052 1527
rect 5118 1493 5152 1527
rect 5218 1493 5252 1527
rect 5318 1493 5352 1527
rect 5418 1493 5452 1527
rect 5518 1493 5552 1527
rect 5718 1493 5752 1527
rect 5812 1493 5846 1527
rect 4924 1353 4958 1387
rect 5018 1353 5052 1387
rect 5112 1353 5146 1387
rect 6024 1633 6058 1667
rect 6112 1633 6146 1667
rect 5924 1493 5958 1527
rect 6012 1493 6046 1527
rect 7024 2333 7058 2367
rect 7118 2333 7152 2367
rect 7212 2333 7246 2367
rect 8324 2703 8358 2737
rect 8418 2703 8452 2737
rect 8518 2703 8552 2737
rect 8618 2703 8652 2737
rect 8712 2703 8746 2737
rect 8324 2563 8358 2597
rect 8412 2563 8446 2597
rect 8524 2563 8558 2597
rect 8618 2563 8652 2597
rect 8712 2563 8746 2597
rect 7324 2333 7358 2367
rect 7418 2333 7452 2367
rect 7718 2333 7752 2367
rect 7818 2333 7852 2367
rect 8418 2333 8452 2367
rect 8512 2333 8546 2367
rect 7024 2193 7058 2227
rect 7118 2193 7152 2227
rect 7418 2193 7452 2227
rect 7512 2193 7546 2227
rect 7624 2193 7658 2227
rect 7712 2193 7746 2227
rect 10124 3543 10158 3577
rect 10218 3543 10252 3577
rect 10518 3543 10552 3577
rect 10612 3543 10646 3577
rect 11224 3773 11258 3807
rect 11318 3773 11352 3807
rect 11418 3773 11452 3807
rect 11512 3773 11546 3807
rect 11624 3773 11658 3807
rect 11718 3773 11752 3807
rect 11818 3773 11852 3807
rect 11918 3773 11952 3807
rect 12018 3773 12052 3807
rect 12112 3773 12146 3807
rect 10724 3543 10758 3577
rect 10818 3543 10852 3577
rect 10918 3543 10952 3577
rect 11318 3543 11352 3577
rect 11412 3543 11446 3577
rect 9824 3403 9858 3437
rect 9918 3403 9952 3437
rect 10018 3403 10052 3437
rect 10318 3403 10352 3437
rect 10418 3403 10452 3437
rect 10918 3403 10952 3437
rect 11018 3403 11052 3437
rect 11318 3403 11352 3437
rect 11412 3403 11446 3437
rect 9624 3263 9658 3297
rect 9718 3263 9752 3297
rect 9818 3263 9852 3297
rect 10118 3263 10152 3297
rect 10218 3263 10252 3297
rect 10312 3263 10346 3297
rect 8924 3123 8958 3157
rect 9018 3123 9052 3157
rect 9118 3123 9152 3157
rect 9218 3123 9252 3157
rect 9418 3123 9452 3157
rect 9518 3123 9552 3157
rect 9618 3123 9652 3157
rect 9718 3123 9752 3157
rect 9818 3123 9852 3157
rect 9912 3123 9946 3157
rect 8924 2983 8958 3017
rect 9018 2983 9052 3017
rect 9112 2983 9146 3017
rect 9224 2983 9258 3017
rect 9318 2983 9352 3017
rect 9412 2983 9446 3017
rect 10024 3123 10058 3157
rect 10112 3123 10146 3157
rect 10224 3123 10258 3157
rect 10312 3123 10346 3157
rect 10424 3263 10458 3297
rect 10512 3263 10546 3297
rect 12224 3773 12258 3807
rect 12318 3773 12352 3807
rect 12418 3773 12452 3807
rect 12518 3773 12552 3807
rect 12924 3788 12958 3822
rect 13018 3773 13052 3807
rect 13112 3758 13146 3792
rect 13228 3773 13262 3807
rect 13328 3773 13362 3807
rect 13428 3773 13462 3807
rect 13528 3773 13562 3807
rect 13628 3773 13662 3807
rect 11524 3543 11558 3577
rect 11618 3543 11652 3577
rect 11718 3543 11752 3577
rect 12018 3543 12052 3577
rect 12118 3543 12152 3577
rect 12218 3543 12252 3577
rect 12518 3543 12552 3577
rect 12618 3543 12652 3577
rect 12924 3558 12958 3592
rect 13018 3543 13052 3577
rect 13112 3528 13146 3562
rect 13228 3543 13262 3577
rect 13328 3543 13362 3577
rect 13428 3543 13462 3577
rect 13528 3543 13562 3577
rect 13628 3543 13662 3577
rect 11524 3403 11558 3437
rect 11618 3403 11652 3437
rect 11718 3403 11752 3437
rect 11918 3403 11952 3437
rect 12018 3403 12052 3437
rect 12112 3403 12146 3437
rect 12224 3403 12258 3437
rect 12318 3403 12352 3437
rect 12618 3403 12652 3437
rect 12718 3403 12752 3437
rect 12812 3403 12846 3437
rect 12924 3418 12958 3452
rect 13018 3403 13052 3437
rect 13112 3388 13146 3422
rect 13228 3403 13262 3437
rect 13328 3403 13362 3437
rect 13428 3403 13462 3437
rect 13528 3403 13562 3437
rect 13628 3403 13662 3437
rect 10624 3263 10658 3297
rect 10718 3263 10752 3297
rect 10818 3263 10852 3297
rect 10918 3263 10952 3297
rect 11018 3263 11052 3297
rect 11118 3263 11152 3297
rect 11218 3263 11252 3297
rect 11318 3263 11352 3297
rect 11418 3263 11452 3297
rect 11518 3263 11552 3297
rect 11618 3263 11652 3297
rect 11718 3263 11752 3297
rect 11818 3263 11852 3297
rect 12318 3263 12352 3297
rect 12412 3263 12446 3297
rect 10424 3123 10458 3157
rect 10518 3123 10552 3157
rect 10718 3123 10752 3157
rect 10812 3123 10846 3157
rect 10924 3123 10958 3157
rect 11018 3123 11052 3157
rect 11118 3123 11152 3157
rect 11418 3123 11452 3157
rect 11512 3123 11546 3157
rect 9524 2983 9558 3017
rect 9618 2983 9652 3017
rect 9918 2983 9952 3017
rect 10018 2983 10052 3017
rect 10118 2983 10152 3017
rect 10418 2983 10452 3017
rect 10518 2983 10552 3017
rect 10618 2983 10652 3017
rect 11018 2983 11052 3017
rect 11118 2983 11152 3017
rect 11318 2983 11352 3017
rect 11418 2983 11452 3017
rect 11512 2983 11546 3017
rect 8824 2843 8858 2877
rect 8918 2843 8952 2877
rect 9018 2843 9052 2877
rect 9118 2843 9152 2877
rect 9318 2843 9352 2877
rect 9418 2843 9452 2877
rect 9818 2843 9852 2877
rect 9918 2843 9952 2877
rect 10118 2843 10152 2877
rect 10218 2843 10252 2877
rect 10318 2843 10352 2877
rect 10418 2843 10452 2877
rect 10512 2843 10546 2877
rect 8824 2703 8858 2737
rect 8912 2703 8946 2737
rect 9024 2703 9058 2737
rect 9112 2703 9146 2737
rect 8824 2563 8858 2597
rect 8918 2563 8952 2597
rect 9012 2563 9046 2597
rect 9224 2703 9258 2737
rect 9312 2703 9346 2737
rect 9124 2563 9158 2597
rect 9212 2563 9246 2597
rect 9424 2703 9458 2737
rect 9512 2703 9546 2737
rect 9324 2563 9358 2597
rect 9418 2563 9452 2597
rect 9512 2563 9546 2597
rect 9624 2703 9658 2737
rect 9718 2703 9752 2737
rect 9818 2703 9852 2737
rect 9912 2703 9946 2737
rect 9624 2563 9658 2597
rect 9718 2563 9752 2597
rect 9818 2563 9852 2597
rect 9912 2563 9946 2597
rect 8624 2333 8658 2367
rect 8718 2333 8752 2367
rect 8918 2333 8952 2367
rect 9018 2333 9052 2367
rect 9118 2333 9152 2367
rect 9518 2333 9552 2367
rect 9612 2333 9646 2367
rect 7824 2193 7858 2227
rect 7918 2193 7952 2227
rect 8218 2193 8252 2227
rect 8318 2193 8352 2227
rect 8518 2193 8552 2227
rect 8618 2193 8652 2227
rect 8718 2193 8752 2227
rect 8812 2193 8846 2227
rect 6924 2053 6958 2087
rect 7018 2053 7052 2087
rect 7118 2053 7152 2087
rect 7418 2053 7452 2087
rect 7518 2053 7552 2087
rect 8018 2053 8052 2087
rect 8112 2053 8146 2087
rect 6824 1913 6858 1947
rect 6912 1913 6946 1947
rect 8224 2053 8258 2087
rect 8312 2053 8346 2087
rect 8424 2053 8458 2087
rect 8518 2053 8552 2087
rect 8618 2053 8652 2087
rect 8712 2053 8746 2087
rect 8924 2193 8958 2227
rect 9012 2193 9046 2227
rect 8824 2053 8858 2087
rect 8912 2053 8946 2087
rect 9124 2193 9158 2227
rect 9212 2193 9246 2227
rect 9024 2053 9058 2087
rect 9118 2053 9152 2087
rect 9212 2053 9246 2087
rect 9324 2193 9358 2227
rect 9418 2193 9452 2227
rect 9512 2193 9546 2227
rect 10024 2703 10058 2737
rect 10118 2703 10152 2737
rect 10218 2703 10252 2737
rect 10318 2703 10352 2737
rect 10412 2703 10446 2737
rect 10624 2843 10658 2877
rect 10718 2843 10752 2877
rect 10918 2843 10952 2877
rect 11018 2843 11052 2877
rect 11118 2843 11152 2877
rect 11218 2843 11252 2877
rect 11312 2843 11346 2877
rect 10524 2703 10558 2737
rect 10612 2703 10646 2737
rect 12524 3263 12558 3297
rect 12618 3263 12652 3297
rect 12718 3263 12752 3297
rect 12924 3278 12958 3312
rect 13018 3263 13052 3297
rect 13112 3248 13146 3282
rect 13228 3263 13262 3297
rect 13328 3263 13362 3297
rect 13428 3263 13462 3297
rect 13528 3263 13562 3297
rect 13628 3263 13662 3297
rect 11624 3123 11658 3157
rect 11718 3123 11752 3157
rect 11818 3123 11852 3157
rect 12018 3123 12052 3157
rect 12118 3123 12152 3157
rect 12318 3123 12352 3157
rect 12418 3123 12452 3157
rect 12518 3123 12552 3157
rect 12618 3123 12652 3157
rect 12718 3123 12752 3157
rect 12924 3138 12958 3172
rect 13018 3123 13052 3157
rect 13112 3108 13146 3142
rect 13228 3123 13262 3157
rect 13328 3123 13362 3157
rect 13428 3123 13462 3157
rect 13528 3123 13562 3157
rect 13628 3123 13662 3157
rect 11624 2983 11658 3017
rect 11718 2983 11752 3017
rect 11818 2983 11852 3017
rect 11918 2983 11952 3017
rect 12018 2983 12052 3017
rect 12218 2983 12252 3017
rect 12318 2983 12352 3017
rect 12718 2983 12752 3017
rect 12812 2983 12846 3017
rect 12924 2998 12958 3032
rect 13018 2983 13052 3017
rect 13112 2968 13146 3002
rect 13228 2983 13262 3017
rect 13328 2983 13362 3017
rect 13428 2983 13462 3017
rect 13528 2983 13562 3017
rect 13628 2983 13662 3017
rect 11424 2843 11458 2877
rect 11518 2843 11552 2877
rect 11618 2843 11652 2877
rect 11718 2843 11752 2877
rect 11812 2843 11846 2877
rect 10724 2703 10758 2737
rect 10818 2703 10852 2737
rect 10918 2703 10952 2737
rect 11518 2703 11552 2737
rect 11612 2703 11646 2737
rect 10024 2563 10058 2597
rect 10118 2563 10152 2597
rect 10218 2563 10252 2597
rect 10618 2563 10652 2597
rect 10718 2563 10752 2597
rect 10818 2563 10852 2597
rect 10912 2563 10946 2597
rect 11024 2563 11058 2597
rect 11112 2563 11146 2597
rect 11224 2563 11258 2597
rect 11312 2563 11346 2597
rect 11424 2563 11458 2597
rect 11518 2563 11552 2597
rect 11612 2563 11646 2597
rect 11924 2843 11958 2877
rect 12018 2843 12052 2877
rect 12718 2843 12752 2877
rect 12812 2843 12846 2877
rect 12924 2858 12958 2892
rect 13018 2843 13052 2877
rect 13112 2828 13146 2862
rect 13228 2843 13262 2877
rect 13328 2843 13362 2877
rect 13428 2843 13462 2877
rect 13528 2843 13562 2877
rect 13628 2843 13662 2877
rect 11724 2703 11758 2737
rect 11818 2703 11852 2737
rect 11918 2703 11952 2737
rect 12218 2703 12252 2737
rect 12318 2703 12352 2737
rect 12418 2703 12452 2737
rect 12518 2703 12552 2737
rect 12618 2703 12652 2737
rect 12718 2703 12752 2737
rect 12924 2718 12958 2752
rect 13018 2703 13052 2737
rect 13112 2688 13146 2722
rect 13228 2703 13262 2737
rect 13328 2703 13362 2737
rect 13428 2703 13462 2737
rect 13528 2703 13562 2737
rect 13628 2703 13662 2737
rect 11724 2563 11758 2597
rect 11818 2563 11852 2597
rect 12218 2563 12252 2597
rect 12318 2563 12352 2597
rect 12418 2563 12452 2597
rect 12618 2563 12652 2597
rect 12718 2563 12752 2597
rect 12924 2578 12958 2612
rect 13018 2563 13052 2597
rect 13112 2548 13146 2582
rect 13228 2563 13262 2597
rect 13328 2563 13362 2597
rect 13428 2563 13462 2597
rect 13528 2563 13562 2597
rect 13628 2563 13662 2597
rect 9724 2333 9758 2367
rect 9818 2333 9852 2367
rect 10018 2333 10052 2367
rect 10118 2333 10152 2367
rect 10318 2333 10352 2367
rect 10418 2333 10452 2367
rect 10518 2333 10552 2367
rect 10618 2333 10652 2367
rect 10718 2333 10752 2367
rect 10818 2333 10852 2367
rect 10918 2333 10952 2367
rect 11118 2333 11152 2367
rect 11218 2333 11252 2367
rect 11318 2333 11352 2367
rect 11418 2333 11452 2367
rect 11618 2333 11652 2367
rect 11712 2333 11746 2367
rect 9624 2193 9658 2227
rect 9718 2193 9752 2227
rect 9818 2193 9852 2227
rect 10218 2193 10252 2227
rect 10318 2193 10352 2227
rect 10418 2193 10452 2227
rect 10512 2193 10546 2227
rect 11824 2333 11858 2367
rect 11912 2333 11946 2367
rect 12024 2333 12058 2367
rect 12118 2333 12152 2367
rect 12318 2333 12352 2367
rect 12418 2333 12452 2367
rect 12512 2333 12546 2367
rect 10624 2193 10658 2227
rect 10718 2193 10752 2227
rect 10818 2193 10852 2227
rect 10918 2193 10952 2227
rect 11318 2193 11352 2227
rect 11418 2193 11452 2227
rect 11518 2193 11552 2227
rect 11818 2193 11852 2227
rect 11918 2193 11952 2227
rect 12012 2193 12046 2227
rect 9324 2053 9358 2087
rect 9418 2053 9452 2087
rect 10118 2053 10152 2087
rect 10218 2053 10252 2087
rect 10318 2053 10352 2087
rect 10418 2053 10452 2087
rect 10618 2053 10652 2087
rect 10718 2053 10752 2087
rect 10918 2053 10952 2087
rect 11018 2053 11052 2087
rect 11118 2053 11152 2087
rect 11212 2053 11246 2087
rect 7024 1913 7058 1947
rect 7118 1913 7152 1947
rect 7218 1913 7252 1947
rect 7318 1913 7352 1947
rect 8218 1913 8252 1947
rect 8318 1913 8352 1947
rect 8418 1913 8452 1947
rect 9318 1913 9352 1947
rect 9418 1913 9452 1947
rect 9618 1913 9652 1947
rect 9718 1913 9752 1947
rect 9818 1913 9852 1947
rect 9918 1913 9952 1947
rect 10018 1913 10052 1947
rect 10318 1913 10352 1947
rect 10418 1913 10452 1947
rect 10618 1913 10652 1947
rect 10718 1913 10752 1947
rect 10818 1913 10852 1947
rect 10918 1913 10952 1947
rect 11012 1913 11046 1947
rect 6424 1773 6458 1807
rect 6518 1773 6552 1807
rect 6818 1773 6852 1807
rect 6918 1773 6952 1807
rect 7018 1773 7052 1807
rect 7112 1773 7146 1807
rect 6224 1633 6258 1667
rect 6318 1633 6352 1667
rect 6418 1633 6452 1667
rect 6512 1633 6546 1667
rect 6124 1493 6158 1527
rect 6218 1493 6252 1527
rect 6312 1493 6346 1527
rect 5224 1353 5258 1387
rect 5318 1353 5352 1387
rect 5618 1353 5652 1387
rect 5718 1353 5752 1387
rect 5818 1353 5852 1387
rect 6018 1353 6052 1387
rect 6118 1353 6152 1387
rect 6212 1353 6246 1387
rect 4724 1123 4758 1157
rect 4818 1123 4852 1157
rect 5118 1123 5152 1157
rect 5218 1123 5252 1157
rect 5318 1123 5352 1157
rect 5412 1123 5446 1157
rect 3924 983 3958 1017
rect 4018 983 4052 1017
rect 4118 983 4152 1017
rect 4218 983 4252 1017
rect 4318 983 4352 1017
rect 4418 983 4452 1017
rect 4718 983 4752 1017
rect 4812 983 4846 1017
rect 4924 983 4958 1017
rect 5018 983 5052 1017
rect 5218 983 5252 1017
rect 5312 983 5346 1017
rect 7224 1773 7258 1807
rect 7318 1773 7352 1807
rect 7412 1773 7446 1807
rect 7524 1773 7558 1807
rect 7618 1773 7652 1807
rect 7712 1773 7746 1807
rect 7824 1773 7858 1807
rect 7918 1773 7952 1807
rect 8012 1773 8046 1807
rect 8124 1773 8158 1807
rect 8218 1773 8252 1807
rect 8318 1773 8352 1807
rect 8418 1773 8452 1807
rect 8518 1773 8552 1807
rect 8612 1773 8646 1807
rect 8724 1773 8758 1807
rect 8818 1773 8852 1807
rect 8918 1773 8952 1807
rect 9318 1773 9352 1807
rect 9418 1773 9452 1807
rect 9518 1773 9552 1807
rect 9718 1773 9752 1807
rect 9812 1773 9846 1807
rect 6624 1633 6658 1667
rect 6718 1633 6752 1667
rect 6818 1633 6852 1667
rect 7018 1633 7052 1667
rect 7118 1633 7152 1667
rect 7618 1633 7652 1667
rect 7718 1633 7752 1667
rect 7918 1633 7952 1667
rect 8018 1633 8052 1667
rect 8218 1633 8252 1667
rect 8318 1633 8352 1667
rect 8418 1633 8452 1667
rect 8818 1633 8852 1667
rect 8918 1633 8952 1667
rect 9018 1633 9052 1667
rect 9418 1633 9452 1667
rect 9512 1633 9546 1667
rect 6424 1493 6458 1527
rect 6518 1493 6552 1527
rect 6618 1493 6652 1527
rect 7418 1493 7452 1527
rect 7518 1493 7552 1527
rect 7618 1493 7652 1527
rect 7712 1493 7746 1527
rect 6324 1353 6358 1387
rect 6412 1353 6446 1387
rect 6524 1353 6558 1387
rect 6618 1353 6652 1387
rect 6712 1353 6746 1387
rect 6824 1353 6858 1387
rect 6912 1353 6946 1387
rect 5524 1123 5558 1157
rect 5618 1123 5652 1157
rect 5718 1123 5752 1157
rect 5818 1123 5852 1157
rect 6518 1123 6552 1157
rect 6618 1123 6652 1157
rect 6712 1123 6746 1157
rect 5424 983 5458 1017
rect 5518 983 5552 1017
rect 5618 983 5652 1017
rect 5718 983 5752 1017
rect 5818 983 5852 1017
rect 5918 983 5952 1017
rect 6118 983 6152 1017
rect 6218 983 6252 1017
rect 6318 983 6352 1017
rect 6412 983 6446 1017
rect 7824 1493 7858 1527
rect 7912 1493 7946 1527
rect 7024 1353 7058 1387
rect 7118 1353 7152 1387
rect 7218 1353 7252 1387
rect 7318 1353 7352 1387
rect 7418 1353 7452 1387
rect 7518 1353 7552 1387
rect 7818 1353 7852 1387
rect 7912 1353 7946 1387
rect 8024 1493 8058 1527
rect 8118 1493 8152 1527
rect 8418 1493 8452 1527
rect 8512 1493 8546 1527
rect 8624 1493 8658 1527
rect 8718 1493 8752 1527
rect 8918 1493 8952 1527
rect 9018 1493 9052 1527
rect 9118 1493 9152 1527
rect 9218 1493 9252 1527
rect 9312 1493 9346 1527
rect 8024 1353 8058 1387
rect 8118 1353 8152 1387
rect 8218 1353 8252 1387
rect 8318 1353 8352 1387
rect 8718 1353 8752 1387
rect 8818 1353 8852 1387
rect 8918 1353 8952 1387
rect 9118 1353 9152 1387
rect 9218 1353 9252 1387
rect 9312 1353 9346 1387
rect 9924 1773 9958 1807
rect 10012 1773 10046 1807
rect 10124 1773 10158 1807
rect 10212 1773 10246 1807
rect 10324 1773 10358 1807
rect 10412 1773 10446 1807
rect 10524 1773 10558 1807
rect 10618 1773 10652 1807
rect 10712 1773 10746 1807
rect 11124 1913 11158 1947
rect 11212 1913 11246 1947
rect 11324 2053 11358 2087
rect 11412 2053 11446 2087
rect 12124 2193 12158 2227
rect 12218 2193 12252 2227
rect 12312 2193 12346 2227
rect 12624 2333 12658 2367
rect 12718 2333 12752 2367
rect 12924 2348 12958 2382
rect 13018 2333 13052 2367
rect 13112 2318 13146 2352
rect 13228 2333 13262 2367
rect 13328 2333 13362 2367
rect 13428 2333 13462 2367
rect 13528 2333 13562 2367
rect 13628 2333 13662 2367
rect 12424 2193 12458 2227
rect 12518 2193 12552 2227
rect 12612 2193 12646 2227
rect 11524 2053 11558 2087
rect 11618 2053 11652 2087
rect 11718 2053 11752 2087
rect 11818 2053 11852 2087
rect 11918 2053 11952 2087
rect 12118 2053 12152 2087
rect 12218 2053 12252 2087
rect 12318 2053 12352 2087
rect 12518 2053 12552 2087
rect 12612 2053 12646 2087
rect 11324 1913 11358 1947
rect 11418 1913 11452 1947
rect 11918 1913 11952 1947
rect 12018 1913 12052 1947
rect 12118 1913 12152 1947
rect 12218 1913 12252 1947
rect 12318 1913 12352 1947
rect 12518 1913 12552 1947
rect 12612 1913 12646 1947
rect 10824 1773 10858 1807
rect 10918 1773 10952 1807
rect 11018 1773 11052 1807
rect 11118 1773 11152 1807
rect 11218 1773 11252 1807
rect 11418 1773 11452 1807
rect 11518 1773 11552 1807
rect 11612 1773 11646 1807
rect 9624 1633 9658 1667
rect 9718 1633 9752 1667
rect 9818 1633 9852 1667
rect 10018 1633 10052 1667
rect 10118 1633 10152 1667
rect 10218 1633 10252 1667
rect 10318 1633 10352 1667
rect 10418 1633 10452 1667
rect 10618 1633 10652 1667
rect 10718 1633 10752 1667
rect 10818 1633 10852 1667
rect 10912 1633 10946 1667
rect 9424 1493 9458 1527
rect 9518 1493 9552 1527
rect 9618 1493 9652 1527
rect 9818 1493 9852 1527
rect 9918 1493 9952 1527
rect 10118 1493 10152 1527
rect 10218 1493 10252 1527
rect 10518 1493 10552 1527
rect 10618 1493 10652 1527
rect 10718 1493 10752 1527
rect 10818 1493 10852 1527
rect 10912 1493 10946 1527
rect 9424 1353 9458 1387
rect 9518 1353 9552 1387
rect 9818 1353 9852 1387
rect 9918 1353 9952 1387
rect 10018 1353 10052 1387
rect 10118 1353 10152 1387
rect 10212 1353 10246 1387
rect 6824 1123 6858 1157
rect 6918 1123 6952 1157
rect 7318 1123 7352 1157
rect 7418 1123 7452 1157
rect 7718 1123 7752 1157
rect 7818 1123 7852 1157
rect 8018 1123 8052 1157
rect 8118 1123 8152 1157
rect 8318 1123 8352 1157
rect 8418 1123 8452 1157
rect 8518 1123 8552 1157
rect 8718 1123 8752 1157
rect 8818 1123 8852 1157
rect 8918 1123 8952 1157
rect 9218 1123 9252 1157
rect 9318 1123 9352 1157
rect 9518 1123 9552 1157
rect 9612 1123 9646 1157
rect 6524 983 6558 1017
rect 6618 983 6652 1017
rect 6718 983 6752 1017
rect 6818 983 6852 1017
rect 6912 983 6946 1017
rect 3924 843 3958 877
rect 4018 843 4052 877
rect 4118 843 4152 877
rect 4218 843 4252 877
rect 4318 843 4352 877
rect 4418 843 4452 877
rect 4718 843 4752 877
rect 4818 843 4852 877
rect 4918 843 4952 877
rect 5018 843 5052 877
rect 5118 843 5152 877
rect 5318 843 5352 877
rect 5418 843 5452 877
rect 5518 843 5552 877
rect 5618 843 5652 877
rect 5918 843 5952 877
rect 6018 843 6052 877
rect 6118 843 6152 877
rect 6218 843 6252 877
rect 6418 843 6452 877
rect 6518 843 6552 877
rect 6612 843 6646 877
rect 3724 703 3758 737
rect 3818 703 3852 737
rect 3918 703 3952 737
rect 4018 703 4052 737
rect 4418 703 4452 737
rect 4518 703 4552 737
rect 4612 703 4646 737
rect 2824 563 2858 597
rect 2918 563 2952 597
rect 3418 563 3452 597
rect 3518 563 3552 597
rect 3618 563 3652 597
rect 3718 563 3752 597
rect 3818 563 3852 597
rect 3912 563 3946 597
rect 4024 563 4058 597
rect 4112 563 4146 597
rect 4724 703 4758 737
rect 4818 703 4852 737
rect 5018 703 5052 737
rect 5112 703 5146 737
rect 4224 563 4258 597
rect 4318 563 4352 597
rect 4618 563 4652 597
rect 4718 563 4752 597
rect 4812 563 4846 597
rect 2724 423 2758 457
rect 2818 423 2852 457
rect 2918 423 2952 457
rect 3118 423 3152 457
rect 3218 423 3252 457
rect 3618 423 3652 457
rect 3718 423 3752 457
rect 3818 423 3852 457
rect 3918 423 3952 457
rect 4018 423 4052 457
rect 4318 423 4352 457
rect 4412 423 4446 457
rect 1824 283 1858 317
rect 1918 283 1952 317
rect 2318 283 2352 317
rect 2418 283 2452 317
rect 2718 283 2752 317
rect 2812 283 2846 317
rect 1724 143 1758 177
rect 1812 143 1846 177
rect 2924 283 2958 317
rect 3012 283 3046 317
rect 4924 563 4958 597
rect 5012 563 5046 597
rect 5224 703 5258 737
rect 5318 703 5352 737
rect 5618 703 5652 737
rect 5712 703 5746 737
rect 5124 563 5158 597
rect 5212 563 5246 597
rect 4524 423 4558 457
rect 4618 423 4652 457
rect 4718 423 4752 457
rect 4818 423 4852 457
rect 5018 423 5052 457
rect 5112 423 5146 457
rect 3124 283 3158 317
rect 3218 283 3252 317
rect 3318 283 3352 317
rect 3518 283 3552 317
rect 3618 283 3652 317
rect 3818 283 3852 317
rect 3918 283 3952 317
rect 4018 283 4052 317
rect 4118 283 4152 317
rect 4218 283 4252 317
rect 4318 283 4352 317
rect 4418 283 4452 317
rect 4512 283 4546 317
rect 4624 283 4658 317
rect 4718 283 4752 317
rect 4812 283 4846 317
rect 4924 283 4958 317
rect 5012 283 5046 317
rect 5824 703 5858 737
rect 5918 703 5952 737
rect 6118 703 6152 737
rect 6212 703 6246 737
rect 6324 703 6358 737
rect 6412 703 6446 737
rect 7024 983 7058 1017
rect 7112 983 7146 1017
rect 7224 983 7258 1017
rect 7312 983 7346 1017
rect 6724 843 6758 877
rect 6818 843 6852 877
rect 7018 843 7052 877
rect 7118 843 7152 877
rect 7218 843 7252 877
rect 7312 843 7346 877
rect 6524 703 6558 737
rect 6618 703 6652 737
rect 6918 703 6952 737
rect 7012 703 7046 737
rect 7424 983 7458 1017
rect 7518 983 7552 1017
rect 7618 983 7652 1017
rect 7718 983 7752 1017
rect 7818 983 7852 1017
rect 8218 983 8252 1017
rect 8318 983 8352 1017
rect 8418 983 8452 1017
rect 8518 983 8552 1017
rect 8612 983 8646 1017
rect 7424 843 7458 877
rect 7512 843 7546 877
rect 7624 843 7658 877
rect 7712 843 7746 877
rect 7824 843 7858 877
rect 7912 843 7946 877
rect 8024 843 8058 877
rect 8118 843 8152 877
rect 8318 843 8352 877
rect 8418 843 8452 877
rect 8518 843 8552 877
rect 8612 843 8646 877
rect 8724 983 8758 1017
rect 8812 983 8846 1017
rect 8724 843 8758 877
rect 8812 843 8846 877
rect 8924 983 8958 1017
rect 9018 983 9052 1017
rect 9118 983 9152 1017
rect 9418 983 9452 1017
rect 9512 983 9546 1017
rect 11724 1773 11758 1807
rect 11818 1773 11852 1807
rect 11912 1773 11946 1807
rect 11024 1633 11058 1667
rect 11118 1633 11152 1667
rect 11218 1633 11252 1667
rect 11618 1633 11652 1667
rect 11712 1633 11746 1667
rect 11024 1493 11058 1527
rect 11112 1493 11146 1527
rect 10324 1353 10358 1387
rect 10418 1353 10452 1387
rect 10918 1353 10952 1387
rect 11018 1353 11052 1387
rect 11112 1353 11146 1387
rect 12724 2193 12758 2227
rect 12812 2193 12846 2227
rect 12924 2208 12958 2242
rect 13018 2193 13052 2227
rect 13112 2178 13146 2212
rect 13228 2193 13262 2227
rect 13328 2193 13362 2227
rect 13428 2193 13462 2227
rect 13528 2193 13562 2227
rect 13628 2193 13662 2227
rect 12724 2053 12758 2087
rect 12812 2053 12846 2087
rect 12924 2068 12958 2102
rect 13018 2053 13052 2087
rect 13112 2038 13146 2072
rect 13228 2053 13262 2087
rect 13328 2053 13362 2087
rect 13428 2053 13462 2087
rect 13528 2053 13562 2087
rect 13628 2053 13662 2087
rect 12724 1913 12758 1947
rect 12812 1913 12846 1947
rect 12924 1928 12958 1962
rect 13018 1913 13052 1947
rect 13112 1898 13146 1932
rect 13228 1913 13262 1947
rect 13328 1913 13362 1947
rect 13428 1913 13462 1947
rect 13528 1913 13562 1947
rect 13628 1913 13662 1947
rect 12024 1773 12058 1807
rect 12118 1773 12152 1807
rect 12218 1773 12252 1807
rect 12618 1773 12652 1807
rect 12718 1773 12752 1807
rect 12812 1773 12846 1807
rect 12924 1788 12958 1822
rect 13018 1773 13052 1807
rect 13112 1758 13146 1792
rect 13228 1773 13262 1807
rect 13328 1773 13362 1807
rect 13428 1773 13462 1807
rect 13528 1773 13562 1807
rect 13628 1773 13662 1807
rect 11824 1633 11858 1667
rect 11918 1633 11952 1667
rect 12118 1633 12152 1667
rect 12218 1633 12252 1667
rect 12318 1633 12352 1667
rect 12418 1633 12452 1667
rect 12518 1633 12552 1667
rect 12618 1633 12652 1667
rect 12718 1633 12752 1667
rect 12924 1648 12958 1682
rect 13018 1633 13052 1667
rect 13112 1618 13146 1652
rect 13228 1633 13262 1667
rect 13328 1633 13362 1667
rect 13428 1633 13462 1667
rect 13528 1633 13562 1667
rect 13628 1633 13662 1667
rect 11224 1493 11258 1527
rect 11318 1493 11352 1527
rect 11518 1493 11552 1527
rect 11618 1493 11652 1527
rect 11918 1493 11952 1527
rect 12012 1493 12046 1527
rect 11224 1353 11258 1387
rect 11318 1353 11352 1387
rect 11518 1353 11552 1387
rect 11618 1353 11652 1387
rect 11712 1353 11746 1387
rect 9724 1123 9758 1157
rect 9818 1123 9852 1157
rect 9918 1123 9952 1157
rect 10018 1123 10052 1157
rect 10518 1123 10552 1157
rect 10618 1123 10652 1157
rect 10718 1123 10752 1157
rect 10918 1123 10952 1157
rect 11012 1123 11046 1157
rect 9624 983 9658 1017
rect 9718 983 9752 1017
rect 9818 983 9852 1017
rect 9912 983 9946 1017
rect 8924 843 8958 877
rect 9018 843 9052 877
rect 9118 843 9152 877
rect 9418 843 9452 877
rect 9518 843 9552 877
rect 9718 843 9752 877
rect 9818 843 9852 877
rect 9912 843 9946 877
rect 7124 703 7158 737
rect 7218 703 7252 737
rect 7318 703 7352 737
rect 7418 703 7452 737
rect 7518 703 7552 737
rect 7618 703 7652 737
rect 7718 703 7752 737
rect 7918 703 7952 737
rect 8018 703 8052 737
rect 8118 703 8152 737
rect 8218 703 8252 737
rect 8318 703 8352 737
rect 8418 703 8452 737
rect 8618 703 8652 737
rect 8718 703 8752 737
rect 8818 703 8852 737
rect 9018 703 9052 737
rect 9112 703 9146 737
rect 5324 563 5358 597
rect 5418 563 5452 597
rect 5518 563 5552 597
rect 5918 563 5952 597
rect 6018 563 6052 597
rect 6118 563 6152 597
rect 6318 563 6352 597
rect 6418 563 6452 597
rect 6718 563 6752 597
rect 6818 563 6852 597
rect 6918 563 6952 597
rect 7218 563 7252 597
rect 7318 563 7352 597
rect 7518 563 7552 597
rect 7618 563 7652 597
rect 7718 563 7752 597
rect 7818 563 7852 597
rect 8118 563 8152 597
rect 8218 563 8252 597
rect 8312 563 8346 597
rect 5224 423 5258 457
rect 5312 423 5346 457
rect 5424 423 5458 457
rect 5518 423 5552 457
rect 5618 423 5652 457
rect 5718 423 5752 457
rect 5818 423 5852 457
rect 6018 423 6052 457
rect 6112 423 6146 457
rect 5124 283 5158 317
rect 5218 283 5252 317
rect 5318 283 5352 317
rect 5718 283 5752 317
rect 5812 283 5846 317
rect 5924 283 5958 317
rect 6012 283 6046 317
rect 6224 423 6258 457
rect 6318 423 6352 457
rect 6412 423 6446 457
rect 6124 283 6158 317
rect 6212 283 6246 317
rect 6324 283 6358 317
rect 6412 283 6446 317
rect 6524 423 6558 457
rect 6618 423 6652 457
rect 6918 423 6952 457
rect 7018 423 7052 457
rect 7112 423 7146 457
rect 6524 283 6558 317
rect 6612 283 6646 317
rect 6724 283 6758 317
rect 6812 283 6846 317
rect 7224 423 7258 457
rect 7312 423 7346 457
rect 7424 423 7458 457
rect 7512 423 7546 457
rect 7624 423 7658 457
rect 7718 423 7752 457
rect 7818 423 7852 457
rect 8218 423 8252 457
rect 8312 423 8346 457
rect 6924 283 6958 317
rect 7018 283 7052 317
rect 7218 283 7252 317
rect 7318 283 7352 317
rect 7418 283 7452 317
rect 7718 283 7752 317
rect 7812 283 7846 317
rect 1924 143 1958 177
rect 2018 143 2052 177
rect 2218 143 2252 177
rect 2318 143 2352 177
rect 2518 143 2552 177
rect 2618 143 2652 177
rect 2918 143 2952 177
rect 3018 143 3052 177
rect 3318 143 3352 177
rect 3418 143 3452 177
rect 3718 143 3752 177
rect 3818 143 3852 177
rect 3918 143 3952 177
rect 4018 143 4052 177
rect 4118 143 4152 177
rect 4218 143 4252 177
rect 4318 143 4352 177
rect 4718 143 4752 177
rect 4818 143 4852 177
rect 4918 143 4952 177
rect 5018 143 5052 177
rect 5518 143 5552 177
rect 5618 143 5652 177
rect 5818 143 5852 177
rect 5918 143 5952 177
rect 6018 143 6052 177
rect 6118 143 6152 177
rect 6218 143 6252 177
rect 6318 143 6352 177
rect 6418 143 6452 177
rect 6918 143 6952 177
rect 7012 143 7046 177
rect 7924 283 7958 317
rect 8012 283 8046 317
rect 9224 703 9258 737
rect 9312 703 9346 737
rect 9424 703 9458 737
rect 9518 703 9552 737
rect 9612 703 9646 737
rect 9724 703 9758 737
rect 9812 703 9846 737
rect 10024 983 10058 1017
rect 10118 983 10152 1017
rect 10218 983 10252 1017
rect 10312 983 10346 1017
rect 11124 1123 11158 1157
rect 11212 1123 11246 1157
rect 11324 1123 11358 1157
rect 11412 1123 11446 1157
rect 10424 983 10458 1017
rect 10518 983 10552 1017
rect 10818 983 10852 1017
rect 10918 983 10952 1017
rect 11018 983 11052 1017
rect 11118 983 11152 1017
rect 11218 983 11252 1017
rect 11312 983 11346 1017
rect 10024 843 10058 877
rect 10118 843 10152 877
rect 10518 843 10552 877
rect 10618 843 10652 877
rect 10712 843 10746 877
rect 9924 703 9958 737
rect 10018 703 10052 737
rect 10112 703 10146 737
rect 10824 843 10858 877
rect 10912 843 10946 877
rect 10224 703 10258 737
rect 10318 703 10352 737
rect 10718 703 10752 737
rect 10818 703 10852 737
rect 10912 703 10946 737
rect 8424 563 8458 597
rect 8518 563 8552 597
rect 8718 563 8752 597
rect 8818 563 8852 597
rect 8918 563 8952 597
rect 9018 563 9052 597
rect 9218 563 9252 597
rect 9318 563 9352 597
rect 9518 563 9552 597
rect 9618 563 9652 597
rect 9918 563 9952 597
rect 10018 563 10052 597
rect 10118 563 10152 597
rect 10212 563 10246 597
rect 8424 423 8458 457
rect 8518 423 8552 457
rect 8718 423 8752 457
rect 8818 423 8852 457
rect 8918 423 8952 457
rect 9018 423 9052 457
rect 9118 423 9152 457
rect 9218 423 9252 457
rect 9418 423 9452 457
rect 9518 423 9552 457
rect 9618 423 9652 457
rect 9718 423 9752 457
rect 9818 423 9852 457
rect 9912 423 9946 457
rect 8124 283 8158 317
rect 8218 283 8252 317
rect 8318 283 8352 317
rect 8418 283 8452 317
rect 8518 283 8552 317
rect 8618 283 8652 317
rect 8712 283 8746 317
rect 8824 283 8858 317
rect 8918 283 8952 317
rect 9012 283 9046 317
rect 9124 283 9158 317
rect 9212 283 9246 317
rect 10024 423 10058 457
rect 10118 423 10152 457
rect 10212 423 10246 457
rect 9324 283 9358 317
rect 9418 283 9452 317
rect 9518 283 9552 317
rect 9618 283 9652 317
rect 10018 283 10052 317
rect 10112 283 10146 317
rect 10324 563 10358 597
rect 10412 563 10446 597
rect 12124 1493 12158 1527
rect 12218 1493 12252 1527
rect 12318 1493 12352 1527
rect 12412 1493 12446 1527
rect 11824 1353 11858 1387
rect 11918 1353 11952 1387
rect 12018 1353 12052 1387
rect 12318 1353 12352 1387
rect 12412 1353 12446 1387
rect 11524 1123 11558 1157
rect 11618 1123 11652 1157
rect 11918 1123 11952 1157
rect 12012 1123 12046 1157
rect 11424 983 11458 1017
rect 11518 983 11552 1017
rect 11612 983 11646 1017
rect 11724 983 11758 1017
rect 11818 983 11852 1017
rect 11912 983 11946 1017
rect 11024 843 11058 877
rect 11118 843 11152 877
rect 11218 843 11252 877
rect 11318 843 11352 877
rect 11718 843 11752 877
rect 11818 843 11852 877
rect 11912 843 11946 877
rect 11024 703 11058 737
rect 11118 703 11152 737
rect 11218 703 11252 737
rect 11318 703 11352 737
rect 11518 703 11552 737
rect 11618 703 11652 737
rect 11712 703 11746 737
rect 10524 563 10558 597
rect 10618 563 10652 597
rect 10718 563 10752 597
rect 10818 563 10852 597
rect 11118 563 11152 597
rect 11212 563 11246 597
rect 10324 423 10358 457
rect 10418 423 10452 457
rect 10518 423 10552 457
rect 10618 423 10652 457
rect 10718 423 10752 457
rect 10812 423 10846 457
rect 10924 423 10958 457
rect 11018 423 11052 457
rect 11112 423 11146 457
rect 12524 1493 12558 1527
rect 12618 1493 12652 1527
rect 12718 1493 12752 1527
rect 12924 1508 12958 1542
rect 13018 1493 13052 1527
rect 13112 1478 13146 1512
rect 13228 1493 13262 1527
rect 13328 1493 13362 1527
rect 13428 1493 13462 1527
rect 13528 1493 13562 1527
rect 13628 1493 13662 1527
rect 12524 1353 12558 1387
rect 12618 1353 12652 1387
rect 12924 1368 12958 1402
rect 13018 1353 13052 1387
rect 13112 1338 13146 1372
rect 13228 1353 13262 1387
rect 13328 1353 13362 1387
rect 13428 1353 13462 1387
rect 13528 1353 13562 1387
rect 13628 1353 13662 1387
rect 12124 1123 12158 1157
rect 12218 1123 12252 1157
rect 12518 1123 12552 1157
rect 12612 1123 12646 1157
rect 12724 1123 12758 1157
rect 12812 1123 12846 1157
rect 12924 1138 12958 1172
rect 13018 1123 13052 1157
rect 13112 1108 13146 1142
rect 13228 1123 13262 1157
rect 13328 1123 13362 1157
rect 13428 1123 13462 1157
rect 13528 1123 13562 1157
rect 13628 1123 13662 1157
rect 12024 983 12058 1017
rect 12118 983 12152 1017
rect 12218 983 12252 1017
rect 12618 983 12652 1017
rect 12718 983 12752 1017
rect 12812 983 12846 1017
rect 12924 998 12958 1032
rect 13018 983 13052 1017
rect 13112 968 13146 1002
rect 13228 983 13262 1017
rect 13328 983 13362 1017
rect 13428 983 13462 1017
rect 13528 983 13562 1017
rect 13628 983 13662 1017
rect 12024 843 12058 877
rect 12118 843 12152 877
rect 12218 843 12252 877
rect 12312 843 12346 877
rect 11824 703 11858 737
rect 11918 703 11952 737
rect 12018 703 12052 737
rect 12112 703 12146 737
rect 12424 843 12458 877
rect 12512 843 12546 877
rect 12624 843 12658 877
rect 12718 843 12752 877
rect 12924 858 12958 892
rect 13018 843 13052 877
rect 13112 828 13146 862
rect 13228 843 13262 877
rect 13328 843 13362 877
rect 13428 843 13462 877
rect 13528 843 13562 877
rect 13628 843 13662 877
rect 12224 703 12258 737
rect 12318 703 12352 737
rect 12518 703 12552 737
rect 12618 703 12652 737
rect 12924 718 12958 752
rect 13018 703 13052 737
rect 13112 688 13146 722
rect 13228 703 13262 737
rect 13328 703 13362 737
rect 13428 703 13462 737
rect 13528 703 13562 737
rect 13628 703 13662 737
rect 11324 563 11358 597
rect 11418 563 11452 597
rect 11518 563 11552 597
rect 11618 563 11652 597
rect 11718 563 11752 597
rect 11818 563 11852 597
rect 11918 563 11952 597
rect 12118 563 12152 597
rect 12218 563 12252 597
rect 12318 563 12352 597
rect 12418 563 12452 597
rect 12518 563 12552 597
rect 12618 563 12652 597
rect 12718 563 12752 597
rect 12812 563 12846 597
rect 12924 578 12958 612
rect 13018 563 13052 597
rect 13112 548 13146 582
rect 13228 563 13262 597
rect 13328 563 13362 597
rect 13428 563 13462 597
rect 13528 563 13562 597
rect 13628 563 13662 597
rect 11224 423 11258 457
rect 11312 423 11346 457
rect 11424 423 11458 457
rect 11518 423 11552 457
rect 12018 423 12052 457
rect 12118 423 12152 457
rect 12218 423 12252 457
rect 12312 423 12346 457
rect 10224 283 10258 317
rect 10318 283 10352 317
rect 10418 283 10452 317
rect 10718 283 10752 317
rect 10818 283 10852 317
rect 10918 283 10952 317
rect 11318 283 11352 317
rect 11412 283 11446 317
rect 7124 143 7158 177
rect 7218 143 7252 177
rect 7318 143 7352 177
rect 7618 143 7652 177
rect 7718 143 7752 177
rect 7918 143 7952 177
rect 8018 143 8052 177
rect 8318 143 8352 177
rect 8418 143 8452 177
rect 8718 143 8752 177
rect 8818 143 8852 177
rect 8918 143 8952 177
rect 9018 143 9052 177
rect 9118 143 9152 177
rect 9318 143 9352 177
rect 9418 143 9452 177
rect 9618 143 9652 177
rect 9718 143 9752 177
rect 9818 143 9852 177
rect 9918 143 9952 177
rect 10018 143 10052 177
rect 10118 143 10152 177
rect 10218 143 10252 177
rect 10618 143 10652 177
rect 10718 143 10752 177
rect 10918 143 10952 177
rect 11018 143 11052 177
rect 11118 143 11152 177
rect 11318 143 11352 177
rect 11412 143 11446 177
rect 11524 283 11558 317
rect 11618 283 11652 317
rect 11718 283 11752 317
rect 11818 283 11852 317
rect 12018 283 12052 317
rect 12118 283 12152 317
rect 12212 283 12246 317
rect 12424 423 12458 457
rect 12518 423 12552 457
rect 12718 423 12752 457
rect 12812 423 12846 457
rect 12924 438 12958 472
rect 13018 423 13052 457
rect 13112 408 13146 442
rect 13228 423 13262 457
rect 13328 423 13362 457
rect 13428 423 13462 457
rect 13528 423 13562 457
rect 13628 423 13662 457
rect 12324 283 12358 317
rect 12418 283 12452 317
rect 12518 283 12552 317
rect 12618 283 12652 317
rect 12924 298 12958 332
rect 13018 283 13052 317
rect 13112 268 13146 302
rect 13228 283 13262 317
rect 13328 283 13362 317
rect 13428 283 13462 317
rect 13528 283 13562 317
rect 13628 283 13662 317
rect 11524 143 11558 177
rect 11618 143 11652 177
rect 11818 143 11852 177
rect 11918 143 11952 177
rect 12018 143 12052 177
rect 12118 143 12152 177
rect 12418 143 12452 177
rect 12518 143 12552 177
rect 12618 143 12652 177
rect 12718 143 12752 177
rect 12924 158 12958 192
rect 13018 143 13052 177
rect 13112 128 13146 162
rect 13228 143 13262 177
rect 13328 143 13362 177
rect 13428 143 13462 177
rect 13528 143 13562 177
rect 13628 143 13662 177
rect -82 -183 -48 -149
rect 18 -183 52 -149
rect 118 -183 152 -149
rect 218 -183 252 -149
rect 318 -183 352 -149
rect 418 -183 452 -149
rect 518 -183 552 -149
rect 618 -183 652 -149
rect 718 -183 752 -149
rect 818 -183 852 -149
rect 918 -183 952 -149
rect 1018 -183 1052 -149
rect 1118 -183 1152 -149
rect 1218 -183 1252 -149
rect 1318 -183 1352 -149
rect 1418 -183 1452 -149
rect 1518 -183 1552 -149
rect 1618 -183 1652 -149
rect 1718 -183 1752 -149
rect 1818 -183 1852 -149
rect 1918 -183 1952 -149
rect 2018 -183 2052 -149
rect 2118 -183 2152 -149
rect 2218 -183 2252 -149
rect 2318 -183 2352 -149
rect 2418 -183 2452 -149
rect 2518 -183 2552 -149
rect 2618 -183 2652 -149
rect 2718 -183 2752 -149
rect 2818 -183 2852 -149
rect 2918 -183 2952 -149
rect 3018 -183 3052 -149
rect 3118 -183 3152 -149
rect 3218 -183 3252 -149
rect 3318 -183 3352 -149
rect 3418 -183 3452 -149
rect 3518 -183 3552 -149
rect 3618 -183 3652 -149
rect 3718 -183 3752 -149
rect 3818 -183 3852 -149
rect 3918 -183 3952 -149
rect 4018 -183 4052 -149
rect 4118 -183 4152 -149
rect 4218 -183 4252 -149
rect 4318 -183 4352 -149
rect 4418 -183 4452 -149
rect 4518 -183 4552 -149
rect 4618 -183 4652 -149
rect 4718 -183 4752 -149
rect 4818 -183 4852 -149
rect 4918 -183 4952 -149
rect 5018 -183 5052 -149
rect 5118 -183 5152 -149
rect 5218 -183 5252 -149
rect 5318 -183 5352 -149
rect 5418 -183 5452 -149
rect 5518 -183 5552 -149
rect 5618 -183 5652 -149
rect 5718 -183 5752 -149
rect 5818 -183 5852 -149
rect 5918 -183 5952 -149
rect 6018 -183 6052 -149
rect 6118 -183 6152 -149
rect 6218 -183 6252 -149
rect 6318 -183 6352 -149
rect 6418 -183 6452 -149
rect 6518 -183 6552 -149
rect 6618 -183 6652 -149
rect 6718 -183 6752 -149
rect 6818 -183 6852 -149
rect 6918 -183 6952 -149
rect 7018 -183 7052 -149
rect 7118 -183 7152 -149
rect 7218 -183 7252 -149
rect 7318 -183 7352 -149
rect 7418 -183 7452 -149
rect 7518 -183 7552 -149
rect 7618 -183 7652 -149
rect 7718 -183 7752 -149
rect 7818 -183 7852 -149
rect 7918 -183 7952 -149
rect 8018 -183 8052 -149
rect 8118 -183 8152 -149
rect 8218 -183 8252 -149
rect 8318 -183 8352 -149
rect 8418 -183 8452 -149
rect 8518 -183 8552 -149
rect 8618 -183 8652 -149
rect 8718 -183 8752 -149
rect 8818 -183 8852 -149
rect 8918 -183 8952 -149
rect 9018 -183 9052 -149
rect 9118 -183 9152 -149
rect 9218 -183 9252 -149
rect 9318 -183 9352 -149
rect 9418 -183 9452 -149
rect 9518 -183 9552 -149
rect 9618 -183 9652 -149
rect 9718 -183 9752 -149
rect 9818 -183 9852 -149
rect 9918 -183 9952 -149
rect 10018 -183 10052 -149
rect 10118 -183 10152 -149
rect 10218 -183 10252 -149
rect 10318 -183 10352 -149
rect 10418 -183 10452 -149
rect 10518 -183 10552 -149
rect 10618 -183 10652 -149
rect 10718 -183 10752 -149
rect 10818 -183 10852 -149
rect 10918 -183 10952 -149
rect 11018 -183 11052 -149
rect 11118 -183 11152 -149
rect 11218 -183 11252 -149
rect 11318 -183 11352 -149
rect 11418 -183 11452 -149
rect 11518 -183 11552 -149
rect 11618 -183 11652 -149
rect 11718 -183 11752 -149
rect 11818 -183 11852 -149
rect 11918 -183 11952 -149
rect 12018 -183 12052 -149
rect 12118 -183 12152 -149
rect 12218 -183 12252 -149
rect 12318 -183 12352 -149
rect 12418 -183 12452 -149
rect 12518 -183 12552 -149
rect 12618 -183 12652 -149
rect 12718 -183 12752 -149
rect 14562 -242 14596 -208
rect 14630 -242 14664 -208
rect 15678 -242 15712 -208
rect 15746 -242 15780 -208
rect 14562 -342 14596 -308
rect 14630 -342 14664 -308
rect 15678 -342 15712 -308
rect 15746 -342 15780 -308
rect 14562 -442 14596 -408
rect 14630 -442 14664 -408
rect 15678 -442 15712 -408
rect 15746 -442 15780 -408
rect 14562 -542 14596 -508
rect 14630 -542 14664 -508
rect 15678 -542 15712 -508
rect 15746 -542 15780 -508
rect 14562 -642 14596 -608
rect 14630 -642 14664 -608
rect 15678 -642 15712 -608
rect 15746 -642 15780 -608
rect 14562 -742 14596 -708
rect 14630 -742 14664 -708
rect 15678 -742 15712 -708
rect 15746 -742 15780 -708
rect 14562 -842 14596 -808
rect 14630 -842 14664 -808
rect -2 -892 32 -858
rect 66 -892 100 -858
rect 170 -892 204 -858
rect 238 -892 272 -858
rect 398 -892 432 -858
rect 466 -892 500 -858
rect 570 -892 604 -858
rect 638 -892 672 -858
rect 798 -892 832 -858
rect 866 -892 900 -858
rect -2 -992 32 -958
rect 66 -992 100 -958
rect 170 -992 204 -958
rect 238 -992 272 -958
rect 398 -992 432 -958
rect 466 -992 500 -958
rect 970 -892 1004 -858
rect 1038 -892 1072 -858
rect 1198 -892 1232 -858
rect 1266 -892 1300 -858
rect 1370 -892 1404 -858
rect 1438 -892 1472 -858
rect 1598 -892 1632 -858
rect 1666 -892 1700 -858
rect 570 -992 604 -958
rect 638 -992 672 -958
rect 798 -992 832 -958
rect 866 -992 900 -958
rect -2 -1092 32 -1058
rect 66 -1092 100 -1058
rect 170 -1092 204 -1058
rect 238 -1092 272 -1058
rect 398 -1092 432 -1058
rect 466 -1092 500 -1058
rect 970 -992 1004 -958
rect 1038 -992 1072 -958
rect 1198 -992 1232 -958
rect 1266 -992 1300 -958
rect 1770 -892 1804 -858
rect 1838 -892 1872 -858
rect 1998 -892 2032 -858
rect 2066 -892 2100 -858
rect 2170 -892 2204 -858
rect 2238 -892 2272 -858
rect 2398 -892 2432 -858
rect 2466 -892 2500 -858
rect 1370 -992 1404 -958
rect 1438 -992 1472 -958
rect 1598 -992 1632 -958
rect 1666 -992 1700 -958
rect 570 -1092 604 -1058
rect 638 -1092 672 -1058
rect 798 -1092 832 -1058
rect 866 -1092 900 -1058
rect -2 -1192 32 -1158
rect 66 -1192 100 -1158
rect 170 -1192 204 -1158
rect 238 -1192 272 -1158
rect 398 -1192 432 -1158
rect 466 -1192 500 -1158
rect 970 -1092 1004 -1058
rect 1038 -1092 1072 -1058
rect 1198 -1092 1232 -1058
rect 1266 -1092 1300 -1058
rect 1770 -992 1804 -958
rect 1838 -992 1872 -958
rect 1998 -992 2032 -958
rect 2066 -992 2100 -958
rect 2570 -892 2604 -858
rect 2638 -892 2672 -858
rect 2798 -892 2832 -858
rect 2866 -892 2900 -858
rect 2970 -892 3004 -858
rect 3038 -892 3072 -858
rect 3198 -892 3232 -858
rect 3266 -892 3300 -858
rect 2170 -992 2204 -958
rect 2238 -992 2272 -958
rect 2398 -992 2432 -958
rect 2466 -992 2500 -958
rect 1370 -1092 1404 -1058
rect 1438 -1092 1472 -1058
rect 1598 -1092 1632 -1058
rect 1666 -1092 1700 -1058
rect 570 -1192 604 -1158
rect 638 -1192 672 -1158
rect 798 -1192 832 -1158
rect 866 -1192 900 -1158
rect -2 -1292 32 -1258
rect 66 -1292 100 -1258
rect 170 -1292 204 -1258
rect 238 -1292 272 -1258
rect 398 -1292 432 -1258
rect 466 -1292 500 -1258
rect 970 -1192 1004 -1158
rect 1038 -1192 1072 -1158
rect 1198 -1192 1232 -1158
rect 1266 -1192 1300 -1158
rect 1770 -1092 1804 -1058
rect 1838 -1092 1872 -1058
rect 1998 -1092 2032 -1058
rect 2066 -1092 2100 -1058
rect 2570 -992 2604 -958
rect 2638 -992 2672 -958
rect 2798 -992 2832 -958
rect 2866 -992 2900 -958
rect 3370 -892 3404 -858
rect 3438 -892 3472 -858
rect 3598 -892 3632 -858
rect 3666 -892 3700 -858
rect 3770 -892 3804 -858
rect 3838 -892 3872 -858
rect 3998 -892 4032 -858
rect 4066 -892 4100 -858
rect 2970 -992 3004 -958
rect 3038 -992 3072 -958
rect 3198 -992 3232 -958
rect 3266 -992 3300 -958
rect 2170 -1092 2204 -1058
rect 2238 -1092 2272 -1058
rect 2398 -1092 2432 -1058
rect 2466 -1092 2500 -1058
rect 1370 -1192 1404 -1158
rect 1438 -1192 1472 -1158
rect 1598 -1192 1632 -1158
rect 1666 -1192 1700 -1158
rect 570 -1292 604 -1258
rect 638 -1292 672 -1258
rect 798 -1292 832 -1258
rect 866 -1292 900 -1258
rect -2 -1392 32 -1358
rect 66 -1392 100 -1358
rect 170 -1392 204 -1358
rect 238 -1392 272 -1358
rect 398 -1392 432 -1358
rect 466 -1392 500 -1358
rect 970 -1292 1004 -1258
rect 1038 -1292 1072 -1258
rect 1198 -1292 1232 -1258
rect 1266 -1292 1300 -1258
rect 1770 -1192 1804 -1158
rect 1838 -1192 1872 -1158
rect 1998 -1192 2032 -1158
rect 2066 -1192 2100 -1158
rect 2570 -1092 2604 -1058
rect 2638 -1092 2672 -1058
rect 2798 -1092 2832 -1058
rect 2866 -1092 2900 -1058
rect 3370 -992 3404 -958
rect 3438 -992 3472 -958
rect 3598 -992 3632 -958
rect 3666 -992 3700 -958
rect 4170 -892 4204 -858
rect 4238 -892 4272 -858
rect 4398 -892 4432 -858
rect 4466 -892 4500 -858
rect 4570 -892 4604 -858
rect 4638 -892 4672 -858
rect 4798 -892 4832 -858
rect 4866 -892 4900 -858
rect 3770 -992 3804 -958
rect 3838 -992 3872 -958
rect 3998 -992 4032 -958
rect 4066 -992 4100 -958
rect 2970 -1092 3004 -1058
rect 3038 -1092 3072 -1058
rect 3198 -1092 3232 -1058
rect 3266 -1092 3300 -1058
rect 2170 -1192 2204 -1158
rect 2238 -1192 2272 -1158
rect 2398 -1192 2432 -1158
rect 2466 -1192 2500 -1158
rect 1370 -1292 1404 -1258
rect 1438 -1292 1472 -1258
rect 1598 -1292 1632 -1258
rect 1666 -1292 1700 -1258
rect 570 -1392 604 -1358
rect 638 -1392 672 -1358
rect 798 -1392 832 -1358
rect 866 -1392 900 -1358
rect -2 -1492 32 -1458
rect 66 -1492 100 -1458
rect 170 -1492 204 -1458
rect 238 -1492 272 -1458
rect 398 -1492 432 -1458
rect 466 -1492 500 -1458
rect 970 -1392 1004 -1358
rect 1038 -1392 1072 -1358
rect 1198 -1392 1232 -1358
rect 1266 -1392 1300 -1358
rect 1770 -1292 1804 -1258
rect 1838 -1292 1872 -1258
rect 1998 -1292 2032 -1258
rect 2066 -1292 2100 -1258
rect 2570 -1192 2604 -1158
rect 2638 -1192 2672 -1158
rect 2798 -1192 2832 -1158
rect 2866 -1192 2900 -1158
rect 3370 -1092 3404 -1058
rect 3438 -1092 3472 -1058
rect 3598 -1092 3632 -1058
rect 3666 -1092 3700 -1058
rect 4170 -992 4204 -958
rect 4238 -992 4272 -958
rect 4398 -992 4432 -958
rect 4466 -992 4500 -958
rect 4970 -892 5004 -858
rect 5038 -892 5072 -858
rect 5198 -892 5232 -858
rect 5266 -892 5300 -858
rect 5370 -892 5404 -858
rect 5438 -892 5472 -858
rect 5598 -892 5632 -858
rect 5666 -892 5700 -858
rect 4570 -992 4604 -958
rect 4638 -992 4672 -958
rect 4798 -992 4832 -958
rect 4866 -992 4900 -958
rect 3770 -1092 3804 -1058
rect 3838 -1092 3872 -1058
rect 3998 -1092 4032 -1058
rect 4066 -1092 4100 -1058
rect 2970 -1192 3004 -1158
rect 3038 -1192 3072 -1158
rect 3198 -1192 3232 -1158
rect 3266 -1192 3300 -1158
rect 2170 -1292 2204 -1258
rect 2238 -1292 2272 -1258
rect 2398 -1292 2432 -1258
rect 2466 -1292 2500 -1258
rect 1370 -1392 1404 -1358
rect 1438 -1392 1472 -1358
rect 1598 -1392 1632 -1358
rect 1666 -1392 1700 -1358
rect 570 -1492 604 -1458
rect 638 -1492 672 -1458
rect 798 -1492 832 -1458
rect 866 -1492 900 -1458
rect -2 -1592 32 -1558
rect 66 -1592 100 -1558
rect 170 -1592 204 -1558
rect 238 -1592 272 -1558
rect 398 -1592 432 -1558
rect 466 -1592 500 -1558
rect 970 -1492 1004 -1458
rect 1038 -1492 1072 -1458
rect 1198 -1492 1232 -1458
rect 1266 -1492 1300 -1458
rect 1770 -1392 1804 -1358
rect 1838 -1392 1872 -1358
rect 1998 -1392 2032 -1358
rect 2066 -1392 2100 -1358
rect 2570 -1292 2604 -1258
rect 2638 -1292 2672 -1258
rect 2798 -1292 2832 -1258
rect 2866 -1292 2900 -1258
rect 3370 -1192 3404 -1158
rect 3438 -1192 3472 -1158
rect 3598 -1192 3632 -1158
rect 3666 -1192 3700 -1158
rect 4170 -1092 4204 -1058
rect 4238 -1092 4272 -1058
rect 4398 -1092 4432 -1058
rect 4466 -1092 4500 -1058
rect 4970 -992 5004 -958
rect 5038 -992 5072 -958
rect 5198 -992 5232 -958
rect 5266 -992 5300 -958
rect 5770 -892 5804 -858
rect 5838 -892 5872 -858
rect 5998 -892 6032 -858
rect 6066 -892 6100 -858
rect 6170 -892 6204 -858
rect 6238 -892 6272 -858
rect 6398 -892 6432 -858
rect 6466 -892 6500 -858
rect 5370 -992 5404 -958
rect 5438 -992 5472 -958
rect 5598 -992 5632 -958
rect 5666 -992 5700 -958
rect 4570 -1092 4604 -1058
rect 4638 -1092 4672 -1058
rect 4798 -1092 4832 -1058
rect 4866 -1092 4900 -1058
rect 3770 -1192 3804 -1158
rect 3838 -1192 3872 -1158
rect 3998 -1192 4032 -1158
rect 4066 -1192 4100 -1158
rect 2970 -1292 3004 -1258
rect 3038 -1292 3072 -1258
rect 3198 -1292 3232 -1258
rect 3266 -1292 3300 -1258
rect 2170 -1392 2204 -1358
rect 2238 -1392 2272 -1358
rect 2398 -1392 2432 -1358
rect 2466 -1392 2500 -1358
rect 1370 -1492 1404 -1458
rect 1438 -1492 1472 -1458
rect 1598 -1492 1632 -1458
rect 1666 -1492 1700 -1458
rect 570 -1592 604 -1558
rect 638 -1592 672 -1558
rect 798 -1592 832 -1558
rect 866 -1592 900 -1558
rect -2 -1692 32 -1658
rect 66 -1692 100 -1658
rect 170 -1692 204 -1658
rect 238 -1692 272 -1658
rect 398 -1692 432 -1658
rect 466 -1692 500 -1658
rect 970 -1592 1004 -1558
rect 1038 -1592 1072 -1558
rect 1198 -1592 1232 -1558
rect 1266 -1592 1300 -1558
rect 1770 -1492 1804 -1458
rect 1838 -1492 1872 -1458
rect 1998 -1492 2032 -1458
rect 2066 -1492 2100 -1458
rect 2570 -1392 2604 -1358
rect 2638 -1392 2672 -1358
rect 2798 -1392 2832 -1358
rect 2866 -1392 2900 -1358
rect 3370 -1292 3404 -1258
rect 3438 -1292 3472 -1258
rect 3598 -1292 3632 -1258
rect 3666 -1292 3700 -1258
rect 4170 -1192 4204 -1158
rect 4238 -1192 4272 -1158
rect 4398 -1192 4432 -1158
rect 4466 -1192 4500 -1158
rect 4970 -1092 5004 -1058
rect 5038 -1092 5072 -1058
rect 5198 -1092 5232 -1058
rect 5266 -1092 5300 -1058
rect 5770 -992 5804 -958
rect 5838 -992 5872 -958
rect 5998 -992 6032 -958
rect 6066 -992 6100 -958
rect 6570 -892 6604 -858
rect 6638 -892 6672 -858
rect 6798 -892 6832 -858
rect 6866 -892 6900 -858
rect 6970 -892 7004 -858
rect 7038 -892 7072 -858
rect 7198 -892 7232 -858
rect 7266 -892 7300 -858
rect 6170 -992 6204 -958
rect 6238 -992 6272 -958
rect 6398 -992 6432 -958
rect 6466 -992 6500 -958
rect 5370 -1092 5404 -1058
rect 5438 -1092 5472 -1058
rect 5598 -1092 5632 -1058
rect 5666 -1092 5700 -1058
rect 4570 -1192 4604 -1158
rect 4638 -1192 4672 -1158
rect 4798 -1192 4832 -1158
rect 4866 -1192 4900 -1158
rect 3770 -1292 3804 -1258
rect 3838 -1292 3872 -1258
rect 3998 -1292 4032 -1258
rect 4066 -1292 4100 -1258
rect 2970 -1392 3004 -1358
rect 3038 -1392 3072 -1358
rect 3198 -1392 3232 -1358
rect 3266 -1392 3300 -1358
rect 2170 -1492 2204 -1458
rect 2238 -1492 2272 -1458
rect 2398 -1492 2432 -1458
rect 2466 -1492 2500 -1458
rect 1370 -1592 1404 -1558
rect 1438 -1592 1472 -1558
rect 1598 -1592 1632 -1558
rect 1666 -1592 1700 -1558
rect 570 -1692 604 -1658
rect 638 -1692 672 -1658
rect 798 -1692 832 -1658
rect 866 -1692 900 -1658
rect -2 -1792 32 -1758
rect 66 -1792 100 -1758
rect 170 -1792 204 -1758
rect 238 -1792 272 -1758
rect 398 -1792 432 -1758
rect 466 -1792 500 -1758
rect 970 -1692 1004 -1658
rect 1038 -1692 1072 -1658
rect 1198 -1692 1232 -1658
rect 1266 -1692 1300 -1658
rect 1770 -1592 1804 -1558
rect 1838 -1592 1872 -1558
rect 1998 -1592 2032 -1558
rect 2066 -1592 2100 -1558
rect 2570 -1492 2604 -1458
rect 2638 -1492 2672 -1458
rect 2798 -1492 2832 -1458
rect 2866 -1492 2900 -1458
rect 3370 -1392 3404 -1358
rect 3438 -1392 3472 -1358
rect 3598 -1392 3632 -1358
rect 3666 -1392 3700 -1358
rect 4170 -1292 4204 -1258
rect 4238 -1292 4272 -1258
rect 4398 -1292 4432 -1258
rect 4466 -1292 4500 -1258
rect 4970 -1192 5004 -1158
rect 5038 -1192 5072 -1158
rect 5198 -1192 5232 -1158
rect 5266 -1192 5300 -1158
rect 5770 -1092 5804 -1058
rect 5838 -1092 5872 -1058
rect 5998 -1092 6032 -1058
rect 6066 -1092 6100 -1058
rect 6570 -992 6604 -958
rect 6638 -992 6672 -958
rect 6798 -992 6832 -958
rect 6866 -992 6900 -958
rect 7370 -892 7404 -858
rect 7438 -892 7472 -858
rect 7598 -892 7632 -858
rect 7666 -892 7700 -858
rect 7770 -892 7804 -858
rect 7838 -892 7872 -858
rect 7998 -892 8032 -858
rect 8066 -892 8100 -858
rect 6970 -992 7004 -958
rect 7038 -992 7072 -958
rect 7198 -992 7232 -958
rect 7266 -992 7300 -958
rect 6170 -1092 6204 -1058
rect 6238 -1092 6272 -1058
rect 6398 -1092 6432 -1058
rect 6466 -1092 6500 -1058
rect 5370 -1192 5404 -1158
rect 5438 -1192 5472 -1158
rect 5598 -1192 5632 -1158
rect 5666 -1192 5700 -1158
rect 4570 -1292 4604 -1258
rect 4638 -1292 4672 -1258
rect 4798 -1292 4832 -1258
rect 4866 -1292 4900 -1258
rect 3770 -1392 3804 -1358
rect 3838 -1392 3872 -1358
rect 3998 -1392 4032 -1358
rect 4066 -1392 4100 -1358
rect 2970 -1492 3004 -1458
rect 3038 -1492 3072 -1458
rect 3198 -1492 3232 -1458
rect 3266 -1492 3300 -1458
rect 2170 -1592 2204 -1558
rect 2238 -1592 2272 -1558
rect 2398 -1592 2432 -1558
rect 2466 -1592 2500 -1558
rect 1370 -1692 1404 -1658
rect 1438 -1692 1472 -1658
rect 1598 -1692 1632 -1658
rect 1666 -1692 1700 -1658
rect 570 -1792 604 -1758
rect 638 -1792 672 -1758
rect 798 -1792 832 -1758
rect 866 -1792 900 -1758
rect -2 -1892 32 -1858
rect 66 -1892 100 -1858
rect 170 -1892 204 -1858
rect 238 -1892 272 -1858
rect 398 -1892 432 -1858
rect 466 -1892 500 -1858
rect 970 -1792 1004 -1758
rect 1038 -1792 1072 -1758
rect 1198 -1792 1232 -1758
rect 1266 -1792 1300 -1758
rect 1770 -1692 1804 -1658
rect 1838 -1692 1872 -1658
rect 1998 -1692 2032 -1658
rect 2066 -1692 2100 -1658
rect 2570 -1592 2604 -1558
rect 2638 -1592 2672 -1558
rect 2798 -1592 2832 -1558
rect 2866 -1592 2900 -1558
rect 3370 -1492 3404 -1458
rect 3438 -1492 3472 -1458
rect 3598 -1492 3632 -1458
rect 3666 -1492 3700 -1458
rect 4170 -1392 4204 -1358
rect 4238 -1392 4272 -1358
rect 4398 -1392 4432 -1358
rect 4466 -1392 4500 -1358
rect 4970 -1292 5004 -1258
rect 5038 -1292 5072 -1258
rect 5198 -1292 5232 -1258
rect 5266 -1292 5300 -1258
rect 5770 -1192 5804 -1158
rect 5838 -1192 5872 -1158
rect 5998 -1192 6032 -1158
rect 6066 -1192 6100 -1158
rect 6570 -1092 6604 -1058
rect 6638 -1092 6672 -1058
rect 6798 -1092 6832 -1058
rect 6866 -1092 6900 -1058
rect 7370 -992 7404 -958
rect 7438 -992 7472 -958
rect 7598 -992 7632 -958
rect 7666 -992 7700 -958
rect 8170 -892 8204 -858
rect 8238 -892 8272 -858
rect 8398 -892 8432 -858
rect 8466 -892 8500 -858
rect 8570 -892 8604 -858
rect 8638 -892 8672 -858
rect 8798 -892 8832 -858
rect 8866 -892 8900 -858
rect 7770 -992 7804 -958
rect 7838 -992 7872 -958
rect 7998 -992 8032 -958
rect 8066 -992 8100 -958
rect 6970 -1092 7004 -1058
rect 7038 -1092 7072 -1058
rect 7198 -1092 7232 -1058
rect 7266 -1092 7300 -1058
rect 6170 -1192 6204 -1158
rect 6238 -1192 6272 -1158
rect 6398 -1192 6432 -1158
rect 6466 -1192 6500 -1158
rect 5370 -1292 5404 -1258
rect 5438 -1292 5472 -1258
rect 5598 -1292 5632 -1258
rect 5666 -1292 5700 -1258
rect 4570 -1392 4604 -1358
rect 4638 -1392 4672 -1358
rect 4798 -1392 4832 -1358
rect 4866 -1392 4900 -1358
rect 3770 -1492 3804 -1458
rect 3838 -1492 3872 -1458
rect 3998 -1492 4032 -1458
rect 4066 -1492 4100 -1458
rect 2970 -1592 3004 -1558
rect 3038 -1592 3072 -1558
rect 3198 -1592 3232 -1558
rect 3266 -1592 3300 -1558
rect 2170 -1692 2204 -1658
rect 2238 -1692 2272 -1658
rect 2398 -1692 2432 -1658
rect 2466 -1692 2500 -1658
rect 1370 -1792 1404 -1758
rect 1438 -1792 1472 -1758
rect 1598 -1792 1632 -1758
rect 1666 -1792 1700 -1758
rect 570 -1892 604 -1858
rect 638 -1892 672 -1858
rect 798 -1892 832 -1858
rect 866 -1892 900 -1858
rect -2 -1992 32 -1958
rect 66 -1992 100 -1958
rect 170 -1992 204 -1958
rect 238 -1992 272 -1958
rect 398 -1992 432 -1958
rect 466 -1992 500 -1958
rect 970 -1892 1004 -1858
rect 1038 -1892 1072 -1858
rect 1198 -1892 1232 -1858
rect 1266 -1892 1300 -1858
rect 1770 -1792 1804 -1758
rect 1838 -1792 1872 -1758
rect 1998 -1792 2032 -1758
rect 2066 -1792 2100 -1758
rect 2570 -1692 2604 -1658
rect 2638 -1692 2672 -1658
rect 2798 -1692 2832 -1658
rect 2866 -1692 2900 -1658
rect 3370 -1592 3404 -1558
rect 3438 -1592 3472 -1558
rect 3598 -1592 3632 -1558
rect 3666 -1592 3700 -1558
rect 4170 -1492 4204 -1458
rect 4238 -1492 4272 -1458
rect 4398 -1492 4432 -1458
rect 4466 -1492 4500 -1458
rect 4970 -1392 5004 -1358
rect 5038 -1392 5072 -1358
rect 5198 -1392 5232 -1358
rect 5266 -1392 5300 -1358
rect 5770 -1292 5804 -1258
rect 5838 -1292 5872 -1258
rect 5998 -1292 6032 -1258
rect 6066 -1292 6100 -1258
rect 6570 -1192 6604 -1158
rect 6638 -1192 6672 -1158
rect 6798 -1192 6832 -1158
rect 6866 -1192 6900 -1158
rect 7370 -1092 7404 -1058
rect 7438 -1092 7472 -1058
rect 7598 -1092 7632 -1058
rect 7666 -1092 7700 -1058
rect 8170 -992 8204 -958
rect 8238 -992 8272 -958
rect 8398 -992 8432 -958
rect 8466 -992 8500 -958
rect 8970 -892 9004 -858
rect 9038 -892 9072 -858
rect 9198 -892 9232 -858
rect 9266 -892 9300 -858
rect 9370 -892 9404 -858
rect 9438 -892 9472 -858
rect 9598 -892 9632 -858
rect 9666 -892 9700 -858
rect 8570 -992 8604 -958
rect 8638 -992 8672 -958
rect 8798 -992 8832 -958
rect 8866 -992 8900 -958
rect 7770 -1092 7804 -1058
rect 7838 -1092 7872 -1058
rect 7998 -1092 8032 -1058
rect 8066 -1092 8100 -1058
rect 6970 -1192 7004 -1158
rect 7038 -1192 7072 -1158
rect 7198 -1192 7232 -1158
rect 7266 -1192 7300 -1158
rect 6170 -1292 6204 -1258
rect 6238 -1292 6272 -1258
rect 6398 -1292 6432 -1258
rect 6466 -1292 6500 -1258
rect 5370 -1392 5404 -1358
rect 5438 -1392 5472 -1358
rect 5598 -1392 5632 -1358
rect 5666 -1392 5700 -1358
rect 4570 -1492 4604 -1458
rect 4638 -1492 4672 -1458
rect 4798 -1492 4832 -1458
rect 4866 -1492 4900 -1458
rect 3770 -1592 3804 -1558
rect 3838 -1592 3872 -1558
rect 3998 -1592 4032 -1558
rect 4066 -1592 4100 -1558
rect 2970 -1692 3004 -1658
rect 3038 -1692 3072 -1658
rect 3198 -1692 3232 -1658
rect 3266 -1692 3300 -1658
rect 2170 -1792 2204 -1758
rect 2238 -1792 2272 -1758
rect 2398 -1792 2432 -1758
rect 2466 -1792 2500 -1758
rect 1370 -1892 1404 -1858
rect 1438 -1892 1472 -1858
rect 1598 -1892 1632 -1858
rect 1666 -1892 1700 -1858
rect 570 -1992 604 -1958
rect 638 -1992 672 -1958
rect 798 -1992 832 -1958
rect 866 -1992 900 -1958
rect -2 -2092 32 -2058
rect 66 -2092 100 -2058
rect 170 -2092 204 -2058
rect 238 -2092 272 -2058
rect 398 -2092 432 -2058
rect 466 -2092 500 -2058
rect 970 -1992 1004 -1958
rect 1038 -1992 1072 -1958
rect 1198 -1992 1232 -1958
rect 1266 -1992 1300 -1958
rect 1770 -1892 1804 -1858
rect 1838 -1892 1872 -1858
rect 1998 -1892 2032 -1858
rect 2066 -1892 2100 -1858
rect 2570 -1792 2604 -1758
rect 2638 -1792 2672 -1758
rect 2798 -1792 2832 -1758
rect 2866 -1792 2900 -1758
rect 3370 -1692 3404 -1658
rect 3438 -1692 3472 -1658
rect 3598 -1692 3632 -1658
rect 3666 -1692 3700 -1658
rect 4170 -1592 4204 -1558
rect 4238 -1592 4272 -1558
rect 4398 -1592 4432 -1558
rect 4466 -1592 4500 -1558
rect 4970 -1492 5004 -1458
rect 5038 -1492 5072 -1458
rect 5198 -1492 5232 -1458
rect 5266 -1492 5300 -1458
rect 5770 -1392 5804 -1358
rect 5838 -1392 5872 -1358
rect 5998 -1392 6032 -1358
rect 6066 -1392 6100 -1358
rect 6570 -1292 6604 -1258
rect 6638 -1292 6672 -1258
rect 6798 -1292 6832 -1258
rect 6866 -1292 6900 -1258
rect 7370 -1192 7404 -1158
rect 7438 -1192 7472 -1158
rect 7598 -1192 7632 -1158
rect 7666 -1192 7700 -1158
rect 8170 -1092 8204 -1058
rect 8238 -1092 8272 -1058
rect 8398 -1092 8432 -1058
rect 8466 -1092 8500 -1058
rect 8970 -992 9004 -958
rect 9038 -992 9072 -958
rect 9198 -992 9232 -958
rect 9266 -992 9300 -958
rect 9770 -892 9804 -858
rect 9838 -892 9872 -858
rect 9998 -892 10032 -858
rect 10066 -892 10100 -858
rect 10170 -892 10204 -858
rect 10238 -892 10272 -858
rect 10398 -892 10432 -858
rect 10466 -892 10500 -858
rect 9370 -992 9404 -958
rect 9438 -992 9472 -958
rect 9598 -992 9632 -958
rect 9666 -992 9700 -958
rect 8570 -1092 8604 -1058
rect 8638 -1092 8672 -1058
rect 8798 -1092 8832 -1058
rect 8866 -1092 8900 -1058
rect 7770 -1192 7804 -1158
rect 7838 -1192 7872 -1158
rect 7998 -1192 8032 -1158
rect 8066 -1192 8100 -1158
rect 6970 -1292 7004 -1258
rect 7038 -1292 7072 -1258
rect 7198 -1292 7232 -1258
rect 7266 -1292 7300 -1258
rect 6170 -1392 6204 -1358
rect 6238 -1392 6272 -1358
rect 6398 -1392 6432 -1358
rect 6466 -1392 6500 -1358
rect 5370 -1492 5404 -1458
rect 5438 -1492 5472 -1458
rect 5598 -1492 5632 -1458
rect 5666 -1492 5700 -1458
rect 4570 -1592 4604 -1558
rect 4638 -1592 4672 -1558
rect 4798 -1592 4832 -1558
rect 4866 -1592 4900 -1558
rect 3770 -1692 3804 -1658
rect 3838 -1692 3872 -1658
rect 3998 -1692 4032 -1658
rect 4066 -1692 4100 -1658
rect 2970 -1792 3004 -1758
rect 3038 -1792 3072 -1758
rect 3198 -1792 3232 -1758
rect 3266 -1792 3300 -1758
rect 2170 -1892 2204 -1858
rect 2238 -1892 2272 -1858
rect 2398 -1892 2432 -1858
rect 2466 -1892 2500 -1858
rect 1370 -1992 1404 -1958
rect 1438 -1992 1472 -1958
rect 1598 -1992 1632 -1958
rect 1666 -1992 1700 -1958
rect 570 -2092 604 -2058
rect 638 -2092 672 -2058
rect 798 -2092 832 -2058
rect 866 -2092 900 -2058
rect 970 -2092 1004 -2058
rect 1038 -2092 1072 -2058
rect 1198 -2092 1232 -2058
rect 1266 -2092 1300 -2058
rect 1770 -1992 1804 -1958
rect 1838 -1992 1872 -1958
rect 1998 -1992 2032 -1958
rect 2066 -1992 2100 -1958
rect 2570 -1892 2604 -1858
rect 2638 -1892 2672 -1858
rect 2798 -1892 2832 -1858
rect 2866 -1892 2900 -1858
rect 3370 -1792 3404 -1758
rect 3438 -1792 3472 -1758
rect 3598 -1792 3632 -1758
rect 3666 -1792 3700 -1758
rect 4170 -1692 4204 -1658
rect 4238 -1692 4272 -1658
rect 4398 -1692 4432 -1658
rect 4466 -1692 4500 -1658
rect 4970 -1592 5004 -1558
rect 5038 -1592 5072 -1558
rect 5198 -1592 5232 -1558
rect 5266 -1592 5300 -1558
rect 5770 -1492 5804 -1458
rect 5838 -1492 5872 -1458
rect 5998 -1492 6032 -1458
rect 6066 -1492 6100 -1458
rect 6570 -1392 6604 -1358
rect 6638 -1392 6672 -1358
rect 6798 -1392 6832 -1358
rect 6866 -1392 6900 -1358
rect 7370 -1292 7404 -1258
rect 7438 -1292 7472 -1258
rect 7598 -1292 7632 -1258
rect 7666 -1292 7700 -1258
rect 8170 -1192 8204 -1158
rect 8238 -1192 8272 -1158
rect 8398 -1192 8432 -1158
rect 8466 -1192 8500 -1158
rect 8970 -1092 9004 -1058
rect 9038 -1092 9072 -1058
rect 9198 -1092 9232 -1058
rect 9266 -1092 9300 -1058
rect 9770 -992 9804 -958
rect 9838 -992 9872 -958
rect 9998 -992 10032 -958
rect 10066 -992 10100 -958
rect 10570 -892 10604 -858
rect 10638 -892 10672 -858
rect 10798 -892 10832 -858
rect 10866 -892 10900 -858
rect 10970 -892 11004 -858
rect 11038 -892 11072 -858
rect 11198 -892 11232 -858
rect 11266 -892 11300 -858
rect 10170 -992 10204 -958
rect 10238 -992 10272 -958
rect 10398 -992 10432 -958
rect 10466 -992 10500 -958
rect 9370 -1092 9404 -1058
rect 9438 -1092 9472 -1058
rect 9598 -1092 9632 -1058
rect 9666 -1092 9700 -1058
rect 8570 -1192 8604 -1158
rect 8638 -1192 8672 -1158
rect 8798 -1192 8832 -1158
rect 8866 -1192 8900 -1158
rect 7770 -1292 7804 -1258
rect 7838 -1292 7872 -1258
rect 7998 -1292 8032 -1258
rect 8066 -1292 8100 -1258
rect 6970 -1392 7004 -1358
rect 7038 -1392 7072 -1358
rect 7198 -1392 7232 -1358
rect 7266 -1392 7300 -1358
rect 6170 -1492 6204 -1458
rect 6238 -1492 6272 -1458
rect 6398 -1492 6432 -1458
rect 6466 -1492 6500 -1458
rect 5370 -1592 5404 -1558
rect 5438 -1592 5472 -1558
rect 5598 -1592 5632 -1558
rect 5666 -1592 5700 -1558
rect 4570 -1692 4604 -1658
rect 4638 -1692 4672 -1658
rect 4798 -1692 4832 -1658
rect 4866 -1692 4900 -1658
rect 3770 -1792 3804 -1758
rect 3838 -1792 3872 -1758
rect 3998 -1792 4032 -1758
rect 4066 -1792 4100 -1758
rect 2970 -1892 3004 -1858
rect 3038 -1892 3072 -1858
rect 3198 -1892 3232 -1858
rect 3266 -1892 3300 -1858
rect 2170 -1992 2204 -1958
rect 2238 -1992 2272 -1958
rect 2398 -1992 2432 -1958
rect 2466 -1992 2500 -1958
rect 1370 -2092 1404 -2058
rect 1438 -2092 1472 -2058
rect 1598 -2092 1632 -2058
rect 1666 -2092 1700 -2058
rect 1770 -2092 1804 -2058
rect 1838 -2092 1872 -2058
rect 1998 -2092 2032 -2058
rect 2066 -2092 2100 -2058
rect 2570 -1992 2604 -1958
rect 2638 -1992 2672 -1958
rect 2798 -1992 2832 -1958
rect 2866 -1992 2900 -1958
rect 3370 -1892 3404 -1858
rect 3438 -1892 3472 -1858
rect 3598 -1892 3632 -1858
rect 3666 -1892 3700 -1858
rect 4170 -1792 4204 -1758
rect 4238 -1792 4272 -1758
rect 4398 -1792 4432 -1758
rect 4466 -1792 4500 -1758
rect 4970 -1692 5004 -1658
rect 5038 -1692 5072 -1658
rect 5198 -1692 5232 -1658
rect 5266 -1692 5300 -1658
rect 5770 -1592 5804 -1558
rect 5838 -1592 5872 -1558
rect 5998 -1592 6032 -1558
rect 6066 -1592 6100 -1558
rect 6570 -1492 6604 -1458
rect 6638 -1492 6672 -1458
rect 6798 -1492 6832 -1458
rect 6866 -1492 6900 -1458
rect 7370 -1392 7404 -1358
rect 7438 -1392 7472 -1358
rect 7598 -1392 7632 -1358
rect 7666 -1392 7700 -1358
rect 8170 -1292 8204 -1258
rect 8238 -1292 8272 -1258
rect 8398 -1292 8432 -1258
rect 8466 -1292 8500 -1258
rect 8970 -1192 9004 -1158
rect 9038 -1192 9072 -1158
rect 9198 -1192 9232 -1158
rect 9266 -1192 9300 -1158
rect 9770 -1092 9804 -1058
rect 9838 -1092 9872 -1058
rect 9998 -1092 10032 -1058
rect 10066 -1092 10100 -1058
rect 10570 -992 10604 -958
rect 10638 -992 10672 -958
rect 10798 -992 10832 -958
rect 10866 -992 10900 -958
rect 11370 -892 11404 -858
rect 11438 -892 11472 -858
rect 11598 -892 11632 -858
rect 11666 -892 11700 -858
rect 11770 -892 11804 -858
rect 11838 -892 11872 -858
rect 11998 -892 12032 -858
rect 12066 -892 12100 -858
rect 10970 -992 11004 -958
rect 11038 -992 11072 -958
rect 11198 -992 11232 -958
rect 11266 -992 11300 -958
rect 10170 -1092 10204 -1058
rect 10238 -1092 10272 -1058
rect 10398 -1092 10432 -1058
rect 10466 -1092 10500 -1058
rect 9370 -1192 9404 -1158
rect 9438 -1192 9472 -1158
rect 9598 -1192 9632 -1158
rect 9666 -1192 9700 -1158
rect 8570 -1292 8604 -1258
rect 8638 -1292 8672 -1258
rect 8798 -1292 8832 -1258
rect 8866 -1292 8900 -1258
rect 7770 -1392 7804 -1358
rect 7838 -1392 7872 -1358
rect 7998 -1392 8032 -1358
rect 8066 -1392 8100 -1358
rect 6970 -1492 7004 -1458
rect 7038 -1492 7072 -1458
rect 7198 -1492 7232 -1458
rect 7266 -1492 7300 -1458
rect 6170 -1592 6204 -1558
rect 6238 -1592 6272 -1558
rect 6398 -1592 6432 -1558
rect 6466 -1592 6500 -1558
rect 5370 -1692 5404 -1658
rect 5438 -1692 5472 -1658
rect 5598 -1692 5632 -1658
rect 5666 -1692 5700 -1658
rect 4570 -1792 4604 -1758
rect 4638 -1792 4672 -1758
rect 4798 -1792 4832 -1758
rect 4866 -1792 4900 -1758
rect 3770 -1892 3804 -1858
rect 3838 -1892 3872 -1858
rect 3998 -1892 4032 -1858
rect 4066 -1892 4100 -1858
rect 2970 -1992 3004 -1958
rect 3038 -1992 3072 -1958
rect 3198 -1992 3232 -1958
rect 3266 -1992 3300 -1958
rect 2170 -2092 2204 -2058
rect 2238 -2092 2272 -2058
rect 2398 -2092 2432 -2058
rect 2466 -2092 2500 -2058
rect 2570 -2092 2604 -2058
rect 2638 -2092 2672 -2058
rect 2798 -2092 2832 -2058
rect 2866 -2092 2900 -2058
rect 3370 -1992 3404 -1958
rect 3438 -1992 3472 -1958
rect 3598 -1992 3632 -1958
rect 3666 -1992 3700 -1958
rect 4170 -1892 4204 -1858
rect 4238 -1892 4272 -1858
rect 4398 -1892 4432 -1858
rect 4466 -1892 4500 -1858
rect 4970 -1792 5004 -1758
rect 5038 -1792 5072 -1758
rect 5198 -1792 5232 -1758
rect 5266 -1792 5300 -1758
rect 5770 -1692 5804 -1658
rect 5838 -1692 5872 -1658
rect 5998 -1692 6032 -1658
rect 6066 -1692 6100 -1658
rect 6570 -1592 6604 -1558
rect 6638 -1592 6672 -1558
rect 6798 -1592 6832 -1558
rect 6866 -1592 6900 -1558
rect 7370 -1492 7404 -1458
rect 7438 -1492 7472 -1458
rect 7598 -1492 7632 -1458
rect 7666 -1492 7700 -1458
rect 8170 -1392 8204 -1358
rect 8238 -1392 8272 -1358
rect 8398 -1392 8432 -1358
rect 8466 -1392 8500 -1358
rect 8970 -1292 9004 -1258
rect 9038 -1292 9072 -1258
rect 9198 -1292 9232 -1258
rect 9266 -1292 9300 -1258
rect 9770 -1192 9804 -1158
rect 9838 -1192 9872 -1158
rect 9998 -1192 10032 -1158
rect 10066 -1192 10100 -1158
rect 10570 -1092 10604 -1058
rect 10638 -1092 10672 -1058
rect 10798 -1092 10832 -1058
rect 10866 -1092 10900 -1058
rect 11370 -992 11404 -958
rect 11438 -992 11472 -958
rect 11598 -992 11632 -958
rect 11666 -992 11700 -958
rect 12170 -892 12204 -858
rect 12238 -892 12272 -858
rect 12398 -892 12432 -858
rect 12466 -892 12500 -858
rect 12570 -892 12604 -858
rect 12638 -892 12672 -858
rect 15678 -842 15712 -808
rect 15746 -842 15780 -808
rect 11770 -992 11804 -958
rect 11838 -992 11872 -958
rect 11998 -992 12032 -958
rect 12066 -992 12100 -958
rect 10970 -1092 11004 -1058
rect 11038 -1092 11072 -1058
rect 11198 -1092 11232 -1058
rect 11266 -1092 11300 -1058
rect 10170 -1192 10204 -1158
rect 10238 -1192 10272 -1158
rect 10398 -1192 10432 -1158
rect 10466 -1192 10500 -1158
rect 9370 -1292 9404 -1258
rect 9438 -1292 9472 -1258
rect 9598 -1292 9632 -1258
rect 9666 -1292 9700 -1258
rect 8570 -1392 8604 -1358
rect 8638 -1392 8672 -1358
rect 8798 -1392 8832 -1358
rect 8866 -1392 8900 -1358
rect 7770 -1492 7804 -1458
rect 7838 -1492 7872 -1458
rect 7998 -1492 8032 -1458
rect 8066 -1492 8100 -1458
rect 6970 -1592 7004 -1558
rect 7038 -1592 7072 -1558
rect 7198 -1592 7232 -1558
rect 7266 -1592 7300 -1558
rect 6170 -1692 6204 -1658
rect 6238 -1692 6272 -1658
rect 6398 -1692 6432 -1658
rect 6466 -1692 6500 -1658
rect 5370 -1792 5404 -1758
rect 5438 -1792 5472 -1758
rect 5598 -1792 5632 -1758
rect 5666 -1792 5700 -1758
rect 4570 -1892 4604 -1858
rect 4638 -1892 4672 -1858
rect 4798 -1892 4832 -1858
rect 4866 -1892 4900 -1858
rect 3770 -1992 3804 -1958
rect 3838 -1992 3872 -1958
rect 3998 -1992 4032 -1958
rect 4066 -1992 4100 -1958
rect 2970 -2092 3004 -2058
rect 3038 -2092 3072 -2058
rect 3198 -2092 3232 -2058
rect 3266 -2092 3300 -2058
rect 3370 -2092 3404 -2058
rect 3438 -2092 3472 -2058
rect 3598 -2092 3632 -2058
rect 3666 -2092 3700 -2058
rect 4170 -1992 4204 -1958
rect 4238 -1992 4272 -1958
rect 4398 -1992 4432 -1958
rect 4466 -1992 4500 -1958
rect 4970 -1892 5004 -1858
rect 5038 -1892 5072 -1858
rect 5198 -1892 5232 -1858
rect 5266 -1892 5300 -1858
rect 5770 -1792 5804 -1758
rect 5838 -1792 5872 -1758
rect 5998 -1792 6032 -1758
rect 6066 -1792 6100 -1758
rect 6570 -1692 6604 -1658
rect 6638 -1692 6672 -1658
rect 6798 -1692 6832 -1658
rect 6866 -1692 6900 -1658
rect 7370 -1592 7404 -1558
rect 7438 -1592 7472 -1558
rect 7598 -1592 7632 -1558
rect 7666 -1592 7700 -1558
rect 8170 -1492 8204 -1458
rect 8238 -1492 8272 -1458
rect 8398 -1492 8432 -1458
rect 8466 -1492 8500 -1458
rect 8970 -1392 9004 -1358
rect 9038 -1392 9072 -1358
rect 9198 -1392 9232 -1358
rect 9266 -1392 9300 -1358
rect 9770 -1292 9804 -1258
rect 9838 -1292 9872 -1258
rect 9998 -1292 10032 -1258
rect 10066 -1292 10100 -1258
rect 10570 -1192 10604 -1158
rect 10638 -1192 10672 -1158
rect 10798 -1192 10832 -1158
rect 10866 -1192 10900 -1158
rect 11370 -1092 11404 -1058
rect 11438 -1092 11472 -1058
rect 11598 -1092 11632 -1058
rect 11666 -1092 11700 -1058
rect 12170 -992 12204 -958
rect 12238 -992 12272 -958
rect 12398 -992 12432 -958
rect 12466 -992 12500 -958
rect 14562 -942 14596 -908
rect 14630 -942 14664 -908
rect 12570 -992 12604 -958
rect 12638 -992 12672 -958
rect 15678 -942 15712 -908
rect 15746 -942 15780 -908
rect 11770 -1092 11804 -1058
rect 11838 -1092 11872 -1058
rect 11998 -1092 12032 -1058
rect 12066 -1092 12100 -1058
rect 10970 -1192 11004 -1158
rect 11038 -1192 11072 -1158
rect 11198 -1192 11232 -1158
rect 11266 -1192 11300 -1158
rect 10170 -1292 10204 -1258
rect 10238 -1292 10272 -1258
rect 10398 -1292 10432 -1258
rect 10466 -1292 10500 -1258
rect 9370 -1392 9404 -1358
rect 9438 -1392 9472 -1358
rect 9598 -1392 9632 -1358
rect 9666 -1392 9700 -1358
rect 8570 -1492 8604 -1458
rect 8638 -1492 8672 -1458
rect 8798 -1492 8832 -1458
rect 8866 -1492 8900 -1458
rect 7770 -1592 7804 -1558
rect 7838 -1592 7872 -1558
rect 7998 -1592 8032 -1558
rect 8066 -1592 8100 -1558
rect 6970 -1692 7004 -1658
rect 7038 -1692 7072 -1658
rect 7198 -1692 7232 -1658
rect 7266 -1692 7300 -1658
rect 6170 -1792 6204 -1758
rect 6238 -1792 6272 -1758
rect 6398 -1792 6432 -1758
rect 6466 -1792 6500 -1758
rect 5370 -1892 5404 -1858
rect 5438 -1892 5472 -1858
rect 5598 -1892 5632 -1858
rect 5666 -1892 5700 -1858
rect 4570 -1992 4604 -1958
rect 4638 -1992 4672 -1958
rect 4798 -1992 4832 -1958
rect 4866 -1992 4900 -1958
rect 3770 -2092 3804 -2058
rect 3838 -2092 3872 -2058
rect 3998 -2092 4032 -2058
rect 4066 -2092 4100 -2058
rect 4170 -2092 4204 -2058
rect 4238 -2092 4272 -2058
rect 4398 -2092 4432 -2058
rect 4466 -2092 4500 -2058
rect 4970 -1992 5004 -1958
rect 5038 -1992 5072 -1958
rect 5198 -1992 5232 -1958
rect 5266 -1992 5300 -1958
rect 5770 -1892 5804 -1858
rect 5838 -1892 5872 -1858
rect 5998 -1892 6032 -1858
rect 6066 -1892 6100 -1858
rect 6570 -1792 6604 -1758
rect 6638 -1792 6672 -1758
rect 6798 -1792 6832 -1758
rect 6866 -1792 6900 -1758
rect 7370 -1692 7404 -1658
rect 7438 -1692 7472 -1658
rect 7598 -1692 7632 -1658
rect 7666 -1692 7700 -1658
rect 8170 -1592 8204 -1558
rect 8238 -1592 8272 -1558
rect 8398 -1592 8432 -1558
rect 8466 -1592 8500 -1558
rect 8970 -1492 9004 -1458
rect 9038 -1492 9072 -1458
rect 9198 -1492 9232 -1458
rect 9266 -1492 9300 -1458
rect 9770 -1392 9804 -1358
rect 9838 -1392 9872 -1358
rect 9998 -1392 10032 -1358
rect 10066 -1392 10100 -1358
rect 10570 -1292 10604 -1258
rect 10638 -1292 10672 -1258
rect 10798 -1292 10832 -1258
rect 10866 -1292 10900 -1258
rect 11370 -1192 11404 -1158
rect 11438 -1192 11472 -1158
rect 11598 -1192 11632 -1158
rect 11666 -1192 11700 -1158
rect 12170 -1092 12204 -1058
rect 12238 -1092 12272 -1058
rect 12398 -1092 12432 -1058
rect 12466 -1092 12500 -1058
rect 14562 -1042 14596 -1008
rect 14630 -1042 14664 -1008
rect 12570 -1092 12604 -1058
rect 12638 -1092 12672 -1058
rect 15678 -1042 15712 -1008
rect 15746 -1042 15780 -1008
rect 11770 -1192 11804 -1158
rect 11838 -1192 11872 -1158
rect 11998 -1192 12032 -1158
rect 12066 -1192 12100 -1158
rect 10970 -1292 11004 -1258
rect 11038 -1292 11072 -1258
rect 11198 -1292 11232 -1258
rect 11266 -1292 11300 -1258
rect 10170 -1392 10204 -1358
rect 10238 -1392 10272 -1358
rect 10398 -1392 10432 -1358
rect 10466 -1392 10500 -1358
rect 9370 -1492 9404 -1458
rect 9438 -1492 9472 -1458
rect 9598 -1492 9632 -1458
rect 9666 -1492 9700 -1458
rect 8570 -1592 8604 -1558
rect 8638 -1592 8672 -1558
rect 8798 -1592 8832 -1558
rect 8866 -1592 8900 -1558
rect 7770 -1692 7804 -1658
rect 7838 -1692 7872 -1658
rect 7998 -1692 8032 -1658
rect 8066 -1692 8100 -1658
rect 6970 -1792 7004 -1758
rect 7038 -1792 7072 -1758
rect 7198 -1792 7232 -1758
rect 7266 -1792 7300 -1758
rect 6170 -1892 6204 -1858
rect 6238 -1892 6272 -1858
rect 6398 -1892 6432 -1858
rect 6466 -1892 6500 -1858
rect 5370 -1992 5404 -1958
rect 5438 -1992 5472 -1958
rect 5598 -1992 5632 -1958
rect 5666 -1992 5700 -1958
rect 4570 -2092 4604 -2058
rect 4638 -2092 4672 -2058
rect 4798 -2092 4832 -2058
rect 4866 -2092 4900 -2058
rect 4970 -2092 5004 -2058
rect 5038 -2092 5072 -2058
rect 5198 -2092 5232 -2058
rect 5266 -2092 5300 -2058
rect 5770 -1992 5804 -1958
rect 5838 -1992 5872 -1958
rect 5998 -1992 6032 -1958
rect 6066 -1992 6100 -1958
rect 6570 -1892 6604 -1858
rect 6638 -1892 6672 -1858
rect 6798 -1892 6832 -1858
rect 6866 -1892 6900 -1858
rect 7370 -1792 7404 -1758
rect 7438 -1792 7472 -1758
rect 7598 -1792 7632 -1758
rect 7666 -1792 7700 -1758
rect 8170 -1692 8204 -1658
rect 8238 -1692 8272 -1658
rect 8398 -1692 8432 -1658
rect 8466 -1692 8500 -1658
rect 8970 -1592 9004 -1558
rect 9038 -1592 9072 -1558
rect 9198 -1592 9232 -1558
rect 9266 -1592 9300 -1558
rect 9770 -1492 9804 -1458
rect 9838 -1492 9872 -1458
rect 9998 -1492 10032 -1458
rect 10066 -1492 10100 -1458
rect 10570 -1392 10604 -1358
rect 10638 -1392 10672 -1358
rect 10798 -1392 10832 -1358
rect 10866 -1392 10900 -1358
rect 11370 -1292 11404 -1258
rect 11438 -1292 11472 -1258
rect 11598 -1292 11632 -1258
rect 11666 -1292 11700 -1258
rect 12170 -1192 12204 -1158
rect 12238 -1192 12272 -1158
rect 12398 -1192 12432 -1158
rect 12466 -1192 12500 -1158
rect 14562 -1142 14596 -1108
rect 14630 -1142 14664 -1108
rect 12570 -1192 12604 -1158
rect 12638 -1192 12672 -1158
rect 15678 -1142 15712 -1108
rect 15746 -1142 15780 -1108
rect 11770 -1292 11804 -1258
rect 11838 -1292 11872 -1258
rect 11998 -1292 12032 -1258
rect 12066 -1292 12100 -1258
rect 10970 -1392 11004 -1358
rect 11038 -1392 11072 -1358
rect 11198 -1392 11232 -1358
rect 11266 -1392 11300 -1358
rect 10170 -1492 10204 -1458
rect 10238 -1492 10272 -1458
rect 10398 -1492 10432 -1458
rect 10466 -1492 10500 -1458
rect 9370 -1592 9404 -1558
rect 9438 -1592 9472 -1558
rect 9598 -1592 9632 -1558
rect 9666 -1592 9700 -1558
rect 8570 -1692 8604 -1658
rect 8638 -1692 8672 -1658
rect 8798 -1692 8832 -1658
rect 8866 -1692 8900 -1658
rect 7770 -1792 7804 -1758
rect 7838 -1792 7872 -1758
rect 7998 -1792 8032 -1758
rect 8066 -1792 8100 -1758
rect 6970 -1892 7004 -1858
rect 7038 -1892 7072 -1858
rect 7198 -1892 7232 -1858
rect 7266 -1892 7300 -1858
rect 6170 -1992 6204 -1958
rect 6238 -1992 6272 -1958
rect 6398 -1992 6432 -1958
rect 6466 -1992 6500 -1958
rect 5370 -2092 5404 -2058
rect 5438 -2092 5472 -2058
rect 5598 -2092 5632 -2058
rect 5666 -2092 5700 -2058
rect 5770 -2092 5804 -2058
rect 5838 -2092 5872 -2058
rect 5998 -2092 6032 -2058
rect 6066 -2092 6100 -2058
rect 6570 -1992 6604 -1958
rect 6638 -1992 6672 -1958
rect 6798 -1992 6832 -1958
rect 6866 -1992 6900 -1958
rect 7370 -1892 7404 -1858
rect 7438 -1892 7472 -1858
rect 7598 -1892 7632 -1858
rect 7666 -1892 7700 -1858
rect 8170 -1792 8204 -1758
rect 8238 -1792 8272 -1758
rect 8398 -1792 8432 -1758
rect 8466 -1792 8500 -1758
rect 8970 -1692 9004 -1658
rect 9038 -1692 9072 -1658
rect 9198 -1692 9232 -1658
rect 9266 -1692 9300 -1658
rect 9770 -1592 9804 -1558
rect 9838 -1592 9872 -1558
rect 9998 -1592 10032 -1558
rect 10066 -1592 10100 -1558
rect 10570 -1492 10604 -1458
rect 10638 -1492 10672 -1458
rect 10798 -1492 10832 -1458
rect 10866 -1492 10900 -1458
rect 11370 -1392 11404 -1358
rect 11438 -1392 11472 -1358
rect 11598 -1392 11632 -1358
rect 11666 -1392 11700 -1358
rect 12170 -1292 12204 -1258
rect 12238 -1292 12272 -1258
rect 12398 -1292 12432 -1258
rect 12466 -1292 12500 -1258
rect 14562 -1242 14596 -1208
rect 14630 -1242 14664 -1208
rect 12570 -1292 12604 -1258
rect 12638 -1292 12672 -1258
rect 15678 -1242 15712 -1208
rect 15746 -1242 15780 -1208
rect 11770 -1392 11804 -1358
rect 11838 -1392 11872 -1358
rect 11998 -1392 12032 -1358
rect 12066 -1392 12100 -1358
rect 10970 -1492 11004 -1458
rect 11038 -1492 11072 -1458
rect 11198 -1492 11232 -1458
rect 11266 -1492 11300 -1458
rect 10170 -1592 10204 -1558
rect 10238 -1592 10272 -1558
rect 10398 -1592 10432 -1558
rect 10466 -1592 10500 -1558
rect 9370 -1692 9404 -1658
rect 9438 -1692 9472 -1658
rect 9598 -1692 9632 -1658
rect 9666 -1692 9700 -1658
rect 8570 -1792 8604 -1758
rect 8638 -1792 8672 -1758
rect 8798 -1792 8832 -1758
rect 8866 -1792 8900 -1758
rect 7770 -1892 7804 -1858
rect 7838 -1892 7872 -1858
rect 7998 -1892 8032 -1858
rect 8066 -1892 8100 -1858
rect 6970 -1992 7004 -1958
rect 7038 -1992 7072 -1958
rect 7198 -1992 7232 -1958
rect 7266 -1992 7300 -1958
rect 6170 -2092 6204 -2058
rect 6238 -2092 6272 -2058
rect 6398 -2092 6432 -2058
rect 6466 -2092 6500 -2058
rect 6570 -2092 6604 -2058
rect 6638 -2092 6672 -2058
rect 6798 -2092 6832 -2058
rect 6866 -2092 6900 -2058
rect 7370 -1992 7404 -1958
rect 7438 -1992 7472 -1958
rect 7598 -1992 7632 -1958
rect 7666 -1992 7700 -1958
rect 8170 -1892 8204 -1858
rect 8238 -1892 8272 -1858
rect 8398 -1892 8432 -1858
rect 8466 -1892 8500 -1858
rect 8970 -1792 9004 -1758
rect 9038 -1792 9072 -1758
rect 9198 -1792 9232 -1758
rect 9266 -1792 9300 -1758
rect 9770 -1692 9804 -1658
rect 9838 -1692 9872 -1658
rect 9998 -1692 10032 -1658
rect 10066 -1692 10100 -1658
rect 10570 -1592 10604 -1558
rect 10638 -1592 10672 -1558
rect 10798 -1592 10832 -1558
rect 10866 -1592 10900 -1558
rect 11370 -1492 11404 -1458
rect 11438 -1492 11472 -1458
rect 11598 -1492 11632 -1458
rect 11666 -1492 11700 -1458
rect 12170 -1392 12204 -1358
rect 12238 -1392 12272 -1358
rect 12398 -1392 12432 -1358
rect 12466 -1392 12500 -1358
rect 14562 -1342 14596 -1308
rect 14630 -1342 14664 -1308
rect 12570 -1392 12604 -1358
rect 12638 -1392 12672 -1358
rect 15678 -1342 15712 -1308
rect 15746 -1342 15780 -1308
rect 11770 -1492 11804 -1458
rect 11838 -1492 11872 -1458
rect 11998 -1492 12032 -1458
rect 12066 -1492 12100 -1458
rect 10970 -1592 11004 -1558
rect 11038 -1592 11072 -1558
rect 11198 -1592 11232 -1558
rect 11266 -1592 11300 -1558
rect 10170 -1692 10204 -1658
rect 10238 -1692 10272 -1658
rect 10398 -1692 10432 -1658
rect 10466 -1692 10500 -1658
rect 9370 -1792 9404 -1758
rect 9438 -1792 9472 -1758
rect 9598 -1792 9632 -1758
rect 9666 -1792 9700 -1758
rect 8570 -1892 8604 -1858
rect 8638 -1892 8672 -1858
rect 8798 -1892 8832 -1858
rect 8866 -1892 8900 -1858
rect 7770 -1992 7804 -1958
rect 7838 -1992 7872 -1958
rect 7998 -1992 8032 -1958
rect 8066 -1992 8100 -1958
rect 6970 -2092 7004 -2058
rect 7038 -2092 7072 -2058
rect 7198 -2092 7232 -2058
rect 7266 -2092 7300 -2058
rect 7370 -2092 7404 -2058
rect 7438 -2092 7472 -2058
rect 7598 -2092 7632 -2058
rect 7666 -2092 7700 -2058
rect 8170 -1992 8204 -1958
rect 8238 -1992 8272 -1958
rect 8398 -1992 8432 -1958
rect 8466 -1992 8500 -1958
rect 8970 -1892 9004 -1858
rect 9038 -1892 9072 -1858
rect 9198 -1892 9232 -1858
rect 9266 -1892 9300 -1858
rect 9770 -1792 9804 -1758
rect 9838 -1792 9872 -1758
rect 9998 -1792 10032 -1758
rect 10066 -1792 10100 -1758
rect 10570 -1692 10604 -1658
rect 10638 -1692 10672 -1658
rect 10798 -1692 10832 -1658
rect 10866 -1692 10900 -1658
rect 11370 -1592 11404 -1558
rect 11438 -1592 11472 -1558
rect 11598 -1592 11632 -1558
rect 11666 -1592 11700 -1558
rect 12170 -1492 12204 -1458
rect 12238 -1492 12272 -1458
rect 12398 -1492 12432 -1458
rect 12466 -1492 12500 -1458
rect 14562 -1442 14596 -1408
rect 14630 -1442 14664 -1408
rect 12570 -1492 12604 -1458
rect 12638 -1492 12672 -1458
rect 15678 -1442 15712 -1408
rect 15746 -1442 15780 -1408
rect 11770 -1592 11804 -1558
rect 11838 -1592 11872 -1558
rect 11998 -1592 12032 -1558
rect 12066 -1592 12100 -1558
rect 10970 -1692 11004 -1658
rect 11038 -1692 11072 -1658
rect 11198 -1692 11232 -1658
rect 11266 -1692 11300 -1658
rect 10170 -1792 10204 -1758
rect 10238 -1792 10272 -1758
rect 10398 -1792 10432 -1758
rect 10466 -1792 10500 -1758
rect 9370 -1892 9404 -1858
rect 9438 -1892 9472 -1858
rect 9598 -1892 9632 -1858
rect 9666 -1892 9700 -1858
rect 8570 -1992 8604 -1958
rect 8638 -1992 8672 -1958
rect 8798 -1992 8832 -1958
rect 8866 -1992 8900 -1958
rect 7770 -2092 7804 -2058
rect 7838 -2092 7872 -2058
rect 7998 -2092 8032 -2058
rect 8066 -2092 8100 -2058
rect 8170 -2092 8204 -2058
rect 8238 -2092 8272 -2058
rect 8398 -2092 8432 -2058
rect 8466 -2092 8500 -2058
rect 8970 -1992 9004 -1958
rect 9038 -1992 9072 -1958
rect 9198 -1992 9232 -1958
rect 9266 -1992 9300 -1958
rect 9770 -1892 9804 -1858
rect 9838 -1892 9872 -1858
rect 9998 -1892 10032 -1858
rect 10066 -1892 10100 -1858
rect 10570 -1792 10604 -1758
rect 10638 -1792 10672 -1758
rect 10798 -1792 10832 -1758
rect 10866 -1792 10900 -1758
rect 11370 -1692 11404 -1658
rect 11438 -1692 11472 -1658
rect 11598 -1692 11632 -1658
rect 11666 -1692 11700 -1658
rect 12170 -1592 12204 -1558
rect 12238 -1592 12272 -1558
rect 12398 -1592 12432 -1558
rect 12466 -1592 12500 -1558
rect 14562 -1542 14596 -1508
rect 14630 -1542 14664 -1508
rect 12570 -1592 12604 -1558
rect 12638 -1592 12672 -1558
rect 15678 -1542 15712 -1508
rect 15746 -1542 15780 -1508
rect 11770 -1692 11804 -1658
rect 11838 -1692 11872 -1658
rect 11998 -1692 12032 -1658
rect 12066 -1692 12100 -1658
rect 10970 -1792 11004 -1758
rect 11038 -1792 11072 -1758
rect 11198 -1792 11232 -1758
rect 11266 -1792 11300 -1758
rect 10170 -1892 10204 -1858
rect 10238 -1892 10272 -1858
rect 10398 -1892 10432 -1858
rect 10466 -1892 10500 -1858
rect 9370 -1992 9404 -1958
rect 9438 -1992 9472 -1958
rect 9598 -1992 9632 -1958
rect 9666 -1992 9700 -1958
rect 8570 -2092 8604 -2058
rect 8638 -2092 8672 -2058
rect 8798 -2092 8832 -2058
rect 8866 -2092 8900 -2058
rect 8970 -2092 9004 -2058
rect 9038 -2092 9072 -2058
rect 9198 -2092 9232 -2058
rect 9266 -2092 9300 -2058
rect 9770 -1992 9804 -1958
rect 9838 -1992 9872 -1958
rect 9998 -1992 10032 -1958
rect 10066 -1992 10100 -1958
rect 10570 -1892 10604 -1858
rect 10638 -1892 10672 -1858
rect 10798 -1892 10832 -1858
rect 10866 -1892 10900 -1858
rect 11370 -1792 11404 -1758
rect 11438 -1792 11472 -1758
rect 11598 -1792 11632 -1758
rect 11666 -1792 11700 -1758
rect 12170 -1692 12204 -1658
rect 12238 -1692 12272 -1658
rect 12398 -1692 12432 -1658
rect 12466 -1692 12500 -1658
rect 14562 -1642 14596 -1608
rect 14630 -1642 14664 -1608
rect 12570 -1692 12604 -1658
rect 12638 -1692 12672 -1658
rect 15678 -1642 15712 -1608
rect 15746 -1642 15780 -1608
rect 11770 -1792 11804 -1758
rect 11838 -1792 11872 -1758
rect 11998 -1792 12032 -1758
rect 12066 -1792 12100 -1758
rect 10970 -1892 11004 -1858
rect 11038 -1892 11072 -1858
rect 11198 -1892 11232 -1858
rect 11266 -1892 11300 -1858
rect 10170 -1992 10204 -1958
rect 10238 -1992 10272 -1958
rect 10398 -1992 10432 -1958
rect 10466 -1992 10500 -1958
rect 9370 -2092 9404 -2058
rect 9438 -2092 9472 -2058
rect 9598 -2092 9632 -2058
rect 9666 -2092 9700 -2058
rect 9770 -2092 9804 -2058
rect 9838 -2092 9872 -2058
rect 9998 -2092 10032 -2058
rect 10066 -2092 10100 -2058
rect 10570 -1992 10604 -1958
rect 10638 -1992 10672 -1958
rect 10798 -1992 10832 -1958
rect 10866 -1992 10900 -1958
rect 11370 -1892 11404 -1858
rect 11438 -1892 11472 -1858
rect 11598 -1892 11632 -1858
rect 11666 -1892 11700 -1858
rect 12170 -1792 12204 -1758
rect 12238 -1792 12272 -1758
rect 12398 -1792 12432 -1758
rect 12466 -1792 12500 -1758
rect 14562 -1742 14596 -1708
rect 14630 -1742 14664 -1708
rect 12570 -1792 12604 -1758
rect 12638 -1792 12672 -1758
rect 15678 -1742 15712 -1708
rect 15746 -1742 15780 -1708
rect 11770 -1892 11804 -1858
rect 11838 -1892 11872 -1858
rect 11998 -1892 12032 -1858
rect 12066 -1892 12100 -1858
rect 10970 -1992 11004 -1958
rect 11038 -1992 11072 -1958
rect 11198 -1992 11232 -1958
rect 11266 -1992 11300 -1958
rect 10170 -2092 10204 -2058
rect 10238 -2092 10272 -2058
rect 10398 -2092 10432 -2058
rect 10466 -2092 10500 -2058
rect 10570 -2092 10604 -2058
rect 10638 -2092 10672 -2058
rect 10798 -2092 10832 -2058
rect 10866 -2092 10900 -2058
rect 11370 -1992 11404 -1958
rect 11438 -1992 11472 -1958
rect 11598 -1992 11632 -1958
rect 11666 -1992 11700 -1958
rect 12170 -1892 12204 -1858
rect 12238 -1892 12272 -1858
rect 12398 -1892 12432 -1858
rect 12466 -1892 12500 -1858
rect 14562 -1842 14596 -1808
rect 14630 -1842 14664 -1808
rect 12570 -1892 12604 -1858
rect 12638 -1892 12672 -1858
rect 15678 -1842 15712 -1808
rect 15746 -1842 15780 -1808
rect 11770 -1992 11804 -1958
rect 11838 -1992 11872 -1958
rect 11998 -1992 12032 -1958
rect 12066 -1992 12100 -1958
rect 10970 -2092 11004 -2058
rect 11038 -2092 11072 -2058
rect 11198 -2092 11232 -2058
rect 11266 -2092 11300 -2058
rect 11370 -2092 11404 -2058
rect 11438 -2092 11472 -2058
rect 11598 -2092 11632 -2058
rect 11666 -2092 11700 -2058
rect 12170 -1992 12204 -1958
rect 12238 -1992 12272 -1958
rect 12398 -1992 12432 -1958
rect 12466 -1992 12500 -1958
rect 14562 -1942 14596 -1908
rect 14630 -1942 14664 -1908
rect 12570 -1992 12604 -1958
rect 12638 -1992 12672 -1958
rect 15678 -1942 15712 -1908
rect 15746 -1942 15780 -1908
rect 11770 -2092 11804 -2058
rect 11838 -2092 11872 -2058
rect 11998 -2092 12032 -2058
rect 12066 -2092 12100 -2058
rect 12170 -2092 12204 -2058
rect 12238 -2092 12272 -2058
rect 12398 -2092 12432 -2058
rect 12466 -2092 12500 -2058
rect 14562 -2042 14596 -2008
rect 14630 -2042 14664 -2008
rect 12570 -2092 12604 -2058
rect 12638 -2092 12672 -2058
rect 15678 -2042 15712 -2008
rect 15746 -2042 15780 -2008
<< pdiffc >>
rect 14847 -242 14881 -208
rect 14915 -242 14949 -208
rect 14983 -242 15017 -208
rect 15051 -242 15085 -208
rect 15257 -242 15291 -208
rect 15325 -242 15359 -208
rect 15393 -242 15427 -208
rect 15461 -242 15495 -208
rect -82 -397 -48 -363
rect -82 -465 -48 -431
rect 18 -397 52 -363
rect 18 -465 52 -431
rect 118 -397 152 -363
rect 118 -465 152 -431
rect 218 -397 252 -363
rect 218 -465 252 -431
rect 318 -397 352 -363
rect 318 -465 352 -431
rect 418 -397 452 -363
rect 418 -465 452 -431
rect 518 -397 552 -363
rect 518 -465 552 -431
rect 618 -397 652 -363
rect 618 -465 652 -431
rect 718 -397 752 -363
rect 718 -465 752 -431
rect 818 -397 852 -363
rect 818 -465 852 -431
rect 918 -397 952 -363
rect 918 -465 952 -431
rect 1018 -397 1052 -363
rect 1018 -465 1052 -431
rect 1118 -397 1152 -363
rect 1118 -465 1152 -431
rect 1218 -397 1252 -363
rect 1218 -465 1252 -431
rect 1318 -397 1352 -363
rect 1318 -465 1352 -431
rect 1418 -397 1452 -363
rect 1418 -465 1452 -431
rect 1518 -397 1552 -363
rect 1518 -465 1552 -431
rect 1618 -397 1652 -363
rect 1618 -465 1652 -431
rect 1718 -397 1752 -363
rect 1718 -465 1752 -431
rect 1818 -397 1852 -363
rect 1818 -465 1852 -431
rect 1918 -397 1952 -363
rect 1918 -465 1952 -431
rect 2018 -397 2052 -363
rect 2018 -465 2052 -431
rect 2118 -397 2152 -363
rect 2118 -465 2152 -431
rect 2218 -397 2252 -363
rect 2218 -465 2252 -431
rect 2318 -397 2352 -363
rect 2318 -465 2352 -431
rect 2418 -397 2452 -363
rect 2418 -465 2452 -431
rect 2518 -397 2552 -363
rect 2518 -465 2552 -431
rect 2618 -397 2652 -363
rect 2618 -465 2652 -431
rect 2718 -397 2752 -363
rect 2718 -465 2752 -431
rect 2818 -397 2852 -363
rect 2818 -465 2852 -431
rect 2918 -397 2952 -363
rect 2918 -465 2952 -431
rect 3018 -397 3052 -363
rect 3018 -465 3052 -431
rect 3118 -397 3152 -363
rect 3118 -465 3152 -431
rect 3218 -397 3252 -363
rect 3218 -465 3252 -431
rect 3318 -397 3352 -363
rect 3318 -465 3352 -431
rect 3418 -397 3452 -363
rect 3418 -465 3452 -431
rect 3518 -397 3552 -363
rect 3518 -465 3552 -431
rect 3618 -397 3652 -363
rect 3618 -465 3652 -431
rect 3718 -397 3752 -363
rect 3718 -465 3752 -431
rect 3818 -397 3852 -363
rect 3818 -465 3852 -431
rect 3918 -397 3952 -363
rect 3918 -465 3952 -431
rect 4018 -397 4052 -363
rect 4018 -465 4052 -431
rect 4118 -397 4152 -363
rect 4118 -465 4152 -431
rect 4218 -397 4252 -363
rect 4218 -465 4252 -431
rect 4318 -397 4352 -363
rect 4318 -465 4352 -431
rect 4418 -397 4452 -363
rect 4418 -465 4452 -431
rect 4518 -397 4552 -363
rect 4518 -465 4552 -431
rect 4618 -397 4652 -363
rect 4618 -465 4652 -431
rect 4718 -397 4752 -363
rect 4718 -465 4752 -431
rect 4818 -397 4852 -363
rect 4818 -465 4852 -431
rect 4918 -397 4952 -363
rect 4918 -465 4952 -431
rect 5018 -397 5052 -363
rect 5018 -465 5052 -431
rect 5118 -397 5152 -363
rect 5118 -465 5152 -431
rect 5218 -397 5252 -363
rect 5218 -465 5252 -431
rect 5318 -397 5352 -363
rect 5318 -465 5352 -431
rect 5418 -397 5452 -363
rect 5418 -465 5452 -431
rect 5518 -397 5552 -363
rect 5518 -465 5552 -431
rect 5618 -397 5652 -363
rect 5618 -465 5652 -431
rect 5718 -397 5752 -363
rect 5718 -465 5752 -431
rect 5818 -397 5852 -363
rect 5818 -465 5852 -431
rect 5918 -397 5952 -363
rect 5918 -465 5952 -431
rect 6018 -397 6052 -363
rect 6018 -465 6052 -431
rect 6118 -397 6152 -363
rect 6118 -465 6152 -431
rect 6218 -397 6252 -363
rect 6218 -465 6252 -431
rect 6318 -397 6352 -363
rect 6318 -465 6352 -431
rect 6418 -397 6452 -363
rect 6418 -465 6452 -431
rect 6518 -397 6552 -363
rect 6518 -465 6552 -431
rect 6618 -397 6652 -363
rect 6618 -465 6652 -431
rect 6718 -397 6752 -363
rect 6718 -465 6752 -431
rect 6818 -397 6852 -363
rect 6818 -465 6852 -431
rect 6918 -397 6952 -363
rect 6918 -465 6952 -431
rect 7018 -397 7052 -363
rect 7018 -465 7052 -431
rect 7118 -397 7152 -363
rect 7118 -465 7152 -431
rect 7218 -397 7252 -363
rect 7218 -465 7252 -431
rect 7318 -397 7352 -363
rect 7318 -465 7352 -431
rect 7418 -397 7452 -363
rect 7418 -465 7452 -431
rect 7518 -397 7552 -363
rect 7518 -465 7552 -431
rect 7618 -397 7652 -363
rect 7618 -465 7652 -431
rect 7718 -397 7752 -363
rect 7718 -465 7752 -431
rect 7818 -397 7852 -363
rect 7818 -465 7852 -431
rect 7918 -397 7952 -363
rect 7918 -465 7952 -431
rect 8018 -397 8052 -363
rect 8018 -465 8052 -431
rect 8118 -397 8152 -363
rect 8118 -465 8152 -431
rect 8218 -397 8252 -363
rect 8218 -465 8252 -431
rect 8318 -397 8352 -363
rect 8318 -465 8352 -431
rect 8418 -397 8452 -363
rect 8418 -465 8452 -431
rect 8518 -397 8552 -363
rect 8518 -465 8552 -431
rect 8618 -397 8652 -363
rect 8618 -465 8652 -431
rect 8718 -397 8752 -363
rect 8718 -465 8752 -431
rect 8818 -397 8852 -363
rect 8818 -465 8852 -431
rect 8918 -397 8952 -363
rect 8918 -465 8952 -431
rect 9018 -397 9052 -363
rect 9018 -465 9052 -431
rect 9118 -397 9152 -363
rect 9118 -465 9152 -431
rect 9218 -397 9252 -363
rect 9218 -465 9252 -431
rect 9318 -397 9352 -363
rect 9318 -465 9352 -431
rect 9418 -397 9452 -363
rect 9418 -465 9452 -431
rect 9518 -397 9552 -363
rect 9518 -465 9552 -431
rect 9618 -397 9652 -363
rect 9618 -465 9652 -431
rect 9718 -397 9752 -363
rect 9718 -465 9752 -431
rect 9818 -397 9852 -363
rect 9818 -465 9852 -431
rect 9918 -397 9952 -363
rect 9918 -465 9952 -431
rect 10018 -397 10052 -363
rect 10018 -465 10052 -431
rect 10118 -397 10152 -363
rect 10118 -465 10152 -431
rect 10218 -397 10252 -363
rect 10218 -465 10252 -431
rect 10318 -397 10352 -363
rect 10318 -465 10352 -431
rect 10418 -397 10452 -363
rect 10418 -465 10452 -431
rect 10518 -397 10552 -363
rect 10518 -465 10552 -431
rect 10618 -397 10652 -363
rect 10618 -465 10652 -431
rect 10718 -397 10752 -363
rect 10718 -465 10752 -431
rect 10818 -397 10852 -363
rect 10818 -465 10852 -431
rect 10918 -397 10952 -363
rect 10918 -465 10952 -431
rect 11018 -397 11052 -363
rect 11018 -465 11052 -431
rect 11118 -397 11152 -363
rect 11118 -465 11152 -431
rect 11218 -397 11252 -363
rect 11218 -465 11252 -431
rect 11318 -397 11352 -363
rect 11318 -465 11352 -431
rect 11418 -397 11452 -363
rect 11418 -465 11452 -431
rect 11518 -397 11552 -363
rect 11518 -465 11552 -431
rect 11618 -397 11652 -363
rect 11618 -465 11652 -431
rect 11718 -397 11752 -363
rect 11718 -465 11752 -431
rect 11818 -397 11852 -363
rect 11818 -465 11852 -431
rect 11918 -397 11952 -363
rect 11918 -465 11952 -431
rect 12018 -397 12052 -363
rect 12018 -465 12052 -431
rect 12118 -397 12152 -363
rect 12118 -465 12152 -431
rect 12218 -397 12252 -363
rect 12218 -465 12252 -431
rect 12318 -397 12352 -363
rect 12318 -465 12352 -431
rect 12418 -397 12452 -363
rect 12418 -465 12452 -431
rect 12518 -397 12552 -363
rect 12518 -465 12552 -431
rect 12618 -397 12652 -363
rect 12618 -465 12652 -431
rect 14847 -342 14881 -308
rect 14915 -342 14949 -308
rect 14983 -342 15017 -308
rect 15051 -342 15085 -308
rect 15257 -342 15291 -308
rect 15325 -342 15359 -308
rect 15393 -342 15427 -308
rect 15461 -342 15495 -308
rect 12718 -397 12752 -363
rect 12718 -465 12752 -431
rect 14847 -442 14881 -408
rect 14915 -442 14949 -408
rect 14983 -442 15017 -408
rect 15051 -442 15085 -408
rect 15257 -442 15291 -408
rect 15325 -442 15359 -408
rect 15393 -442 15427 -408
rect 15461 -442 15495 -408
rect 14847 -542 14881 -508
rect 14915 -542 14949 -508
rect 14983 -542 15017 -508
rect 15051 -542 15085 -508
rect 15257 -542 15291 -508
rect 15325 -542 15359 -508
rect 15393 -542 15427 -508
rect 15461 -542 15495 -508
rect -30 -717 4 -683
rect 118 -717 152 -683
rect 266 -717 300 -683
rect 370 -717 404 -683
rect 518 -717 552 -683
rect 666 -717 700 -683
rect 770 -717 804 -683
rect 918 -717 952 -683
rect 1066 -717 1100 -683
rect 1170 -717 1204 -683
rect 1318 -717 1352 -683
rect 1466 -717 1500 -683
rect 1570 -717 1604 -683
rect 1718 -717 1752 -683
rect 1866 -717 1900 -683
rect 1970 -717 2004 -683
rect 2118 -717 2152 -683
rect 2266 -717 2300 -683
rect 2370 -717 2404 -683
rect 2518 -717 2552 -683
rect 2666 -717 2700 -683
rect 2770 -717 2804 -683
rect 2918 -717 2952 -683
rect 3066 -717 3100 -683
rect 3170 -717 3204 -683
rect 3318 -717 3352 -683
rect 3466 -717 3500 -683
rect 3570 -717 3604 -683
rect 3718 -717 3752 -683
rect 3866 -717 3900 -683
rect 3970 -717 4004 -683
rect 4118 -717 4152 -683
rect 4266 -717 4300 -683
rect 4370 -717 4404 -683
rect 4518 -717 4552 -683
rect 4666 -717 4700 -683
rect 4770 -717 4804 -683
rect 4918 -717 4952 -683
rect 5066 -717 5100 -683
rect 5170 -717 5204 -683
rect 5318 -717 5352 -683
rect 5466 -717 5500 -683
rect 5570 -717 5604 -683
rect 5718 -717 5752 -683
rect 5866 -717 5900 -683
rect 5970 -717 6004 -683
rect 6118 -717 6152 -683
rect 6266 -717 6300 -683
rect 6370 -717 6404 -683
rect 6518 -717 6552 -683
rect 6666 -717 6700 -683
rect 6770 -717 6804 -683
rect 6918 -717 6952 -683
rect 7066 -717 7100 -683
rect 7170 -717 7204 -683
rect 7318 -717 7352 -683
rect 7466 -717 7500 -683
rect 7570 -717 7604 -683
rect 7718 -717 7752 -683
rect 7866 -717 7900 -683
rect 7970 -717 8004 -683
rect 8118 -717 8152 -683
rect 8266 -717 8300 -683
rect 8370 -717 8404 -683
rect 8518 -717 8552 -683
rect 8666 -717 8700 -683
rect 8770 -717 8804 -683
rect 8918 -717 8952 -683
rect 9066 -717 9100 -683
rect 9170 -717 9204 -683
rect 9318 -717 9352 -683
rect 9466 -717 9500 -683
rect 9570 -717 9604 -683
rect 9718 -717 9752 -683
rect 9866 -717 9900 -683
rect 9970 -717 10004 -683
rect 10118 -717 10152 -683
rect 10266 -717 10300 -683
rect 10370 -717 10404 -683
rect 10518 -717 10552 -683
rect 10666 -717 10700 -683
rect 10770 -717 10804 -683
rect 10918 -717 10952 -683
rect 11066 -717 11100 -683
rect 11170 -717 11204 -683
rect 11318 -717 11352 -683
rect 11466 -717 11500 -683
rect 11570 -717 11604 -683
rect 11718 -717 11752 -683
rect 11866 -717 11900 -683
rect 11970 -717 12004 -683
rect 12118 -717 12152 -683
rect 12266 -717 12300 -683
rect 12370 -717 12404 -683
rect 12518 -717 12552 -683
rect 14847 -642 14881 -608
rect 14915 -642 14949 -608
rect 14983 -642 15017 -608
rect 15051 -642 15085 -608
rect 15257 -642 15291 -608
rect 15325 -642 15359 -608
rect 15393 -642 15427 -608
rect 15461 -642 15495 -608
rect 12666 -717 12700 -683
rect 14847 -742 14881 -708
rect 14915 -742 14949 -708
rect 14983 -742 15017 -708
rect 15051 -742 15085 -708
rect 15257 -742 15291 -708
rect 15325 -742 15359 -708
rect 15393 -742 15427 -708
rect 15461 -742 15495 -708
rect 14847 -842 14881 -808
rect 14915 -842 14949 -808
rect 14983 -842 15017 -808
rect 15051 -842 15085 -808
rect 15257 -842 15291 -808
rect 15325 -842 15359 -808
rect 15393 -842 15427 -808
rect 15461 -842 15495 -808
rect 14847 -942 14881 -908
rect 14915 -942 14949 -908
rect 14983 -942 15017 -908
rect 15051 -942 15085 -908
rect 15257 -942 15291 -908
rect 15325 -942 15359 -908
rect 15393 -942 15427 -908
rect 15461 -942 15495 -908
rect 14847 -1042 14881 -1008
rect 14915 -1042 14949 -1008
rect 14983 -1042 15017 -1008
rect 15051 -1042 15085 -1008
rect 15257 -1042 15291 -1008
rect 15325 -1042 15359 -1008
rect 15393 -1042 15427 -1008
rect 15461 -1042 15495 -1008
rect 14847 -1142 14881 -1108
rect 14915 -1142 14949 -1108
rect 14983 -1142 15017 -1108
rect 15051 -1142 15085 -1108
rect 15257 -1142 15291 -1108
rect 15325 -1142 15359 -1108
rect 15393 -1142 15427 -1108
rect 15461 -1142 15495 -1108
rect 14847 -1242 14881 -1208
rect 14915 -1242 14949 -1208
rect 14983 -1242 15017 -1208
rect 15051 -1242 15085 -1208
rect 15257 -1242 15291 -1208
rect 15325 -1242 15359 -1208
rect 15393 -1242 15427 -1208
rect 15461 -1242 15495 -1208
rect 14847 -1342 14881 -1308
rect 14915 -1342 14949 -1308
rect 14983 -1342 15017 -1308
rect 15051 -1342 15085 -1308
rect 15257 -1342 15291 -1308
rect 15325 -1342 15359 -1308
rect 15393 -1342 15427 -1308
rect 15461 -1342 15495 -1308
rect 14847 -1442 14881 -1408
rect 14915 -1442 14949 -1408
rect 14983 -1442 15017 -1408
rect 15051 -1442 15085 -1408
rect 15257 -1442 15291 -1408
rect 15325 -1442 15359 -1408
rect 15393 -1442 15427 -1408
rect 15461 -1442 15495 -1408
rect 14847 -1542 14881 -1508
rect 14915 -1542 14949 -1508
rect 14983 -1542 15017 -1508
rect 15051 -1542 15085 -1508
rect 15257 -1542 15291 -1508
rect 15325 -1542 15359 -1508
rect 15393 -1542 15427 -1508
rect 15461 -1542 15495 -1508
rect 14847 -1642 14881 -1608
rect 14915 -1642 14949 -1608
rect 14983 -1642 15017 -1608
rect 15051 -1642 15085 -1608
rect 15257 -1642 15291 -1608
rect 15325 -1642 15359 -1608
rect 15393 -1642 15427 -1608
rect 15461 -1642 15495 -1608
rect 14847 -1742 14881 -1708
rect 14915 -1742 14949 -1708
rect 14983 -1742 15017 -1708
rect 15051 -1742 15085 -1708
rect 15257 -1742 15291 -1708
rect 15325 -1742 15359 -1708
rect 15393 -1742 15427 -1708
rect 15461 -1742 15495 -1708
rect 14847 -1842 14881 -1808
rect 14915 -1842 14949 -1808
rect 14983 -1842 15017 -1808
rect 15051 -1842 15085 -1808
rect 15257 -1842 15291 -1808
rect 15325 -1842 15359 -1808
rect 15393 -1842 15427 -1808
rect 15461 -1842 15495 -1808
rect 14847 -1942 14881 -1908
rect 14915 -1942 14949 -1908
rect 14983 -1942 15017 -1908
rect 15051 -1942 15085 -1908
rect 15257 -1942 15291 -1908
rect 15325 -1942 15359 -1908
rect 15393 -1942 15427 -1908
rect 15461 -1942 15495 -1908
rect 14847 -2042 14881 -2008
rect 14915 -2042 14949 -2008
rect 14983 -2042 15017 -2008
rect 15051 -2042 15085 -2008
rect 15257 -2042 15291 -2008
rect 15325 -2042 15359 -2008
rect 15393 -2042 15427 -2008
rect 15461 -2042 15495 -2008
<< psubdiff >>
rect 116 5017 154 5041
rect 116 4983 118 5017
rect 152 4983 154 5017
rect 116 4959 154 4983
rect 316 5017 354 5041
rect 316 4983 318 5017
rect 352 4983 354 5017
rect 316 4959 354 4983
rect 516 5017 554 5041
rect 516 4983 518 5017
rect 552 4983 554 5017
rect 516 4959 554 4983
rect 716 5017 754 5041
rect 716 4983 718 5017
rect 752 4983 754 5017
rect 716 4959 754 4983
rect 916 5017 954 5041
rect 916 4983 918 5017
rect 952 4983 954 5017
rect 916 4959 954 4983
rect 1116 5017 1154 5041
rect 1116 4983 1118 5017
rect 1152 4983 1154 5017
rect 1116 4959 1154 4983
rect 1316 5017 1354 5041
rect 1316 4983 1318 5017
rect 1352 4983 1354 5017
rect 1316 4959 1354 4983
rect 1516 5017 1554 5041
rect 1516 4983 1518 5017
rect 1552 4983 1554 5017
rect 1516 4959 1554 4983
rect 1716 5017 1754 5041
rect 1716 4983 1718 5017
rect 1752 4983 1754 5017
rect 1716 4959 1754 4983
rect 1916 5017 1954 5041
rect 1916 4983 1918 5017
rect 1952 4983 1954 5017
rect 1916 4959 1954 4983
rect 2116 5017 2154 5041
rect 2116 4983 2118 5017
rect 2152 4983 2154 5017
rect 2116 4959 2154 4983
rect 2316 5017 2354 5041
rect 2316 4983 2318 5017
rect 2352 4983 2354 5017
rect 2316 4959 2354 4983
rect 2516 5017 2554 5041
rect 2516 4983 2518 5017
rect 2552 4983 2554 5017
rect 2516 4959 2554 4983
rect 2716 5017 2754 5041
rect 2716 4983 2718 5017
rect 2752 4983 2754 5017
rect 2716 4959 2754 4983
rect 2916 5017 2954 5041
rect 2916 4983 2918 5017
rect 2952 4983 2954 5017
rect 2916 4959 2954 4983
rect 3116 5017 3154 5041
rect 3116 4983 3118 5017
rect 3152 4983 3154 5017
rect 3116 4959 3154 4983
rect 3316 5017 3354 5041
rect 3316 4983 3318 5017
rect 3352 4983 3354 5017
rect 3316 4959 3354 4983
rect 3516 5017 3554 5041
rect 3516 4983 3518 5017
rect 3552 4983 3554 5017
rect 3516 4959 3554 4983
rect 3716 5017 3754 5041
rect 3716 4983 3718 5017
rect 3752 4983 3754 5017
rect 3716 4959 3754 4983
rect 3916 5017 3954 5041
rect 3916 4983 3918 5017
rect 3952 4983 3954 5017
rect 3916 4959 3954 4983
rect 4116 5017 4154 5041
rect 4116 4983 4118 5017
rect 4152 4983 4154 5017
rect 4116 4959 4154 4983
rect 4316 5017 4354 5041
rect 4316 4983 4318 5017
rect 4352 4983 4354 5017
rect 4316 4959 4354 4983
rect 4516 5017 4554 5041
rect 4516 4983 4518 5017
rect 4552 4983 4554 5017
rect 4516 4959 4554 4983
rect 4716 5017 4754 5041
rect 4716 4983 4718 5017
rect 4752 4983 4754 5017
rect 4716 4959 4754 4983
rect 4916 5017 4954 5041
rect 4916 4983 4918 5017
rect 4952 4983 4954 5017
rect 4916 4959 4954 4983
rect 5116 5017 5154 5041
rect 5116 4983 5118 5017
rect 5152 4983 5154 5017
rect 5116 4959 5154 4983
rect 5316 5017 5354 5041
rect 5316 4983 5318 5017
rect 5352 4983 5354 5017
rect 5316 4959 5354 4983
rect 5516 5017 5554 5041
rect 5516 4983 5518 5017
rect 5552 4983 5554 5017
rect 5516 4959 5554 4983
rect 5716 5017 5754 5041
rect 5716 4983 5718 5017
rect 5752 4983 5754 5017
rect 5716 4959 5754 4983
rect 5916 5017 5954 5041
rect 5916 4983 5918 5017
rect 5952 4983 5954 5017
rect 5916 4959 5954 4983
rect 6116 5017 6154 5041
rect 6116 4983 6118 5017
rect 6152 4983 6154 5017
rect 6116 4959 6154 4983
rect 6316 5017 6354 5041
rect 6316 4983 6318 5017
rect 6352 4983 6354 5017
rect 6316 4959 6354 4983
rect 6516 5017 6554 5041
rect 6516 4983 6518 5017
rect 6552 4983 6554 5017
rect 6516 4959 6554 4983
rect 6716 5017 6754 5041
rect 6716 4983 6718 5017
rect 6752 4983 6754 5017
rect 6716 4959 6754 4983
rect 6916 5017 6954 5041
rect 6916 4983 6918 5017
rect 6952 4983 6954 5017
rect 6916 4959 6954 4983
rect 7116 5017 7154 5041
rect 7116 4983 7118 5017
rect 7152 4983 7154 5017
rect 7116 4959 7154 4983
rect 7316 5017 7354 5041
rect 7316 4983 7318 5017
rect 7352 4983 7354 5017
rect 7316 4959 7354 4983
rect 7516 5017 7554 5041
rect 7516 4983 7518 5017
rect 7552 4983 7554 5017
rect 7516 4959 7554 4983
rect 7716 5017 7754 5041
rect 7716 4983 7718 5017
rect 7752 4983 7754 5017
rect 7716 4959 7754 4983
rect 7916 5017 7954 5041
rect 7916 4983 7918 5017
rect 7952 4983 7954 5017
rect 7916 4959 7954 4983
rect 8116 5017 8154 5041
rect 8116 4983 8118 5017
rect 8152 4983 8154 5017
rect 8116 4959 8154 4983
rect 8316 5017 8354 5041
rect 8316 4983 8318 5017
rect 8352 4983 8354 5017
rect 8316 4959 8354 4983
rect 8516 5017 8554 5041
rect 8516 4983 8518 5017
rect 8552 4983 8554 5017
rect 8516 4959 8554 4983
rect 8716 5017 8754 5041
rect 8716 4983 8718 5017
rect 8752 4983 8754 5017
rect 8716 4959 8754 4983
rect 8916 5017 8954 5041
rect 8916 4983 8918 5017
rect 8952 4983 8954 5017
rect 8916 4959 8954 4983
rect 9116 5017 9154 5041
rect 9116 4983 9118 5017
rect 9152 4983 9154 5017
rect 9116 4959 9154 4983
rect 9316 5017 9354 5041
rect 9316 4983 9318 5017
rect 9352 4983 9354 5017
rect 9316 4959 9354 4983
rect 9516 5017 9554 5041
rect 9516 4983 9518 5017
rect 9552 4983 9554 5017
rect 9516 4959 9554 4983
rect 9716 5017 9754 5041
rect 9716 4983 9718 5017
rect 9752 4983 9754 5017
rect 9716 4959 9754 4983
rect 9916 5017 9954 5041
rect 9916 4983 9918 5017
rect 9952 4983 9954 5017
rect 9916 4959 9954 4983
rect 10116 5017 10154 5041
rect 10116 4983 10118 5017
rect 10152 4983 10154 5017
rect 10116 4959 10154 4983
rect 10316 5017 10354 5041
rect 10316 4983 10318 5017
rect 10352 4983 10354 5017
rect 10316 4959 10354 4983
rect 10516 5017 10554 5041
rect 10516 4983 10518 5017
rect 10552 4983 10554 5017
rect 10516 4959 10554 4983
rect 10716 5017 10754 5041
rect 10716 4983 10718 5017
rect 10752 4983 10754 5017
rect 10716 4959 10754 4983
rect 10916 5017 10954 5041
rect 10916 4983 10918 5017
rect 10952 4983 10954 5017
rect 10916 4959 10954 4983
rect 11116 5017 11154 5041
rect 11116 4983 11118 5017
rect 11152 4983 11154 5017
rect 11116 4959 11154 4983
rect 11316 5017 11354 5041
rect 11316 4983 11318 5017
rect 11352 4983 11354 5017
rect 11316 4959 11354 4983
rect 11516 5017 11554 5041
rect 11516 4983 11518 5017
rect 11552 4983 11554 5017
rect 11516 4959 11554 4983
rect 11716 5017 11754 5041
rect 11716 4983 11718 5017
rect 11752 4983 11754 5017
rect 11716 4959 11754 4983
rect 11916 5017 11954 5041
rect 11916 4983 11918 5017
rect 11952 4983 11954 5017
rect 11916 4959 11954 4983
rect 12116 5017 12154 5041
rect 12116 4983 12118 5017
rect 12152 4983 12154 5017
rect 12116 4959 12154 4983
rect 12316 5017 12354 5041
rect 12316 4983 12318 5017
rect 12352 4983 12354 5017
rect 12316 4959 12354 4983
rect 12516 5017 12554 5041
rect 12516 4983 12518 5017
rect 12552 4983 12554 5017
rect 12516 4959 12554 4983
rect 12716 5017 12754 5041
rect 12716 4983 12718 5017
rect 12752 4983 12754 5017
rect 12716 4959 12754 4983
rect -140 -61 -116 -27
rect -82 -61 -48 -27
rect -14 -61 84 -27
rect 118 -61 152 -27
rect 186 -61 284 -27
rect 318 -61 352 -27
rect 386 -61 484 -27
rect 518 -61 552 -27
rect 586 -61 684 -27
rect 718 -61 752 -27
rect 786 -61 884 -27
rect 918 -61 952 -27
rect 986 -61 1084 -27
rect 1118 -61 1152 -27
rect 1186 -61 1284 -27
rect 1318 -61 1352 -27
rect 1386 -61 1484 -27
rect 1518 -61 1552 -27
rect 1586 -61 1684 -27
rect 1718 -61 1752 -27
rect 1786 -61 1884 -27
rect 1918 -61 1952 -27
rect 1986 -61 2084 -27
rect 2118 -61 2152 -27
rect 2186 -61 2284 -27
rect 2318 -61 2352 -27
rect 2386 -61 2484 -27
rect 2518 -61 2552 -27
rect 2586 -61 2684 -27
rect 2718 -61 2752 -27
rect 2786 -61 2884 -27
rect 2918 -61 2952 -27
rect 2986 -61 3084 -27
rect 3118 -61 3152 -27
rect 3186 -61 3284 -27
rect 3318 -61 3352 -27
rect 3386 -61 3484 -27
rect 3518 -61 3552 -27
rect 3586 -61 3684 -27
rect 3718 -61 3752 -27
rect 3786 -61 3884 -27
rect 3918 -61 3952 -27
rect 3986 -61 4084 -27
rect 4118 -61 4152 -27
rect 4186 -61 4284 -27
rect 4318 -61 4352 -27
rect 4386 -61 4484 -27
rect 4518 -61 4552 -27
rect 4586 -61 4684 -27
rect 4718 -61 4752 -27
rect 4786 -61 4884 -27
rect 4918 -61 4952 -27
rect 4986 -61 5084 -27
rect 5118 -61 5152 -27
rect 5186 -61 5284 -27
rect 5318 -61 5352 -27
rect 5386 -61 5484 -27
rect 5518 -61 5552 -27
rect 5586 -61 5684 -27
rect 5718 -61 5752 -27
rect 5786 -61 5884 -27
rect 5918 -61 5952 -27
rect 5986 -61 6084 -27
rect 6118 -61 6152 -27
rect 6186 -61 6284 -27
rect 6318 -61 6352 -27
rect 6386 -61 6484 -27
rect 6518 -61 6552 -27
rect 6586 -61 6684 -27
rect 6718 -61 6752 -27
rect 6786 -61 6884 -27
rect 6918 -61 6952 -27
rect 6986 -61 7084 -27
rect 7118 -61 7152 -27
rect 7186 -61 7284 -27
rect 7318 -61 7352 -27
rect 7386 -61 7484 -27
rect 7518 -61 7552 -27
rect 7586 -61 7684 -27
rect 7718 -61 7752 -27
rect 7786 -61 7884 -27
rect 7918 -61 7952 -27
rect 7986 -61 8084 -27
rect 8118 -61 8152 -27
rect 8186 -61 8284 -27
rect 8318 -61 8352 -27
rect 8386 -61 8484 -27
rect 8518 -61 8552 -27
rect 8586 -61 8684 -27
rect 8718 -61 8752 -27
rect 8786 -61 8884 -27
rect 8918 -61 8952 -27
rect 8986 -61 9084 -27
rect 9118 -61 9152 -27
rect 9186 -61 9284 -27
rect 9318 -61 9352 -27
rect 9386 -61 9484 -27
rect 9518 -61 9552 -27
rect 9586 -61 9684 -27
rect 9718 -61 9752 -27
rect 9786 -61 9884 -27
rect 9918 -61 9952 -27
rect 9986 -61 10084 -27
rect 10118 -61 10152 -27
rect 10186 -61 10284 -27
rect 10318 -61 10352 -27
rect 10386 -61 10484 -27
rect 10518 -61 10552 -27
rect 10586 -61 10684 -27
rect 10718 -61 10752 -27
rect 10786 -61 10884 -27
rect 10918 -61 10952 -27
rect 10986 -61 11084 -27
rect 11118 -61 11152 -27
rect 11186 -61 11284 -27
rect 11318 -61 11352 -27
rect 11386 -61 11484 -27
rect 11518 -61 11552 -27
rect 11586 -61 11684 -27
rect 11718 -61 11752 -27
rect 11786 -61 11884 -27
rect 11918 -61 11952 -27
rect 11986 -61 12084 -27
rect 12118 -61 12152 -27
rect 12186 -61 12284 -27
rect 12318 -61 12352 -27
rect 12386 -61 12484 -27
rect 12518 -61 12552 -27
rect 12586 -61 12684 -27
rect 12718 -61 12752 -27
rect 12786 -61 12810 -27
rect 14540 -115 14690 -113
rect 14540 -149 14564 -115
rect 14598 -149 14632 -115
rect 14666 -149 14690 -115
rect 14540 -171 14690 -149
rect 15652 -115 15802 -113
rect 15652 -149 15676 -115
rect 15710 -149 15744 -115
rect 15778 -149 15802 -115
rect 15652 -171 15802 -149
rect -10 -2151 108 -2129
rect -10 -2185 32 -2151
rect 66 -2185 108 -2151
rect -10 -2187 108 -2185
rect 162 -2151 280 -2129
rect 162 -2185 204 -2151
rect 238 -2185 280 -2151
rect 162 -2187 280 -2185
rect 390 -2151 508 -2129
rect 390 -2185 432 -2151
rect 466 -2185 508 -2151
rect 390 -2187 508 -2185
rect 562 -2151 680 -2129
rect 562 -2185 604 -2151
rect 638 -2185 680 -2151
rect 562 -2187 680 -2185
rect 790 -2151 908 -2129
rect 790 -2185 832 -2151
rect 866 -2185 908 -2151
rect 790 -2187 908 -2185
rect 962 -2151 1080 -2129
rect 962 -2185 1004 -2151
rect 1038 -2185 1080 -2151
rect 962 -2187 1080 -2185
rect 1190 -2151 1308 -2129
rect 1190 -2185 1232 -2151
rect 1266 -2185 1308 -2151
rect 1190 -2187 1308 -2185
rect 1362 -2151 1480 -2129
rect 1362 -2185 1404 -2151
rect 1438 -2185 1480 -2151
rect 1362 -2187 1480 -2185
rect 1590 -2151 1708 -2129
rect 1590 -2185 1632 -2151
rect 1666 -2185 1708 -2151
rect 1590 -2187 1708 -2185
rect 1762 -2151 1880 -2129
rect 1762 -2185 1804 -2151
rect 1838 -2185 1880 -2151
rect 1762 -2187 1880 -2185
rect 1990 -2151 2108 -2129
rect 1990 -2185 2032 -2151
rect 2066 -2185 2108 -2151
rect 1990 -2187 2108 -2185
rect 2162 -2151 2280 -2129
rect 2162 -2185 2204 -2151
rect 2238 -2185 2280 -2151
rect 2162 -2187 2280 -2185
rect 2390 -2151 2508 -2129
rect 2390 -2185 2432 -2151
rect 2466 -2185 2508 -2151
rect 2390 -2187 2508 -2185
rect 2562 -2151 2680 -2129
rect 2562 -2185 2604 -2151
rect 2638 -2185 2680 -2151
rect 2562 -2187 2680 -2185
rect 2790 -2151 2908 -2129
rect 2790 -2185 2832 -2151
rect 2866 -2185 2908 -2151
rect 2790 -2187 2908 -2185
rect 2962 -2151 3080 -2129
rect 2962 -2185 3004 -2151
rect 3038 -2185 3080 -2151
rect 2962 -2187 3080 -2185
rect 3190 -2151 3308 -2129
rect 3190 -2185 3232 -2151
rect 3266 -2185 3308 -2151
rect 3190 -2187 3308 -2185
rect 3362 -2151 3480 -2129
rect 3362 -2185 3404 -2151
rect 3438 -2185 3480 -2151
rect 3362 -2187 3480 -2185
rect 3590 -2151 3708 -2129
rect 3590 -2185 3632 -2151
rect 3666 -2185 3708 -2151
rect 3590 -2187 3708 -2185
rect 3762 -2151 3880 -2129
rect 3762 -2185 3804 -2151
rect 3838 -2185 3880 -2151
rect 3762 -2187 3880 -2185
rect 3990 -2151 4108 -2129
rect 3990 -2185 4032 -2151
rect 4066 -2185 4108 -2151
rect 3990 -2187 4108 -2185
rect 4162 -2151 4280 -2129
rect 4162 -2185 4204 -2151
rect 4238 -2185 4280 -2151
rect 4162 -2187 4280 -2185
rect 4390 -2151 4508 -2129
rect 4390 -2185 4432 -2151
rect 4466 -2185 4508 -2151
rect 4390 -2187 4508 -2185
rect 4562 -2151 4680 -2129
rect 4562 -2185 4604 -2151
rect 4638 -2185 4680 -2151
rect 4562 -2187 4680 -2185
rect 4790 -2151 4908 -2129
rect 4790 -2185 4832 -2151
rect 4866 -2185 4908 -2151
rect 4790 -2187 4908 -2185
rect 4962 -2151 5080 -2129
rect 4962 -2185 5004 -2151
rect 5038 -2185 5080 -2151
rect 4962 -2187 5080 -2185
rect 5190 -2151 5308 -2129
rect 5190 -2185 5232 -2151
rect 5266 -2185 5308 -2151
rect 5190 -2187 5308 -2185
rect 5362 -2151 5480 -2129
rect 5362 -2185 5404 -2151
rect 5438 -2185 5480 -2151
rect 5362 -2187 5480 -2185
rect 5590 -2151 5708 -2129
rect 5590 -2185 5632 -2151
rect 5666 -2185 5708 -2151
rect 5590 -2187 5708 -2185
rect 5762 -2151 5880 -2129
rect 5762 -2185 5804 -2151
rect 5838 -2185 5880 -2151
rect 5762 -2187 5880 -2185
rect 5990 -2151 6108 -2129
rect 5990 -2185 6032 -2151
rect 6066 -2185 6108 -2151
rect 5990 -2187 6108 -2185
rect 6162 -2151 6280 -2129
rect 6162 -2185 6204 -2151
rect 6238 -2185 6280 -2151
rect 6162 -2187 6280 -2185
rect 6390 -2151 6508 -2129
rect 6390 -2185 6432 -2151
rect 6466 -2185 6508 -2151
rect 6390 -2187 6508 -2185
rect 6562 -2151 6680 -2129
rect 6562 -2185 6604 -2151
rect 6638 -2185 6680 -2151
rect 6562 -2187 6680 -2185
rect 6790 -2151 6908 -2129
rect 6790 -2185 6832 -2151
rect 6866 -2185 6908 -2151
rect 6790 -2187 6908 -2185
rect 6962 -2151 7080 -2129
rect 6962 -2185 7004 -2151
rect 7038 -2185 7080 -2151
rect 6962 -2187 7080 -2185
rect 7190 -2151 7308 -2129
rect 7190 -2185 7232 -2151
rect 7266 -2185 7308 -2151
rect 7190 -2187 7308 -2185
rect 7362 -2151 7480 -2129
rect 7362 -2185 7404 -2151
rect 7438 -2185 7480 -2151
rect 7362 -2187 7480 -2185
rect 7590 -2151 7708 -2129
rect 7590 -2185 7632 -2151
rect 7666 -2185 7708 -2151
rect 7590 -2187 7708 -2185
rect 7762 -2151 7880 -2129
rect 7762 -2185 7804 -2151
rect 7838 -2185 7880 -2151
rect 7762 -2187 7880 -2185
rect 7990 -2151 8108 -2129
rect 7990 -2185 8032 -2151
rect 8066 -2185 8108 -2151
rect 7990 -2187 8108 -2185
rect 8162 -2151 8280 -2129
rect 8162 -2185 8204 -2151
rect 8238 -2185 8280 -2151
rect 8162 -2187 8280 -2185
rect 8390 -2151 8508 -2129
rect 8390 -2185 8432 -2151
rect 8466 -2185 8508 -2151
rect 8390 -2187 8508 -2185
rect 8562 -2151 8680 -2129
rect 8562 -2185 8604 -2151
rect 8638 -2185 8680 -2151
rect 8562 -2187 8680 -2185
rect 8790 -2151 8908 -2129
rect 8790 -2185 8832 -2151
rect 8866 -2185 8908 -2151
rect 8790 -2187 8908 -2185
rect 8962 -2151 9080 -2129
rect 8962 -2185 9004 -2151
rect 9038 -2185 9080 -2151
rect 8962 -2187 9080 -2185
rect 9190 -2151 9308 -2129
rect 9190 -2185 9232 -2151
rect 9266 -2185 9308 -2151
rect 9190 -2187 9308 -2185
rect 9362 -2151 9480 -2129
rect 9362 -2185 9404 -2151
rect 9438 -2185 9480 -2151
rect 9362 -2187 9480 -2185
rect 9590 -2151 9708 -2129
rect 9590 -2185 9632 -2151
rect 9666 -2185 9708 -2151
rect 9590 -2187 9708 -2185
rect 9762 -2151 9880 -2129
rect 9762 -2185 9804 -2151
rect 9838 -2185 9880 -2151
rect 9762 -2187 9880 -2185
rect 9990 -2151 10108 -2129
rect 9990 -2185 10032 -2151
rect 10066 -2185 10108 -2151
rect 9990 -2187 10108 -2185
rect 10162 -2151 10280 -2129
rect 10162 -2185 10204 -2151
rect 10238 -2185 10280 -2151
rect 10162 -2187 10280 -2185
rect 10390 -2151 10508 -2129
rect 10390 -2185 10432 -2151
rect 10466 -2185 10508 -2151
rect 10390 -2187 10508 -2185
rect 10562 -2151 10680 -2129
rect 10562 -2185 10604 -2151
rect 10638 -2185 10680 -2151
rect 10562 -2187 10680 -2185
rect 10790 -2151 10908 -2129
rect 10790 -2185 10832 -2151
rect 10866 -2185 10908 -2151
rect 10790 -2187 10908 -2185
rect 10962 -2151 11080 -2129
rect 10962 -2185 11004 -2151
rect 11038 -2185 11080 -2151
rect 10962 -2187 11080 -2185
rect 11190 -2151 11308 -2129
rect 11190 -2185 11232 -2151
rect 11266 -2185 11308 -2151
rect 11190 -2187 11308 -2185
rect 11362 -2151 11480 -2129
rect 11362 -2185 11404 -2151
rect 11438 -2185 11480 -2151
rect 11362 -2187 11480 -2185
rect 11590 -2151 11708 -2129
rect 11590 -2185 11632 -2151
rect 11666 -2185 11708 -2151
rect 11590 -2187 11708 -2185
rect 11762 -2151 11880 -2129
rect 11762 -2185 11804 -2151
rect 11838 -2185 11880 -2151
rect 11762 -2187 11880 -2185
rect 11990 -2151 12108 -2129
rect 11990 -2185 12032 -2151
rect 12066 -2185 12108 -2151
rect 11990 -2187 12108 -2185
rect 12162 -2151 12280 -2129
rect 12162 -2185 12204 -2151
rect 12238 -2185 12280 -2151
rect 12162 -2187 12280 -2185
rect 12390 -2151 12508 -2129
rect 12390 -2185 12432 -2151
rect 12466 -2185 12508 -2151
rect 12390 -2187 12508 -2185
rect 12562 -2151 12680 -2129
rect 14540 -2101 14690 -2079
rect 14540 -2135 14564 -2101
rect 14598 -2135 14632 -2101
rect 14666 -2135 14690 -2101
rect 14540 -2137 14690 -2135
rect 15652 -2101 15802 -2079
rect 15652 -2135 15676 -2101
rect 15710 -2135 15744 -2101
rect 15778 -2135 15802 -2101
rect 15652 -2137 15802 -2135
rect 12562 -2185 12604 -2151
rect 12638 -2185 12680 -2151
rect 12562 -2187 12680 -2185
<< nsubdiff >>
rect 14816 -115 15116 -113
rect 14816 -149 14847 -115
rect 14881 -149 14915 -115
rect 14949 -149 14983 -115
rect 15017 -149 15051 -115
rect 15085 -149 15116 -115
rect 14816 -171 15116 -149
rect 15226 -115 15526 -113
rect 15226 -149 15257 -115
rect 15291 -149 15325 -115
rect 15359 -149 15393 -115
rect 15427 -149 15461 -115
rect 15495 -149 15526 -115
rect 15226 -171 15526 -149
rect -133 -595 -82 -561
rect -48 -595 3 -561
rect 267 -595 318 -561
rect 352 -595 403 -561
rect 667 -595 718 -561
rect 752 -595 803 -561
rect 1067 -595 1118 -561
rect 1152 -595 1203 -561
rect 1467 -595 1518 -561
rect 1552 -595 1603 -561
rect 1867 -595 1918 -561
rect 1952 -595 2003 -561
rect 2267 -595 2318 -561
rect 2352 -595 2403 -561
rect 2667 -595 2718 -561
rect 2752 -595 2803 -561
rect 3067 -595 3118 -561
rect 3152 -595 3203 -561
rect 3467 -595 3518 -561
rect 3552 -595 3603 -561
rect 3867 -595 3918 -561
rect 3952 -595 4003 -561
rect 4267 -595 4318 -561
rect 4352 -595 4403 -561
rect 4667 -595 4718 -561
rect 4752 -595 4803 -561
rect 5067 -595 5118 -561
rect 5152 -595 5203 -561
rect 5467 -595 5518 -561
rect 5552 -595 5603 -561
rect 5867 -595 5918 -561
rect 5952 -595 6003 -561
rect 6267 -595 6318 -561
rect 6352 -595 6403 -561
rect 6667 -595 6718 -561
rect 6752 -595 6803 -561
rect 7067 -595 7118 -561
rect 7152 -595 7203 -561
rect 7467 -595 7518 -561
rect 7552 -595 7603 -561
rect 7867 -595 7918 -561
rect 7952 -595 8003 -561
rect 8267 -595 8318 -561
rect 8352 -595 8403 -561
rect 8667 -595 8718 -561
rect 8752 -595 8803 -561
rect 9067 -595 9118 -561
rect 9152 -595 9203 -561
rect 9467 -595 9518 -561
rect 9552 -595 9603 -561
rect 9867 -595 9918 -561
rect 9952 -595 10003 -561
rect 10267 -595 10318 -561
rect 10352 -595 10403 -561
rect 10667 -595 10718 -561
rect 10752 -595 10803 -561
rect 11067 -595 11118 -561
rect 11152 -595 11203 -561
rect 11467 -595 11518 -561
rect 11552 -595 11603 -561
rect 11867 -595 11918 -561
rect 11952 -595 12003 -561
rect 12267 -595 12318 -561
rect 12352 -595 12403 -561
rect 12667 -595 12718 -561
rect 12752 -595 12803 -561
rect 14816 -2101 15116 -2079
rect 14816 -2135 14847 -2101
rect 14881 -2135 14915 -2101
rect 14949 -2135 14983 -2101
rect 15017 -2135 15051 -2101
rect 15085 -2135 15116 -2101
rect 14816 -2137 15116 -2135
rect 15226 -2101 15526 -2079
rect 15226 -2135 15257 -2101
rect 15291 -2135 15325 -2101
rect 15359 -2135 15393 -2101
rect 15427 -2135 15461 -2101
rect 15495 -2135 15526 -2101
rect 15226 -2137 15526 -2135
<< psubdiffcont >>
rect 118 4983 152 5017
rect 318 4983 352 5017
rect 518 4983 552 5017
rect 718 4983 752 5017
rect 918 4983 952 5017
rect 1118 4983 1152 5017
rect 1318 4983 1352 5017
rect 1518 4983 1552 5017
rect 1718 4983 1752 5017
rect 1918 4983 1952 5017
rect 2118 4983 2152 5017
rect 2318 4983 2352 5017
rect 2518 4983 2552 5017
rect 2718 4983 2752 5017
rect 2918 4983 2952 5017
rect 3118 4983 3152 5017
rect 3318 4983 3352 5017
rect 3518 4983 3552 5017
rect 3718 4983 3752 5017
rect 3918 4983 3952 5017
rect 4118 4983 4152 5017
rect 4318 4983 4352 5017
rect 4518 4983 4552 5017
rect 4718 4983 4752 5017
rect 4918 4983 4952 5017
rect 5118 4983 5152 5017
rect 5318 4983 5352 5017
rect 5518 4983 5552 5017
rect 5718 4983 5752 5017
rect 5918 4983 5952 5017
rect 6118 4983 6152 5017
rect 6318 4983 6352 5017
rect 6518 4983 6552 5017
rect 6718 4983 6752 5017
rect 6918 4983 6952 5017
rect 7118 4983 7152 5017
rect 7318 4983 7352 5017
rect 7518 4983 7552 5017
rect 7718 4983 7752 5017
rect 7918 4983 7952 5017
rect 8118 4983 8152 5017
rect 8318 4983 8352 5017
rect 8518 4983 8552 5017
rect 8718 4983 8752 5017
rect 8918 4983 8952 5017
rect 9118 4983 9152 5017
rect 9318 4983 9352 5017
rect 9518 4983 9552 5017
rect 9718 4983 9752 5017
rect 9918 4983 9952 5017
rect 10118 4983 10152 5017
rect 10318 4983 10352 5017
rect 10518 4983 10552 5017
rect 10718 4983 10752 5017
rect 10918 4983 10952 5017
rect 11118 4983 11152 5017
rect 11318 4983 11352 5017
rect 11518 4983 11552 5017
rect 11718 4983 11752 5017
rect 11918 4983 11952 5017
rect 12118 4983 12152 5017
rect 12318 4983 12352 5017
rect 12518 4983 12552 5017
rect 12718 4983 12752 5017
rect -116 -61 -82 -27
rect -48 -61 -14 -27
rect 84 -61 118 -27
rect 152 -61 186 -27
rect 284 -61 318 -27
rect 352 -61 386 -27
rect 484 -61 518 -27
rect 552 -61 586 -27
rect 684 -61 718 -27
rect 752 -61 786 -27
rect 884 -61 918 -27
rect 952 -61 986 -27
rect 1084 -61 1118 -27
rect 1152 -61 1186 -27
rect 1284 -61 1318 -27
rect 1352 -61 1386 -27
rect 1484 -61 1518 -27
rect 1552 -61 1586 -27
rect 1684 -61 1718 -27
rect 1752 -61 1786 -27
rect 1884 -61 1918 -27
rect 1952 -61 1986 -27
rect 2084 -61 2118 -27
rect 2152 -61 2186 -27
rect 2284 -61 2318 -27
rect 2352 -61 2386 -27
rect 2484 -61 2518 -27
rect 2552 -61 2586 -27
rect 2684 -61 2718 -27
rect 2752 -61 2786 -27
rect 2884 -61 2918 -27
rect 2952 -61 2986 -27
rect 3084 -61 3118 -27
rect 3152 -61 3186 -27
rect 3284 -61 3318 -27
rect 3352 -61 3386 -27
rect 3484 -61 3518 -27
rect 3552 -61 3586 -27
rect 3684 -61 3718 -27
rect 3752 -61 3786 -27
rect 3884 -61 3918 -27
rect 3952 -61 3986 -27
rect 4084 -61 4118 -27
rect 4152 -61 4186 -27
rect 4284 -61 4318 -27
rect 4352 -61 4386 -27
rect 4484 -61 4518 -27
rect 4552 -61 4586 -27
rect 4684 -61 4718 -27
rect 4752 -61 4786 -27
rect 4884 -61 4918 -27
rect 4952 -61 4986 -27
rect 5084 -61 5118 -27
rect 5152 -61 5186 -27
rect 5284 -61 5318 -27
rect 5352 -61 5386 -27
rect 5484 -61 5518 -27
rect 5552 -61 5586 -27
rect 5684 -61 5718 -27
rect 5752 -61 5786 -27
rect 5884 -61 5918 -27
rect 5952 -61 5986 -27
rect 6084 -61 6118 -27
rect 6152 -61 6186 -27
rect 6284 -61 6318 -27
rect 6352 -61 6386 -27
rect 6484 -61 6518 -27
rect 6552 -61 6586 -27
rect 6684 -61 6718 -27
rect 6752 -61 6786 -27
rect 6884 -61 6918 -27
rect 6952 -61 6986 -27
rect 7084 -61 7118 -27
rect 7152 -61 7186 -27
rect 7284 -61 7318 -27
rect 7352 -61 7386 -27
rect 7484 -61 7518 -27
rect 7552 -61 7586 -27
rect 7684 -61 7718 -27
rect 7752 -61 7786 -27
rect 7884 -61 7918 -27
rect 7952 -61 7986 -27
rect 8084 -61 8118 -27
rect 8152 -61 8186 -27
rect 8284 -61 8318 -27
rect 8352 -61 8386 -27
rect 8484 -61 8518 -27
rect 8552 -61 8586 -27
rect 8684 -61 8718 -27
rect 8752 -61 8786 -27
rect 8884 -61 8918 -27
rect 8952 -61 8986 -27
rect 9084 -61 9118 -27
rect 9152 -61 9186 -27
rect 9284 -61 9318 -27
rect 9352 -61 9386 -27
rect 9484 -61 9518 -27
rect 9552 -61 9586 -27
rect 9684 -61 9718 -27
rect 9752 -61 9786 -27
rect 9884 -61 9918 -27
rect 9952 -61 9986 -27
rect 10084 -61 10118 -27
rect 10152 -61 10186 -27
rect 10284 -61 10318 -27
rect 10352 -61 10386 -27
rect 10484 -61 10518 -27
rect 10552 -61 10586 -27
rect 10684 -61 10718 -27
rect 10752 -61 10786 -27
rect 10884 -61 10918 -27
rect 10952 -61 10986 -27
rect 11084 -61 11118 -27
rect 11152 -61 11186 -27
rect 11284 -61 11318 -27
rect 11352 -61 11386 -27
rect 11484 -61 11518 -27
rect 11552 -61 11586 -27
rect 11684 -61 11718 -27
rect 11752 -61 11786 -27
rect 11884 -61 11918 -27
rect 11952 -61 11986 -27
rect 12084 -61 12118 -27
rect 12152 -61 12186 -27
rect 12284 -61 12318 -27
rect 12352 -61 12386 -27
rect 12484 -61 12518 -27
rect 12552 -61 12586 -27
rect 12684 -61 12718 -27
rect 12752 -61 12786 -27
rect 14564 -149 14598 -115
rect 14632 -149 14666 -115
rect 15676 -149 15710 -115
rect 15744 -149 15778 -115
rect 32 -2185 66 -2151
rect 204 -2185 238 -2151
rect 432 -2185 466 -2151
rect 604 -2185 638 -2151
rect 832 -2185 866 -2151
rect 1004 -2185 1038 -2151
rect 1232 -2185 1266 -2151
rect 1404 -2185 1438 -2151
rect 1632 -2185 1666 -2151
rect 1804 -2185 1838 -2151
rect 2032 -2185 2066 -2151
rect 2204 -2185 2238 -2151
rect 2432 -2185 2466 -2151
rect 2604 -2185 2638 -2151
rect 2832 -2185 2866 -2151
rect 3004 -2185 3038 -2151
rect 3232 -2185 3266 -2151
rect 3404 -2185 3438 -2151
rect 3632 -2185 3666 -2151
rect 3804 -2185 3838 -2151
rect 4032 -2185 4066 -2151
rect 4204 -2185 4238 -2151
rect 4432 -2185 4466 -2151
rect 4604 -2185 4638 -2151
rect 4832 -2185 4866 -2151
rect 5004 -2185 5038 -2151
rect 5232 -2185 5266 -2151
rect 5404 -2185 5438 -2151
rect 5632 -2185 5666 -2151
rect 5804 -2185 5838 -2151
rect 6032 -2185 6066 -2151
rect 6204 -2185 6238 -2151
rect 6432 -2185 6466 -2151
rect 6604 -2185 6638 -2151
rect 6832 -2185 6866 -2151
rect 7004 -2185 7038 -2151
rect 7232 -2185 7266 -2151
rect 7404 -2185 7438 -2151
rect 7632 -2185 7666 -2151
rect 7804 -2185 7838 -2151
rect 8032 -2185 8066 -2151
rect 8204 -2185 8238 -2151
rect 8432 -2185 8466 -2151
rect 8604 -2185 8638 -2151
rect 8832 -2185 8866 -2151
rect 9004 -2185 9038 -2151
rect 9232 -2185 9266 -2151
rect 9404 -2185 9438 -2151
rect 9632 -2185 9666 -2151
rect 9804 -2185 9838 -2151
rect 10032 -2185 10066 -2151
rect 10204 -2185 10238 -2151
rect 10432 -2185 10466 -2151
rect 10604 -2185 10638 -2151
rect 10832 -2185 10866 -2151
rect 11004 -2185 11038 -2151
rect 11232 -2185 11266 -2151
rect 11404 -2185 11438 -2151
rect 11632 -2185 11666 -2151
rect 11804 -2185 11838 -2151
rect 12032 -2185 12066 -2151
rect 12204 -2185 12238 -2151
rect 12432 -2185 12466 -2151
rect 14564 -2135 14598 -2101
rect 14632 -2135 14666 -2101
rect 15676 -2135 15710 -2101
rect 15744 -2135 15778 -2101
rect 12604 -2185 12638 -2151
<< nsubdiffcont >>
rect 14847 -149 14881 -115
rect 14915 -149 14949 -115
rect 14983 -149 15017 -115
rect 15051 -149 15085 -115
rect 15257 -149 15291 -115
rect 15325 -149 15359 -115
rect 15393 -149 15427 -115
rect 15461 -149 15495 -115
rect -82 -595 -48 -561
rect 318 -595 352 -561
rect 718 -595 752 -561
rect 1118 -595 1152 -561
rect 1518 -595 1552 -561
rect 1918 -595 1952 -561
rect 2318 -595 2352 -561
rect 2718 -595 2752 -561
rect 3118 -595 3152 -561
rect 3518 -595 3552 -561
rect 3918 -595 3952 -561
rect 4318 -595 4352 -561
rect 4718 -595 4752 -561
rect 5118 -595 5152 -561
rect 5518 -595 5552 -561
rect 5918 -595 5952 -561
rect 6318 -595 6352 -561
rect 6718 -595 6752 -561
rect 7118 -595 7152 -561
rect 7518 -595 7552 -561
rect 7918 -595 7952 -561
rect 8318 -595 8352 -561
rect 8718 -595 8752 -561
rect 9118 -595 9152 -561
rect 9518 -595 9552 -561
rect 9918 -595 9952 -561
rect 10318 -595 10352 -561
rect 10718 -595 10752 -561
rect 11118 -595 11152 -561
rect 11518 -595 11552 -561
rect 11918 -595 11952 -561
rect 12318 -595 12352 -561
rect 12718 -595 12752 -561
rect 14847 -2135 14881 -2101
rect 14915 -2135 14949 -2101
rect 14983 -2135 15017 -2101
rect 15051 -2135 15085 -2101
rect 15257 -2135 15291 -2101
rect 15325 -2135 15359 -2101
rect 15393 -2135 15427 -2101
rect 15461 -2135 15495 -2101
<< poly >>
rect 70 4904 100 5070
rect 170 4904 200 5070
rect 70 4894 200 4904
rect 70 4860 118 4894
rect 152 4860 200 4894
rect 70 4850 200 4860
rect 70 4813 100 4850
rect 170 4813 200 4850
rect 270 4920 300 5070
rect 370 4920 400 5070
rect 270 4910 400 4920
rect 270 4876 318 4910
rect 352 4876 400 4910
rect 270 4866 400 4876
rect 270 4813 300 4866
rect 70 4673 100 4727
rect 170 4673 200 4727
rect 270 4673 300 4727
rect 370 4673 400 4866
rect 470 4904 500 5070
rect 570 4904 600 5070
rect 470 4894 600 4904
rect 470 4860 518 4894
rect 552 4860 600 4894
rect 470 4850 600 4860
rect 470 4813 500 4850
rect 570 4813 600 4850
rect 670 4920 700 5070
rect 770 4920 800 5070
rect 670 4910 800 4920
rect 670 4876 718 4910
rect 752 4876 800 4910
rect 670 4866 800 4876
rect 670 4813 700 4866
rect 770 4813 800 4866
rect 870 4904 900 5070
rect 970 4904 1000 5070
rect 870 4894 1000 4904
rect 870 4860 918 4894
rect 952 4860 1000 4894
rect 870 4850 1000 4860
rect 870 4813 900 4850
rect 970 4813 1000 4850
rect 1070 4920 1100 5070
rect 1170 4920 1200 5070
rect 1070 4910 1200 4920
rect 1070 4876 1118 4910
rect 1152 4876 1200 4910
rect 1070 4866 1200 4876
rect 1070 4813 1100 4866
rect 470 4673 500 4727
rect 570 4673 600 4727
rect 670 4673 700 4727
rect 770 4673 800 4727
rect 870 4673 900 4727
rect 970 4673 1000 4727
rect 1070 4673 1100 4727
rect 70 4533 100 4587
rect 170 4533 200 4587
rect 270 4533 300 4587
rect 70 4393 100 4447
rect 170 4393 200 4447
rect 270 4393 300 4447
rect 370 4393 400 4587
rect 470 4533 500 4587
rect 570 4533 600 4587
rect 670 4533 700 4587
rect 770 4533 800 4587
rect 870 4533 900 4587
rect 970 4533 1000 4587
rect 1070 4533 1100 4587
rect 1170 4533 1200 4866
rect 1270 4904 1300 5070
rect 1370 4904 1400 5070
rect 1270 4894 1400 4904
rect 1270 4860 1318 4894
rect 1352 4860 1400 4894
rect 1270 4850 1400 4860
rect 1270 4813 1300 4850
rect 1370 4813 1400 4850
rect 1470 4920 1500 5070
rect 1570 4920 1600 5070
rect 1470 4910 1600 4920
rect 1470 4876 1518 4910
rect 1552 4876 1600 4910
rect 1470 4866 1600 4876
rect 1470 4813 1500 4866
rect 1570 4813 1600 4866
rect 1670 4904 1700 5070
rect 1770 4904 1800 5070
rect 1670 4894 1800 4904
rect 1670 4860 1718 4894
rect 1752 4860 1800 4894
rect 1670 4850 1800 4860
rect 1670 4813 1700 4850
rect 1770 4813 1800 4850
rect 1870 4920 1900 5070
rect 1970 4920 2000 5070
rect 1870 4910 2000 4920
rect 1870 4876 1918 4910
rect 1952 4876 2000 4910
rect 1870 4866 2000 4876
rect 1870 4813 1900 4866
rect 1970 4813 2000 4866
rect 2070 4904 2100 5070
rect 2170 4904 2200 5070
rect 2070 4894 2200 4904
rect 2070 4860 2118 4894
rect 2152 4860 2200 4894
rect 2070 4850 2200 4860
rect 2070 4813 2100 4850
rect 2170 4813 2200 4850
rect 2270 4920 2300 5070
rect 2370 4920 2400 5070
rect 2270 4910 2400 4920
rect 2270 4876 2318 4910
rect 2352 4876 2400 4910
rect 2270 4866 2400 4876
rect 2270 4813 2300 4866
rect 1270 4673 1300 4727
rect 1370 4673 1400 4727
rect 1470 4673 1500 4727
rect 1570 4673 1600 4727
rect 1670 4673 1700 4727
rect 1770 4673 1800 4727
rect 1870 4673 1900 4727
rect 1970 4673 2000 4727
rect 2070 4673 2100 4727
rect 2170 4673 2200 4727
rect 2270 4673 2300 4727
rect 2370 4673 2400 4866
rect 2470 4904 2500 5070
rect 2570 4904 2600 5070
rect 2470 4894 2600 4904
rect 2470 4860 2518 4894
rect 2552 4860 2600 4894
rect 2470 4850 2600 4860
rect 2470 4813 2500 4850
rect 2570 4813 2600 4850
rect 2670 4920 2700 5070
rect 2770 4920 2800 5070
rect 2670 4910 2800 4920
rect 2670 4876 2718 4910
rect 2752 4876 2800 4910
rect 2670 4866 2800 4876
rect 2670 4813 2700 4866
rect 2770 4813 2800 4866
rect 2870 4904 2900 5070
rect 2970 4904 3000 5070
rect 2870 4894 3000 4904
rect 2870 4860 2918 4894
rect 2952 4860 3000 4894
rect 2870 4850 3000 4860
rect 2870 4813 2900 4850
rect 2970 4813 3000 4850
rect 3070 4920 3100 5070
rect 3170 4920 3200 5070
rect 3070 4910 3200 4920
rect 3070 4876 3118 4910
rect 3152 4876 3200 4910
rect 3070 4866 3200 4876
rect 3070 4813 3100 4866
rect 2470 4673 2500 4727
rect 2570 4673 2600 4727
rect 2670 4673 2700 4727
rect 2770 4673 2800 4727
rect 2870 4673 2900 4727
rect 1270 4533 1300 4587
rect 1370 4533 1400 4587
rect 1470 4533 1500 4587
rect 1570 4533 1600 4587
rect 470 4393 500 4447
rect 570 4393 600 4447
rect 670 4393 700 4447
rect 770 4393 800 4447
rect 870 4393 900 4447
rect 970 4393 1000 4447
rect 1070 4393 1100 4447
rect 1170 4393 1200 4447
rect 70 4253 100 4307
rect 170 4253 200 4307
rect 270 4253 300 4307
rect 370 4253 400 4307
rect 470 4253 500 4307
rect 70 4113 100 4167
rect 170 4113 200 4167
rect 70 3973 100 4027
rect 170 3973 200 4027
rect 270 3973 300 4167
rect 370 4113 400 4167
rect 370 3973 400 4027
rect 470 3973 500 4167
rect 570 4113 600 4307
rect 670 4253 700 4307
rect 770 4253 800 4307
rect 870 4253 900 4307
rect 970 4253 1000 4307
rect 1070 4253 1100 4307
rect 670 4113 700 4167
rect 770 4113 800 4167
rect 870 4113 900 4167
rect 970 4113 1000 4167
rect 1070 4113 1100 4167
rect 1170 4113 1200 4307
rect 1270 4253 1300 4447
rect 1370 4393 1400 4447
rect 1470 4393 1500 4447
rect 1570 4393 1600 4447
rect 1670 4393 1700 4587
rect 1770 4533 1800 4587
rect 1770 4393 1800 4447
rect 1870 4393 1900 4587
rect 1970 4533 2000 4587
rect 2070 4533 2100 4587
rect 2170 4533 2200 4587
rect 2270 4533 2300 4587
rect 1370 4253 1400 4307
rect 1470 4253 1500 4307
rect 1570 4253 1600 4307
rect 1670 4253 1700 4307
rect 1770 4253 1800 4307
rect 1870 4253 1900 4307
rect 1270 4113 1300 4167
rect 570 3973 600 4027
rect 670 3973 700 4027
rect 770 3973 800 4027
rect 870 3973 900 4027
rect 970 3973 1000 4027
rect 1070 3973 1100 4027
rect 1170 3973 1200 4027
rect 1270 3973 1300 4027
rect 1370 3973 1400 4167
rect 1470 4113 1500 4167
rect 1570 4113 1600 4167
rect 1470 3973 1500 4027
rect 1570 3973 1600 4027
rect 1670 3973 1700 4167
rect 1770 4113 1800 4167
rect 1870 4113 1900 4167
rect 1970 4113 2000 4447
rect 2070 4393 2100 4447
rect 2170 4393 2200 4447
rect 2270 4393 2300 4447
rect 2370 4393 2400 4587
rect 2470 4533 2500 4587
rect 2570 4533 2600 4587
rect 2470 4393 2500 4447
rect 2570 4393 2600 4447
rect 2670 4393 2700 4587
rect 2770 4533 2800 4587
rect 2770 4393 2800 4447
rect 2870 4393 2900 4587
rect 2970 4533 3000 4727
rect 3070 4673 3100 4727
rect 3170 4673 3200 4866
rect 3270 4904 3300 5070
rect 3370 4904 3400 5070
rect 3270 4894 3400 4904
rect 3270 4860 3318 4894
rect 3352 4860 3400 4894
rect 3270 4850 3400 4860
rect 3270 4813 3300 4850
rect 3370 4813 3400 4850
rect 3470 4920 3500 5070
rect 3570 4920 3600 5070
rect 3470 4910 3600 4920
rect 3470 4876 3518 4910
rect 3552 4876 3600 4910
rect 3470 4866 3600 4876
rect 3270 4673 3300 4727
rect 3370 4673 3400 4727
rect 3470 4673 3500 4866
rect 3570 4813 3600 4866
rect 3670 4904 3700 5070
rect 3770 4904 3800 5070
rect 3670 4894 3800 4904
rect 3670 4860 3718 4894
rect 3752 4860 3800 4894
rect 3670 4850 3800 4860
rect 3670 4813 3700 4850
rect 3770 4813 3800 4850
rect 3870 4920 3900 5070
rect 3970 4920 4000 5070
rect 3870 4910 4000 4920
rect 3870 4876 3918 4910
rect 3952 4876 4000 4910
rect 3870 4866 4000 4876
rect 3870 4813 3900 4866
rect 3970 4813 4000 4866
rect 4070 4904 4100 5070
rect 4170 4904 4200 5070
rect 4070 4894 4200 4904
rect 4070 4860 4118 4894
rect 4152 4860 4200 4894
rect 4070 4850 4200 4860
rect 4070 4813 4100 4850
rect 4170 4813 4200 4850
rect 4270 4920 4300 5070
rect 4370 4920 4400 5070
rect 4270 4910 4400 4920
rect 4270 4876 4318 4910
rect 4352 4876 4400 4910
rect 4270 4866 4400 4876
rect 3570 4673 3600 4727
rect 3070 4533 3100 4587
rect 3170 4533 3200 4587
rect 3270 4533 3300 4587
rect 3370 4533 3400 4587
rect 3470 4533 3500 4587
rect 3570 4533 3600 4587
rect 3670 4533 3700 4727
rect 3770 4673 3800 4727
rect 3870 4673 3900 4727
rect 3970 4673 4000 4727
rect 4070 4673 4100 4727
rect 4170 4673 4200 4727
rect 4270 4673 4300 4866
rect 4370 4813 4400 4866
rect 4470 4904 4500 5070
rect 4570 4904 4600 5070
rect 4470 4894 4600 4904
rect 4470 4860 4518 4894
rect 4552 4860 4600 4894
rect 4470 4850 4600 4860
rect 4470 4813 4500 4850
rect 4570 4813 4600 4850
rect 4670 4920 4700 5070
rect 4770 4920 4800 5070
rect 4670 4910 4800 4920
rect 4670 4876 4718 4910
rect 4752 4876 4800 4910
rect 4670 4866 4800 4876
rect 4670 4813 4700 4866
rect 4770 4813 4800 4866
rect 4870 4904 4900 5070
rect 4970 4904 5000 5070
rect 4870 4894 5000 4904
rect 4870 4860 4918 4894
rect 4952 4860 5000 4894
rect 4870 4850 5000 4860
rect 4870 4813 4900 4850
rect 4970 4813 5000 4850
rect 5070 4920 5100 5070
rect 5170 4920 5200 5070
rect 5070 4910 5200 4920
rect 5070 4876 5118 4910
rect 5152 4876 5200 4910
rect 5070 4866 5200 4876
rect 5070 4813 5100 4866
rect 5170 4813 5200 4866
rect 5270 4904 5300 5070
rect 5370 4904 5400 5070
rect 5270 4894 5400 4904
rect 5270 4860 5318 4894
rect 5352 4860 5400 4894
rect 5270 4850 5400 4860
rect 5270 4813 5300 4850
rect 5370 4813 5400 4850
rect 5470 4920 5500 5070
rect 5570 4920 5600 5070
rect 5470 4910 5600 4920
rect 5470 4876 5518 4910
rect 5552 4876 5600 4910
rect 5470 4866 5600 4876
rect 5470 4813 5500 4866
rect 5570 4813 5600 4866
rect 5670 4904 5700 5070
rect 5770 4904 5800 5070
rect 5670 4894 5800 4904
rect 5670 4860 5718 4894
rect 5752 4860 5800 4894
rect 5670 4850 5800 4860
rect 5670 4813 5700 4850
rect 5770 4813 5800 4850
rect 5870 4920 5900 5070
rect 5970 4920 6000 5070
rect 5870 4910 6000 4920
rect 5870 4876 5918 4910
rect 5952 4876 6000 4910
rect 5870 4866 6000 4876
rect 5870 4813 5900 4866
rect 5970 4813 6000 4866
rect 6070 4904 6100 5070
rect 6170 4904 6200 5070
rect 6070 4894 6200 4904
rect 6070 4860 6118 4894
rect 6152 4860 6200 4894
rect 6070 4850 6200 4860
rect 6070 4813 6100 4850
rect 6170 4813 6200 4850
rect 6270 4920 6300 5070
rect 6370 4920 6400 5070
rect 6270 4910 6400 4920
rect 6270 4876 6318 4910
rect 6352 4876 6400 4910
rect 6270 4866 6400 4876
rect 6270 4813 6300 4866
rect 6370 4813 6400 4866
rect 6470 4904 6500 5070
rect 6570 4904 6600 5070
rect 6470 4894 6600 4904
rect 6470 4860 6518 4894
rect 6552 4860 6600 4894
rect 6470 4850 6600 4860
rect 4370 4673 4400 4727
rect 4470 4673 4500 4727
rect 4570 4673 4600 4727
rect 4670 4673 4700 4727
rect 2970 4393 3000 4447
rect 3070 4393 3100 4447
rect 3170 4393 3200 4447
rect 3270 4393 3300 4447
rect 3370 4393 3400 4447
rect 3470 4393 3500 4447
rect 3570 4393 3600 4447
rect 3670 4393 3700 4447
rect 2070 4253 2100 4307
rect 2170 4253 2200 4307
rect 2270 4253 2300 4307
rect 2370 4253 2400 4307
rect 2470 4253 2500 4307
rect 2570 4253 2600 4307
rect 2670 4253 2700 4307
rect 2770 4253 2800 4307
rect 2870 4253 2900 4307
rect 2970 4253 3000 4307
rect 3070 4253 3100 4307
rect 3170 4253 3200 4307
rect 3270 4253 3300 4307
rect 3370 4253 3400 4307
rect 3470 4253 3500 4307
rect 3570 4253 3600 4307
rect 3670 4253 3700 4307
rect 3770 4253 3800 4587
rect 3870 4533 3900 4587
rect 3970 4533 4000 4587
rect 4070 4533 4100 4587
rect 4170 4533 4200 4587
rect 4270 4533 4300 4587
rect 4370 4533 4400 4587
rect 4470 4533 4500 4587
rect 4570 4533 4600 4587
rect 4670 4533 4700 4587
rect 4770 4533 4800 4727
rect 4870 4673 4900 4727
rect 4970 4673 5000 4727
rect 4870 4533 4900 4587
rect 4970 4533 5000 4587
rect 3870 4393 3900 4447
rect 3970 4393 4000 4447
rect 4070 4393 4100 4447
rect 4170 4393 4200 4447
rect 4270 4393 4300 4447
rect 4370 4393 4400 4447
rect 4470 4393 4500 4447
rect 4570 4393 4600 4447
rect 4670 4393 4700 4447
rect 4770 4393 4800 4447
rect 4870 4393 4900 4447
rect 4970 4393 5000 4447
rect 5070 4393 5100 4727
rect 5170 4673 5200 4727
rect 5270 4673 5300 4727
rect 5370 4673 5400 4727
rect 5470 4673 5500 4727
rect 5570 4673 5600 4727
rect 5670 4673 5700 4727
rect 5770 4673 5800 4727
rect 5170 4533 5200 4587
rect 5270 4533 5300 4587
rect 5170 4393 5200 4447
rect 5270 4393 5300 4447
rect 5370 4393 5400 4587
rect 5470 4533 5500 4587
rect 5570 4533 5600 4587
rect 5670 4533 5700 4587
rect 5770 4533 5800 4587
rect 5870 4533 5900 4727
rect 5970 4673 6000 4727
rect 6070 4673 6100 4727
rect 6170 4673 6200 4727
rect 6270 4673 6300 4727
rect 6370 4673 6400 4727
rect 5970 4533 6000 4587
rect 5470 4393 5500 4447
rect 5570 4393 5600 4447
rect 5670 4393 5700 4447
rect 5770 4393 5800 4447
rect 5870 4393 5900 4447
rect 5970 4393 6000 4447
rect 3870 4253 3900 4307
rect 3970 4253 4000 4307
rect 2070 4113 2100 4167
rect 2170 4113 2200 4167
rect 1770 3973 1800 4027
rect 1870 3973 1900 4027
rect 70 3833 100 3887
rect 170 3833 200 3887
rect 270 3833 300 3887
rect 370 3833 400 3887
rect 470 3833 500 3887
rect 570 3833 600 3887
rect 670 3833 700 3887
rect 770 3833 800 3887
rect 870 3833 900 3887
rect 970 3833 1000 3887
rect 1070 3833 1100 3887
rect 1170 3833 1200 3887
rect 1270 3833 1300 3887
rect 1370 3833 1400 3887
rect 1470 3833 1500 3887
rect 1570 3833 1600 3887
rect 1670 3833 1700 3887
rect 1770 3833 1800 3887
rect 1870 3833 1900 3887
rect 1970 3833 2000 4027
rect 2070 3973 2100 4027
rect 2170 3973 2200 4027
rect 2270 3973 2300 4167
rect 2370 4113 2400 4167
rect 2470 4113 2500 4167
rect 2570 4113 2600 4167
rect 2370 3973 2400 4027
rect 2470 3973 2500 4027
rect 2570 3973 2600 4027
rect 2670 3973 2700 4167
rect 2770 4113 2800 4167
rect 2870 4113 2900 4167
rect 2770 3973 2800 4027
rect 2870 3973 2900 4027
rect 2970 3973 3000 4167
rect 3070 4113 3100 4167
rect 3170 4113 3200 4167
rect 3070 3973 3100 4027
rect 3170 3973 3200 4027
rect 3270 3973 3300 4167
rect 3370 4113 3400 4167
rect 3470 4113 3500 4167
rect 3570 4113 3600 4167
rect 3670 4113 3700 4167
rect 3770 4113 3800 4167
rect 3870 4113 3900 4167
rect 3970 4113 4000 4167
rect 4070 4113 4100 4307
rect 4170 4253 4200 4307
rect 3370 3973 3400 4027
rect 3470 3973 3500 4027
rect 3570 3973 3600 4027
rect 3670 3973 3700 4027
rect 3770 3973 3800 4027
rect 3870 3973 3900 4027
rect 2070 3833 2100 3887
rect 70 3694 100 3747
rect 170 3694 200 3747
rect 70 3684 200 3694
rect 70 3650 118 3684
rect 152 3650 200 3684
rect 70 3640 200 3650
rect 70 3603 100 3640
rect 170 3603 200 3640
rect 270 3710 300 3747
rect 370 3710 400 3747
rect 270 3700 400 3710
rect 270 3666 318 3700
rect 352 3666 400 3700
rect 270 3656 400 3666
rect 270 3603 300 3656
rect 370 3603 400 3656
rect 470 3694 500 3747
rect 570 3694 600 3747
rect 470 3684 600 3694
rect 470 3650 518 3684
rect 552 3650 600 3684
rect 470 3640 600 3650
rect 470 3603 500 3640
rect 570 3603 600 3640
rect 670 3710 700 3747
rect 770 3710 800 3747
rect 670 3700 800 3710
rect 670 3666 718 3700
rect 752 3666 800 3700
rect 670 3656 800 3666
rect 670 3603 700 3656
rect 770 3603 800 3656
rect 870 3694 900 3747
rect 970 3694 1000 3747
rect 870 3684 1000 3694
rect 870 3650 918 3684
rect 952 3650 1000 3684
rect 870 3640 1000 3650
rect 70 3463 100 3517
rect 170 3463 200 3517
rect 270 3463 300 3517
rect 70 3323 100 3377
rect 170 3323 200 3377
rect 270 3323 300 3377
rect 370 3323 400 3517
rect 470 3463 500 3517
rect 470 3323 500 3377
rect 570 3323 600 3517
rect 670 3463 700 3517
rect 670 3323 700 3377
rect 70 3183 100 3237
rect 70 3043 100 3097
rect 170 3043 200 3237
rect 270 3183 300 3237
rect 370 3183 400 3237
rect 470 3183 500 3237
rect 570 3183 600 3237
rect 670 3183 700 3237
rect 770 3183 800 3517
rect 870 3463 900 3640
rect 970 3603 1000 3640
rect 1070 3710 1100 3747
rect 1170 3710 1200 3747
rect 1070 3700 1200 3710
rect 1070 3666 1118 3700
rect 1152 3666 1200 3700
rect 1070 3656 1200 3666
rect 870 3323 900 3377
rect 870 3183 900 3237
rect 970 3183 1000 3517
rect 1070 3463 1100 3656
rect 1170 3603 1200 3656
rect 1270 3694 1300 3747
rect 1370 3694 1400 3747
rect 1270 3684 1400 3694
rect 1270 3650 1318 3684
rect 1352 3650 1400 3684
rect 1270 3640 1400 3650
rect 1270 3603 1300 3640
rect 1370 3603 1400 3640
rect 1470 3710 1500 3747
rect 1570 3710 1600 3747
rect 1470 3700 1600 3710
rect 1470 3666 1518 3700
rect 1552 3666 1600 3700
rect 1470 3656 1600 3666
rect 1470 3603 1500 3656
rect 1570 3603 1600 3656
rect 1670 3694 1700 3747
rect 1770 3694 1800 3747
rect 1670 3684 1800 3694
rect 1670 3650 1718 3684
rect 1752 3650 1800 3684
rect 1670 3640 1800 3650
rect 1670 3603 1700 3640
rect 1770 3603 1800 3640
rect 1870 3710 1900 3747
rect 1970 3710 2000 3747
rect 1870 3700 2000 3710
rect 1870 3666 1918 3700
rect 1952 3666 2000 3700
rect 1870 3656 2000 3666
rect 1870 3603 1900 3656
rect 1970 3603 2000 3656
rect 2070 3694 2100 3747
rect 2170 3694 2200 3887
rect 2270 3833 2300 3887
rect 2370 3833 2400 3887
rect 2470 3833 2500 3887
rect 2070 3684 2200 3694
rect 2070 3650 2118 3684
rect 2152 3650 2200 3684
rect 2070 3640 2200 3650
rect 2070 3603 2100 3640
rect 2170 3603 2200 3640
rect 2270 3710 2300 3747
rect 2370 3710 2400 3747
rect 2270 3700 2400 3710
rect 2270 3666 2318 3700
rect 2352 3666 2400 3700
rect 2270 3656 2400 3666
rect 2270 3603 2300 3656
rect 2370 3603 2400 3656
rect 2470 3694 2500 3747
rect 2570 3694 2600 3887
rect 2670 3833 2700 3887
rect 2470 3684 2600 3694
rect 2470 3650 2518 3684
rect 2552 3650 2600 3684
rect 2470 3640 2600 3650
rect 2470 3603 2500 3640
rect 1170 3463 1200 3517
rect 1270 3463 1300 3517
rect 1370 3463 1400 3517
rect 1470 3463 1500 3517
rect 1570 3463 1600 3517
rect 1670 3463 1700 3517
rect 1770 3463 1800 3517
rect 1870 3463 1900 3517
rect 1970 3463 2000 3517
rect 2070 3463 2100 3517
rect 2170 3463 2200 3517
rect 2270 3463 2300 3517
rect 2370 3463 2400 3517
rect 2470 3463 2500 3517
rect 2570 3463 2600 3640
rect 2670 3710 2700 3747
rect 2770 3710 2800 3887
rect 2870 3833 2900 3887
rect 2970 3833 3000 3887
rect 3070 3833 3100 3887
rect 2670 3700 2800 3710
rect 2670 3666 2718 3700
rect 2752 3666 2800 3700
rect 2670 3656 2800 3666
rect 2670 3603 2700 3656
rect 2770 3603 2800 3656
rect 2870 3694 2900 3747
rect 2970 3694 3000 3747
rect 2870 3684 3000 3694
rect 2870 3650 2918 3684
rect 2952 3650 3000 3684
rect 2870 3640 3000 3650
rect 2870 3603 2900 3640
rect 2970 3603 3000 3640
rect 3070 3710 3100 3747
rect 3170 3710 3200 3887
rect 3270 3833 3300 3887
rect 3370 3833 3400 3887
rect 3470 3833 3500 3887
rect 3570 3833 3600 3887
rect 3670 3833 3700 3887
rect 3770 3833 3800 3887
rect 3870 3833 3900 3887
rect 3970 3833 4000 4027
rect 4070 3973 4100 4027
rect 4070 3833 4100 3887
rect 4170 3833 4200 4167
rect 4270 4113 4300 4307
rect 4370 4253 4400 4307
rect 4270 3973 4300 4027
rect 4370 3973 4400 4167
rect 4470 4113 4500 4307
rect 4570 4253 4600 4307
rect 4470 3973 4500 4027
rect 4570 3973 4600 4167
rect 4670 4113 4700 4307
rect 4770 4253 4800 4307
rect 4670 3973 4700 4027
rect 4770 3973 4800 4167
rect 4870 4113 4900 4307
rect 4970 4253 5000 4307
rect 5070 4253 5100 4307
rect 5170 4253 5200 4307
rect 5270 4253 5300 4307
rect 5370 4253 5400 4307
rect 5470 4253 5500 4307
rect 4870 3973 4900 4027
rect 4970 3973 5000 4167
rect 5070 4113 5100 4167
rect 5170 4113 5200 4167
rect 4270 3833 4300 3887
rect 4370 3833 4400 3887
rect 4470 3833 4500 3887
rect 3070 3700 3200 3710
rect 3070 3666 3118 3700
rect 3152 3666 3200 3700
rect 3070 3656 3200 3666
rect 3070 3603 3100 3656
rect 2670 3463 2700 3517
rect 2770 3463 2800 3517
rect 2870 3463 2900 3517
rect 2970 3463 3000 3517
rect 3070 3463 3100 3517
rect 3170 3463 3200 3656
rect 3270 3694 3300 3747
rect 3370 3694 3400 3747
rect 3270 3684 3400 3694
rect 3270 3650 3318 3684
rect 3352 3650 3400 3684
rect 3270 3640 3400 3650
rect 3270 3603 3300 3640
rect 3370 3603 3400 3640
rect 3470 3710 3500 3747
rect 3570 3710 3600 3747
rect 3470 3700 3600 3710
rect 3470 3666 3518 3700
rect 3552 3666 3600 3700
rect 3470 3656 3600 3666
rect 3470 3603 3500 3656
rect 3570 3603 3600 3656
rect 3670 3694 3700 3747
rect 3770 3694 3800 3747
rect 3670 3684 3800 3694
rect 3670 3650 3718 3684
rect 3752 3650 3800 3684
rect 3670 3640 3800 3650
rect 3670 3603 3700 3640
rect 3770 3603 3800 3640
rect 3870 3710 3900 3747
rect 3970 3710 4000 3747
rect 3870 3700 4000 3710
rect 3870 3666 3918 3700
rect 3952 3666 4000 3700
rect 3870 3656 4000 3666
rect 3870 3603 3900 3656
rect 3970 3603 4000 3656
rect 4070 3694 4100 3747
rect 4170 3694 4200 3747
rect 4070 3684 4200 3694
rect 4070 3650 4118 3684
rect 4152 3650 4200 3684
rect 4070 3640 4200 3650
rect 4070 3603 4100 3640
rect 4170 3603 4200 3640
rect 4270 3710 4300 3747
rect 4370 3710 4400 3747
rect 4270 3700 4400 3710
rect 4270 3666 4318 3700
rect 4352 3666 4400 3700
rect 4270 3656 4400 3666
rect 4270 3603 4300 3656
rect 4370 3603 4400 3656
rect 4470 3694 4500 3747
rect 4570 3694 4600 3887
rect 4670 3833 4700 3887
rect 4770 3833 4800 3887
rect 4870 3833 4900 3887
rect 4970 3833 5000 3887
rect 5070 3833 5100 4027
rect 5170 3973 5200 4027
rect 5170 3833 5200 3887
rect 5270 3833 5300 4167
rect 5370 4113 5400 4167
rect 5470 4113 5500 4167
rect 5570 4113 5600 4307
rect 5670 4253 5700 4307
rect 5770 4253 5800 4307
rect 5870 4253 5900 4307
rect 5970 4253 6000 4307
rect 5370 3973 5400 4027
rect 5470 3973 5500 4027
rect 5370 3833 5400 3887
rect 4470 3684 4600 3694
rect 4470 3650 4518 3684
rect 4552 3650 4600 3684
rect 4470 3640 4600 3650
rect 3270 3463 3300 3517
rect 3370 3463 3400 3517
rect 3470 3463 3500 3517
rect 3570 3463 3600 3517
rect 3670 3463 3700 3517
rect 3770 3463 3800 3517
rect 1070 3323 1100 3377
rect 1170 3323 1200 3377
rect 1270 3323 1300 3377
rect 1370 3323 1400 3377
rect 1470 3323 1500 3377
rect 1570 3323 1600 3377
rect 1670 3323 1700 3377
rect 1770 3323 1800 3377
rect 1870 3323 1900 3377
rect 1970 3323 2000 3377
rect 2070 3323 2100 3377
rect 2170 3323 2200 3377
rect 2270 3323 2300 3377
rect 2370 3323 2400 3377
rect 2470 3323 2500 3377
rect 2570 3323 2600 3377
rect 2670 3323 2700 3377
rect 1070 3183 1100 3237
rect 1170 3183 1200 3237
rect 1270 3183 1300 3237
rect 270 3043 300 3097
rect 370 3043 400 3097
rect 470 3043 500 3097
rect 570 3043 600 3097
rect 70 2903 100 2957
rect 170 2903 200 2957
rect 270 2903 300 2957
rect 370 2903 400 2957
rect 470 2903 500 2957
rect 570 2903 600 2957
rect 670 2903 700 3097
rect 770 3043 800 3097
rect 870 3043 900 3097
rect 970 3043 1000 3097
rect 1070 3043 1100 3097
rect 1170 3043 1200 3097
rect 1270 3043 1300 3097
rect 1370 3043 1400 3237
rect 1470 3183 1500 3237
rect 1570 3183 1600 3237
rect 1670 3183 1700 3237
rect 1770 3183 1800 3237
rect 1870 3183 1900 3237
rect 1970 3183 2000 3237
rect 2070 3183 2100 3237
rect 2170 3183 2200 3237
rect 2270 3183 2300 3237
rect 2370 3183 2400 3237
rect 2470 3183 2500 3237
rect 1470 3043 1500 3097
rect 1570 3043 1600 3097
rect 1670 3043 1700 3097
rect 1770 3043 1800 3097
rect 1870 3043 1900 3097
rect 1970 3043 2000 3097
rect 770 2903 800 2957
rect 70 2763 100 2817
rect 170 2763 200 2817
rect 270 2763 300 2817
rect 370 2763 400 2817
rect 470 2763 500 2817
rect 570 2763 600 2817
rect 670 2763 700 2817
rect 770 2763 800 2817
rect 870 2763 900 2957
rect 970 2903 1000 2957
rect 1070 2903 1100 2957
rect 1170 2903 1200 2957
rect 1270 2903 1300 2957
rect 1370 2903 1400 2957
rect 1470 2903 1500 2957
rect 1570 2903 1600 2957
rect 1670 2903 1700 2957
rect 1770 2903 1800 2957
rect 1870 2903 1900 2957
rect 1970 2903 2000 2957
rect 2070 2903 2100 3097
rect 2170 3043 2200 3097
rect 2270 3043 2300 3097
rect 2370 3043 2400 3097
rect 2470 3043 2500 3097
rect 2570 3043 2600 3237
rect 2670 3183 2700 3237
rect 2770 3183 2800 3377
rect 2870 3323 2900 3377
rect 2970 3323 3000 3377
rect 3070 3323 3100 3377
rect 3170 3323 3200 3377
rect 2870 3183 2900 3237
rect 2970 3183 3000 3237
rect 3070 3183 3100 3237
rect 3170 3183 3200 3237
rect 2670 3043 2700 3097
rect 2770 3043 2800 3097
rect 2870 3043 2900 3097
rect 2970 3043 3000 3097
rect 2170 2903 2200 2957
rect 2270 2903 2300 2957
rect 2370 2903 2400 2957
rect 2470 2903 2500 2957
rect 2570 2903 2600 2957
rect 970 2763 1000 2817
rect 1070 2763 1100 2817
rect 70 2623 100 2677
rect 170 2623 200 2677
rect 270 2623 300 2677
rect 370 2623 400 2677
rect 470 2623 500 2677
rect 570 2623 600 2677
rect 670 2623 700 2677
rect 770 2623 800 2677
rect 870 2623 900 2677
rect 970 2623 1000 2677
rect 1070 2623 1100 2677
rect 1170 2623 1200 2817
rect 1270 2763 1300 2817
rect 1370 2763 1400 2817
rect 1470 2763 1500 2817
rect 1570 2763 1600 2817
rect 1670 2763 1700 2817
rect 1770 2763 1800 2817
rect 1870 2763 1900 2817
rect 1970 2763 2000 2817
rect 2070 2763 2100 2817
rect 2170 2763 2200 2817
rect 2270 2763 2300 2817
rect 1270 2623 1300 2677
rect 1370 2623 1400 2677
rect 1470 2623 1500 2677
rect 1570 2623 1600 2677
rect 1670 2623 1700 2677
rect 1770 2623 1800 2677
rect 1870 2623 1900 2677
rect 1970 2623 2000 2677
rect 2070 2623 2100 2677
rect 2170 2623 2200 2677
rect 2270 2623 2300 2677
rect 2370 2623 2400 2817
rect 2470 2763 2500 2817
rect 2570 2763 2600 2817
rect 2670 2763 2700 2957
rect 2770 2903 2800 2957
rect 2870 2903 2900 2957
rect 2770 2763 2800 2817
rect 2870 2763 2900 2817
rect 2970 2763 3000 2957
rect 3070 2903 3100 3097
rect 3170 3043 3200 3097
rect 3270 3043 3300 3377
rect 3370 3323 3400 3377
rect 3370 3183 3400 3237
rect 3470 3183 3500 3377
rect 3570 3323 3600 3377
rect 3670 3323 3700 3377
rect 3770 3323 3800 3377
rect 3870 3323 3900 3517
rect 3970 3463 4000 3517
rect 4070 3463 4100 3517
rect 4170 3463 4200 3517
rect 4270 3463 4300 3517
rect 4370 3463 4400 3517
rect 3970 3323 4000 3377
rect 4070 3323 4100 3377
rect 4170 3323 4200 3377
rect 4270 3323 4300 3377
rect 4370 3323 4400 3377
rect 4470 3323 4500 3640
rect 4570 3603 4600 3640
rect 4670 3710 4700 3747
rect 4770 3710 4800 3747
rect 4670 3700 4800 3710
rect 4670 3666 4718 3700
rect 4752 3666 4800 3700
rect 4670 3656 4800 3666
rect 4670 3603 4700 3656
rect 4770 3603 4800 3656
rect 4870 3694 4900 3747
rect 4970 3694 5000 3747
rect 4870 3684 5000 3694
rect 4870 3650 4918 3684
rect 4952 3650 5000 3684
rect 4870 3640 5000 3650
rect 4870 3603 4900 3640
rect 4970 3603 5000 3640
rect 5070 3710 5100 3747
rect 5170 3710 5200 3747
rect 5070 3700 5200 3710
rect 5070 3666 5118 3700
rect 5152 3666 5200 3700
rect 5070 3656 5200 3666
rect 5070 3603 5100 3656
rect 5170 3603 5200 3656
rect 5270 3694 5300 3747
rect 5370 3694 5400 3747
rect 5270 3684 5400 3694
rect 5270 3650 5318 3684
rect 5352 3650 5400 3684
rect 5270 3640 5400 3650
rect 5270 3603 5300 3640
rect 5370 3603 5400 3640
rect 5470 3710 5500 3887
rect 5570 3833 5600 4027
rect 5670 3973 5700 4167
rect 5770 4113 5800 4167
rect 5870 4113 5900 4167
rect 5970 4113 6000 4167
rect 6070 4113 6100 4587
rect 6170 4533 6200 4587
rect 6270 4533 6300 4587
rect 6370 4533 6400 4587
rect 6470 4533 6500 4850
rect 6570 4813 6600 4850
rect 6670 4920 6700 5070
rect 6770 4920 6800 5070
rect 6670 4910 6800 4920
rect 6670 4876 6718 4910
rect 6752 4876 6800 4910
rect 6670 4866 6800 4876
rect 6670 4813 6700 4866
rect 6770 4813 6800 4866
rect 6870 4904 6900 5070
rect 6970 4904 7000 5070
rect 6870 4894 7000 4904
rect 6870 4860 6918 4894
rect 6952 4860 7000 4894
rect 6870 4850 7000 4860
rect 6870 4813 6900 4850
rect 6970 4813 7000 4850
rect 7070 4920 7100 5070
rect 7170 4920 7200 5070
rect 7070 4910 7200 4920
rect 7070 4876 7118 4910
rect 7152 4876 7200 4910
rect 7070 4866 7200 4876
rect 7070 4813 7100 4866
rect 7170 4813 7200 4866
rect 7270 4904 7300 5070
rect 7370 4904 7400 5070
rect 7270 4894 7400 4904
rect 7270 4860 7318 4894
rect 7352 4860 7400 4894
rect 7270 4850 7400 4860
rect 7270 4813 7300 4850
rect 7370 4813 7400 4850
rect 7470 4920 7500 5070
rect 7570 4920 7600 5070
rect 7470 4910 7600 4920
rect 7470 4876 7518 4910
rect 7552 4876 7600 4910
rect 7470 4866 7600 4876
rect 7470 4813 7500 4866
rect 7570 4813 7600 4866
rect 7670 4904 7700 5070
rect 7770 4904 7800 5070
rect 7670 4894 7800 4904
rect 7670 4860 7718 4894
rect 7752 4860 7800 4894
rect 7670 4850 7800 4860
rect 7670 4813 7700 4850
rect 7770 4813 7800 4850
rect 7870 4920 7900 5070
rect 7970 4920 8000 5070
rect 7870 4910 8000 4920
rect 7870 4876 7918 4910
rect 7952 4876 8000 4910
rect 7870 4866 8000 4876
rect 7870 4813 7900 4866
rect 7970 4813 8000 4866
rect 8070 4904 8100 5070
rect 8170 4904 8200 5070
rect 8070 4894 8200 4904
rect 8070 4860 8118 4894
rect 8152 4860 8200 4894
rect 8070 4850 8200 4860
rect 8070 4813 8100 4850
rect 8170 4813 8200 4850
rect 8270 4920 8300 5070
rect 8370 4920 8400 5070
rect 8270 4910 8400 4920
rect 8270 4876 8318 4910
rect 8352 4876 8400 4910
rect 8270 4866 8400 4876
rect 8270 4813 8300 4866
rect 8370 4813 8400 4866
rect 8470 4904 8500 5070
rect 8570 4904 8600 5070
rect 8470 4894 8600 4904
rect 8470 4860 8518 4894
rect 8552 4860 8600 4894
rect 8470 4850 8600 4860
rect 8470 4813 8500 4850
rect 8570 4813 8600 4850
rect 8670 4920 8700 5070
rect 8770 4920 8800 5070
rect 8670 4910 8800 4920
rect 8670 4876 8718 4910
rect 8752 4876 8800 4910
rect 8670 4866 8800 4876
rect 8670 4813 8700 4866
rect 8770 4813 8800 4866
rect 8870 4904 8900 5070
rect 8970 4904 9000 5070
rect 8870 4894 9000 4904
rect 8870 4860 8918 4894
rect 8952 4860 9000 4894
rect 8870 4850 9000 4860
rect 8870 4813 8900 4850
rect 8970 4813 9000 4850
rect 9070 4920 9100 5070
rect 9170 4920 9200 5070
rect 9070 4910 9200 4920
rect 9070 4876 9118 4910
rect 9152 4876 9200 4910
rect 9070 4866 9200 4876
rect 9070 4813 9100 4866
rect 9170 4813 9200 4866
rect 9270 4904 9300 5070
rect 9370 4904 9400 5070
rect 9270 4894 9400 4904
rect 9270 4860 9318 4894
rect 9352 4860 9400 4894
rect 9270 4850 9400 4860
rect 9270 4813 9300 4850
rect 9370 4813 9400 4850
rect 9470 4920 9500 5070
rect 9570 4920 9600 5070
rect 9470 4910 9600 4920
rect 9470 4876 9518 4910
rect 9552 4876 9600 4910
rect 9470 4866 9600 4876
rect 9470 4813 9500 4866
rect 9570 4813 9600 4866
rect 9670 4904 9700 5070
rect 9770 4904 9800 5070
rect 9670 4894 9800 4904
rect 9670 4860 9718 4894
rect 9752 4860 9800 4894
rect 9670 4850 9800 4860
rect 9670 4813 9700 4850
rect 9770 4813 9800 4850
rect 9870 4920 9900 5070
rect 9970 4920 10000 5070
rect 9870 4910 10000 4920
rect 9870 4876 9918 4910
rect 9952 4876 10000 4910
rect 9870 4866 10000 4876
rect 6570 4673 6600 4727
rect 6670 4673 6700 4727
rect 6770 4673 6800 4727
rect 6870 4673 6900 4727
rect 6970 4673 7000 4727
rect 7070 4673 7100 4727
rect 7170 4673 7200 4727
rect 7270 4673 7300 4727
rect 7370 4673 7400 4727
rect 7470 4673 7500 4727
rect 7570 4673 7600 4727
rect 7670 4673 7700 4727
rect 7770 4673 7800 4727
rect 7870 4673 7900 4727
rect 7970 4673 8000 4727
rect 8070 4673 8100 4727
rect 8170 4673 8200 4727
rect 8270 4673 8300 4727
rect 8370 4673 8400 4727
rect 8470 4673 8500 4727
rect 8570 4673 8600 4727
rect 8670 4673 8700 4727
rect 6570 4533 6600 4587
rect 6670 4533 6700 4587
rect 6770 4533 6800 4587
rect 6870 4533 6900 4587
rect 6970 4533 7000 4587
rect 7070 4533 7100 4587
rect 7170 4533 7200 4587
rect 7270 4533 7300 4587
rect 7370 4533 7400 4587
rect 7470 4533 7500 4587
rect 7570 4533 7600 4587
rect 7670 4533 7700 4587
rect 7770 4533 7800 4587
rect 7870 4533 7900 4587
rect 7970 4533 8000 4587
rect 6170 4393 6200 4447
rect 6270 4393 6300 4447
rect 6370 4393 6400 4447
rect 6470 4393 6500 4447
rect 6570 4393 6600 4447
rect 6170 4253 6200 4307
rect 6170 4113 6200 4167
rect 6270 4113 6300 4307
rect 6370 4253 6400 4307
rect 6370 4113 6400 4167
rect 6470 4113 6500 4307
rect 6570 4253 6600 4307
rect 6570 4113 6600 4167
rect 6670 4113 6700 4447
rect 6770 4393 6800 4447
rect 6870 4393 6900 4447
rect 6970 4393 7000 4447
rect 7070 4393 7100 4447
rect 7170 4393 7200 4447
rect 7270 4393 7300 4447
rect 6770 4253 6800 4307
rect 6870 4253 6900 4307
rect 6970 4253 7000 4307
rect 7070 4253 7100 4307
rect 6770 4113 6800 4167
rect 6870 4113 6900 4167
rect 6970 4113 7000 4167
rect 7070 4113 7100 4167
rect 7170 4113 7200 4307
rect 7270 4253 7300 4307
rect 7370 4253 7400 4447
rect 7470 4393 7500 4447
rect 7570 4393 7600 4447
rect 7670 4393 7700 4447
rect 7770 4393 7800 4447
rect 7870 4393 7900 4447
rect 7970 4393 8000 4447
rect 8070 4393 8100 4587
rect 8170 4533 8200 4587
rect 8270 4533 8300 4587
rect 8170 4393 8200 4447
rect 8270 4393 8300 4447
rect 8370 4393 8400 4587
rect 8470 4533 8500 4587
rect 8570 4533 8600 4587
rect 8670 4533 8700 4587
rect 8770 4533 8800 4727
rect 8870 4673 8900 4727
rect 8970 4673 9000 4727
rect 9070 4673 9100 4727
rect 9170 4673 9200 4727
rect 9270 4673 9300 4727
rect 9370 4673 9400 4727
rect 9470 4673 9500 4727
rect 9570 4673 9600 4727
rect 9670 4673 9700 4727
rect 9770 4673 9800 4727
rect 9870 4673 9900 4866
rect 9970 4813 10000 4866
rect 10070 4904 10100 5070
rect 10170 4904 10200 5070
rect 10070 4894 10200 4904
rect 10070 4860 10118 4894
rect 10152 4860 10200 4894
rect 10070 4850 10200 4860
rect 10070 4813 10100 4850
rect 10170 4813 10200 4850
rect 10270 4920 10300 5070
rect 10370 4920 10400 5070
rect 10270 4910 10400 4920
rect 10270 4876 10318 4910
rect 10352 4876 10400 4910
rect 10270 4866 10400 4876
rect 10270 4813 10300 4866
rect 10370 4813 10400 4866
rect 10470 4904 10500 5070
rect 10570 4904 10600 5070
rect 10470 4894 10600 4904
rect 10470 4860 10518 4894
rect 10552 4860 10600 4894
rect 10470 4850 10600 4860
rect 10470 4813 10500 4850
rect 10570 4813 10600 4850
rect 10670 4920 10700 5070
rect 10770 4920 10800 5070
rect 10670 4910 10800 4920
rect 10670 4876 10718 4910
rect 10752 4876 10800 4910
rect 10670 4866 10800 4876
rect 10670 4813 10700 4866
rect 9970 4673 10000 4727
rect 10070 4673 10100 4727
rect 10170 4673 10200 4727
rect 10270 4673 10300 4727
rect 10370 4673 10400 4727
rect 10470 4673 10500 4727
rect 10570 4673 10600 4727
rect 10670 4673 10700 4727
rect 10770 4673 10800 4866
rect 10870 4904 10900 5070
rect 10970 4904 11000 5070
rect 10870 4894 11000 4904
rect 10870 4860 10918 4894
rect 10952 4860 11000 4894
rect 10870 4850 11000 4860
rect 10870 4813 10900 4850
rect 10970 4813 11000 4850
rect 11070 4920 11100 5070
rect 11170 4920 11200 5070
rect 11070 4910 11200 4920
rect 11070 4876 11118 4910
rect 11152 4876 11200 4910
rect 11070 4866 11200 4876
rect 11070 4813 11100 4866
rect 11170 4813 11200 4866
rect 11270 4904 11300 5070
rect 11370 4904 11400 5070
rect 11270 4894 11400 4904
rect 11270 4860 11318 4894
rect 11352 4860 11400 4894
rect 11270 4850 11400 4860
rect 11270 4813 11300 4850
rect 11370 4813 11400 4850
rect 11470 4920 11500 5070
rect 11570 4920 11600 5070
rect 11470 4910 11600 4920
rect 11470 4876 11518 4910
rect 11552 4876 11600 4910
rect 11470 4866 11600 4876
rect 11470 4813 11500 4866
rect 11570 4813 11600 4866
rect 11670 4904 11700 5070
rect 11770 4904 11800 5070
rect 11670 4894 11800 4904
rect 11670 4860 11718 4894
rect 11752 4860 11800 4894
rect 11670 4850 11800 4860
rect 10870 4673 10900 4727
rect 10970 4673 11000 4727
rect 11070 4673 11100 4727
rect 11170 4673 11200 4727
rect 11270 4673 11300 4727
rect 11370 4673 11400 4727
rect 11470 4673 11500 4727
rect 11570 4673 11600 4727
rect 11670 4673 11700 4850
rect 11770 4813 11800 4850
rect 11870 4920 11900 5070
rect 11970 4920 12000 5070
rect 11870 4910 12000 4920
rect 11870 4876 11918 4910
rect 11952 4876 12000 4910
rect 11870 4866 12000 4876
rect 11870 4813 11900 4866
rect 11970 4813 12000 4866
rect 12070 4904 12100 5070
rect 12170 4904 12200 5070
rect 12070 4894 12200 4904
rect 12070 4860 12118 4894
rect 12152 4860 12200 4894
rect 12070 4850 12200 4860
rect 12070 4813 12100 4850
rect 12170 4813 12200 4850
rect 12270 4920 12300 5070
rect 12370 4920 12400 5070
rect 12270 4910 12400 4920
rect 12270 4876 12318 4910
rect 12352 4876 12400 4910
rect 12270 4866 12400 4876
rect 12270 4813 12300 4866
rect 12370 4813 12400 4866
rect 12470 4904 12500 5070
rect 12570 4904 12600 5070
rect 12470 4894 12600 4904
rect 12470 4860 12518 4894
rect 12552 4860 12600 4894
rect 12470 4850 12600 4860
rect 11770 4673 11800 4727
rect 11870 4673 11900 4727
rect 11970 4673 12000 4727
rect 12070 4673 12100 4727
rect 12170 4673 12200 4727
rect 12270 4673 12300 4727
rect 12370 4673 12400 4727
rect 12470 4673 12500 4850
rect 12570 4813 12600 4850
rect 12670 4920 12700 5070
rect 12770 4920 12800 5070
rect 12970 4924 13000 5070
rect 13070 4924 13100 5070
rect 13280 4924 13310 5070
rect 13380 4924 13410 5070
rect 13480 4924 13510 5070
rect 13580 4924 13610 5070
rect 12670 4910 12800 4920
rect 12670 4876 12718 4910
rect 12752 4876 12800 4910
rect 12670 4866 12800 4876
rect 12670 4813 12700 4866
rect 12770 4813 12800 4866
rect 12958 4908 13012 4924
rect 12958 4874 12968 4908
rect 13002 4874 13012 4908
rect 12958 4858 13012 4874
rect 13058 4908 13112 4924
rect 13058 4874 13068 4908
rect 13102 4874 13112 4908
rect 13058 4858 13112 4874
rect 13268 4908 13322 4924
rect 13268 4874 13278 4908
rect 13312 4874 13322 4908
rect 13268 4858 13322 4874
rect 13368 4908 13422 4924
rect 13368 4874 13378 4908
rect 13412 4874 13422 4908
rect 13368 4858 13422 4874
rect 13468 4908 13522 4924
rect 13468 4874 13478 4908
rect 13512 4874 13522 4908
rect 13468 4858 13522 4874
rect 13568 4908 13622 4924
rect 13568 4874 13578 4908
rect 13612 4874 13622 4908
rect 13568 4858 13622 4874
rect 12970 4813 13000 4858
rect 13070 4813 13100 4858
rect 13280 4813 13310 4858
rect 13380 4813 13410 4858
rect 13480 4813 13510 4858
rect 13580 4813 13610 4858
rect 12570 4673 12600 4727
rect 8470 4393 8500 4447
rect 8570 4393 8600 4447
rect 8670 4393 8700 4447
rect 8770 4393 8800 4447
rect 8870 4393 8900 4587
rect 8970 4533 9000 4587
rect 8970 4393 9000 4447
rect 9070 4393 9100 4587
rect 9170 4533 9200 4587
rect 9270 4533 9300 4587
rect 9170 4393 9200 4447
rect 9270 4393 9300 4447
rect 9370 4393 9400 4587
rect 9470 4533 9500 4587
rect 9570 4533 9600 4587
rect 9470 4393 9500 4447
rect 9570 4393 9600 4447
rect 9670 4393 9700 4587
rect 9770 4533 9800 4587
rect 9870 4533 9900 4587
rect 9770 4393 9800 4447
rect 9870 4393 9900 4447
rect 9970 4393 10000 4587
rect 10070 4533 10100 4587
rect 10170 4533 10200 4587
rect 10070 4393 10100 4447
rect 10170 4393 10200 4447
rect 10270 4393 10300 4587
rect 10370 4533 10400 4587
rect 10470 4533 10500 4587
rect 10370 4393 10400 4447
rect 10470 4393 10500 4447
rect 10570 4393 10600 4587
rect 10670 4533 10700 4587
rect 10670 4393 10700 4447
rect 10770 4393 10800 4587
rect 10870 4533 10900 4587
rect 7470 4253 7500 4307
rect 7570 4253 7600 4307
rect 7670 4253 7700 4307
rect 7770 4253 7800 4307
rect 7870 4253 7900 4307
rect 7970 4253 8000 4307
rect 8070 4253 8100 4307
rect 7270 4113 7300 4167
rect 5770 3973 5800 4027
rect 5870 3973 5900 4027
rect 5670 3833 5700 3887
rect 5770 3833 5800 3887
rect 5870 3833 5900 3887
rect 5570 3710 5600 3747
rect 5470 3700 5600 3710
rect 5470 3666 5518 3700
rect 5552 3666 5600 3700
rect 5470 3656 5600 3666
rect 5470 3603 5500 3656
rect 5570 3603 5600 3656
rect 5670 3694 5700 3747
rect 5770 3694 5800 3747
rect 5670 3684 5800 3694
rect 5670 3650 5718 3684
rect 5752 3650 5800 3684
rect 5670 3640 5800 3650
rect 5670 3603 5700 3640
rect 4570 3463 4600 3517
rect 4670 3463 4700 3517
rect 4770 3463 4800 3517
rect 4570 3323 4600 3377
rect 4670 3323 4700 3377
rect 4770 3323 4800 3377
rect 4870 3323 4900 3517
rect 4970 3463 5000 3517
rect 4970 3323 5000 3377
rect 5070 3323 5100 3517
rect 5170 3463 5200 3517
rect 5270 3463 5300 3517
rect 5370 3463 5400 3517
rect 5470 3463 5500 3517
rect 5570 3463 5600 3517
rect 5670 3463 5700 3517
rect 5770 3463 5800 3640
rect 5870 3710 5900 3747
rect 5970 3710 6000 4027
rect 6070 3973 6100 4027
rect 6170 3973 6200 4027
rect 6270 3973 6300 4027
rect 6370 3973 6400 4027
rect 6470 3973 6500 4027
rect 6570 3973 6600 4027
rect 6670 3973 6700 4027
rect 6770 3973 6800 4027
rect 6870 3973 6900 4027
rect 6070 3833 6100 3887
rect 6170 3833 6200 3887
rect 6270 3833 6300 3887
rect 6370 3833 6400 3887
rect 6470 3833 6500 3887
rect 6570 3833 6600 3887
rect 6670 3833 6700 3887
rect 6770 3833 6800 3887
rect 6870 3833 6900 3887
rect 6970 3833 7000 4027
rect 7070 3973 7100 4027
rect 7070 3833 7100 3887
rect 7170 3833 7200 4027
rect 7270 3973 7300 4027
rect 7370 3973 7400 4167
rect 7470 4113 7500 4167
rect 7570 4113 7600 4167
rect 7470 3973 7500 4027
rect 7570 3973 7600 4027
rect 7670 3973 7700 4167
rect 7770 4113 7800 4167
rect 7770 3973 7800 4027
rect 7870 3973 7900 4167
rect 7970 4113 8000 4167
rect 8070 4113 8100 4167
rect 8170 4113 8200 4307
rect 8270 4253 8300 4307
rect 8270 4113 8300 4167
rect 8370 4113 8400 4307
rect 8470 4253 8500 4307
rect 8470 4113 8500 4167
rect 8570 4113 8600 4307
rect 8670 4253 8700 4307
rect 8670 4113 8700 4167
rect 7970 3973 8000 4027
rect 8070 3973 8100 4027
rect 8170 3973 8200 4027
rect 8270 3973 8300 4027
rect 8370 3973 8400 4027
rect 8470 3973 8500 4027
rect 8570 3973 8600 4027
rect 8670 3973 8700 4027
rect 7270 3833 7300 3887
rect 7370 3833 7400 3887
rect 7470 3833 7500 3887
rect 7570 3833 7600 3887
rect 5870 3700 6000 3710
rect 5870 3666 5918 3700
rect 5952 3666 6000 3700
rect 5870 3656 6000 3666
rect 5870 3603 5900 3656
rect 5970 3603 6000 3656
rect 6070 3694 6100 3747
rect 6170 3694 6200 3747
rect 6070 3684 6200 3694
rect 6070 3650 6118 3684
rect 6152 3650 6200 3684
rect 6070 3640 6200 3650
rect 6070 3603 6100 3640
rect 6170 3603 6200 3640
rect 6270 3710 6300 3747
rect 6370 3710 6400 3747
rect 6270 3700 6400 3710
rect 6270 3666 6318 3700
rect 6352 3666 6400 3700
rect 6270 3656 6400 3666
rect 6270 3603 6300 3656
rect 6370 3603 6400 3656
rect 6470 3694 6500 3747
rect 6570 3694 6600 3747
rect 6470 3684 6600 3694
rect 6470 3650 6518 3684
rect 6552 3650 6600 3684
rect 6470 3640 6600 3650
rect 6470 3603 6500 3640
rect 6570 3603 6600 3640
rect 6670 3710 6700 3747
rect 6770 3710 6800 3747
rect 6670 3700 6800 3710
rect 6670 3666 6718 3700
rect 6752 3666 6800 3700
rect 6670 3656 6800 3666
rect 6670 3603 6700 3656
rect 6770 3603 6800 3656
rect 6870 3694 6900 3747
rect 6970 3694 7000 3747
rect 6870 3684 7000 3694
rect 6870 3650 6918 3684
rect 6952 3650 7000 3684
rect 6870 3640 7000 3650
rect 6870 3603 6900 3640
rect 6970 3603 7000 3640
rect 7070 3710 7100 3747
rect 7170 3710 7200 3747
rect 7070 3700 7200 3710
rect 7070 3666 7118 3700
rect 7152 3666 7200 3700
rect 7070 3656 7200 3666
rect 7070 3603 7100 3656
rect 7170 3603 7200 3656
rect 7270 3694 7300 3747
rect 7370 3694 7400 3747
rect 7270 3684 7400 3694
rect 7270 3650 7318 3684
rect 7352 3650 7400 3684
rect 7270 3640 7400 3650
rect 7270 3603 7300 3640
rect 7370 3603 7400 3640
rect 7470 3710 7500 3747
rect 7570 3710 7600 3747
rect 7470 3700 7600 3710
rect 7470 3666 7518 3700
rect 7552 3666 7600 3700
rect 7470 3656 7600 3666
rect 7470 3603 7500 3656
rect 7570 3603 7600 3656
rect 7670 3694 7700 3887
rect 7770 3833 7800 3887
rect 7870 3833 7900 3887
rect 7970 3833 8000 3887
rect 8070 3833 8100 3887
rect 8170 3833 8200 3887
rect 8270 3833 8300 3887
rect 8370 3833 8400 3887
rect 8470 3833 8500 3887
rect 8570 3833 8600 3887
rect 8670 3833 8700 3887
rect 8770 3833 8800 4307
rect 8870 4253 8900 4307
rect 8870 4113 8900 4167
rect 8870 3973 8900 4027
rect 8970 3973 9000 4307
rect 9070 4253 9100 4307
rect 9170 4253 9200 4307
rect 9270 4253 9300 4307
rect 9070 4113 9100 4167
rect 9170 4113 9200 4167
rect 9270 4113 9300 4167
rect 9370 4113 9400 4307
rect 9470 4253 9500 4307
rect 9470 4113 9500 4167
rect 9070 3973 9100 4027
rect 9170 3973 9200 4027
rect 9270 3973 9300 4027
rect 9370 3973 9400 4027
rect 9470 3973 9500 4027
rect 8870 3833 8900 3887
rect 8970 3833 9000 3887
rect 9070 3833 9100 3887
rect 9170 3833 9200 3887
rect 9270 3833 9300 3887
rect 9370 3833 9400 3887
rect 7770 3694 7800 3747
rect 7670 3684 7800 3694
rect 7670 3650 7718 3684
rect 7752 3650 7800 3684
rect 7670 3640 7800 3650
rect 7670 3603 7700 3640
rect 7770 3603 7800 3640
rect 7870 3710 7900 3747
rect 7970 3710 8000 3747
rect 7870 3700 8000 3710
rect 7870 3666 7918 3700
rect 7952 3666 8000 3700
rect 7870 3656 8000 3666
rect 7870 3603 7900 3656
rect 7970 3603 8000 3656
rect 8070 3694 8100 3747
rect 8170 3694 8200 3747
rect 8070 3684 8200 3694
rect 8070 3650 8118 3684
rect 8152 3650 8200 3684
rect 8070 3640 8200 3650
rect 8070 3603 8100 3640
rect 8170 3603 8200 3640
rect 8270 3710 8300 3747
rect 8370 3710 8400 3747
rect 8270 3700 8400 3710
rect 8270 3666 8318 3700
rect 8352 3666 8400 3700
rect 8270 3656 8400 3666
rect 8270 3603 8300 3656
rect 8370 3603 8400 3656
rect 8470 3694 8500 3747
rect 8570 3694 8600 3747
rect 8470 3684 8600 3694
rect 8470 3650 8518 3684
rect 8552 3650 8600 3684
rect 8470 3640 8600 3650
rect 8470 3603 8500 3640
rect 8570 3603 8600 3640
rect 8670 3710 8700 3747
rect 8770 3710 8800 3747
rect 8670 3700 8800 3710
rect 8670 3666 8718 3700
rect 8752 3666 8800 3700
rect 8670 3656 8800 3666
rect 8670 3603 8700 3656
rect 8770 3603 8800 3656
rect 8870 3694 8900 3747
rect 8970 3694 9000 3747
rect 8870 3684 9000 3694
rect 8870 3650 8918 3684
rect 8952 3650 9000 3684
rect 8870 3640 9000 3650
rect 8870 3603 8900 3640
rect 5870 3463 5900 3517
rect 5970 3463 6000 3517
rect 5170 3323 5200 3377
rect 5270 3323 5300 3377
rect 5370 3323 5400 3377
rect 5470 3323 5500 3377
rect 5570 3323 5600 3377
rect 5670 3323 5700 3377
rect 5770 3323 5800 3377
rect 5870 3323 5900 3377
rect 5970 3323 6000 3377
rect 6070 3323 6100 3517
rect 6170 3463 6200 3517
rect 6270 3463 6300 3517
rect 6370 3463 6400 3517
rect 6170 3323 6200 3377
rect 6270 3323 6300 3377
rect 6370 3323 6400 3377
rect 6470 3323 6500 3517
rect 6570 3463 6600 3517
rect 6670 3463 6700 3517
rect 6570 3323 6600 3377
rect 6670 3323 6700 3377
rect 6770 3323 6800 3517
rect 6870 3463 6900 3517
rect 6970 3463 7000 3517
rect 7070 3463 7100 3517
rect 7170 3463 7200 3517
rect 7270 3463 7300 3517
rect 7370 3463 7400 3517
rect 7470 3463 7500 3517
rect 7570 3463 7600 3517
rect 7670 3463 7700 3517
rect 7770 3463 7800 3517
rect 7870 3463 7900 3517
rect 7970 3463 8000 3517
rect 8070 3463 8100 3517
rect 8170 3463 8200 3517
rect 8270 3463 8300 3517
rect 8370 3463 8400 3517
rect 8470 3463 8500 3517
rect 8570 3463 8600 3517
rect 8670 3463 8700 3517
rect 8770 3463 8800 3517
rect 8870 3463 8900 3517
rect 8970 3463 9000 3640
rect 9070 3710 9100 3747
rect 9170 3710 9200 3747
rect 9070 3700 9200 3710
rect 9070 3666 9118 3700
rect 9152 3666 9200 3700
rect 9070 3656 9200 3666
rect 9070 3603 9100 3656
rect 9070 3463 9100 3517
rect 9170 3463 9200 3656
rect 9270 3694 9300 3747
rect 9370 3694 9400 3747
rect 9270 3684 9400 3694
rect 9270 3650 9318 3684
rect 9352 3650 9400 3684
rect 9270 3640 9400 3650
rect 9270 3603 9300 3640
rect 9270 3463 9300 3517
rect 9370 3463 9400 3640
rect 9470 3710 9500 3887
rect 9570 3833 9600 4307
rect 9670 4253 9700 4307
rect 9670 4113 9700 4167
rect 9770 4113 9800 4307
rect 9870 4253 9900 4307
rect 9970 4253 10000 4307
rect 9870 4113 9900 4167
rect 9970 4113 10000 4167
rect 10070 4113 10100 4307
rect 10170 4253 10200 4307
rect 10270 4253 10300 4307
rect 10370 4253 10400 4307
rect 10470 4253 10500 4307
rect 10570 4253 10600 4307
rect 10670 4253 10700 4307
rect 10770 4253 10800 4307
rect 10870 4253 10900 4447
rect 10970 4393 11000 4587
rect 11070 4533 11100 4587
rect 11170 4533 11200 4587
rect 11070 4393 11100 4447
rect 10170 4113 10200 4167
rect 10270 4113 10300 4167
rect 10370 4113 10400 4167
rect 10470 4113 10500 4167
rect 10570 4113 10600 4167
rect 9670 3973 9700 4027
rect 9770 3973 9800 4027
rect 9870 3973 9900 4027
rect 9970 3973 10000 4027
rect 10070 3973 10100 4027
rect 10170 3973 10200 4027
rect 10270 3973 10300 4027
rect 10370 3973 10400 4027
rect 10470 3973 10500 4027
rect 10570 3973 10600 4027
rect 10670 3973 10700 4167
rect 10770 4113 10800 4167
rect 10770 3973 10800 4027
rect 10870 3973 10900 4167
rect 10970 4113 11000 4307
rect 11070 4253 11100 4307
rect 11170 4253 11200 4447
rect 11270 4393 11300 4587
rect 11370 4533 11400 4587
rect 11470 4533 11500 4587
rect 11570 4533 11600 4587
rect 11670 4533 11700 4587
rect 11770 4533 11800 4587
rect 11870 4533 11900 4587
rect 11970 4533 12000 4587
rect 12070 4533 12100 4587
rect 12170 4533 12200 4587
rect 12270 4533 12300 4587
rect 12370 4533 12400 4587
rect 11370 4393 11400 4447
rect 11470 4393 11500 4447
rect 11570 4393 11600 4447
rect 11670 4393 11700 4447
rect 11770 4393 11800 4447
rect 11870 4393 11900 4447
rect 11270 4253 11300 4307
rect 11070 4113 11100 4167
rect 11170 4113 11200 4167
rect 11270 4113 11300 4167
rect 10970 3973 11000 4027
rect 9670 3833 9700 3887
rect 9770 3833 9800 3887
rect 9870 3833 9900 3887
rect 9970 3833 10000 3887
rect 9570 3710 9600 3747
rect 9470 3700 9600 3710
rect 9470 3666 9518 3700
rect 9552 3666 9600 3700
rect 9470 3656 9600 3666
rect 9470 3603 9500 3656
rect 9570 3603 9600 3656
rect 9670 3694 9700 3747
rect 9770 3694 9800 3747
rect 9670 3684 9800 3694
rect 9670 3650 9718 3684
rect 9752 3650 9800 3684
rect 9670 3640 9800 3650
rect 9670 3603 9700 3640
rect 9770 3603 9800 3640
rect 9870 3710 9900 3747
rect 9970 3710 10000 3747
rect 9870 3700 10000 3710
rect 9870 3666 9918 3700
rect 9952 3666 10000 3700
rect 9870 3656 10000 3666
rect 9870 3603 9900 3656
rect 9970 3603 10000 3656
rect 10070 3694 10100 3887
rect 10170 3833 10200 3887
rect 10270 3833 10300 3887
rect 10370 3833 10400 3887
rect 10470 3833 10500 3887
rect 10570 3833 10600 3887
rect 10670 3833 10700 3887
rect 10770 3833 10800 3887
rect 10870 3833 10900 3887
rect 10970 3833 11000 3887
rect 11070 3833 11100 4027
rect 11170 3973 11200 4027
rect 11270 3973 11300 4027
rect 11370 3973 11400 4307
rect 11470 4253 11500 4307
rect 11470 4113 11500 4167
rect 11470 3973 11500 4027
rect 11570 3973 11600 4307
rect 11670 4253 11700 4307
rect 11770 4253 11800 4307
rect 11870 4253 11900 4307
rect 11970 4253 12000 4447
rect 12070 4393 12100 4447
rect 12170 4393 12200 4447
rect 12270 4393 12300 4447
rect 12370 4393 12400 4447
rect 12470 4393 12500 4587
rect 12570 4533 12600 4587
rect 12670 4533 12700 4727
rect 12770 4673 12800 4727
rect 12970 4673 13000 4727
rect 13070 4673 13100 4727
rect 13280 4673 13310 4727
rect 13380 4673 13410 4727
rect 13480 4673 13510 4727
rect 13580 4673 13610 4727
rect 12770 4533 12800 4587
rect 12970 4533 13000 4587
rect 13070 4533 13100 4587
rect 13280 4533 13310 4587
rect 13380 4533 13410 4587
rect 13480 4533 13510 4587
rect 13580 4533 13610 4587
rect 12570 4393 12600 4447
rect 12670 4393 12700 4447
rect 12770 4393 12800 4447
rect 12970 4393 13000 4447
rect 13070 4393 13100 4447
rect 13280 4393 13310 4447
rect 13380 4393 13410 4447
rect 13480 4393 13510 4447
rect 13580 4393 13610 4447
rect 12070 4253 12100 4307
rect 12170 4253 12200 4307
rect 12270 4253 12300 4307
rect 12370 4253 12400 4307
rect 12470 4253 12500 4307
rect 12570 4253 12600 4307
rect 12670 4253 12700 4307
rect 12770 4253 12800 4307
rect 12970 4253 13000 4307
rect 13070 4253 13100 4307
rect 13280 4253 13310 4307
rect 13380 4253 13410 4307
rect 13480 4253 13510 4307
rect 13580 4253 13610 4307
rect 11670 4113 11700 4167
rect 11770 4113 11800 4167
rect 11670 3973 11700 4027
rect 11770 3973 11800 4027
rect 11870 3973 11900 4167
rect 11970 4113 12000 4167
rect 12070 4113 12100 4167
rect 12170 4113 12200 4167
rect 12270 4113 12300 4167
rect 12370 4113 12400 4167
rect 12470 4113 12500 4167
rect 12570 4113 12600 4167
rect 11970 3973 12000 4027
rect 12070 3973 12100 4027
rect 12170 3973 12200 4027
rect 12270 3973 12300 4027
rect 12370 3973 12400 4027
rect 12470 3973 12500 4027
rect 12570 3973 12600 4027
rect 12670 3973 12700 4167
rect 12770 4113 12800 4167
rect 12970 4113 13000 4167
rect 13070 4113 13100 4167
rect 13280 4113 13310 4167
rect 13380 4113 13410 4167
rect 13480 4113 13510 4167
rect 13580 4113 13610 4167
rect 12770 3973 12800 4027
rect 12970 3973 13000 4027
rect 13070 3973 13100 4027
rect 13280 3973 13310 4027
rect 13380 3973 13410 4027
rect 13480 3973 13510 4027
rect 13580 3973 13610 4027
rect 10170 3694 10200 3747
rect 10070 3684 10200 3694
rect 10070 3650 10118 3684
rect 10152 3650 10200 3684
rect 10070 3640 10200 3650
rect 6870 3323 6900 3377
rect 6970 3323 7000 3377
rect 7070 3323 7100 3377
rect 7170 3323 7200 3377
rect 7270 3323 7300 3377
rect 3570 3183 3600 3237
rect 3370 3043 3400 3097
rect 3470 3043 3500 3097
rect 3570 3043 3600 3097
rect 3670 3043 3700 3237
rect 3770 3183 3800 3237
rect 3870 3183 3900 3237
rect 3970 3183 4000 3237
rect 4070 3183 4100 3237
rect 4170 3183 4200 3237
rect 4270 3183 4300 3237
rect 4370 3183 4400 3237
rect 4470 3183 4500 3237
rect 4570 3183 4600 3237
rect 4670 3183 4700 3237
rect 4770 3183 4800 3237
rect 4870 3183 4900 3237
rect 4970 3183 5000 3237
rect 5070 3183 5100 3237
rect 5170 3183 5200 3237
rect 5270 3183 5300 3237
rect 5370 3183 5400 3237
rect 3770 3043 3800 3097
rect 3170 2903 3200 2957
rect 3270 2903 3300 2957
rect 3070 2763 3100 2817
rect 3170 2763 3200 2817
rect 3270 2763 3300 2817
rect 3370 2763 3400 2957
rect 3470 2903 3500 2957
rect 3570 2903 3600 2957
rect 3670 2903 3700 2957
rect 3770 2903 3800 2957
rect 3870 2903 3900 3097
rect 3970 3043 4000 3097
rect 4070 3043 4100 3097
rect 4170 3043 4200 3097
rect 4270 3043 4300 3097
rect 4370 3043 4400 3097
rect 4470 3043 4500 3097
rect 3470 2763 3500 2817
rect 3570 2763 3600 2817
rect 3670 2763 3700 2817
rect 3770 2763 3800 2817
rect 3870 2763 3900 2817
rect 3970 2763 4000 2957
rect 4070 2903 4100 2957
rect 4170 2903 4200 2957
rect 4270 2903 4300 2957
rect 4370 2903 4400 2957
rect 4470 2903 4500 2957
rect 4570 2903 4600 3097
rect 4670 3043 4700 3097
rect 4770 3043 4800 3097
rect 4870 3043 4900 3097
rect 4670 2903 4700 2957
rect 4770 2903 4800 2957
rect 4870 2903 4900 2957
rect 4970 2903 5000 3097
rect 5070 3043 5100 3097
rect 5170 3043 5200 3097
rect 5270 3043 5300 3097
rect 5370 3043 5400 3097
rect 5470 3043 5500 3237
rect 5570 3183 5600 3237
rect 5570 3043 5600 3097
rect 5670 3043 5700 3237
rect 5770 3183 5800 3237
rect 5770 3043 5800 3097
rect 5870 3043 5900 3237
rect 5970 3183 6000 3237
rect 6070 3183 6100 3237
rect 6170 3183 6200 3237
rect 6270 3183 6300 3237
rect 5070 2903 5100 2957
rect 5170 2903 5200 2957
rect 5270 2903 5300 2957
rect 4070 2763 4100 2817
rect 2470 2623 2500 2677
rect 70 2484 100 2537
rect 170 2484 200 2537
rect 70 2474 200 2484
rect 70 2440 118 2474
rect 152 2440 200 2474
rect 70 2430 200 2440
rect 70 2393 100 2430
rect 70 2253 100 2307
rect 170 2253 200 2430
rect 270 2500 300 2537
rect 370 2500 400 2537
rect 270 2490 400 2500
rect 270 2456 318 2490
rect 352 2456 400 2490
rect 270 2446 400 2456
rect 270 2393 300 2446
rect 370 2393 400 2446
rect 470 2484 500 2537
rect 570 2484 600 2537
rect 470 2474 600 2484
rect 470 2440 518 2474
rect 552 2440 600 2474
rect 470 2430 600 2440
rect 270 2253 300 2307
rect 370 2253 400 2307
rect 470 2253 500 2430
rect 570 2393 600 2430
rect 670 2500 700 2537
rect 770 2500 800 2537
rect 670 2490 800 2500
rect 670 2456 718 2490
rect 752 2456 800 2490
rect 670 2446 800 2456
rect 570 2253 600 2307
rect 670 2253 700 2446
rect 770 2393 800 2446
rect 870 2484 900 2537
rect 970 2484 1000 2537
rect 870 2474 1000 2484
rect 870 2440 918 2474
rect 952 2440 1000 2474
rect 870 2430 1000 2440
rect 870 2393 900 2430
rect 970 2393 1000 2430
rect 1070 2500 1100 2537
rect 1170 2500 1200 2537
rect 1070 2490 1200 2500
rect 1070 2456 1118 2490
rect 1152 2456 1200 2490
rect 1070 2446 1200 2456
rect 1070 2393 1100 2446
rect 1170 2393 1200 2446
rect 1270 2484 1300 2537
rect 1370 2484 1400 2537
rect 1270 2474 1400 2484
rect 1270 2440 1318 2474
rect 1352 2440 1400 2474
rect 1270 2430 1400 2440
rect 1270 2393 1300 2430
rect 1370 2393 1400 2430
rect 1470 2500 1500 2537
rect 1570 2500 1600 2537
rect 1470 2490 1600 2500
rect 1470 2456 1518 2490
rect 1552 2456 1600 2490
rect 1470 2446 1600 2456
rect 1470 2393 1500 2446
rect 1570 2393 1600 2446
rect 1670 2484 1700 2537
rect 1770 2484 1800 2537
rect 1670 2474 1800 2484
rect 1670 2440 1718 2474
rect 1752 2440 1800 2474
rect 1670 2430 1800 2440
rect 1670 2393 1700 2430
rect 1770 2393 1800 2430
rect 1870 2500 1900 2537
rect 1970 2500 2000 2537
rect 1870 2490 2000 2500
rect 1870 2456 1918 2490
rect 1952 2456 2000 2490
rect 1870 2446 2000 2456
rect 1870 2393 1900 2446
rect 1970 2393 2000 2446
rect 2070 2484 2100 2537
rect 2170 2484 2200 2537
rect 2070 2474 2200 2484
rect 2070 2440 2118 2474
rect 2152 2440 2200 2474
rect 2070 2430 2200 2440
rect 2070 2393 2100 2430
rect 2170 2393 2200 2430
rect 2270 2500 2300 2537
rect 2370 2500 2400 2537
rect 2270 2490 2400 2500
rect 2270 2456 2318 2490
rect 2352 2456 2400 2490
rect 2270 2446 2400 2456
rect 2270 2393 2300 2446
rect 770 2253 800 2307
rect 70 2113 100 2167
rect 170 2113 200 2167
rect 270 2113 300 2167
rect 370 2113 400 2167
rect 470 2113 500 2167
rect 570 2113 600 2167
rect 670 2113 700 2167
rect 70 1973 100 2027
rect 170 1973 200 2027
rect 270 1973 300 2027
rect 370 1973 400 2027
rect 470 1973 500 2027
rect 570 1973 600 2027
rect 670 1973 700 2027
rect 770 1973 800 2167
rect 870 2113 900 2307
rect 970 2253 1000 2307
rect 970 2113 1000 2167
rect 1070 2113 1100 2307
rect 1170 2253 1200 2307
rect 1270 2253 1300 2307
rect 1370 2253 1400 2307
rect 1470 2253 1500 2307
rect 1570 2253 1600 2307
rect 1670 2253 1700 2307
rect 1770 2253 1800 2307
rect 1870 2253 1900 2307
rect 1970 2253 2000 2307
rect 2070 2253 2100 2307
rect 2170 2253 2200 2307
rect 2270 2253 2300 2307
rect 2370 2253 2400 2446
rect 2470 2484 2500 2537
rect 2570 2484 2600 2677
rect 2670 2623 2700 2677
rect 2770 2623 2800 2677
rect 2870 2623 2900 2677
rect 2970 2623 3000 2677
rect 3070 2623 3100 2677
rect 3170 2623 3200 2677
rect 3270 2623 3300 2677
rect 2470 2474 2600 2484
rect 2470 2440 2518 2474
rect 2552 2440 2600 2474
rect 2470 2430 2600 2440
rect 2470 2393 2500 2430
rect 2570 2393 2600 2430
rect 2670 2500 2700 2537
rect 2770 2500 2800 2537
rect 2670 2490 2800 2500
rect 2670 2456 2718 2490
rect 2752 2456 2800 2490
rect 2670 2446 2800 2456
rect 2470 2253 2500 2307
rect 2570 2253 2600 2307
rect 1170 2113 1200 2167
rect 1270 2113 1300 2167
rect 1370 2113 1400 2167
rect 870 1973 900 2027
rect 70 1833 100 1887
rect 170 1833 200 1887
rect 270 1833 300 1887
rect 370 1833 400 1887
rect 470 1833 500 1887
rect 570 1833 600 1887
rect 670 1833 700 1887
rect 770 1833 800 1887
rect 870 1833 900 1887
rect 970 1833 1000 2027
rect 1070 1973 1100 2027
rect 1170 1973 1200 2027
rect 1270 1973 1300 2027
rect 1370 1973 1400 2027
rect 1470 1973 1500 2167
rect 1570 2113 1600 2167
rect 1670 2113 1700 2167
rect 1770 2113 1800 2167
rect 1870 2113 1900 2167
rect 1970 2113 2000 2167
rect 2070 2113 2100 2167
rect 2170 2113 2200 2167
rect 2270 2113 2300 2167
rect 2370 2113 2400 2167
rect 2470 2113 2500 2167
rect 2570 2113 2600 2167
rect 2670 2113 2700 2446
rect 2770 2393 2800 2446
rect 2870 2484 2900 2537
rect 2970 2484 3000 2537
rect 2870 2474 3000 2484
rect 2870 2440 2918 2474
rect 2952 2440 3000 2474
rect 2870 2430 3000 2440
rect 2870 2393 2900 2430
rect 2970 2393 3000 2430
rect 3070 2500 3100 2537
rect 3170 2500 3200 2537
rect 3070 2490 3200 2500
rect 3070 2456 3118 2490
rect 3152 2456 3200 2490
rect 3070 2446 3200 2456
rect 3070 2393 3100 2446
rect 3170 2393 3200 2446
rect 3270 2484 3300 2537
rect 3370 2484 3400 2677
rect 3470 2623 3500 2677
rect 3570 2623 3600 2677
rect 3670 2623 3700 2677
rect 3770 2623 3800 2677
rect 3870 2623 3900 2677
rect 3270 2474 3400 2484
rect 3270 2440 3318 2474
rect 3352 2440 3400 2474
rect 3270 2430 3400 2440
rect 3270 2393 3300 2430
rect 3370 2393 3400 2430
rect 3470 2500 3500 2537
rect 3570 2500 3600 2537
rect 3470 2490 3600 2500
rect 3470 2456 3518 2490
rect 3552 2456 3600 2490
rect 3470 2446 3600 2456
rect 3470 2393 3500 2446
rect 3570 2393 3600 2446
rect 3670 2484 3700 2537
rect 3770 2484 3800 2537
rect 3670 2474 3800 2484
rect 3670 2440 3718 2474
rect 3752 2440 3800 2474
rect 3670 2430 3800 2440
rect 3670 2393 3700 2430
rect 3770 2393 3800 2430
rect 3870 2500 3900 2537
rect 3970 2500 4000 2677
rect 4070 2623 4100 2677
rect 3870 2490 4000 2500
rect 3870 2456 3918 2490
rect 3952 2456 4000 2490
rect 3870 2446 4000 2456
rect 3870 2393 3900 2446
rect 3970 2393 4000 2446
rect 4070 2484 4100 2537
rect 4170 2484 4200 2817
rect 4270 2763 4300 2817
rect 4370 2763 4400 2817
rect 4470 2763 4500 2817
rect 4570 2763 4600 2817
rect 4670 2763 4700 2817
rect 4270 2623 4300 2677
rect 4070 2474 4200 2484
rect 4070 2440 4118 2474
rect 4152 2440 4200 2474
rect 4070 2430 4200 2440
rect 4070 2393 4100 2430
rect 4170 2393 4200 2430
rect 4270 2500 4300 2537
rect 4370 2500 4400 2677
rect 4470 2623 4500 2677
rect 4570 2623 4600 2677
rect 4670 2623 4700 2677
rect 4270 2490 4400 2500
rect 4270 2456 4318 2490
rect 4352 2456 4400 2490
rect 4270 2446 4400 2456
rect 4270 2393 4300 2446
rect 4370 2393 4400 2446
rect 4470 2484 4500 2537
rect 4570 2484 4600 2537
rect 4470 2474 4600 2484
rect 4470 2440 4518 2474
rect 4552 2440 4600 2474
rect 4470 2430 4600 2440
rect 4470 2393 4500 2430
rect 4570 2393 4600 2430
rect 4670 2500 4700 2537
rect 4770 2500 4800 2817
rect 4870 2763 4900 2817
rect 4970 2763 5000 2817
rect 5070 2763 5100 2817
rect 4870 2623 4900 2677
rect 4970 2623 5000 2677
rect 5070 2623 5100 2677
rect 5170 2623 5200 2817
rect 5270 2763 5300 2817
rect 5270 2623 5300 2677
rect 5370 2623 5400 2957
rect 5470 2903 5500 2957
rect 5570 2903 5600 2957
rect 5670 2903 5700 2957
rect 5770 2903 5800 2957
rect 5870 2903 5900 2957
rect 5970 2903 6000 3097
rect 6070 3043 6100 3097
rect 6170 3043 6200 3097
rect 6270 3043 6300 3097
rect 6370 3043 6400 3237
rect 6470 3183 6500 3237
rect 6470 3043 6500 3097
rect 6570 3043 6600 3237
rect 6670 3183 6700 3237
rect 6770 3183 6800 3237
rect 6870 3183 6900 3237
rect 6970 3183 7000 3237
rect 6670 3043 6700 3097
rect 6770 3043 6800 3097
rect 6870 3043 6900 3097
rect 6970 3043 7000 3097
rect 7070 3043 7100 3237
rect 7170 3183 7200 3237
rect 7270 3183 7300 3237
rect 7370 3183 7400 3377
rect 7470 3323 7500 3377
rect 7570 3323 7600 3377
rect 7670 3323 7700 3377
rect 7770 3323 7800 3377
rect 7870 3323 7900 3377
rect 7970 3323 8000 3377
rect 8070 3323 8100 3377
rect 8170 3323 8200 3377
rect 8270 3323 8300 3377
rect 8370 3323 8400 3377
rect 8470 3323 8500 3377
rect 8570 3323 8600 3377
rect 8670 3323 8700 3377
rect 8770 3323 8800 3377
rect 8870 3323 8900 3377
rect 8970 3323 9000 3377
rect 9070 3323 9100 3377
rect 9170 3323 9200 3377
rect 9270 3323 9300 3377
rect 9370 3323 9400 3377
rect 9470 3323 9500 3517
rect 9570 3463 9600 3517
rect 9670 3463 9700 3517
rect 7470 3183 7500 3237
rect 7570 3183 7600 3237
rect 7670 3183 7700 3237
rect 7770 3183 7800 3237
rect 7870 3183 7900 3237
rect 7970 3183 8000 3237
rect 8070 3183 8100 3237
rect 7170 3043 7200 3097
rect 7270 3043 7300 3097
rect 7370 3043 7400 3097
rect 7470 3043 7500 3097
rect 7570 3043 7600 3097
rect 7670 3043 7700 3097
rect 7770 3043 7800 3097
rect 7870 3043 7900 3097
rect 7970 3043 8000 3097
rect 5470 2763 5500 2817
rect 5570 2763 5600 2817
rect 5670 2763 5700 2817
rect 5770 2763 5800 2817
rect 5870 2763 5900 2817
rect 5970 2763 6000 2817
rect 5470 2623 5500 2677
rect 5570 2623 5600 2677
rect 5670 2623 5700 2677
rect 5770 2623 5800 2677
rect 5870 2623 5900 2677
rect 5970 2623 6000 2677
rect 6070 2623 6100 2957
rect 6170 2903 6200 2957
rect 6270 2903 6300 2957
rect 6370 2903 6400 2957
rect 6470 2903 6500 2957
rect 6570 2903 6600 2957
rect 6670 2903 6700 2957
rect 6770 2903 6800 2957
rect 6870 2903 6900 2957
rect 6170 2763 6200 2817
rect 6170 2623 6200 2677
rect 4670 2490 4800 2500
rect 4670 2456 4718 2490
rect 4752 2456 4800 2490
rect 4670 2446 4800 2456
rect 4670 2393 4700 2446
rect 4770 2393 4800 2446
rect 4870 2484 4900 2537
rect 4970 2484 5000 2537
rect 4870 2474 5000 2484
rect 4870 2440 4918 2474
rect 4952 2440 5000 2474
rect 4870 2430 5000 2440
rect 4870 2393 4900 2430
rect 4970 2393 5000 2430
rect 5070 2500 5100 2537
rect 5170 2500 5200 2537
rect 5070 2490 5200 2500
rect 5070 2456 5118 2490
rect 5152 2456 5200 2490
rect 5070 2446 5200 2456
rect 5070 2393 5100 2446
rect 5170 2393 5200 2446
rect 5270 2484 5300 2537
rect 5370 2484 5400 2537
rect 5270 2474 5400 2484
rect 5270 2440 5318 2474
rect 5352 2440 5400 2474
rect 5270 2430 5400 2440
rect 5270 2393 5300 2430
rect 5370 2393 5400 2430
rect 5470 2500 5500 2537
rect 5570 2500 5600 2537
rect 5470 2490 5600 2500
rect 5470 2456 5518 2490
rect 5552 2456 5600 2490
rect 5470 2446 5600 2456
rect 5470 2393 5500 2446
rect 5570 2393 5600 2446
rect 5670 2484 5700 2537
rect 5770 2484 5800 2537
rect 5670 2474 5800 2484
rect 5670 2440 5718 2474
rect 5752 2440 5800 2474
rect 5670 2430 5800 2440
rect 5670 2393 5700 2430
rect 5770 2393 5800 2430
rect 5870 2500 5900 2537
rect 5970 2500 6000 2537
rect 5870 2490 6000 2500
rect 5870 2456 5918 2490
rect 5952 2456 6000 2490
rect 5870 2446 6000 2456
rect 5870 2393 5900 2446
rect 5970 2393 6000 2446
rect 6070 2484 6100 2537
rect 6170 2484 6200 2537
rect 6070 2474 6200 2484
rect 6070 2440 6118 2474
rect 6152 2440 6200 2474
rect 6070 2430 6200 2440
rect 6070 2393 6100 2430
rect 6170 2393 6200 2430
rect 6270 2500 6300 2817
rect 6370 2763 6400 2817
rect 6470 2763 6500 2817
rect 6370 2623 6400 2677
rect 6470 2623 6500 2677
rect 6570 2623 6600 2817
rect 6670 2763 6700 2817
rect 6770 2763 6800 2817
rect 6870 2763 6900 2817
rect 6970 2763 7000 2957
rect 7070 2903 7100 2957
rect 7170 2903 7200 2957
rect 7270 2903 7300 2957
rect 7070 2763 7100 2817
rect 7170 2763 7200 2817
rect 7270 2763 7300 2817
rect 7370 2763 7400 2957
rect 7470 2903 7500 2957
rect 7570 2903 7600 2957
rect 7670 2903 7700 2957
rect 7770 2903 7800 2957
rect 7870 2903 7900 2957
rect 7470 2763 7500 2817
rect 7570 2763 7600 2817
rect 7670 2763 7700 2817
rect 7770 2763 7800 2817
rect 7870 2763 7900 2817
rect 7970 2763 8000 2957
rect 8070 2903 8100 3097
rect 8170 3043 8200 3237
rect 8270 3183 8300 3237
rect 8370 3183 8400 3237
rect 8470 3183 8500 3237
rect 8570 3183 8600 3237
rect 8670 3183 8700 3237
rect 8770 3183 8800 3237
rect 8270 3043 8300 3097
rect 8370 3043 8400 3097
rect 8470 3043 8500 3097
rect 8570 3043 8600 3097
rect 8670 3043 8700 3097
rect 8770 3043 8800 3097
rect 8170 2903 8200 2957
rect 8270 2903 8300 2957
rect 8370 2903 8400 2957
rect 8470 2903 8500 2957
rect 8570 2903 8600 2957
rect 8670 2903 8700 2957
rect 8070 2763 8100 2817
rect 8170 2763 8200 2817
rect 6670 2623 6700 2677
rect 6370 2500 6400 2537
rect 6270 2490 6400 2500
rect 6270 2456 6318 2490
rect 6352 2456 6400 2490
rect 6270 2446 6400 2456
rect 6270 2393 6300 2446
rect 6370 2393 6400 2446
rect 6470 2484 6500 2537
rect 6570 2484 6600 2537
rect 6470 2474 6600 2484
rect 6470 2440 6518 2474
rect 6552 2440 6600 2474
rect 6470 2430 6600 2440
rect 6470 2393 6500 2430
rect 6570 2393 6600 2430
rect 6670 2500 6700 2537
rect 6770 2500 6800 2677
rect 6870 2623 6900 2677
rect 6970 2623 7000 2677
rect 7070 2623 7100 2677
rect 7170 2623 7200 2677
rect 7270 2623 7300 2677
rect 7370 2623 7400 2677
rect 7470 2623 7500 2677
rect 7570 2623 7600 2677
rect 7670 2623 7700 2677
rect 7770 2623 7800 2677
rect 7870 2623 7900 2677
rect 7970 2623 8000 2677
rect 8070 2623 8100 2677
rect 8170 2623 8200 2677
rect 6670 2490 6800 2500
rect 6670 2456 6718 2490
rect 6752 2456 6800 2490
rect 6670 2446 6800 2456
rect 6670 2393 6700 2446
rect 6770 2393 6800 2446
rect 6870 2484 6900 2537
rect 6970 2484 7000 2537
rect 6870 2474 7000 2484
rect 6870 2440 6918 2474
rect 6952 2440 7000 2474
rect 6870 2430 7000 2440
rect 6870 2393 6900 2430
rect 2770 2253 2800 2307
rect 1070 1833 1100 1887
rect 1170 1833 1200 1887
rect 1270 1833 1300 1887
rect 1370 1833 1400 1887
rect 1470 1833 1500 1887
rect 1570 1833 1600 2027
rect 1670 1973 1700 2027
rect 1770 1973 1800 2027
rect 1870 1973 1900 2027
rect 1970 1973 2000 2027
rect 2070 1973 2100 2027
rect 2170 1973 2200 2027
rect 2270 1973 2300 2027
rect 2370 1973 2400 2027
rect 2470 1973 2500 2027
rect 2570 1973 2600 2027
rect 2670 1973 2700 2027
rect 2770 1973 2800 2167
rect 2870 2113 2900 2307
rect 2970 2253 3000 2307
rect 2870 1973 2900 2027
rect 2970 1973 3000 2167
rect 3070 2113 3100 2307
rect 3170 2253 3200 2307
rect 3270 2253 3300 2307
rect 3170 2113 3200 2167
rect 3270 2113 3300 2167
rect 3370 2113 3400 2307
rect 3470 2253 3500 2307
rect 3570 2253 3600 2307
rect 3470 2113 3500 2167
rect 3070 1973 3100 2027
rect 3170 1973 3200 2027
rect 3270 1973 3300 2027
rect 3370 1973 3400 2027
rect 3470 1973 3500 2027
rect 3570 1973 3600 2167
rect 3670 2113 3700 2307
rect 3770 2253 3800 2307
rect 3770 2113 3800 2167
rect 3870 2113 3900 2307
rect 3970 2253 4000 2307
rect 4070 2253 4100 2307
rect 4170 2253 4200 2307
rect 4270 2253 4300 2307
rect 3970 2113 4000 2167
rect 4070 2113 4100 2167
rect 4170 2113 4200 2167
rect 4270 2113 4300 2167
rect 4370 2113 4400 2307
rect 4470 2253 4500 2307
rect 4570 2253 4600 2307
rect 4670 2253 4700 2307
rect 4770 2253 4800 2307
rect 4870 2253 4900 2307
rect 4970 2253 5000 2307
rect 5070 2253 5100 2307
rect 5170 2253 5200 2307
rect 5270 2253 5300 2307
rect 5370 2253 5400 2307
rect 5470 2253 5500 2307
rect 5570 2253 5600 2307
rect 5670 2253 5700 2307
rect 5770 2253 5800 2307
rect 5870 2253 5900 2307
rect 5970 2253 6000 2307
rect 6070 2253 6100 2307
rect 4470 2113 4500 2167
rect 4570 2113 4600 2167
rect 1670 1833 1700 1887
rect 1770 1833 1800 1887
rect 1870 1833 1900 1887
rect 1970 1833 2000 1887
rect 2070 1833 2100 1887
rect 2170 1833 2200 1887
rect 2270 1833 2300 1887
rect 2370 1833 2400 1887
rect 2470 1833 2500 1887
rect 2570 1833 2600 1887
rect 2670 1833 2700 1887
rect 2770 1833 2800 1887
rect 2870 1833 2900 1887
rect 2970 1833 3000 1887
rect 3070 1833 3100 1887
rect 70 1693 100 1747
rect 170 1693 200 1747
rect 270 1693 300 1747
rect 370 1693 400 1747
rect 470 1693 500 1747
rect 570 1693 600 1747
rect 70 1553 100 1607
rect 170 1553 200 1607
rect 270 1553 300 1607
rect 370 1553 400 1607
rect 70 1413 100 1467
rect 170 1413 200 1467
rect 270 1413 300 1467
rect 370 1413 400 1467
rect 470 1413 500 1607
rect 570 1553 600 1607
rect 670 1553 700 1747
rect 770 1693 800 1747
rect 870 1693 900 1747
rect 970 1693 1000 1747
rect 770 1553 800 1607
rect 870 1553 900 1607
rect 970 1553 1000 1607
rect 1070 1553 1100 1747
rect 1170 1693 1200 1747
rect 1170 1553 1200 1607
rect 1270 1553 1300 1747
rect 1370 1693 1400 1747
rect 1470 1693 1500 1747
rect 1370 1553 1400 1607
rect 1470 1553 1500 1607
rect 1570 1553 1600 1747
rect 1670 1693 1700 1747
rect 1770 1693 1800 1747
rect 1870 1693 1900 1747
rect 1970 1693 2000 1747
rect 2070 1693 2100 1747
rect 2170 1693 2200 1747
rect 2270 1693 2300 1747
rect 2370 1693 2400 1747
rect 2470 1693 2500 1747
rect 2570 1693 2600 1747
rect 1670 1553 1700 1607
rect 1770 1553 1800 1607
rect 1870 1553 1900 1607
rect 1970 1553 2000 1607
rect 2070 1553 2100 1607
rect 2170 1553 2200 1607
rect 2270 1553 2300 1607
rect 2370 1553 2400 1607
rect 2470 1553 2500 1607
rect 570 1413 600 1467
rect 670 1413 700 1467
rect 770 1413 800 1467
rect 70 1274 100 1327
rect 170 1274 200 1327
rect 70 1264 200 1274
rect 70 1230 118 1264
rect 152 1230 200 1264
rect 70 1220 200 1230
rect 70 1183 100 1220
rect 170 1183 200 1220
rect 270 1290 300 1327
rect 370 1290 400 1327
rect 270 1280 400 1290
rect 270 1246 318 1280
rect 352 1246 400 1280
rect 270 1236 400 1246
rect 270 1183 300 1236
rect 370 1183 400 1236
rect 470 1274 500 1327
rect 570 1274 600 1327
rect 470 1264 600 1274
rect 470 1230 518 1264
rect 552 1230 600 1264
rect 470 1220 600 1230
rect 470 1183 500 1220
rect 570 1183 600 1220
rect 670 1290 700 1327
rect 770 1290 800 1327
rect 670 1280 800 1290
rect 670 1246 718 1280
rect 752 1246 800 1280
rect 670 1236 800 1246
rect 670 1183 700 1236
rect 770 1183 800 1236
rect 870 1274 900 1467
rect 970 1413 1000 1467
rect 1070 1413 1100 1467
rect 1170 1413 1200 1467
rect 1270 1413 1300 1467
rect 1370 1413 1400 1467
rect 1470 1413 1500 1467
rect 1570 1413 1600 1467
rect 1670 1413 1700 1467
rect 1770 1413 1800 1467
rect 1870 1413 1900 1467
rect 1970 1413 2000 1467
rect 2070 1413 2100 1467
rect 2170 1413 2200 1467
rect 2270 1413 2300 1467
rect 2370 1413 2400 1467
rect 2470 1413 2500 1467
rect 2570 1413 2600 1607
rect 2670 1553 2700 1747
rect 2770 1693 2800 1747
rect 2870 1693 2900 1747
rect 2970 1693 3000 1747
rect 3070 1693 3100 1747
rect 3170 1693 3200 1887
rect 3270 1833 3300 1887
rect 3270 1693 3300 1747
rect 3370 1693 3400 1887
rect 3470 1833 3500 1887
rect 3570 1833 3600 1887
rect 3670 1833 3700 2027
rect 3770 1973 3800 2027
rect 3870 1973 3900 2027
rect 3970 1973 4000 2027
rect 4070 1973 4100 2027
rect 4170 1973 4200 2027
rect 3770 1833 3800 1887
rect 3870 1833 3900 1887
rect 3470 1693 3500 1747
rect 3570 1693 3600 1747
rect 3670 1693 3700 1747
rect 2770 1553 2800 1607
rect 2870 1553 2900 1607
rect 2970 1553 3000 1607
rect 3070 1553 3100 1607
rect 2670 1413 2700 1467
rect 2770 1413 2800 1467
rect 970 1274 1000 1327
rect 870 1264 1000 1274
rect 870 1230 918 1264
rect 952 1230 1000 1264
rect 870 1220 1000 1230
rect 870 1183 900 1220
rect 970 1183 1000 1220
rect 1070 1290 1100 1327
rect 1170 1290 1200 1327
rect 1070 1280 1200 1290
rect 1070 1246 1118 1280
rect 1152 1246 1200 1280
rect 1070 1236 1200 1246
rect 1070 1183 1100 1236
rect 1170 1183 1200 1236
rect 1270 1274 1300 1327
rect 1370 1274 1400 1327
rect 1270 1264 1400 1274
rect 1270 1230 1318 1264
rect 1352 1230 1400 1264
rect 1270 1220 1400 1230
rect 1270 1183 1300 1220
rect 1370 1183 1400 1220
rect 1470 1290 1500 1327
rect 1570 1290 1600 1327
rect 1470 1280 1600 1290
rect 1470 1246 1518 1280
rect 1552 1246 1600 1280
rect 1470 1236 1600 1246
rect 1470 1183 1500 1236
rect 1570 1183 1600 1236
rect 1670 1274 1700 1327
rect 1770 1274 1800 1327
rect 1670 1264 1800 1274
rect 1670 1230 1718 1264
rect 1752 1230 1800 1264
rect 1670 1220 1800 1230
rect 1670 1183 1700 1220
rect 70 1043 100 1097
rect 70 903 100 957
rect 70 763 100 817
rect 170 763 200 1097
rect 270 1043 300 1097
rect 370 1043 400 1097
rect 470 1043 500 1097
rect 570 1043 600 1097
rect 270 903 300 957
rect 370 903 400 957
rect 470 903 500 957
rect 570 903 600 957
rect 670 903 700 1097
rect 770 1043 800 1097
rect 870 1043 900 1097
rect 970 1043 1000 1097
rect 1070 1043 1100 1097
rect 1170 1043 1200 1097
rect 770 903 800 957
rect 870 903 900 957
rect 970 903 1000 957
rect 1070 903 1100 957
rect 1170 903 1200 957
rect 1270 903 1300 1097
rect 1370 1043 1400 1097
rect 1470 1043 1500 1097
rect 1570 1043 1600 1097
rect 1670 1043 1700 1097
rect 1770 1043 1800 1220
rect 1870 1290 1900 1327
rect 1970 1290 2000 1327
rect 1870 1280 2000 1290
rect 1870 1246 1918 1280
rect 1952 1246 2000 1280
rect 1870 1236 2000 1246
rect 1870 1183 1900 1236
rect 1970 1183 2000 1236
rect 2070 1274 2100 1327
rect 2170 1274 2200 1327
rect 2070 1264 2200 1274
rect 2070 1230 2118 1264
rect 2152 1230 2200 1264
rect 2070 1220 2200 1230
rect 1870 1043 1900 1097
rect 1970 1043 2000 1097
rect 2070 1043 2100 1220
rect 2170 1183 2200 1220
rect 2270 1290 2300 1327
rect 2370 1290 2400 1327
rect 2270 1280 2400 1290
rect 2270 1246 2318 1280
rect 2352 1246 2400 1280
rect 2270 1236 2400 1246
rect 2270 1183 2300 1236
rect 2370 1183 2400 1236
rect 2470 1274 2500 1327
rect 2570 1274 2600 1327
rect 2470 1264 2600 1274
rect 2470 1230 2518 1264
rect 2552 1230 2600 1264
rect 2470 1220 2600 1230
rect 2470 1183 2500 1220
rect 2570 1183 2600 1220
rect 2670 1290 2700 1327
rect 2770 1290 2800 1327
rect 2670 1280 2800 1290
rect 2670 1246 2718 1280
rect 2752 1246 2800 1280
rect 2670 1236 2800 1246
rect 2670 1183 2700 1236
rect 2770 1183 2800 1236
rect 2870 1274 2900 1467
rect 2970 1413 3000 1467
rect 3070 1413 3100 1467
rect 3170 1413 3200 1607
rect 3270 1553 3300 1607
rect 3370 1553 3400 1607
rect 3470 1553 3500 1607
rect 3270 1413 3300 1467
rect 3370 1413 3400 1467
rect 3470 1413 3500 1467
rect 3570 1413 3600 1607
rect 3670 1553 3700 1607
rect 3770 1553 3800 1747
rect 3870 1693 3900 1747
rect 3870 1553 3900 1607
rect 3970 1553 4000 1887
rect 4070 1833 4100 1887
rect 4070 1693 4100 1747
rect 3670 1413 3700 1467
rect 3770 1413 3800 1467
rect 3870 1413 3900 1467
rect 3970 1413 4000 1467
rect 4070 1413 4100 1607
rect 4170 1553 4200 1887
rect 4270 1833 4300 2027
rect 4370 1973 4400 2027
rect 4370 1833 4400 1887
rect 4470 1833 4500 2027
rect 4570 1973 4600 2027
rect 4570 1833 4600 1887
rect 4670 1833 4700 2167
rect 4770 2113 4800 2167
rect 4870 2113 4900 2167
rect 4770 1973 4800 2027
rect 4870 1973 4900 2027
rect 4970 1973 5000 2167
rect 5070 2113 5100 2167
rect 5170 2113 5200 2167
rect 5270 2113 5300 2167
rect 5370 2113 5400 2167
rect 5470 2113 5500 2167
rect 5570 2113 5600 2167
rect 5670 2113 5700 2167
rect 5070 1973 5100 2027
rect 4770 1833 4800 1887
rect 4270 1693 4300 1747
rect 4370 1693 4400 1747
rect 4270 1553 4300 1607
rect 4370 1553 4400 1607
rect 4470 1553 4500 1747
rect 4570 1693 4600 1747
rect 4670 1693 4700 1747
rect 4770 1693 4800 1747
rect 4870 1693 4900 1887
rect 4970 1833 5000 1887
rect 5070 1833 5100 1887
rect 5170 1833 5200 2027
rect 5270 1973 5300 2027
rect 5370 1973 5400 2027
rect 5470 1973 5500 2027
rect 5570 1973 5600 2027
rect 5670 1973 5700 2027
rect 5270 1833 5300 1887
rect 5370 1833 5400 1887
rect 5470 1833 5500 1887
rect 5570 1833 5600 1887
rect 5670 1833 5700 1887
rect 5770 1833 5800 2167
rect 5870 2113 5900 2167
rect 5970 2113 6000 2167
rect 6070 2113 6100 2167
rect 6170 2113 6200 2307
rect 6270 2253 6300 2307
rect 6370 2253 6400 2307
rect 6270 2113 6300 2167
rect 6370 2113 6400 2167
rect 6470 2113 6500 2307
rect 6570 2253 6600 2307
rect 6670 2253 6700 2307
rect 6570 2113 6600 2167
rect 5870 1973 5900 2027
rect 5970 1973 6000 2027
rect 6070 1973 6100 2027
rect 6170 1973 6200 2027
rect 6270 1973 6300 2027
rect 6370 1973 6400 2027
rect 6470 1973 6500 2027
rect 6570 1973 6600 2027
rect 6670 1973 6700 2167
rect 6770 2113 6800 2307
rect 6870 2253 6900 2307
rect 5870 1833 5900 1887
rect 5970 1833 6000 1887
rect 6070 1833 6100 1887
rect 6170 1833 6200 1887
rect 6270 1833 6300 1887
rect 4570 1553 4600 1607
rect 4670 1553 4700 1607
rect 4770 1553 4800 1607
rect 4170 1413 4200 1467
rect 4270 1413 4300 1467
rect 4370 1413 4400 1467
rect 4470 1413 4500 1467
rect 4570 1413 4600 1467
rect 2970 1274 3000 1327
rect 2870 1264 3000 1274
rect 2870 1230 2918 1264
rect 2952 1230 3000 1264
rect 2870 1220 3000 1230
rect 2870 1183 2900 1220
rect 2970 1183 3000 1220
rect 3070 1290 3100 1327
rect 3170 1290 3200 1327
rect 3070 1280 3200 1290
rect 3070 1246 3118 1280
rect 3152 1246 3200 1280
rect 3070 1236 3200 1246
rect 2170 1043 2200 1097
rect 2270 1043 2300 1097
rect 2370 1043 2400 1097
rect 2470 1043 2500 1097
rect 2570 1043 2600 1097
rect 1370 903 1400 957
rect 1470 903 1500 957
rect 1570 903 1600 957
rect 1670 903 1700 957
rect 1770 903 1800 957
rect 1870 903 1900 957
rect 1970 903 2000 957
rect 2070 903 2100 957
rect 2170 903 2200 957
rect 2270 903 2300 957
rect 2370 903 2400 957
rect 2470 903 2500 957
rect 2570 903 2600 957
rect 2670 903 2700 1097
rect 2770 1043 2800 1097
rect 2770 903 2800 957
rect 2870 903 2900 1097
rect 2970 1043 3000 1097
rect 3070 1043 3100 1236
rect 3170 1183 3200 1236
rect 3270 1274 3300 1327
rect 3370 1274 3400 1327
rect 3270 1264 3400 1274
rect 3270 1230 3318 1264
rect 3352 1230 3400 1264
rect 3270 1220 3400 1230
rect 270 763 300 817
rect 370 763 400 817
rect 470 763 500 817
rect 70 623 100 677
rect 170 623 200 677
rect 270 623 300 677
rect 370 623 400 677
rect 470 623 500 677
rect 570 623 600 817
rect 670 763 700 817
rect 670 623 700 677
rect 70 483 100 537
rect 170 483 200 537
rect 270 483 300 537
rect 70 343 100 397
rect 170 343 200 397
rect 270 343 300 397
rect 370 343 400 537
rect 470 483 500 537
rect 570 483 600 537
rect 670 483 700 537
rect 770 483 800 817
rect 870 763 900 817
rect 970 763 1000 817
rect 1070 763 1100 817
rect 1170 763 1200 817
rect 870 623 900 677
rect 970 623 1000 677
rect 1070 623 1100 677
rect 1170 623 1200 677
rect 870 483 900 537
rect 970 483 1000 537
rect 1070 483 1100 537
rect 470 343 500 397
rect 570 343 600 397
rect 670 343 700 397
rect 770 343 800 397
rect 870 343 900 397
rect 970 343 1000 397
rect 1070 343 1100 397
rect 1170 343 1200 537
rect 1270 483 1300 817
rect 1370 763 1400 817
rect 1370 623 1400 677
rect 1470 623 1500 817
rect 1570 763 1600 817
rect 1670 763 1700 817
rect 1770 763 1800 817
rect 1870 763 1900 817
rect 1970 763 2000 817
rect 1570 623 1600 677
rect 1670 623 1700 677
rect 1770 623 1800 677
rect 1870 623 1900 677
rect 1970 623 2000 677
rect 2070 623 2100 817
rect 2170 763 2200 817
rect 2270 763 2300 817
rect 2370 763 2400 817
rect 1370 483 1400 537
rect 1470 483 1500 537
rect 1570 483 1600 537
rect 1670 483 1700 537
rect 1770 483 1800 537
rect 1270 343 1300 397
rect 1370 343 1400 397
rect 1470 343 1500 397
rect 1570 343 1600 397
rect 1670 343 1700 397
rect 70 203 100 257
rect 170 203 200 257
rect 270 203 300 257
rect 370 203 400 257
rect 470 203 500 257
rect 570 203 600 257
rect 670 203 700 257
rect 770 203 800 257
rect 870 203 900 257
rect 970 203 1000 257
rect 1070 203 1100 257
rect 1170 203 1200 257
rect 1270 203 1300 257
rect 1370 203 1400 257
rect 1470 203 1500 257
rect 1570 203 1600 257
rect 70 64 100 117
rect 170 64 200 117
rect 70 54 200 64
rect 70 20 118 54
rect 152 20 200 54
rect 70 10 200 20
rect 70 0 100 10
rect 170 0 200 10
rect 270 80 300 117
rect 370 80 400 117
rect 270 70 400 80
rect 270 36 318 70
rect 352 36 400 70
rect 270 26 400 36
rect 270 0 300 26
rect 370 0 400 26
rect 470 64 500 117
rect 570 64 600 117
rect 470 54 600 64
rect 470 20 518 54
rect 552 20 600 54
rect 470 10 600 20
rect 470 0 500 10
rect 570 0 600 10
rect 670 80 700 117
rect 770 80 800 117
rect 670 70 800 80
rect 670 36 718 70
rect 752 36 800 70
rect 670 26 800 36
rect 670 0 700 26
rect 770 0 800 26
rect 870 64 900 117
rect 970 64 1000 117
rect 870 54 1000 64
rect 870 20 918 54
rect 952 20 1000 54
rect 870 10 1000 20
rect 870 0 900 10
rect 970 0 1000 10
rect 1070 80 1100 117
rect 1170 80 1200 117
rect 1070 70 1200 80
rect 1070 36 1118 70
rect 1152 36 1200 70
rect 1070 26 1200 36
rect 1070 0 1100 26
rect 1170 0 1200 26
rect 1270 64 1300 117
rect 1370 64 1400 117
rect 1270 54 1400 64
rect 1270 20 1318 54
rect 1352 20 1400 54
rect 1270 10 1400 20
rect 1270 0 1300 10
rect 1370 0 1400 10
rect 1470 80 1500 117
rect 1570 80 1600 117
rect 1470 70 1600 80
rect 1470 36 1518 70
rect 1552 36 1600 70
rect 1470 26 1600 36
rect 1470 0 1500 26
rect 1570 0 1600 26
rect 1670 64 1700 257
rect 1770 203 1800 397
rect 1870 343 1900 537
rect 1970 483 2000 537
rect 2070 483 2100 537
rect 2170 483 2200 677
rect 2270 623 2300 677
rect 2370 623 2400 677
rect 2470 623 2500 817
rect 2570 763 2600 817
rect 2670 763 2700 817
rect 2770 763 2800 817
rect 2570 623 2600 677
rect 2670 623 2700 677
rect 2270 483 2300 537
rect 1970 343 2000 397
rect 2070 343 2100 397
rect 2170 343 2200 397
rect 2270 343 2300 397
rect 2370 343 2400 537
rect 2470 483 2500 537
rect 2570 483 2600 537
rect 2470 343 2500 397
rect 2570 343 2600 397
rect 2670 343 2700 537
rect 2770 483 2800 677
rect 2870 623 2900 817
rect 2970 763 3000 957
rect 3070 903 3100 957
rect 3170 903 3200 1097
rect 3270 1043 3300 1220
rect 3370 1183 3400 1220
rect 3470 1290 3500 1327
rect 3570 1290 3600 1327
rect 3470 1280 3600 1290
rect 3470 1246 3518 1280
rect 3552 1246 3600 1280
rect 3470 1236 3600 1246
rect 3470 1183 3500 1236
rect 3570 1183 3600 1236
rect 3670 1274 3700 1327
rect 3770 1274 3800 1327
rect 3670 1264 3800 1274
rect 3670 1230 3718 1264
rect 3752 1230 3800 1264
rect 3670 1220 3800 1230
rect 3670 1183 3700 1220
rect 3270 903 3300 957
rect 3370 903 3400 1097
rect 3470 1043 3500 1097
rect 3570 1043 3600 1097
rect 3470 903 3500 957
rect 3570 903 3600 957
rect 3670 903 3700 1097
rect 3770 1043 3800 1220
rect 3870 1290 3900 1327
rect 3970 1290 4000 1327
rect 3870 1280 4000 1290
rect 3870 1246 3918 1280
rect 3952 1246 4000 1280
rect 3870 1236 4000 1246
rect 3870 1183 3900 1236
rect 3970 1183 4000 1236
rect 4070 1274 4100 1327
rect 4170 1274 4200 1327
rect 4070 1264 4200 1274
rect 4070 1230 4118 1264
rect 4152 1230 4200 1264
rect 4070 1220 4200 1230
rect 4070 1183 4100 1220
rect 4170 1183 4200 1220
rect 4270 1290 4300 1327
rect 4370 1290 4400 1327
rect 4270 1280 4400 1290
rect 4270 1246 4318 1280
rect 4352 1246 4400 1280
rect 4270 1236 4400 1246
rect 4270 1183 4300 1236
rect 4370 1183 4400 1236
rect 4470 1274 4500 1327
rect 4570 1274 4600 1327
rect 4470 1264 4600 1274
rect 4470 1230 4518 1264
rect 4552 1230 4600 1264
rect 4470 1220 4600 1230
rect 3770 903 3800 957
rect 2970 623 3000 677
rect 3070 623 3100 817
rect 3170 763 3200 817
rect 3270 763 3300 817
rect 3170 623 3200 677
rect 3270 623 3300 677
rect 3370 623 3400 817
rect 3470 763 3500 817
rect 3570 763 3600 817
rect 3470 623 3500 677
rect 3570 623 3600 677
rect 3670 623 3700 817
rect 3770 763 3800 817
rect 3870 763 3900 1097
rect 3970 1043 4000 1097
rect 4070 1043 4100 1097
rect 4170 1043 4200 1097
rect 4270 1043 4300 1097
rect 4370 1043 4400 1097
rect 4470 1043 4500 1220
rect 4570 1183 4600 1220
rect 4670 1290 4700 1467
rect 4770 1413 4800 1467
rect 4770 1290 4800 1327
rect 4670 1280 4800 1290
rect 4670 1246 4718 1280
rect 4752 1246 4800 1280
rect 4670 1236 4800 1246
rect 4570 1043 4600 1097
rect 4670 1043 4700 1236
rect 4770 1183 4800 1236
rect 4870 1274 4900 1607
rect 4970 1553 5000 1747
rect 5070 1693 5100 1747
rect 5170 1693 5200 1747
rect 5070 1553 5100 1607
rect 5170 1553 5200 1607
rect 5270 1553 5300 1747
rect 5370 1693 5400 1747
rect 5470 1693 5500 1747
rect 5570 1693 5600 1747
rect 5370 1553 5400 1607
rect 5470 1553 5500 1607
rect 5570 1553 5600 1607
rect 5670 1553 5700 1747
rect 5770 1693 5800 1747
rect 5870 1693 5900 1747
rect 5770 1553 5800 1607
rect 4970 1413 5000 1467
rect 5070 1413 5100 1467
rect 4970 1274 5000 1327
rect 4870 1264 5000 1274
rect 4870 1230 4918 1264
rect 4952 1230 5000 1264
rect 4870 1220 5000 1230
rect 4870 1183 4900 1220
rect 4970 1183 5000 1220
rect 5070 1290 5100 1327
rect 5170 1290 5200 1467
rect 5270 1413 5300 1467
rect 5370 1413 5400 1467
rect 5470 1413 5500 1467
rect 5570 1413 5600 1467
rect 5670 1413 5700 1467
rect 5770 1413 5800 1467
rect 5870 1413 5900 1607
rect 5970 1553 6000 1747
rect 6070 1693 6100 1747
rect 5970 1413 6000 1467
rect 6070 1413 6100 1607
rect 6170 1553 6200 1747
rect 6270 1693 6300 1747
rect 6370 1693 6400 1887
rect 6470 1833 6500 1887
rect 6570 1833 6600 1887
rect 6670 1833 6700 1887
rect 6770 1833 6800 2027
rect 6870 1973 6900 2167
rect 6970 2113 7000 2430
rect 7070 2500 7100 2537
rect 7170 2500 7200 2537
rect 7070 2490 7200 2500
rect 7070 2456 7118 2490
rect 7152 2456 7200 2490
rect 7070 2446 7200 2456
rect 7070 2393 7100 2446
rect 7170 2393 7200 2446
rect 7270 2484 7300 2537
rect 7370 2484 7400 2537
rect 7270 2474 7400 2484
rect 7270 2440 7318 2474
rect 7352 2440 7400 2474
rect 7270 2430 7400 2440
rect 7070 2253 7100 2307
rect 7170 2253 7200 2307
rect 7270 2253 7300 2430
rect 7370 2393 7400 2430
rect 7470 2500 7500 2537
rect 7570 2500 7600 2537
rect 7470 2490 7600 2500
rect 7470 2456 7518 2490
rect 7552 2456 7600 2490
rect 7470 2446 7600 2456
rect 7470 2393 7500 2446
rect 7570 2393 7600 2446
rect 7670 2484 7700 2537
rect 7770 2484 7800 2537
rect 7670 2474 7800 2484
rect 7670 2440 7718 2474
rect 7752 2440 7800 2474
rect 7670 2430 7800 2440
rect 7670 2393 7700 2430
rect 7770 2393 7800 2430
rect 7870 2500 7900 2537
rect 7970 2500 8000 2537
rect 7870 2490 8000 2500
rect 7870 2456 7918 2490
rect 7952 2456 8000 2490
rect 7870 2446 8000 2456
rect 7870 2393 7900 2446
rect 7970 2393 8000 2446
rect 8070 2484 8100 2537
rect 8170 2484 8200 2537
rect 8070 2474 8200 2484
rect 8070 2440 8118 2474
rect 8152 2440 8200 2474
rect 8070 2430 8200 2440
rect 8070 2393 8100 2430
rect 8170 2393 8200 2430
rect 8270 2500 8300 2817
rect 8370 2763 8400 2817
rect 8470 2763 8500 2817
rect 8570 2763 8600 2817
rect 8670 2763 8700 2817
rect 8370 2623 8400 2677
rect 8370 2500 8400 2537
rect 8270 2490 8400 2500
rect 8270 2456 8318 2490
rect 8352 2456 8400 2490
rect 8270 2446 8400 2456
rect 8270 2393 8300 2446
rect 8370 2393 8400 2446
rect 8470 2484 8500 2677
rect 8570 2623 8600 2677
rect 8670 2623 8700 2677
rect 8570 2484 8600 2537
rect 8470 2474 8600 2484
rect 8470 2440 8518 2474
rect 8552 2440 8600 2474
rect 8470 2430 8600 2440
rect 8470 2393 8500 2430
rect 7370 2253 7400 2307
rect 7470 2253 7500 2307
rect 7070 2113 7100 2167
rect 7170 2113 7200 2167
rect 7270 2113 7300 2167
rect 7370 2113 7400 2167
rect 7470 2113 7500 2167
rect 7570 2113 7600 2307
rect 7670 2253 7700 2307
rect 7670 2113 7700 2167
rect 7770 2113 7800 2307
rect 7870 2253 7900 2307
rect 7970 2253 8000 2307
rect 8070 2253 8100 2307
rect 8170 2253 8200 2307
rect 8270 2253 8300 2307
rect 8370 2253 8400 2307
rect 8470 2253 8500 2307
rect 8570 2253 8600 2430
rect 8670 2500 8700 2537
rect 8770 2500 8800 2957
rect 8870 2903 8900 3237
rect 8970 3183 9000 3237
rect 9070 3183 9100 3237
rect 9170 3183 9200 3237
rect 9270 3183 9300 3237
rect 9370 3183 9400 3237
rect 9470 3183 9500 3237
rect 9570 3183 9600 3377
rect 9670 3323 9700 3377
rect 9770 3323 9800 3517
rect 9870 3463 9900 3517
rect 9970 3463 10000 3517
rect 10070 3463 10100 3640
rect 10170 3603 10200 3640
rect 10270 3710 10300 3747
rect 10370 3710 10400 3747
rect 10270 3700 10400 3710
rect 10270 3666 10318 3700
rect 10352 3666 10400 3700
rect 10270 3656 10400 3666
rect 10270 3603 10300 3656
rect 10370 3603 10400 3656
rect 10470 3694 10500 3747
rect 10570 3694 10600 3747
rect 10470 3684 10600 3694
rect 10470 3650 10518 3684
rect 10552 3650 10600 3684
rect 10470 3640 10600 3650
rect 10470 3603 10500 3640
rect 10570 3603 10600 3640
rect 10670 3710 10700 3747
rect 10770 3710 10800 3747
rect 10670 3700 10800 3710
rect 10670 3666 10718 3700
rect 10752 3666 10800 3700
rect 10670 3656 10800 3666
rect 10170 3463 10200 3517
rect 10270 3463 10300 3517
rect 10370 3463 10400 3517
rect 10470 3463 10500 3517
rect 10570 3463 10600 3517
rect 10670 3463 10700 3656
rect 10770 3603 10800 3656
rect 10870 3694 10900 3747
rect 10970 3694 11000 3747
rect 10870 3684 11000 3694
rect 10870 3650 10918 3684
rect 10952 3650 11000 3684
rect 10870 3640 11000 3650
rect 10870 3603 10900 3640
rect 10970 3603 11000 3640
rect 11070 3710 11100 3747
rect 11170 3710 11200 3887
rect 11270 3833 11300 3887
rect 11370 3833 11400 3887
rect 11470 3833 11500 3887
rect 11070 3700 11200 3710
rect 11070 3666 11118 3700
rect 11152 3666 11200 3700
rect 11070 3656 11200 3666
rect 11070 3603 11100 3656
rect 11170 3603 11200 3656
rect 11270 3694 11300 3747
rect 11370 3694 11400 3747
rect 11270 3684 11400 3694
rect 11270 3650 11318 3684
rect 11352 3650 11400 3684
rect 11270 3640 11400 3650
rect 11270 3603 11300 3640
rect 11370 3603 11400 3640
rect 11470 3710 11500 3747
rect 11570 3710 11600 3887
rect 11670 3833 11700 3887
rect 11770 3833 11800 3887
rect 11870 3833 11900 3887
rect 11970 3833 12000 3887
rect 12070 3833 12100 3887
rect 11470 3700 11600 3710
rect 11470 3666 11518 3700
rect 11552 3666 11600 3700
rect 11470 3656 11600 3666
rect 10770 3463 10800 3517
rect 10870 3463 10900 3517
rect 10970 3463 11000 3517
rect 11070 3463 11100 3517
rect 11170 3463 11200 3517
rect 11270 3463 11300 3517
rect 11370 3463 11400 3517
rect 9870 3323 9900 3377
rect 9970 3323 10000 3377
rect 10070 3323 10100 3377
rect 10170 3323 10200 3377
rect 10270 3323 10300 3377
rect 9670 3183 9700 3237
rect 9770 3183 9800 3237
rect 9870 3183 9900 3237
rect 8970 3043 9000 3097
rect 9070 3043 9100 3097
rect 8970 2903 9000 2957
rect 9070 2903 9100 2957
rect 9170 2903 9200 3097
rect 9270 3043 9300 3097
rect 9370 3043 9400 3097
rect 9270 2903 9300 2957
rect 9370 2903 9400 2957
rect 9470 2903 9500 3097
rect 9570 3043 9600 3097
rect 9670 3043 9700 3097
rect 9770 3043 9800 3097
rect 9870 3043 9900 3097
rect 9970 3043 10000 3237
rect 10070 3183 10100 3237
rect 10070 3043 10100 3097
rect 10170 3043 10200 3237
rect 10270 3183 10300 3237
rect 10270 3043 10300 3097
rect 10370 3043 10400 3377
rect 10470 3323 10500 3377
rect 10470 3183 10500 3237
rect 10570 3183 10600 3377
rect 10670 3323 10700 3377
rect 10770 3323 10800 3377
rect 10870 3323 10900 3377
rect 10970 3323 11000 3377
rect 11070 3323 11100 3377
rect 11170 3323 11200 3377
rect 11270 3323 11300 3377
rect 11370 3323 11400 3377
rect 11470 3323 11500 3656
rect 11570 3603 11600 3656
rect 11670 3694 11700 3747
rect 11770 3694 11800 3747
rect 11670 3684 11800 3694
rect 11670 3650 11718 3684
rect 11752 3650 11800 3684
rect 11670 3640 11800 3650
rect 11670 3603 11700 3640
rect 11770 3603 11800 3640
rect 11870 3710 11900 3747
rect 11970 3710 12000 3747
rect 11870 3700 12000 3710
rect 11870 3666 11918 3700
rect 11952 3666 12000 3700
rect 11870 3656 12000 3666
rect 11870 3603 11900 3656
rect 11970 3603 12000 3656
rect 12070 3694 12100 3747
rect 12170 3694 12200 3887
rect 12270 3833 12300 3887
rect 12370 3833 12400 3887
rect 12470 3833 12500 3887
rect 12570 3833 12600 3887
rect 12670 3833 12700 3887
rect 12770 3833 12800 3887
rect 12970 3833 13000 3887
rect 13070 3833 13100 3887
rect 13280 3833 13310 3887
rect 13380 3833 13410 3887
rect 13480 3833 13510 3887
rect 13580 3833 13610 3887
rect 12070 3684 12200 3694
rect 12070 3650 12118 3684
rect 12152 3650 12200 3684
rect 12070 3640 12200 3650
rect 12070 3603 12100 3640
rect 12170 3603 12200 3640
rect 12270 3710 12300 3747
rect 12370 3710 12400 3747
rect 12270 3700 12400 3710
rect 12270 3666 12318 3700
rect 12352 3666 12400 3700
rect 12270 3656 12400 3666
rect 12270 3603 12300 3656
rect 12370 3603 12400 3656
rect 12470 3694 12500 3747
rect 12570 3694 12600 3747
rect 12470 3684 12600 3694
rect 12470 3650 12518 3684
rect 12552 3650 12600 3684
rect 12470 3640 12600 3650
rect 12470 3603 12500 3640
rect 12570 3603 12600 3640
rect 12670 3710 12700 3747
rect 12770 3710 12800 3747
rect 12970 3714 13000 3747
rect 13070 3714 13100 3747
rect 13280 3714 13310 3747
rect 13380 3714 13410 3747
rect 13480 3714 13510 3747
rect 13580 3714 13610 3747
rect 12670 3700 12800 3710
rect 12670 3666 12718 3700
rect 12752 3666 12800 3700
rect 12670 3656 12800 3666
rect 12670 3603 12700 3656
rect 12770 3603 12800 3656
rect 12958 3698 13012 3714
rect 12958 3664 12968 3698
rect 13002 3664 13012 3698
rect 12958 3648 13012 3664
rect 13058 3698 13112 3714
rect 13058 3664 13068 3698
rect 13102 3664 13112 3698
rect 13058 3648 13112 3664
rect 13268 3698 13322 3714
rect 13268 3664 13278 3698
rect 13312 3664 13322 3698
rect 13268 3648 13322 3664
rect 13368 3698 13422 3714
rect 13368 3664 13378 3698
rect 13412 3664 13422 3698
rect 13368 3648 13422 3664
rect 13468 3698 13522 3714
rect 13468 3664 13478 3698
rect 13512 3664 13522 3698
rect 13468 3648 13522 3664
rect 13568 3698 13622 3714
rect 13568 3664 13578 3698
rect 13612 3664 13622 3698
rect 13568 3648 13622 3664
rect 12970 3603 13000 3648
rect 13070 3603 13100 3648
rect 13280 3603 13310 3648
rect 13380 3603 13410 3648
rect 13480 3603 13510 3648
rect 13580 3603 13610 3648
rect 11570 3463 11600 3517
rect 11670 3463 11700 3517
rect 11770 3463 11800 3517
rect 11870 3463 11900 3517
rect 11970 3463 12000 3517
rect 12070 3463 12100 3517
rect 11570 3323 11600 3377
rect 11670 3323 11700 3377
rect 11770 3323 11800 3377
rect 11870 3323 11900 3377
rect 11970 3323 12000 3377
rect 12070 3323 12100 3377
rect 12170 3323 12200 3517
rect 12270 3463 12300 3517
rect 12370 3463 12400 3517
rect 12470 3463 12500 3517
rect 12570 3463 12600 3517
rect 12670 3463 12700 3517
rect 12770 3463 12800 3517
rect 12970 3463 13000 3517
rect 13070 3463 13100 3517
rect 13280 3463 13310 3517
rect 13380 3463 13410 3517
rect 13480 3463 13510 3517
rect 13580 3463 13610 3517
rect 12270 3323 12300 3377
rect 12370 3323 12400 3377
rect 10670 3183 10700 3237
rect 10770 3183 10800 3237
rect 10470 3043 10500 3097
rect 10570 3043 10600 3097
rect 10670 3043 10700 3097
rect 10770 3043 10800 3097
rect 10870 3043 10900 3237
rect 10970 3183 11000 3237
rect 11070 3183 11100 3237
rect 11170 3183 11200 3237
rect 11270 3183 11300 3237
rect 11370 3183 11400 3237
rect 11470 3183 11500 3237
rect 10970 3043 11000 3097
rect 11070 3043 11100 3097
rect 11170 3043 11200 3097
rect 11270 3043 11300 3097
rect 11370 3043 11400 3097
rect 11470 3043 11500 3097
rect 9570 2903 9600 2957
rect 9670 2903 9700 2957
rect 9770 2903 9800 2957
rect 9870 2903 9900 2957
rect 9970 2903 10000 2957
rect 10070 2903 10100 2957
rect 10170 2903 10200 2957
rect 10270 2903 10300 2957
rect 10370 2903 10400 2957
rect 10470 2903 10500 2957
rect 8870 2763 8900 2817
rect 8870 2623 8900 2677
rect 8970 2623 9000 2817
rect 9070 2763 9100 2817
rect 8670 2490 8800 2500
rect 8670 2456 8718 2490
rect 8752 2456 8800 2490
rect 8670 2446 8800 2456
rect 8670 2393 8700 2446
rect 8770 2393 8800 2446
rect 8870 2484 8900 2537
rect 8970 2484 9000 2537
rect 8870 2474 9000 2484
rect 8870 2440 8918 2474
rect 8952 2440 9000 2474
rect 8870 2430 9000 2440
rect 8870 2393 8900 2430
rect 8970 2393 9000 2430
rect 9070 2500 9100 2677
rect 9170 2623 9200 2817
rect 9270 2763 9300 2817
rect 9170 2500 9200 2537
rect 9070 2490 9200 2500
rect 9070 2456 9118 2490
rect 9152 2456 9200 2490
rect 9070 2446 9200 2456
rect 9070 2393 9100 2446
rect 9170 2393 9200 2446
rect 9270 2484 9300 2677
rect 9370 2623 9400 2817
rect 9470 2763 9500 2817
rect 9470 2623 9500 2677
rect 9370 2484 9400 2537
rect 9270 2474 9400 2484
rect 9270 2440 9318 2474
rect 9352 2440 9400 2474
rect 9270 2430 9400 2440
rect 9270 2393 9300 2430
rect 9370 2393 9400 2430
rect 9470 2500 9500 2537
rect 9570 2500 9600 2817
rect 9670 2763 9700 2817
rect 9770 2763 9800 2817
rect 9870 2763 9900 2817
rect 9670 2623 9700 2677
rect 9770 2623 9800 2677
rect 9870 2623 9900 2677
rect 9470 2490 9600 2500
rect 9470 2456 9518 2490
rect 9552 2456 9600 2490
rect 9470 2446 9600 2456
rect 9470 2393 9500 2446
rect 9570 2393 9600 2446
rect 9670 2484 9700 2537
rect 9770 2484 9800 2537
rect 9670 2474 9800 2484
rect 9670 2440 9718 2474
rect 9752 2440 9800 2474
rect 9670 2430 9800 2440
rect 8670 2253 8700 2307
rect 8770 2253 8800 2307
rect 7870 2113 7900 2167
rect 7970 2113 8000 2167
rect 8070 2113 8100 2167
rect 6870 1833 6900 1887
rect 6970 1833 7000 2027
rect 7070 1973 7100 2027
rect 7170 1973 7200 2027
rect 7270 1973 7300 2027
rect 7370 1973 7400 2027
rect 7470 1973 7500 2027
rect 7570 1973 7600 2027
rect 7670 1973 7700 2027
rect 7770 1973 7800 2027
rect 7870 1973 7900 2027
rect 7970 1973 8000 2027
rect 8070 1973 8100 2027
rect 8170 1973 8200 2167
rect 8270 2113 8300 2167
rect 8270 1973 8300 2027
rect 8370 1973 8400 2167
rect 8470 2113 8500 2167
rect 8570 2113 8600 2167
rect 8670 2113 8700 2167
rect 8470 1973 8500 2027
rect 8570 1973 8600 2027
rect 8670 1973 8700 2027
rect 8770 1973 8800 2167
rect 8870 2113 8900 2307
rect 8970 2253 9000 2307
rect 8870 1973 8900 2027
rect 8970 1973 9000 2167
rect 9070 2113 9100 2307
rect 9170 2253 9200 2307
rect 9170 2113 9200 2167
rect 9070 1973 9100 2027
rect 9170 1973 9200 2027
rect 9270 1973 9300 2307
rect 9370 2253 9400 2307
rect 9470 2253 9500 2307
rect 9370 2113 9400 2167
rect 9470 2113 9500 2167
rect 9570 2113 9600 2307
rect 9670 2253 9700 2430
rect 9770 2393 9800 2430
rect 9870 2500 9900 2537
rect 9970 2500 10000 2817
rect 10070 2763 10100 2817
rect 10170 2763 10200 2817
rect 10270 2763 10300 2817
rect 10370 2763 10400 2817
rect 10070 2623 10100 2677
rect 10170 2623 10200 2677
rect 10270 2623 10300 2677
rect 10370 2623 10400 2677
rect 10470 2623 10500 2817
rect 10570 2763 10600 2957
rect 10670 2903 10700 2957
rect 10770 2903 10800 2957
rect 10870 2903 10900 2957
rect 10970 2903 11000 2957
rect 11070 2903 11100 2957
rect 11170 2903 11200 2957
rect 11270 2903 11300 2957
rect 10570 2623 10600 2677
rect 10670 2623 10700 2817
rect 10770 2763 10800 2817
rect 10870 2763 10900 2817
rect 10970 2763 11000 2817
rect 11070 2763 11100 2817
rect 11170 2763 11200 2817
rect 11270 2763 11300 2817
rect 11370 2763 11400 2957
rect 11470 2903 11500 2957
rect 11570 2903 11600 3237
rect 11670 3183 11700 3237
rect 11770 3183 11800 3237
rect 11870 3183 11900 3237
rect 11970 3183 12000 3237
rect 12070 3183 12100 3237
rect 12170 3183 12200 3237
rect 12270 3183 12300 3237
rect 12370 3183 12400 3237
rect 12470 3183 12500 3377
rect 12570 3323 12600 3377
rect 12670 3323 12700 3377
rect 12770 3323 12800 3377
rect 12970 3323 13000 3377
rect 13070 3323 13100 3377
rect 13280 3323 13310 3377
rect 13380 3323 13410 3377
rect 13480 3323 13510 3377
rect 13580 3323 13610 3377
rect 12570 3183 12600 3237
rect 12670 3183 12700 3237
rect 12770 3183 12800 3237
rect 12970 3183 13000 3237
rect 13070 3183 13100 3237
rect 13280 3183 13310 3237
rect 13380 3183 13410 3237
rect 13480 3183 13510 3237
rect 13580 3183 13610 3237
rect 11670 3043 11700 3097
rect 11770 3043 11800 3097
rect 11870 3043 11900 3097
rect 11970 3043 12000 3097
rect 12070 3043 12100 3097
rect 12170 3043 12200 3097
rect 12270 3043 12300 3097
rect 12370 3043 12400 3097
rect 12470 3043 12500 3097
rect 12570 3043 12600 3097
rect 12670 3043 12700 3097
rect 12770 3043 12800 3097
rect 12970 3043 13000 3097
rect 13070 3043 13100 3097
rect 13280 3043 13310 3097
rect 13380 3043 13410 3097
rect 13480 3043 13510 3097
rect 13580 3043 13610 3097
rect 11670 2903 11700 2957
rect 11770 2903 11800 2957
rect 11470 2763 11500 2817
rect 11570 2763 11600 2817
rect 10770 2623 10800 2677
rect 10870 2623 10900 2677
rect 9870 2490 10000 2500
rect 9870 2456 9918 2490
rect 9952 2456 10000 2490
rect 9870 2446 10000 2456
rect 9870 2393 9900 2446
rect 9970 2393 10000 2446
rect 10070 2484 10100 2537
rect 10170 2484 10200 2537
rect 10070 2474 10200 2484
rect 10070 2440 10118 2474
rect 10152 2440 10200 2474
rect 10070 2430 10200 2440
rect 10070 2393 10100 2430
rect 10170 2393 10200 2430
rect 10270 2500 10300 2537
rect 10370 2500 10400 2537
rect 10270 2490 10400 2500
rect 10270 2456 10318 2490
rect 10352 2456 10400 2490
rect 10270 2446 10400 2456
rect 10270 2393 10300 2446
rect 10370 2393 10400 2446
rect 10470 2484 10500 2537
rect 10570 2484 10600 2537
rect 10470 2474 10600 2484
rect 10470 2440 10518 2474
rect 10552 2440 10600 2474
rect 10470 2430 10600 2440
rect 10470 2393 10500 2430
rect 10570 2393 10600 2430
rect 10670 2500 10700 2537
rect 10770 2500 10800 2537
rect 10670 2490 10800 2500
rect 10670 2456 10718 2490
rect 10752 2456 10800 2490
rect 10670 2446 10800 2456
rect 10670 2393 10700 2446
rect 10770 2393 10800 2446
rect 10870 2484 10900 2537
rect 10970 2484 11000 2677
rect 11070 2623 11100 2677
rect 10870 2474 11000 2484
rect 10870 2440 10918 2474
rect 10952 2440 11000 2474
rect 10870 2430 11000 2440
rect 10870 2393 10900 2430
rect 10970 2393 11000 2430
rect 11070 2500 11100 2537
rect 11170 2500 11200 2677
rect 11270 2623 11300 2677
rect 11070 2490 11200 2500
rect 11070 2456 11118 2490
rect 11152 2456 11200 2490
rect 11070 2446 11200 2456
rect 11070 2393 11100 2446
rect 11170 2393 11200 2446
rect 11270 2484 11300 2537
rect 11370 2484 11400 2677
rect 11470 2623 11500 2677
rect 11570 2623 11600 2677
rect 11270 2474 11400 2484
rect 11270 2440 11318 2474
rect 11352 2440 11400 2474
rect 11270 2430 11400 2440
rect 11270 2393 11300 2430
rect 11370 2393 11400 2430
rect 11470 2500 11500 2537
rect 11570 2500 11600 2537
rect 11470 2490 11600 2500
rect 11470 2456 11518 2490
rect 11552 2456 11600 2490
rect 11470 2446 11600 2456
rect 11470 2393 11500 2446
rect 11570 2393 11600 2446
rect 11670 2484 11700 2817
rect 11770 2763 11800 2817
rect 11870 2763 11900 2957
rect 11970 2903 12000 2957
rect 12070 2903 12100 2957
rect 12170 2903 12200 2957
rect 12270 2903 12300 2957
rect 12370 2903 12400 2957
rect 12470 2903 12500 2957
rect 12570 2903 12600 2957
rect 12670 2903 12700 2957
rect 12770 2903 12800 2957
rect 12970 2903 13000 2957
rect 13070 2903 13100 2957
rect 13280 2903 13310 2957
rect 13380 2903 13410 2957
rect 13480 2903 13510 2957
rect 13580 2903 13610 2957
rect 11970 2763 12000 2817
rect 12070 2763 12100 2817
rect 12170 2763 12200 2817
rect 12270 2763 12300 2817
rect 12370 2763 12400 2817
rect 12470 2763 12500 2817
rect 12570 2763 12600 2817
rect 12670 2763 12700 2817
rect 12770 2763 12800 2817
rect 12970 2763 13000 2817
rect 13070 2763 13100 2817
rect 13280 2763 13310 2817
rect 13380 2763 13410 2817
rect 13480 2763 13510 2817
rect 13580 2763 13610 2817
rect 11770 2623 11800 2677
rect 11870 2623 11900 2677
rect 11970 2623 12000 2677
rect 12070 2623 12100 2677
rect 12170 2623 12200 2677
rect 12270 2623 12300 2677
rect 12370 2623 12400 2677
rect 12470 2623 12500 2677
rect 12570 2623 12600 2677
rect 12670 2623 12700 2677
rect 12770 2623 12800 2677
rect 12970 2623 13000 2677
rect 13070 2623 13100 2677
rect 13280 2623 13310 2677
rect 13380 2623 13410 2677
rect 13480 2623 13510 2677
rect 13580 2623 13610 2677
rect 11770 2484 11800 2537
rect 11670 2474 11800 2484
rect 11670 2440 11718 2474
rect 11752 2440 11800 2474
rect 11670 2430 11800 2440
rect 11670 2393 11700 2430
rect 9770 2253 9800 2307
rect 9870 2253 9900 2307
rect 9970 2253 10000 2307
rect 10070 2253 10100 2307
rect 10170 2253 10200 2307
rect 10270 2253 10300 2307
rect 10370 2253 10400 2307
rect 10470 2253 10500 2307
rect 9670 2113 9700 2167
rect 9770 2113 9800 2167
rect 9870 2113 9900 2167
rect 9970 2113 10000 2167
rect 10070 2113 10100 2167
rect 10170 2113 10200 2167
rect 10270 2113 10300 2167
rect 10370 2113 10400 2167
rect 10470 2113 10500 2167
rect 10570 2113 10600 2307
rect 10670 2253 10700 2307
rect 10770 2253 10800 2307
rect 10870 2253 10900 2307
rect 10970 2253 11000 2307
rect 11070 2253 11100 2307
rect 11170 2253 11200 2307
rect 11270 2253 11300 2307
rect 11370 2253 11400 2307
rect 11470 2253 11500 2307
rect 11570 2253 11600 2307
rect 11670 2253 11700 2307
rect 11770 2253 11800 2430
rect 11870 2500 11900 2537
rect 11970 2500 12000 2537
rect 11870 2490 12000 2500
rect 11870 2456 11918 2490
rect 11952 2456 12000 2490
rect 11870 2446 12000 2456
rect 11870 2393 11900 2446
rect 11870 2253 11900 2307
rect 11970 2253 12000 2446
rect 12070 2484 12100 2537
rect 12170 2484 12200 2537
rect 12070 2474 12200 2484
rect 12070 2440 12118 2474
rect 12152 2440 12200 2474
rect 12070 2430 12200 2440
rect 12070 2393 12100 2430
rect 12170 2393 12200 2430
rect 12270 2500 12300 2537
rect 12370 2500 12400 2537
rect 12270 2490 12400 2500
rect 12270 2456 12318 2490
rect 12352 2456 12400 2490
rect 12270 2446 12400 2456
rect 12270 2393 12300 2446
rect 12370 2393 12400 2446
rect 12470 2484 12500 2537
rect 12570 2484 12600 2537
rect 12470 2474 12600 2484
rect 12470 2440 12518 2474
rect 12552 2440 12600 2474
rect 12470 2430 12600 2440
rect 12470 2393 12500 2430
rect 10670 2113 10700 2167
rect 10770 2113 10800 2167
rect 10870 2113 10900 2167
rect 10970 2113 11000 2167
rect 11070 2113 11100 2167
rect 11170 2113 11200 2167
rect 9370 1973 9400 2027
rect 9470 1973 9500 2027
rect 9570 1973 9600 2027
rect 9670 1973 9700 2027
rect 9770 1973 9800 2027
rect 9870 1973 9900 2027
rect 9970 1973 10000 2027
rect 10070 1973 10100 2027
rect 10170 1973 10200 2027
rect 10270 1973 10300 2027
rect 10370 1973 10400 2027
rect 10470 1973 10500 2027
rect 10570 1973 10600 2027
rect 10670 1973 10700 2027
rect 10770 1973 10800 2027
rect 10870 1973 10900 2027
rect 10970 1973 11000 2027
rect 7070 1833 7100 1887
rect 6470 1693 6500 1747
rect 6270 1553 6300 1607
rect 6170 1413 6200 1467
rect 5070 1280 5200 1290
rect 5070 1246 5118 1280
rect 5152 1246 5200 1280
rect 5070 1236 5200 1246
rect 5070 1183 5100 1236
rect 5170 1183 5200 1236
rect 5270 1274 5300 1327
rect 5370 1274 5400 1327
rect 5270 1264 5400 1274
rect 5270 1230 5318 1264
rect 5352 1230 5400 1264
rect 5270 1220 5400 1230
rect 5270 1183 5300 1220
rect 5370 1183 5400 1220
rect 5470 1290 5500 1327
rect 5570 1290 5600 1327
rect 5470 1280 5600 1290
rect 5470 1246 5518 1280
rect 5552 1246 5600 1280
rect 5470 1236 5600 1246
rect 4770 1043 4800 1097
rect 3970 903 4000 957
rect 4070 903 4100 957
rect 4170 903 4200 957
rect 4270 903 4300 957
rect 4370 903 4400 957
rect 4470 903 4500 957
rect 4570 903 4600 957
rect 4670 903 4700 957
rect 4770 903 4800 957
rect 4870 903 4900 1097
rect 4970 1043 5000 1097
rect 5070 1043 5100 1097
rect 5170 1043 5200 1097
rect 5270 1043 5300 1097
rect 4970 903 5000 957
rect 5070 903 5100 957
rect 5170 903 5200 957
rect 5270 903 5300 957
rect 5370 903 5400 1097
rect 5470 1043 5500 1236
rect 5570 1183 5600 1236
rect 5670 1274 5700 1327
rect 5770 1274 5800 1327
rect 5670 1264 5800 1274
rect 5670 1230 5718 1264
rect 5752 1230 5800 1264
rect 5670 1220 5800 1230
rect 5670 1183 5700 1220
rect 5770 1183 5800 1220
rect 5870 1290 5900 1327
rect 5970 1290 6000 1327
rect 5870 1280 6000 1290
rect 5870 1246 5918 1280
rect 5952 1246 6000 1280
rect 5870 1236 6000 1246
rect 5870 1183 5900 1236
rect 5970 1183 6000 1236
rect 6070 1274 6100 1327
rect 6170 1274 6200 1327
rect 6070 1264 6200 1274
rect 6070 1230 6118 1264
rect 6152 1230 6200 1264
rect 6070 1220 6200 1230
rect 6070 1183 6100 1220
rect 6170 1183 6200 1220
rect 6270 1290 6300 1467
rect 6370 1413 6400 1607
rect 6470 1553 6500 1607
rect 6570 1553 6600 1747
rect 6670 1693 6700 1747
rect 6770 1693 6800 1747
rect 6870 1693 6900 1747
rect 6970 1693 7000 1747
rect 7070 1693 7100 1747
rect 7170 1693 7200 1887
rect 7270 1833 7300 1887
rect 7370 1833 7400 1887
rect 7270 1693 7300 1747
rect 7370 1693 7400 1747
rect 7470 1693 7500 1887
rect 7570 1833 7600 1887
rect 7670 1833 7700 1887
rect 7570 1693 7600 1747
rect 7670 1693 7700 1747
rect 7770 1693 7800 1887
rect 7870 1833 7900 1887
rect 7970 1833 8000 1887
rect 7870 1693 7900 1747
rect 7970 1693 8000 1747
rect 8070 1693 8100 1887
rect 8170 1833 8200 1887
rect 8270 1833 8300 1887
rect 8370 1833 8400 1887
rect 8470 1833 8500 1887
rect 8570 1833 8600 1887
rect 8170 1693 8200 1747
rect 8270 1693 8300 1747
rect 8370 1693 8400 1747
rect 8470 1693 8500 1747
rect 8570 1693 8600 1747
rect 8670 1693 8700 1887
rect 8770 1833 8800 1887
rect 8870 1833 8900 1887
rect 8970 1833 9000 1887
rect 9070 1833 9100 1887
rect 9170 1833 9200 1887
rect 9270 1833 9300 1887
rect 9370 1833 9400 1887
rect 9470 1833 9500 1887
rect 9570 1833 9600 1887
rect 9670 1833 9700 1887
rect 9770 1833 9800 1887
rect 8770 1693 8800 1747
rect 8870 1693 8900 1747
rect 8970 1693 9000 1747
rect 9070 1693 9100 1747
rect 9170 1693 9200 1747
rect 9270 1693 9300 1747
rect 9370 1693 9400 1747
rect 9470 1693 9500 1747
rect 6670 1553 6700 1607
rect 6770 1553 6800 1607
rect 6870 1553 6900 1607
rect 6970 1553 7000 1607
rect 7070 1553 7100 1607
rect 7170 1553 7200 1607
rect 7270 1553 7300 1607
rect 7370 1553 7400 1607
rect 7470 1553 7500 1607
rect 7570 1553 7600 1607
rect 7670 1553 7700 1607
rect 6370 1290 6400 1327
rect 6270 1280 6400 1290
rect 6270 1246 6318 1280
rect 6352 1246 6400 1280
rect 6270 1236 6400 1246
rect 6270 1183 6300 1236
rect 6370 1183 6400 1236
rect 6470 1274 6500 1467
rect 6570 1413 6600 1467
rect 6670 1413 6700 1467
rect 6570 1274 6600 1327
rect 6470 1264 6600 1274
rect 6470 1230 6518 1264
rect 6552 1230 6600 1264
rect 6470 1220 6600 1230
rect 6470 1183 6500 1220
rect 6570 1183 6600 1220
rect 6670 1290 6700 1327
rect 6770 1290 6800 1467
rect 6870 1413 6900 1467
rect 6670 1280 6800 1290
rect 6670 1246 6718 1280
rect 6752 1246 6800 1280
rect 6670 1236 6800 1246
rect 6670 1183 6700 1236
rect 5570 1043 5600 1097
rect 5670 1043 5700 1097
rect 5770 1043 5800 1097
rect 5870 1043 5900 1097
rect 5970 1043 6000 1097
rect 6070 1043 6100 1097
rect 6170 1043 6200 1097
rect 6270 1043 6300 1097
rect 6370 1043 6400 1097
rect 5470 903 5500 957
rect 5570 903 5600 957
rect 5670 903 5700 957
rect 5770 903 5800 957
rect 5870 903 5900 957
rect 5970 903 6000 957
rect 6070 903 6100 957
rect 6170 903 6200 957
rect 6270 903 6300 957
rect 6370 903 6400 957
rect 6470 903 6500 1097
rect 6570 1043 6600 1097
rect 6670 1043 6700 1097
rect 6770 1043 6800 1236
rect 6870 1274 6900 1327
rect 6970 1274 7000 1467
rect 7070 1413 7100 1467
rect 7170 1413 7200 1467
rect 7270 1413 7300 1467
rect 7370 1413 7400 1467
rect 7470 1413 7500 1467
rect 7570 1413 7600 1467
rect 7670 1413 7700 1467
rect 7770 1413 7800 1607
rect 7870 1553 7900 1607
rect 7870 1413 7900 1467
rect 6870 1264 7000 1274
rect 6870 1230 6918 1264
rect 6952 1230 7000 1264
rect 6870 1220 7000 1230
rect 6870 1183 6900 1220
rect 6970 1183 7000 1220
rect 7070 1290 7100 1327
rect 7170 1290 7200 1327
rect 7070 1280 7200 1290
rect 7070 1246 7118 1280
rect 7152 1246 7200 1280
rect 7070 1236 7200 1246
rect 7070 1183 7100 1236
rect 7170 1183 7200 1236
rect 7270 1274 7300 1327
rect 7370 1274 7400 1327
rect 7270 1264 7400 1274
rect 7270 1230 7318 1264
rect 7352 1230 7400 1264
rect 7270 1220 7400 1230
rect 7270 1183 7300 1220
rect 7370 1183 7400 1220
rect 7470 1290 7500 1327
rect 7570 1290 7600 1327
rect 7470 1280 7600 1290
rect 7470 1246 7518 1280
rect 7552 1246 7600 1280
rect 7470 1236 7600 1246
rect 7470 1183 7500 1236
rect 7570 1183 7600 1236
rect 7670 1274 7700 1327
rect 7770 1274 7800 1327
rect 7670 1264 7800 1274
rect 7670 1230 7718 1264
rect 7752 1230 7800 1264
rect 7670 1220 7800 1230
rect 7670 1183 7700 1220
rect 7770 1183 7800 1220
rect 7870 1290 7900 1327
rect 7970 1290 8000 1607
rect 8070 1553 8100 1607
rect 8170 1553 8200 1607
rect 8270 1553 8300 1607
rect 8370 1553 8400 1607
rect 8470 1553 8500 1607
rect 8070 1413 8100 1467
rect 8170 1413 8200 1467
rect 8270 1413 8300 1467
rect 8370 1413 8400 1467
rect 8470 1413 8500 1467
rect 8570 1413 8600 1607
rect 8670 1553 8700 1607
rect 8770 1553 8800 1607
rect 8870 1553 8900 1607
rect 8970 1553 9000 1607
rect 9070 1553 9100 1607
rect 9170 1553 9200 1607
rect 9270 1553 9300 1607
rect 8670 1413 8700 1467
rect 8770 1413 8800 1467
rect 8870 1413 8900 1467
rect 8970 1413 9000 1467
rect 9070 1413 9100 1467
rect 9170 1413 9200 1467
rect 9270 1413 9300 1467
rect 7870 1280 8000 1290
rect 7870 1246 7918 1280
rect 7952 1246 8000 1280
rect 7870 1236 8000 1246
rect 7870 1183 7900 1236
rect 7970 1183 8000 1236
rect 8070 1274 8100 1327
rect 8170 1274 8200 1327
rect 8070 1264 8200 1274
rect 8070 1230 8118 1264
rect 8152 1230 8200 1264
rect 8070 1220 8200 1230
rect 8070 1183 8100 1220
rect 8170 1183 8200 1220
rect 8270 1290 8300 1327
rect 8370 1290 8400 1327
rect 8270 1280 8400 1290
rect 8270 1246 8318 1280
rect 8352 1246 8400 1280
rect 8270 1236 8400 1246
rect 8270 1183 8300 1236
rect 8370 1183 8400 1236
rect 8470 1274 8500 1327
rect 8570 1274 8600 1327
rect 8470 1264 8600 1274
rect 8470 1230 8518 1264
rect 8552 1230 8600 1264
rect 8470 1220 8600 1230
rect 8470 1183 8500 1220
rect 8570 1183 8600 1220
rect 8670 1290 8700 1327
rect 8770 1290 8800 1327
rect 8670 1280 8800 1290
rect 8670 1246 8718 1280
rect 8752 1246 8800 1280
rect 8670 1236 8800 1246
rect 8670 1183 8700 1236
rect 8770 1183 8800 1236
rect 8870 1274 8900 1327
rect 8970 1274 9000 1327
rect 8870 1264 9000 1274
rect 8870 1230 8918 1264
rect 8952 1230 9000 1264
rect 8870 1220 9000 1230
rect 8870 1183 8900 1220
rect 8970 1183 9000 1220
rect 9070 1290 9100 1327
rect 9170 1290 9200 1327
rect 9070 1280 9200 1290
rect 9070 1246 9118 1280
rect 9152 1246 9200 1280
rect 9070 1236 9200 1246
rect 9070 1183 9100 1236
rect 9170 1183 9200 1236
rect 9270 1274 9300 1327
rect 9370 1274 9400 1607
rect 9470 1553 9500 1607
rect 9570 1553 9600 1747
rect 9670 1693 9700 1747
rect 9770 1693 9800 1747
rect 9870 1693 9900 1887
rect 9970 1833 10000 1887
rect 9970 1693 10000 1747
rect 10070 1693 10100 1887
rect 10170 1833 10200 1887
rect 10170 1693 10200 1747
rect 10270 1693 10300 1887
rect 10370 1833 10400 1887
rect 10370 1693 10400 1747
rect 10470 1693 10500 1887
rect 10570 1833 10600 1887
rect 10670 1833 10700 1887
rect 10570 1693 10600 1747
rect 10670 1693 10700 1747
rect 10770 1693 10800 1887
rect 10870 1833 10900 1887
rect 10970 1833 11000 1887
rect 11070 1833 11100 2027
rect 11170 1973 11200 2027
rect 11170 1833 11200 1887
rect 11270 1833 11300 2167
rect 11370 2113 11400 2167
rect 11370 1973 11400 2027
rect 11470 1973 11500 2167
rect 11570 2113 11600 2167
rect 11670 2113 11700 2167
rect 11770 2113 11800 2167
rect 11870 2113 11900 2167
rect 11970 2113 12000 2167
rect 12070 2113 12100 2307
rect 12170 2253 12200 2307
rect 12270 2253 12300 2307
rect 12170 2113 12200 2167
rect 12270 2113 12300 2167
rect 12370 2113 12400 2307
rect 12470 2253 12500 2307
rect 12570 2253 12600 2430
rect 12670 2500 12700 2537
rect 12770 2500 12800 2537
rect 12970 2504 13000 2537
rect 13070 2504 13100 2537
rect 13280 2504 13310 2537
rect 13380 2504 13410 2537
rect 13480 2504 13510 2537
rect 13580 2504 13610 2537
rect 12670 2490 12800 2500
rect 12670 2456 12718 2490
rect 12752 2456 12800 2490
rect 12670 2446 12800 2456
rect 12670 2393 12700 2446
rect 12770 2393 12800 2446
rect 12958 2488 13012 2504
rect 12958 2454 12968 2488
rect 13002 2454 13012 2488
rect 12958 2438 13012 2454
rect 13058 2488 13112 2504
rect 13058 2454 13068 2488
rect 13102 2454 13112 2488
rect 13058 2438 13112 2454
rect 13268 2488 13322 2504
rect 13268 2454 13278 2488
rect 13312 2454 13322 2488
rect 13268 2438 13322 2454
rect 13368 2488 13422 2504
rect 13368 2454 13378 2488
rect 13412 2454 13422 2488
rect 13368 2438 13422 2454
rect 13468 2488 13522 2504
rect 13468 2454 13478 2488
rect 13512 2454 13522 2488
rect 13468 2438 13522 2454
rect 13568 2488 13622 2504
rect 13568 2454 13578 2488
rect 13612 2454 13622 2488
rect 13568 2438 13622 2454
rect 12970 2393 13000 2438
rect 13070 2393 13100 2438
rect 13280 2393 13310 2438
rect 13380 2393 13410 2438
rect 13480 2393 13510 2438
rect 13580 2393 13610 2438
rect 12470 2113 12500 2167
rect 12570 2113 12600 2167
rect 11570 1973 11600 2027
rect 11670 1973 11700 2027
rect 11770 1973 11800 2027
rect 11870 1973 11900 2027
rect 11970 1973 12000 2027
rect 12070 1973 12100 2027
rect 12170 1973 12200 2027
rect 12270 1973 12300 2027
rect 12370 1973 12400 2027
rect 12470 1973 12500 2027
rect 12570 1973 12600 2027
rect 11370 1833 11400 1887
rect 11470 1833 11500 1887
rect 11570 1833 11600 1887
rect 10870 1693 10900 1747
rect 9670 1553 9700 1607
rect 9770 1553 9800 1607
rect 9870 1553 9900 1607
rect 9970 1553 10000 1607
rect 10070 1553 10100 1607
rect 10170 1553 10200 1607
rect 10270 1553 10300 1607
rect 10370 1553 10400 1607
rect 10470 1553 10500 1607
rect 10570 1553 10600 1607
rect 10670 1553 10700 1607
rect 10770 1553 10800 1607
rect 10870 1553 10900 1607
rect 9470 1413 9500 1467
rect 9570 1413 9600 1467
rect 9670 1413 9700 1467
rect 9770 1413 9800 1467
rect 9870 1413 9900 1467
rect 9970 1413 10000 1467
rect 10070 1413 10100 1467
rect 10170 1413 10200 1467
rect 9270 1264 9400 1274
rect 9270 1230 9318 1264
rect 9352 1230 9400 1264
rect 9270 1220 9400 1230
rect 9270 1183 9300 1220
rect 9370 1183 9400 1220
rect 9470 1290 9500 1327
rect 9570 1290 9600 1327
rect 9470 1280 9600 1290
rect 9470 1246 9518 1280
rect 9552 1246 9600 1280
rect 9470 1236 9600 1246
rect 9470 1183 9500 1236
rect 9570 1183 9600 1236
rect 9670 1274 9700 1327
rect 9770 1274 9800 1327
rect 9670 1264 9800 1274
rect 9670 1230 9718 1264
rect 9752 1230 9800 1264
rect 9670 1220 9800 1230
rect 6870 1043 6900 1097
rect 6570 903 6600 957
rect 3970 763 4000 817
rect 4070 763 4100 817
rect 4170 763 4200 817
rect 4270 763 4300 817
rect 4370 763 4400 817
rect 4470 763 4500 817
rect 4570 763 4600 817
rect 3770 623 3800 677
rect 3870 623 3900 677
rect 2870 483 2900 537
rect 2970 483 3000 537
rect 3070 483 3100 537
rect 3170 483 3200 537
rect 3270 483 3300 537
rect 3370 483 3400 537
rect 3470 483 3500 537
rect 3570 483 3600 537
rect 3670 483 3700 537
rect 3770 483 3800 537
rect 3870 483 3900 537
rect 3970 483 4000 677
rect 4070 623 4100 677
rect 4070 483 4100 537
rect 4170 483 4200 677
rect 4270 623 4300 677
rect 4370 623 4400 677
rect 4470 623 4500 677
rect 4570 623 4600 677
rect 4670 623 4700 817
rect 4770 763 4800 817
rect 4870 763 4900 817
rect 4970 763 5000 817
rect 5070 763 5100 817
rect 4770 623 4800 677
rect 4270 483 4300 537
rect 4370 483 4400 537
rect 2770 343 2800 397
rect 1770 64 1800 117
rect 1670 54 1800 64
rect 1670 20 1718 54
rect 1752 20 1800 54
rect 1670 10 1800 20
rect 1670 0 1700 10
rect 1770 0 1800 10
rect 1870 80 1900 257
rect 1970 203 2000 257
rect 2070 203 2100 257
rect 2170 203 2200 257
rect 2270 203 2300 257
rect 2370 203 2400 257
rect 2470 203 2500 257
rect 2570 203 2600 257
rect 2670 203 2700 257
rect 2770 203 2800 257
rect 2870 203 2900 397
rect 2970 343 3000 397
rect 2970 203 3000 257
rect 3070 203 3100 397
rect 3170 343 3200 397
rect 3270 343 3300 397
rect 3370 343 3400 397
rect 3470 343 3500 397
rect 3570 343 3600 397
rect 3670 343 3700 397
rect 3770 343 3800 397
rect 3870 343 3900 397
rect 3970 343 4000 397
rect 4070 343 4100 397
rect 4170 343 4200 397
rect 4270 343 4300 397
rect 4370 343 4400 397
rect 4470 343 4500 537
rect 4570 483 4600 537
rect 4670 483 4700 537
rect 4770 483 4800 537
rect 4870 483 4900 677
rect 4970 623 5000 677
rect 4970 483 5000 537
rect 5070 483 5100 677
rect 5170 623 5200 817
rect 5270 763 5300 817
rect 5370 763 5400 817
rect 5470 763 5500 817
rect 5570 763 5600 817
rect 5670 763 5700 817
rect 3170 203 3200 257
rect 3270 203 3300 257
rect 3370 203 3400 257
rect 3470 203 3500 257
rect 3570 203 3600 257
rect 3670 203 3700 257
rect 3770 203 3800 257
rect 3870 203 3900 257
rect 3970 203 4000 257
rect 4070 203 4100 257
rect 4170 203 4200 257
rect 4270 203 4300 257
rect 4370 203 4400 257
rect 4470 203 4500 257
rect 4570 203 4600 397
rect 4670 343 4700 397
rect 4770 343 4800 397
rect 4670 203 4700 257
rect 4770 203 4800 257
rect 4870 203 4900 397
rect 4970 343 5000 397
rect 4970 203 5000 257
rect 5070 203 5100 397
rect 5170 343 5200 537
rect 5270 483 5300 677
rect 5370 623 5400 677
rect 5470 623 5500 677
rect 5570 623 5600 677
rect 5670 623 5700 677
rect 5770 623 5800 817
rect 5870 763 5900 817
rect 5970 763 6000 817
rect 6070 763 6100 817
rect 6170 763 6200 817
rect 5870 623 5900 677
rect 5970 623 6000 677
rect 6070 623 6100 677
rect 6170 623 6200 677
rect 6270 623 6300 817
rect 6370 763 6400 817
rect 6370 623 6400 677
rect 6470 623 6500 817
rect 6570 763 6600 817
rect 6670 763 6700 957
rect 6770 903 6800 957
rect 6870 903 6900 957
rect 6970 903 7000 1097
rect 7070 1043 7100 1097
rect 7070 903 7100 957
rect 7170 903 7200 1097
rect 7270 1043 7300 1097
rect 7270 903 7300 957
rect 6770 763 6800 817
rect 6870 763 6900 817
rect 6970 763 7000 817
rect 6570 623 6600 677
rect 6670 623 6700 677
rect 6770 623 6800 677
rect 6870 623 6900 677
rect 6970 623 7000 677
rect 7070 623 7100 817
rect 7170 763 7200 817
rect 7270 763 7300 817
rect 7370 763 7400 1097
rect 7470 1043 7500 1097
rect 7570 1043 7600 1097
rect 7670 1043 7700 1097
rect 7770 1043 7800 1097
rect 7870 1043 7900 1097
rect 7970 1043 8000 1097
rect 8070 1043 8100 1097
rect 8170 1043 8200 1097
rect 8270 1043 8300 1097
rect 8370 1043 8400 1097
rect 8470 1043 8500 1097
rect 8570 1043 8600 1097
rect 7470 903 7500 957
rect 7470 763 7500 817
rect 7570 763 7600 957
rect 7670 903 7700 957
rect 7670 763 7700 817
rect 7770 763 7800 957
rect 7870 903 7900 957
rect 7870 763 7900 817
rect 7970 763 8000 957
rect 8070 903 8100 957
rect 8170 903 8200 957
rect 8270 903 8300 957
rect 8370 903 8400 957
rect 8470 903 8500 957
rect 8570 903 8600 957
rect 8070 763 8100 817
rect 8170 763 8200 817
rect 8270 763 8300 817
rect 8370 763 8400 817
rect 8470 763 8500 817
rect 8570 763 8600 817
rect 8670 763 8700 1097
rect 8770 1043 8800 1097
rect 8770 903 8800 957
rect 8770 763 8800 817
rect 8870 763 8900 1097
rect 8970 1043 9000 1097
rect 9070 1043 9100 1097
rect 9170 1043 9200 1097
rect 9270 1043 9300 1097
rect 9370 1043 9400 1097
rect 9470 1043 9500 1097
rect 8970 903 9000 957
rect 9070 903 9100 957
rect 9170 903 9200 957
rect 9270 903 9300 957
rect 9370 903 9400 957
rect 9470 903 9500 957
rect 9570 903 9600 1097
rect 9670 1043 9700 1220
rect 9770 1183 9800 1220
rect 9870 1290 9900 1327
rect 9970 1290 10000 1327
rect 9870 1280 10000 1290
rect 9870 1246 9918 1280
rect 9952 1246 10000 1280
rect 9870 1236 10000 1246
rect 9870 1183 9900 1236
rect 9970 1183 10000 1236
rect 10070 1274 10100 1327
rect 10170 1274 10200 1327
rect 10070 1264 10200 1274
rect 10070 1230 10118 1264
rect 10152 1230 10200 1264
rect 10070 1220 10200 1230
rect 10070 1183 10100 1220
rect 10170 1183 10200 1220
rect 10270 1290 10300 1467
rect 10370 1413 10400 1467
rect 10470 1413 10500 1467
rect 10570 1413 10600 1467
rect 10670 1413 10700 1467
rect 10770 1413 10800 1467
rect 10870 1413 10900 1467
rect 10970 1413 11000 1747
rect 11070 1693 11100 1747
rect 11170 1693 11200 1747
rect 11270 1693 11300 1747
rect 11370 1693 11400 1747
rect 11470 1693 11500 1747
rect 11570 1693 11600 1747
rect 11670 1693 11700 1887
rect 11770 1833 11800 1887
rect 11870 1833 11900 1887
rect 11070 1553 11100 1607
rect 11070 1413 11100 1467
rect 10370 1290 10400 1327
rect 10270 1280 10400 1290
rect 10270 1246 10318 1280
rect 10352 1246 10400 1280
rect 10270 1236 10400 1246
rect 10270 1183 10300 1236
rect 10370 1183 10400 1236
rect 10470 1274 10500 1327
rect 10570 1274 10600 1327
rect 10470 1264 10600 1274
rect 10470 1230 10518 1264
rect 10552 1230 10600 1264
rect 10470 1220 10600 1230
rect 10470 1183 10500 1220
rect 10570 1183 10600 1220
rect 10670 1290 10700 1327
rect 10770 1290 10800 1327
rect 10670 1280 10800 1290
rect 10670 1246 10718 1280
rect 10752 1246 10800 1280
rect 10670 1236 10800 1246
rect 10670 1183 10700 1236
rect 10770 1183 10800 1236
rect 10870 1274 10900 1327
rect 10970 1274 11000 1327
rect 10870 1264 11000 1274
rect 10870 1230 10918 1264
rect 10952 1230 11000 1264
rect 10870 1220 11000 1230
rect 10870 1183 10900 1220
rect 10970 1183 11000 1220
rect 11070 1290 11100 1327
rect 11170 1290 11200 1607
rect 11270 1553 11300 1607
rect 11370 1553 11400 1607
rect 11470 1553 11500 1607
rect 11570 1553 11600 1607
rect 11670 1553 11700 1607
rect 11770 1553 11800 1747
rect 11870 1693 11900 1747
rect 11970 1693 12000 1887
rect 12070 1833 12100 1887
rect 12170 1833 12200 1887
rect 12270 1833 12300 1887
rect 12370 1833 12400 1887
rect 12470 1833 12500 1887
rect 12570 1833 12600 1887
rect 12670 1833 12700 2307
rect 12770 2253 12800 2307
rect 12970 2253 13000 2307
rect 13070 2253 13100 2307
rect 13280 2253 13310 2307
rect 13380 2253 13410 2307
rect 13480 2253 13510 2307
rect 13580 2253 13610 2307
rect 12770 2113 12800 2167
rect 12970 2113 13000 2167
rect 13070 2113 13100 2167
rect 13280 2113 13310 2167
rect 13380 2113 13410 2167
rect 13480 2113 13510 2167
rect 13580 2113 13610 2167
rect 12770 1973 12800 2027
rect 12970 1973 13000 2027
rect 13070 1973 13100 2027
rect 13280 1973 13310 2027
rect 13380 1973 13410 2027
rect 13480 1973 13510 2027
rect 13580 1973 13610 2027
rect 12770 1833 12800 1887
rect 12970 1833 13000 1887
rect 13070 1833 13100 1887
rect 13280 1833 13310 1887
rect 13380 1833 13410 1887
rect 13480 1833 13510 1887
rect 13580 1833 13610 1887
rect 12070 1693 12100 1747
rect 12170 1693 12200 1747
rect 12270 1693 12300 1747
rect 12370 1693 12400 1747
rect 12470 1693 12500 1747
rect 12570 1693 12600 1747
rect 12670 1693 12700 1747
rect 12770 1693 12800 1747
rect 12970 1693 13000 1747
rect 13070 1693 13100 1747
rect 13280 1693 13310 1747
rect 13380 1693 13410 1747
rect 13480 1693 13510 1747
rect 13580 1693 13610 1747
rect 11870 1553 11900 1607
rect 11970 1553 12000 1607
rect 11270 1413 11300 1467
rect 11370 1413 11400 1467
rect 11470 1413 11500 1467
rect 11570 1413 11600 1467
rect 11670 1413 11700 1467
rect 11070 1280 11200 1290
rect 11070 1246 11118 1280
rect 11152 1246 11200 1280
rect 11070 1236 11200 1246
rect 9770 1043 9800 1097
rect 9870 1043 9900 1097
rect 9670 903 9700 957
rect 9770 903 9800 957
rect 9870 903 9900 957
rect 8970 763 9000 817
rect 9070 763 9100 817
rect 7170 623 7200 677
rect 7270 623 7300 677
rect 7370 623 7400 677
rect 7470 623 7500 677
rect 7570 623 7600 677
rect 7670 623 7700 677
rect 7770 623 7800 677
rect 7870 623 7900 677
rect 7970 623 8000 677
rect 8070 623 8100 677
rect 8170 623 8200 677
rect 8270 623 8300 677
rect 5270 343 5300 397
rect 5370 343 5400 537
rect 5470 483 5500 537
rect 5570 483 5600 537
rect 5670 483 5700 537
rect 5770 483 5800 537
rect 5870 483 5900 537
rect 5970 483 6000 537
rect 6070 483 6100 537
rect 5470 343 5500 397
rect 5570 343 5600 397
rect 5670 343 5700 397
rect 5770 343 5800 397
rect 5170 203 5200 257
rect 5270 203 5300 257
rect 5370 203 5400 257
rect 5470 203 5500 257
rect 5570 203 5600 257
rect 5670 203 5700 257
rect 5770 203 5800 257
rect 5870 203 5900 397
rect 5970 343 6000 397
rect 5970 203 6000 257
rect 6070 203 6100 397
rect 6170 343 6200 537
rect 6270 483 6300 537
rect 6370 483 6400 537
rect 6170 203 6200 257
rect 6270 203 6300 397
rect 6370 343 6400 397
rect 6370 203 6400 257
rect 6470 203 6500 537
rect 6570 483 6600 537
rect 6670 483 6700 537
rect 6770 483 6800 537
rect 6870 483 6900 537
rect 6970 483 7000 537
rect 7070 483 7100 537
rect 6570 343 6600 397
rect 6570 203 6600 257
rect 6670 203 6700 397
rect 6770 343 6800 397
rect 6770 203 6800 257
rect 6870 203 6900 397
rect 6970 343 7000 397
rect 7070 343 7100 397
rect 7170 343 7200 537
rect 7270 483 7300 537
rect 7270 343 7300 397
rect 7370 343 7400 537
rect 7470 483 7500 537
rect 7470 343 7500 397
rect 7570 343 7600 537
rect 7670 483 7700 537
rect 7770 483 7800 537
rect 7870 483 7900 537
rect 7970 483 8000 537
rect 8070 483 8100 537
rect 8170 483 8200 537
rect 8270 483 8300 537
rect 7670 343 7700 397
rect 7770 343 7800 397
rect 6970 203 7000 257
rect 1970 80 2000 117
rect 1870 70 2000 80
rect 1870 36 1918 70
rect 1952 36 2000 70
rect 1870 26 2000 36
rect 1870 0 1900 26
rect 1970 0 2000 26
rect 2070 64 2100 117
rect 2170 64 2200 117
rect 2070 54 2200 64
rect 2070 20 2118 54
rect 2152 20 2200 54
rect 2070 10 2200 20
rect 2070 0 2100 10
rect 2170 0 2200 10
rect 2270 80 2300 117
rect 2370 80 2400 117
rect 2270 70 2400 80
rect 2270 36 2318 70
rect 2352 36 2400 70
rect 2270 26 2400 36
rect 2270 0 2300 26
rect 2370 0 2400 26
rect 2470 64 2500 117
rect 2570 64 2600 117
rect 2470 54 2600 64
rect 2470 20 2518 54
rect 2552 20 2600 54
rect 2470 10 2600 20
rect 2470 0 2500 10
rect 2570 0 2600 10
rect 2670 80 2700 117
rect 2770 80 2800 117
rect 2670 70 2800 80
rect 2670 36 2718 70
rect 2752 36 2800 70
rect 2670 26 2800 36
rect 2670 0 2700 26
rect 2770 0 2800 26
rect 2870 64 2900 117
rect 2970 64 3000 117
rect 2870 54 3000 64
rect 2870 20 2918 54
rect 2952 20 3000 54
rect 2870 10 3000 20
rect 2870 0 2900 10
rect 2970 0 3000 10
rect 3070 80 3100 117
rect 3170 80 3200 117
rect 3070 70 3200 80
rect 3070 36 3118 70
rect 3152 36 3200 70
rect 3070 26 3200 36
rect 3070 0 3100 26
rect 3170 0 3200 26
rect 3270 64 3300 117
rect 3370 64 3400 117
rect 3270 54 3400 64
rect 3270 20 3318 54
rect 3352 20 3400 54
rect 3270 10 3400 20
rect 3270 0 3300 10
rect 3370 0 3400 10
rect 3470 80 3500 117
rect 3570 80 3600 117
rect 3470 70 3600 80
rect 3470 36 3518 70
rect 3552 36 3600 70
rect 3470 26 3600 36
rect 3470 0 3500 26
rect 3570 0 3600 26
rect 3670 64 3700 117
rect 3770 64 3800 117
rect 3670 54 3800 64
rect 3670 20 3718 54
rect 3752 20 3800 54
rect 3670 10 3800 20
rect 3670 0 3700 10
rect 3770 0 3800 10
rect 3870 80 3900 117
rect 3970 80 4000 117
rect 3870 70 4000 80
rect 3870 36 3918 70
rect 3952 36 4000 70
rect 3870 26 4000 36
rect 3870 0 3900 26
rect 3970 0 4000 26
rect 4070 64 4100 117
rect 4170 64 4200 117
rect 4070 54 4200 64
rect 4070 20 4118 54
rect 4152 20 4200 54
rect 4070 10 4200 20
rect 4070 0 4100 10
rect 4170 0 4200 10
rect 4270 80 4300 117
rect 4370 80 4400 117
rect 4270 70 4400 80
rect 4270 36 4318 70
rect 4352 36 4400 70
rect 4270 26 4400 36
rect 4270 0 4300 26
rect 4370 0 4400 26
rect 4470 64 4500 117
rect 4570 64 4600 117
rect 4470 54 4600 64
rect 4470 20 4518 54
rect 4552 20 4600 54
rect 4470 10 4600 20
rect 4470 0 4500 10
rect 4570 0 4600 10
rect 4670 80 4700 117
rect 4770 80 4800 117
rect 4670 70 4800 80
rect 4670 36 4718 70
rect 4752 36 4800 70
rect 4670 26 4800 36
rect 4670 0 4700 26
rect 4770 0 4800 26
rect 4870 64 4900 117
rect 4970 64 5000 117
rect 4870 54 5000 64
rect 4870 20 4918 54
rect 4952 20 5000 54
rect 4870 10 5000 20
rect 4870 0 4900 10
rect 4970 0 5000 10
rect 5070 80 5100 117
rect 5170 80 5200 117
rect 5070 70 5200 80
rect 5070 36 5118 70
rect 5152 36 5200 70
rect 5070 26 5200 36
rect 5070 0 5100 26
rect 5170 0 5200 26
rect 5270 64 5300 117
rect 5370 64 5400 117
rect 5270 54 5400 64
rect 5270 20 5318 54
rect 5352 20 5400 54
rect 5270 10 5400 20
rect 5270 0 5300 10
rect 5370 0 5400 10
rect 5470 80 5500 117
rect 5570 80 5600 117
rect 5470 70 5600 80
rect 5470 36 5518 70
rect 5552 36 5600 70
rect 5470 26 5600 36
rect 5470 0 5500 26
rect 5570 0 5600 26
rect 5670 64 5700 117
rect 5770 64 5800 117
rect 5670 54 5800 64
rect 5670 20 5718 54
rect 5752 20 5800 54
rect 5670 10 5800 20
rect 5670 0 5700 10
rect 5770 0 5800 10
rect 5870 80 5900 117
rect 5970 80 6000 117
rect 5870 70 6000 80
rect 5870 36 5918 70
rect 5952 36 6000 70
rect 5870 26 6000 36
rect 5870 0 5900 26
rect 5970 0 6000 26
rect 6070 64 6100 117
rect 6170 64 6200 117
rect 6070 54 6200 64
rect 6070 20 6118 54
rect 6152 20 6200 54
rect 6070 10 6200 20
rect 6070 0 6100 10
rect 6170 0 6200 10
rect 6270 80 6300 117
rect 6370 80 6400 117
rect 6270 70 6400 80
rect 6270 36 6318 70
rect 6352 36 6400 70
rect 6270 26 6400 36
rect 6270 0 6300 26
rect 6370 0 6400 26
rect 6470 64 6500 117
rect 6570 64 6600 117
rect 6470 54 6600 64
rect 6470 20 6518 54
rect 6552 20 6600 54
rect 6470 10 6600 20
rect 6470 0 6500 10
rect 6570 0 6600 10
rect 6670 80 6700 117
rect 6770 80 6800 117
rect 6670 70 6800 80
rect 6670 36 6718 70
rect 6752 36 6800 70
rect 6670 26 6800 36
rect 6670 0 6700 26
rect 6770 0 6800 26
rect 6870 64 6900 117
rect 6970 64 7000 117
rect 6870 54 7000 64
rect 6870 20 6918 54
rect 6952 20 7000 54
rect 6870 10 7000 20
rect 6870 0 6900 10
rect 6970 0 7000 10
rect 7070 80 7100 257
rect 7170 203 7200 257
rect 7270 203 7300 257
rect 7370 203 7400 257
rect 7470 203 7500 257
rect 7570 203 7600 257
rect 7670 203 7700 257
rect 7770 203 7800 257
rect 7870 203 7900 397
rect 7970 343 8000 397
rect 7970 203 8000 257
rect 8070 203 8100 397
rect 8170 343 8200 397
rect 8270 343 8300 397
rect 8370 343 8400 677
rect 8470 623 8500 677
rect 8570 623 8600 677
rect 8670 623 8700 677
rect 8770 623 8800 677
rect 8870 623 8900 677
rect 8970 623 9000 677
rect 9070 623 9100 677
rect 9170 623 9200 817
rect 9270 763 9300 817
rect 9270 623 9300 677
rect 9370 623 9400 817
rect 9470 763 9500 817
rect 9570 763 9600 817
rect 9470 623 9500 677
rect 9570 623 9600 677
rect 9670 623 9700 817
rect 9770 763 9800 817
rect 9770 623 9800 677
rect 9870 623 9900 817
rect 9970 763 10000 1097
rect 10070 1043 10100 1097
rect 10170 1043 10200 1097
rect 10270 1043 10300 1097
rect 10070 903 10100 957
rect 10170 903 10200 957
rect 10270 903 10300 957
rect 10370 903 10400 1097
rect 10470 1043 10500 1097
rect 10570 1043 10600 1097
rect 10670 1043 10700 1097
rect 10770 1043 10800 1097
rect 10870 1043 10900 1097
rect 10970 1043 11000 1097
rect 11070 1043 11100 1236
rect 11170 1183 11200 1236
rect 11270 1274 11300 1327
rect 11370 1274 11400 1327
rect 11270 1264 11400 1274
rect 11270 1230 11318 1264
rect 11352 1230 11400 1264
rect 11270 1220 11400 1230
rect 11170 1043 11200 1097
rect 11270 1043 11300 1220
rect 11370 1183 11400 1220
rect 11470 1290 11500 1327
rect 11570 1290 11600 1327
rect 11470 1280 11600 1290
rect 11470 1246 11518 1280
rect 11552 1246 11600 1280
rect 11470 1236 11600 1246
rect 10470 903 10500 957
rect 10570 903 10600 957
rect 10670 903 10700 957
rect 10070 763 10100 817
rect 9970 623 10000 677
rect 10070 623 10100 677
rect 10170 623 10200 817
rect 10270 763 10300 817
rect 10370 763 10400 817
rect 10470 763 10500 817
rect 10570 763 10600 817
rect 10670 763 10700 817
rect 10770 763 10800 957
rect 10870 903 10900 957
rect 10870 763 10900 817
rect 8470 483 8500 537
rect 8570 483 8600 537
rect 8670 483 8700 537
rect 8770 483 8800 537
rect 8870 483 8900 537
rect 8970 483 9000 537
rect 9070 483 9100 537
rect 9170 483 9200 537
rect 9270 483 9300 537
rect 9370 483 9400 537
rect 9470 483 9500 537
rect 9570 483 9600 537
rect 9670 483 9700 537
rect 9770 483 9800 537
rect 9870 483 9900 537
rect 8470 343 8500 397
rect 8570 343 8600 397
rect 8670 343 8700 397
rect 8170 203 8200 257
rect 8270 203 8300 257
rect 8370 203 8400 257
rect 8470 203 8500 257
rect 8570 203 8600 257
rect 8670 203 8700 257
rect 8770 203 8800 397
rect 8870 343 8900 397
rect 8970 343 9000 397
rect 8870 203 8900 257
rect 8970 203 9000 257
rect 9070 203 9100 397
rect 9170 343 9200 397
rect 9170 203 9200 257
rect 9270 203 9300 397
rect 9370 343 9400 397
rect 9470 343 9500 397
rect 9570 343 9600 397
rect 9670 343 9700 397
rect 9770 343 9800 397
rect 9870 343 9900 397
rect 9970 343 10000 537
rect 10070 483 10100 537
rect 10170 483 10200 537
rect 10070 343 10100 397
rect 9370 203 9400 257
rect 9470 203 9500 257
rect 9570 203 9600 257
rect 9670 203 9700 257
rect 9770 203 9800 257
rect 9870 203 9900 257
rect 9970 203 10000 257
rect 10070 203 10100 257
rect 10170 203 10200 397
rect 10270 343 10300 677
rect 10370 623 10400 677
rect 10370 483 10400 537
rect 10470 483 10500 677
rect 10570 623 10600 677
rect 10670 623 10700 677
rect 10770 623 10800 677
rect 10870 623 10900 677
rect 10970 623 11000 957
rect 11070 903 11100 957
rect 11170 903 11200 957
rect 11270 903 11300 957
rect 11370 903 11400 1097
rect 11470 1043 11500 1236
rect 11570 1183 11600 1236
rect 11670 1274 11700 1327
rect 11770 1274 11800 1467
rect 11870 1413 11900 1467
rect 11970 1413 12000 1467
rect 12070 1413 12100 1607
rect 12170 1553 12200 1607
rect 12270 1553 12300 1607
rect 12370 1553 12400 1607
rect 12170 1413 12200 1467
rect 12270 1413 12300 1467
rect 12370 1413 12400 1467
rect 11670 1264 11800 1274
rect 11670 1230 11718 1264
rect 11752 1230 11800 1264
rect 11670 1220 11800 1230
rect 11670 1183 11700 1220
rect 11770 1183 11800 1220
rect 11870 1290 11900 1327
rect 11970 1290 12000 1327
rect 11870 1280 12000 1290
rect 11870 1246 11918 1280
rect 11952 1246 12000 1280
rect 11870 1236 12000 1246
rect 11870 1183 11900 1236
rect 11970 1183 12000 1236
rect 12070 1274 12100 1327
rect 12170 1274 12200 1327
rect 12070 1264 12200 1274
rect 12070 1230 12118 1264
rect 12152 1230 12200 1264
rect 12070 1220 12200 1230
rect 11570 1043 11600 1097
rect 11470 903 11500 957
rect 11570 903 11600 957
rect 11670 903 11700 1097
rect 11770 1043 11800 1097
rect 11870 1043 11900 1097
rect 11770 903 11800 957
rect 11870 903 11900 957
rect 11070 763 11100 817
rect 11170 763 11200 817
rect 11270 763 11300 817
rect 11370 763 11400 817
rect 11470 763 11500 817
rect 11570 763 11600 817
rect 11670 763 11700 817
rect 11070 623 11100 677
rect 11170 623 11200 677
rect 10570 483 10600 537
rect 10670 483 10700 537
rect 10770 483 10800 537
rect 10370 343 10400 397
rect 10470 343 10500 397
rect 10570 343 10600 397
rect 10670 343 10700 397
rect 10770 343 10800 397
rect 10870 343 10900 537
rect 10970 483 11000 537
rect 11070 483 11100 537
rect 10970 343 11000 397
rect 11070 343 11100 397
rect 11170 343 11200 537
rect 11270 483 11300 677
rect 11370 623 11400 677
rect 11470 623 11500 677
rect 11570 623 11600 677
rect 11670 623 11700 677
rect 11770 623 11800 817
rect 11870 763 11900 817
rect 11970 763 12000 1097
rect 12070 1043 12100 1220
rect 12170 1183 12200 1220
rect 12270 1290 12300 1327
rect 12370 1290 12400 1327
rect 12270 1280 12400 1290
rect 12270 1246 12318 1280
rect 12352 1246 12400 1280
rect 12270 1236 12400 1246
rect 12270 1183 12300 1236
rect 12370 1183 12400 1236
rect 12470 1274 12500 1607
rect 12570 1553 12600 1607
rect 12670 1553 12700 1607
rect 12770 1553 12800 1607
rect 12970 1553 13000 1607
rect 13070 1553 13100 1607
rect 13280 1553 13310 1607
rect 13380 1553 13410 1607
rect 13480 1553 13510 1607
rect 13580 1553 13610 1607
rect 12570 1413 12600 1467
rect 12670 1413 12700 1467
rect 12770 1413 12800 1467
rect 12970 1413 13000 1467
rect 13070 1413 13100 1467
rect 13280 1413 13310 1467
rect 13380 1413 13410 1467
rect 13480 1413 13510 1467
rect 13580 1413 13610 1467
rect 12570 1274 12600 1327
rect 12470 1264 12600 1274
rect 12470 1230 12518 1264
rect 12552 1230 12600 1264
rect 12470 1220 12600 1230
rect 12470 1183 12500 1220
rect 12570 1183 12600 1220
rect 12670 1290 12700 1327
rect 12770 1290 12800 1327
rect 12970 1294 13000 1327
rect 13070 1294 13100 1327
rect 13280 1294 13310 1327
rect 13380 1294 13410 1327
rect 13480 1294 13510 1327
rect 13580 1294 13610 1327
rect 12670 1280 12800 1290
rect 12670 1246 12718 1280
rect 12752 1246 12800 1280
rect 12670 1236 12800 1246
rect 12170 1043 12200 1097
rect 12270 1043 12300 1097
rect 12370 1043 12400 1097
rect 12470 1043 12500 1097
rect 12570 1043 12600 1097
rect 12670 1043 12700 1236
rect 12770 1183 12800 1236
rect 12958 1278 13012 1294
rect 12958 1244 12968 1278
rect 13002 1244 13012 1278
rect 12958 1228 13012 1244
rect 13058 1278 13112 1294
rect 13058 1244 13068 1278
rect 13102 1244 13112 1278
rect 13058 1228 13112 1244
rect 13268 1278 13322 1294
rect 13268 1244 13278 1278
rect 13312 1244 13322 1278
rect 13268 1228 13322 1244
rect 13368 1278 13422 1294
rect 13368 1244 13378 1278
rect 13412 1244 13422 1278
rect 13368 1228 13422 1244
rect 13468 1278 13522 1294
rect 13468 1244 13478 1278
rect 13512 1244 13522 1278
rect 13468 1228 13522 1244
rect 13568 1278 13622 1294
rect 13568 1244 13578 1278
rect 13612 1244 13622 1278
rect 13568 1228 13622 1244
rect 12970 1183 13000 1228
rect 13070 1183 13100 1228
rect 13280 1183 13310 1228
rect 13380 1183 13410 1228
rect 13480 1183 13510 1228
rect 13580 1183 13610 1228
rect 12770 1043 12800 1097
rect 12970 1043 13000 1097
rect 13070 1043 13100 1097
rect 13280 1043 13310 1097
rect 13380 1043 13410 1097
rect 13480 1043 13510 1097
rect 13580 1043 13610 1097
rect 12070 903 12100 957
rect 12170 903 12200 957
rect 12270 903 12300 957
rect 12070 763 12100 817
rect 11870 623 11900 677
rect 11970 623 12000 677
rect 12070 623 12100 677
rect 12170 623 12200 817
rect 12270 763 12300 817
rect 12370 763 12400 957
rect 12470 903 12500 957
rect 12470 763 12500 817
rect 12570 763 12600 957
rect 12670 903 12700 957
rect 12770 903 12800 957
rect 12970 903 13000 957
rect 13070 903 13100 957
rect 13280 903 13310 957
rect 13380 903 13410 957
rect 13480 903 13510 957
rect 13580 903 13610 957
rect 12670 763 12700 817
rect 12770 763 12800 817
rect 12970 763 13000 817
rect 13070 763 13100 817
rect 13280 763 13310 817
rect 13380 763 13410 817
rect 13480 763 13510 817
rect 13580 763 13610 817
rect 12270 623 12300 677
rect 12370 623 12400 677
rect 12470 623 12500 677
rect 12570 623 12600 677
rect 12670 623 12700 677
rect 12770 623 12800 677
rect 12970 623 13000 677
rect 13070 623 13100 677
rect 13280 623 13310 677
rect 13380 623 13410 677
rect 13480 623 13510 677
rect 13580 623 13610 677
rect 11270 343 11300 397
rect 11370 343 11400 537
rect 11470 483 11500 537
rect 11570 483 11600 537
rect 11670 483 11700 537
rect 11770 483 11800 537
rect 11870 483 11900 537
rect 11970 483 12000 537
rect 12070 483 12100 537
rect 12170 483 12200 537
rect 12270 483 12300 537
rect 10270 203 10300 257
rect 10370 203 10400 257
rect 10470 203 10500 257
rect 10570 203 10600 257
rect 10670 203 10700 257
rect 10770 203 10800 257
rect 10870 203 10900 257
rect 10970 203 11000 257
rect 11070 203 11100 257
rect 11170 203 11200 257
rect 11270 203 11300 257
rect 11370 203 11400 257
rect 7170 80 7200 117
rect 7070 70 7200 80
rect 7070 36 7118 70
rect 7152 36 7200 70
rect 7070 26 7200 36
rect 7070 0 7100 26
rect 7170 0 7200 26
rect 7270 64 7300 117
rect 7370 64 7400 117
rect 7270 54 7400 64
rect 7270 20 7318 54
rect 7352 20 7400 54
rect 7270 10 7400 20
rect 7270 0 7300 10
rect 7370 0 7400 10
rect 7470 80 7500 117
rect 7570 80 7600 117
rect 7470 70 7600 80
rect 7470 36 7518 70
rect 7552 36 7600 70
rect 7470 26 7600 36
rect 7470 0 7500 26
rect 7570 0 7600 26
rect 7670 64 7700 117
rect 7770 64 7800 117
rect 7670 54 7800 64
rect 7670 20 7718 54
rect 7752 20 7800 54
rect 7670 10 7800 20
rect 7670 0 7700 10
rect 7770 0 7800 10
rect 7870 80 7900 117
rect 7970 80 8000 117
rect 7870 70 8000 80
rect 7870 36 7918 70
rect 7952 36 8000 70
rect 7870 26 8000 36
rect 7870 0 7900 26
rect 7970 0 8000 26
rect 8070 64 8100 117
rect 8170 64 8200 117
rect 8070 54 8200 64
rect 8070 20 8118 54
rect 8152 20 8200 54
rect 8070 10 8200 20
rect 8070 0 8100 10
rect 8170 0 8200 10
rect 8270 80 8300 117
rect 8370 80 8400 117
rect 8270 70 8400 80
rect 8270 36 8318 70
rect 8352 36 8400 70
rect 8270 26 8400 36
rect 8270 0 8300 26
rect 8370 0 8400 26
rect 8470 64 8500 117
rect 8570 64 8600 117
rect 8470 54 8600 64
rect 8470 20 8518 54
rect 8552 20 8600 54
rect 8470 10 8600 20
rect 8470 0 8500 10
rect 8570 0 8600 10
rect 8670 80 8700 117
rect 8770 80 8800 117
rect 8670 70 8800 80
rect 8670 36 8718 70
rect 8752 36 8800 70
rect 8670 26 8800 36
rect 8670 0 8700 26
rect 8770 0 8800 26
rect 8870 64 8900 117
rect 8970 64 9000 117
rect 8870 54 9000 64
rect 8870 20 8918 54
rect 8952 20 9000 54
rect 8870 10 9000 20
rect 8870 0 8900 10
rect 8970 0 9000 10
rect 9070 80 9100 117
rect 9170 80 9200 117
rect 9070 70 9200 80
rect 9070 36 9118 70
rect 9152 36 9200 70
rect 9070 26 9200 36
rect 9070 0 9100 26
rect 9170 0 9200 26
rect 9270 64 9300 117
rect 9370 64 9400 117
rect 9270 54 9400 64
rect 9270 20 9318 54
rect 9352 20 9400 54
rect 9270 10 9400 20
rect 9270 0 9300 10
rect 9370 0 9400 10
rect 9470 80 9500 117
rect 9570 80 9600 117
rect 9470 70 9600 80
rect 9470 36 9518 70
rect 9552 36 9600 70
rect 9470 26 9600 36
rect 9470 0 9500 26
rect 9570 0 9600 26
rect 9670 64 9700 117
rect 9770 64 9800 117
rect 9670 54 9800 64
rect 9670 20 9718 54
rect 9752 20 9800 54
rect 9670 10 9800 20
rect 9670 0 9700 10
rect 9770 0 9800 10
rect 9870 80 9900 117
rect 9970 80 10000 117
rect 9870 70 10000 80
rect 9870 36 9918 70
rect 9952 36 10000 70
rect 9870 26 10000 36
rect 9870 0 9900 26
rect 9970 0 10000 26
rect 10070 64 10100 117
rect 10170 64 10200 117
rect 10070 54 10200 64
rect 10070 20 10118 54
rect 10152 20 10200 54
rect 10070 10 10200 20
rect 10070 0 10100 10
rect 10170 0 10200 10
rect 10270 80 10300 117
rect 10370 80 10400 117
rect 10270 70 10400 80
rect 10270 36 10318 70
rect 10352 36 10400 70
rect 10270 26 10400 36
rect 10270 0 10300 26
rect 10370 0 10400 26
rect 10470 64 10500 117
rect 10570 64 10600 117
rect 10470 54 10600 64
rect 10470 20 10518 54
rect 10552 20 10600 54
rect 10470 10 10600 20
rect 10470 0 10500 10
rect 10570 0 10600 10
rect 10670 80 10700 117
rect 10770 80 10800 117
rect 10670 70 10800 80
rect 10670 36 10718 70
rect 10752 36 10800 70
rect 10670 26 10800 36
rect 10670 0 10700 26
rect 10770 0 10800 26
rect 10870 64 10900 117
rect 10970 64 11000 117
rect 10870 54 11000 64
rect 10870 20 10918 54
rect 10952 20 11000 54
rect 10870 10 11000 20
rect 10870 0 10900 10
rect 10970 0 11000 10
rect 11070 80 11100 117
rect 11170 80 11200 117
rect 11070 70 11200 80
rect 11070 36 11118 70
rect 11152 36 11200 70
rect 11070 26 11200 36
rect 11070 0 11100 26
rect 11170 0 11200 26
rect 11270 64 11300 117
rect 11370 64 11400 117
rect 11270 54 11400 64
rect 11270 20 11318 54
rect 11352 20 11400 54
rect 11270 10 11400 20
rect 11270 0 11300 10
rect 11370 0 11400 10
rect 11470 80 11500 397
rect 11570 343 11600 397
rect 11670 343 11700 397
rect 11770 343 11800 397
rect 11870 343 11900 397
rect 11970 343 12000 397
rect 12070 343 12100 397
rect 12170 343 12200 397
rect 11570 203 11600 257
rect 11670 203 11700 257
rect 11770 203 11800 257
rect 11870 203 11900 257
rect 11970 203 12000 257
rect 12070 203 12100 257
rect 12170 203 12200 257
rect 12270 203 12300 397
rect 12370 343 12400 537
rect 12470 483 12500 537
rect 12570 483 12600 537
rect 12670 483 12700 537
rect 12770 483 12800 537
rect 12970 483 13000 537
rect 13070 483 13100 537
rect 13280 483 13310 537
rect 13380 483 13410 537
rect 13480 483 13510 537
rect 13580 483 13610 537
rect 12470 343 12500 397
rect 12570 343 12600 397
rect 12670 343 12700 397
rect 12770 343 12800 397
rect 12970 343 13000 397
rect 13070 343 13100 397
rect 13280 343 13310 397
rect 13380 343 13410 397
rect 13480 343 13510 397
rect 13580 343 13610 397
rect 12370 203 12400 257
rect 12470 203 12500 257
rect 12570 203 12600 257
rect 12670 203 12700 257
rect 12770 203 12800 257
rect 12970 203 13000 257
rect 13070 203 13100 257
rect 13280 203 13310 257
rect 13380 203 13410 257
rect 13480 203 13510 257
rect 13580 203 13610 257
rect 11570 80 11600 117
rect 11470 70 11600 80
rect 11470 36 11518 70
rect 11552 36 11600 70
rect 11470 26 11600 36
rect 11470 0 11500 26
rect 11570 0 11600 26
rect 11670 64 11700 117
rect 11770 64 11800 117
rect 11670 54 11800 64
rect 11670 20 11718 54
rect 11752 20 11800 54
rect 11670 10 11800 20
rect 11670 0 11700 10
rect 11770 0 11800 10
rect 11870 80 11900 117
rect 11970 80 12000 117
rect 11870 70 12000 80
rect 11870 36 11918 70
rect 11952 36 12000 70
rect 11870 26 12000 36
rect 11870 0 11900 26
rect 11970 0 12000 26
rect 12070 64 12100 117
rect 12170 64 12200 117
rect 12070 54 12200 64
rect 12070 20 12118 54
rect 12152 20 12200 54
rect 12070 10 12200 20
rect 12070 0 12100 10
rect 12170 0 12200 10
rect 12270 80 12300 117
rect 12370 80 12400 117
rect 12270 70 12400 80
rect 12270 36 12318 70
rect 12352 36 12400 70
rect 12270 26 12400 36
rect 12270 0 12300 26
rect 12370 0 12400 26
rect 12470 64 12500 117
rect 12570 64 12600 117
rect 12470 54 12600 64
rect 12470 20 12518 54
rect 12552 20 12600 54
rect 12470 10 12600 20
rect 12470 0 12500 10
rect 12570 0 12600 10
rect 12670 80 12700 117
rect 12770 80 12800 117
rect 12970 84 13000 117
rect 13070 84 13100 117
rect 13280 84 13310 117
rect 13380 84 13410 117
rect 13480 84 13510 117
rect 13580 84 13610 117
rect 12670 70 12800 80
rect 12670 36 12718 70
rect 12752 36 12800 70
rect 12670 26 12800 36
rect 12670 0 12700 26
rect 12770 0 12800 26
rect 12958 68 13012 84
rect 12958 34 12968 68
rect 13002 34 13012 68
rect 12958 18 13012 34
rect 13058 68 13112 84
rect 13058 34 13068 68
rect 13102 34 13112 68
rect 13058 18 13112 34
rect 13268 68 13322 84
rect 13268 34 13278 68
rect 13312 34 13322 68
rect 13268 18 13322 34
rect 13368 68 13422 84
rect 13368 34 13378 68
rect 13412 34 13422 68
rect 13368 18 13422 34
rect 13468 68 13522 84
rect 13468 34 13478 68
rect 13512 34 13522 68
rect 13468 18 13522 34
rect 13568 68 13622 84
rect 13568 34 13578 68
rect 13612 34 13622 68
rect 13568 18 13622 34
rect 12970 0 13000 18
rect 13070 0 13100 18
rect 13280 0 13310 18
rect 13380 0 13410 18
rect 13480 0 13510 18
rect 13580 0 13610 18
rect -30 -126 0 -100
rect 70 -126 100 -100
rect 170 -126 200 -100
rect 270 -126 300 -100
rect 370 -126 400 -100
rect 470 -126 500 -100
rect 570 -126 600 -100
rect 670 -126 700 -100
rect 770 -126 800 -100
rect 870 -126 900 -100
rect 970 -126 1000 -100
rect 1070 -126 1100 -100
rect 1170 -126 1200 -100
rect 1270 -126 1300 -100
rect 1370 -126 1400 -100
rect 1470 -126 1500 -100
rect 1570 -126 1600 -100
rect 1670 -126 1700 -100
rect 1770 -126 1800 -100
rect 1870 -126 1900 -100
rect 1970 -126 2000 -100
rect 2070 -126 2100 -100
rect 2170 -126 2200 -100
rect 2270 -126 2300 -100
rect 2370 -126 2400 -100
rect 2470 -126 2500 -100
rect 2570 -126 2600 -100
rect 2670 -126 2700 -100
rect 2770 -126 2800 -100
rect 2870 -126 2900 -100
rect 2970 -126 3000 -100
rect 3070 -126 3100 -100
rect 3170 -126 3200 -100
rect 3270 -126 3300 -100
rect 3370 -126 3400 -100
rect 3470 -126 3500 -100
rect 3570 -126 3600 -100
rect 3670 -126 3700 -100
rect 3770 -126 3800 -100
rect 3870 -126 3900 -100
rect 3970 -126 4000 -100
rect 4070 -126 4100 -100
rect 4170 -126 4200 -100
rect 4270 -126 4300 -100
rect 4370 -126 4400 -100
rect 4470 -126 4500 -100
rect 4570 -126 4600 -100
rect 4670 -126 4700 -100
rect 4770 -126 4800 -100
rect 4870 -126 4900 -100
rect 4970 -126 5000 -100
rect 5070 -126 5100 -100
rect 5170 -126 5200 -100
rect 5270 -126 5300 -100
rect 5370 -126 5400 -100
rect 5470 -126 5500 -100
rect 5570 -126 5600 -100
rect 5670 -126 5700 -100
rect 5770 -126 5800 -100
rect 5870 -126 5900 -100
rect 5970 -126 6000 -100
rect 6070 -126 6100 -100
rect 6170 -126 6200 -100
rect 6270 -126 6300 -100
rect 6370 -126 6400 -100
rect 6470 -126 6500 -100
rect 6570 -126 6600 -100
rect 6670 -126 6700 -100
rect 6770 -126 6800 -100
rect 6870 -126 6900 -100
rect 6970 -126 7000 -100
rect 7070 -126 7100 -100
rect 7170 -126 7200 -100
rect 7270 -126 7300 -100
rect 7370 -126 7400 -100
rect 7470 -126 7500 -100
rect 7570 -126 7600 -100
rect 7670 -126 7700 -100
rect 7770 -126 7800 -100
rect 7870 -126 7900 -100
rect 7970 -126 8000 -100
rect 8070 -126 8100 -100
rect 8170 -126 8200 -100
rect 8270 -126 8300 -100
rect 8370 -126 8400 -100
rect 8470 -126 8500 -100
rect 8570 -126 8600 -100
rect 8670 -126 8700 -100
rect 8770 -126 8800 -100
rect 8870 -126 8900 -100
rect 8970 -126 9000 -100
rect 9070 -126 9100 -100
rect 9170 -126 9200 -100
rect 9270 -126 9300 -100
rect 9370 -126 9400 -100
rect 9470 -126 9500 -100
rect 9570 -126 9600 -100
rect 9670 -126 9700 -100
rect 9770 -126 9800 -100
rect 9870 -126 9900 -100
rect 9970 -126 10000 -100
rect 10070 -126 10100 -100
rect 10170 -126 10200 -100
rect 10270 -126 10300 -100
rect 10370 -126 10400 -100
rect 10470 -126 10500 -100
rect 10570 -126 10600 -100
rect 10670 -126 10700 -100
rect 10770 -126 10800 -100
rect 10870 -126 10900 -100
rect 10970 -126 11000 -100
rect 11070 -126 11100 -100
rect 11170 -126 11200 -100
rect 11270 -126 11300 -100
rect 11370 -126 11400 -100
rect 11470 -126 11500 -100
rect 11570 -126 11600 -100
rect 11670 -126 11700 -100
rect 11770 -126 11800 -100
rect 11870 -126 11900 -100
rect 11970 -126 12000 -100
rect 12070 -126 12100 -100
rect 12170 -126 12200 -100
rect 12270 -126 12300 -100
rect 12370 -126 12400 -100
rect 12470 -126 12500 -100
rect 12570 -126 12600 -100
rect 12670 -126 12700 -100
rect -30 -226 0 -210
rect 70 -226 100 -210
rect -30 -248 100 -226
rect -30 -282 18 -248
rect 52 -282 100 -248
rect -30 -314 100 -282
rect -30 -330 0 -314
rect 70 -330 100 -314
rect 170 -226 200 -210
rect 270 -226 300 -210
rect 170 -248 300 -226
rect 170 -282 218 -248
rect 252 -282 300 -248
rect 170 -314 300 -282
rect 170 -330 200 -314
rect 270 -330 300 -314
rect 370 -226 400 -210
rect 470 -226 500 -210
rect 370 -248 500 -226
rect 370 -282 418 -248
rect 452 -282 500 -248
rect 370 -314 500 -282
rect 370 -330 400 -314
rect 470 -330 500 -314
rect 570 -226 600 -210
rect 670 -226 700 -210
rect 570 -248 700 -226
rect 570 -282 618 -248
rect 652 -282 700 -248
rect 570 -314 700 -282
rect 570 -330 600 -314
rect 670 -330 700 -314
rect 770 -226 800 -210
rect 870 -226 900 -210
rect 770 -248 900 -226
rect 770 -282 818 -248
rect 852 -282 900 -248
rect 770 -314 900 -282
rect 770 -330 800 -314
rect 870 -330 900 -314
rect 970 -226 1000 -210
rect 1070 -226 1100 -210
rect 970 -248 1100 -226
rect 970 -282 1018 -248
rect 1052 -282 1100 -248
rect 970 -314 1100 -282
rect 970 -330 1000 -314
rect 1070 -330 1100 -314
rect 1170 -226 1200 -210
rect 1270 -226 1300 -210
rect 1170 -248 1300 -226
rect 1170 -282 1218 -248
rect 1252 -282 1300 -248
rect 1170 -314 1300 -282
rect 1170 -330 1200 -314
rect 1270 -330 1300 -314
rect 1370 -226 1400 -210
rect 1470 -226 1500 -210
rect 1370 -248 1500 -226
rect 1370 -282 1418 -248
rect 1452 -282 1500 -248
rect 1370 -314 1500 -282
rect 1370 -330 1400 -314
rect 1470 -330 1500 -314
rect 1570 -226 1600 -210
rect 1670 -226 1700 -210
rect 1570 -248 1700 -226
rect 1570 -282 1618 -248
rect 1652 -282 1700 -248
rect 1570 -314 1700 -282
rect 1570 -330 1600 -314
rect 1670 -330 1700 -314
rect 1770 -226 1800 -210
rect 1870 -226 1900 -210
rect 1770 -248 1900 -226
rect 1770 -282 1818 -248
rect 1852 -282 1900 -248
rect 1770 -314 1900 -282
rect 1770 -330 1800 -314
rect 1870 -330 1900 -314
rect 1970 -226 2000 -210
rect 2070 -226 2100 -210
rect 1970 -248 2100 -226
rect 1970 -282 2018 -248
rect 2052 -282 2100 -248
rect 1970 -314 2100 -282
rect 1970 -330 2000 -314
rect 2070 -330 2100 -314
rect 2170 -226 2200 -210
rect 2270 -226 2300 -210
rect 2170 -248 2300 -226
rect 2170 -282 2218 -248
rect 2252 -282 2300 -248
rect 2170 -314 2300 -282
rect 2170 -330 2200 -314
rect 2270 -330 2300 -314
rect 2370 -226 2400 -210
rect 2470 -226 2500 -210
rect 2370 -248 2500 -226
rect 2370 -282 2418 -248
rect 2452 -282 2500 -248
rect 2370 -314 2500 -282
rect 2370 -330 2400 -314
rect 2470 -330 2500 -314
rect 2570 -226 2600 -210
rect 2670 -226 2700 -210
rect 2570 -248 2700 -226
rect 2570 -282 2618 -248
rect 2652 -282 2700 -248
rect 2570 -314 2700 -282
rect 2570 -330 2600 -314
rect 2670 -330 2700 -314
rect 2770 -226 2800 -210
rect 2870 -226 2900 -210
rect 2770 -248 2900 -226
rect 2770 -282 2818 -248
rect 2852 -282 2900 -248
rect 2770 -314 2900 -282
rect 2770 -330 2800 -314
rect 2870 -330 2900 -314
rect 2970 -226 3000 -210
rect 3070 -226 3100 -210
rect 2970 -248 3100 -226
rect 2970 -282 3018 -248
rect 3052 -282 3100 -248
rect 2970 -314 3100 -282
rect 2970 -330 3000 -314
rect 3070 -330 3100 -314
rect 3170 -226 3200 -210
rect 3270 -226 3300 -210
rect 3170 -248 3300 -226
rect 3170 -282 3218 -248
rect 3252 -282 3300 -248
rect 3170 -314 3300 -282
rect 3170 -330 3200 -314
rect 3270 -330 3300 -314
rect 3370 -226 3400 -210
rect 3470 -226 3500 -210
rect 3370 -248 3500 -226
rect 3370 -282 3418 -248
rect 3452 -282 3500 -248
rect 3370 -314 3500 -282
rect 3370 -330 3400 -314
rect 3470 -330 3500 -314
rect 3570 -226 3600 -210
rect 3670 -226 3700 -210
rect 3570 -248 3700 -226
rect 3570 -282 3618 -248
rect 3652 -282 3700 -248
rect 3570 -314 3700 -282
rect 3570 -330 3600 -314
rect 3670 -330 3700 -314
rect 3770 -226 3800 -210
rect 3870 -226 3900 -210
rect 3770 -248 3900 -226
rect 3770 -282 3818 -248
rect 3852 -282 3900 -248
rect 3770 -314 3900 -282
rect 3770 -330 3800 -314
rect 3870 -330 3900 -314
rect 3970 -226 4000 -210
rect 4070 -226 4100 -210
rect 3970 -248 4100 -226
rect 3970 -282 4018 -248
rect 4052 -282 4100 -248
rect 3970 -314 4100 -282
rect 3970 -330 4000 -314
rect 4070 -330 4100 -314
rect 4170 -226 4200 -210
rect 4270 -226 4300 -210
rect 4170 -248 4300 -226
rect 4170 -282 4218 -248
rect 4252 -282 4300 -248
rect 4170 -314 4300 -282
rect 4170 -330 4200 -314
rect 4270 -330 4300 -314
rect 4370 -226 4400 -210
rect 4470 -226 4500 -210
rect 4370 -248 4500 -226
rect 4370 -282 4418 -248
rect 4452 -282 4500 -248
rect 4370 -314 4500 -282
rect 4370 -330 4400 -314
rect 4470 -330 4500 -314
rect 4570 -226 4600 -210
rect 4670 -226 4700 -210
rect 4570 -248 4700 -226
rect 4570 -282 4618 -248
rect 4652 -282 4700 -248
rect 4570 -314 4700 -282
rect 4570 -330 4600 -314
rect 4670 -330 4700 -314
rect 4770 -226 4800 -210
rect 4870 -226 4900 -210
rect 4770 -248 4900 -226
rect 4770 -282 4818 -248
rect 4852 -282 4900 -248
rect 4770 -314 4900 -282
rect 4770 -330 4800 -314
rect 4870 -330 4900 -314
rect 4970 -226 5000 -210
rect 5070 -226 5100 -210
rect 4970 -248 5100 -226
rect 4970 -282 5018 -248
rect 5052 -282 5100 -248
rect 4970 -314 5100 -282
rect 4970 -330 5000 -314
rect 5070 -330 5100 -314
rect 5170 -226 5200 -210
rect 5270 -226 5300 -210
rect 5170 -248 5300 -226
rect 5170 -282 5218 -248
rect 5252 -282 5300 -248
rect 5170 -314 5300 -282
rect 5170 -330 5200 -314
rect 5270 -330 5300 -314
rect 5370 -226 5400 -210
rect 5470 -226 5500 -210
rect 5370 -248 5500 -226
rect 5370 -282 5418 -248
rect 5452 -282 5500 -248
rect 5370 -314 5500 -282
rect 5370 -330 5400 -314
rect 5470 -330 5500 -314
rect 5570 -226 5600 -210
rect 5670 -226 5700 -210
rect 5570 -248 5700 -226
rect 5570 -282 5618 -248
rect 5652 -282 5700 -248
rect 5570 -314 5700 -282
rect 5570 -330 5600 -314
rect 5670 -330 5700 -314
rect 5770 -226 5800 -210
rect 5870 -226 5900 -210
rect 5770 -248 5900 -226
rect 5770 -282 5818 -248
rect 5852 -282 5900 -248
rect 5770 -314 5900 -282
rect 5770 -330 5800 -314
rect 5870 -330 5900 -314
rect 5970 -226 6000 -210
rect 6070 -226 6100 -210
rect 5970 -248 6100 -226
rect 5970 -282 6018 -248
rect 6052 -282 6100 -248
rect 5970 -314 6100 -282
rect 5970 -330 6000 -314
rect 6070 -330 6100 -314
rect 6170 -226 6200 -210
rect 6270 -226 6300 -210
rect 6170 -248 6300 -226
rect 6170 -282 6218 -248
rect 6252 -282 6300 -248
rect 6170 -314 6300 -282
rect 6170 -330 6200 -314
rect 6270 -330 6300 -314
rect 6370 -226 6400 -210
rect 6470 -226 6500 -210
rect 6370 -248 6500 -226
rect 6370 -282 6418 -248
rect 6452 -282 6500 -248
rect 6370 -314 6500 -282
rect 6370 -330 6400 -314
rect 6470 -330 6500 -314
rect 6570 -226 6600 -210
rect 6670 -226 6700 -210
rect 6570 -248 6700 -226
rect 6570 -282 6618 -248
rect 6652 -282 6700 -248
rect 6570 -314 6700 -282
rect 6570 -330 6600 -314
rect 6670 -330 6700 -314
rect 6770 -226 6800 -210
rect 6870 -226 6900 -210
rect 6770 -248 6900 -226
rect 6770 -282 6818 -248
rect 6852 -282 6900 -248
rect 6770 -314 6900 -282
rect 6770 -330 6800 -314
rect 6870 -330 6900 -314
rect 6970 -226 7000 -210
rect 7070 -226 7100 -210
rect 6970 -248 7100 -226
rect 6970 -282 7018 -248
rect 7052 -282 7100 -248
rect 6970 -314 7100 -282
rect 6970 -330 7000 -314
rect 7070 -330 7100 -314
rect 7170 -226 7200 -210
rect 7270 -226 7300 -210
rect 7170 -248 7300 -226
rect 7170 -282 7218 -248
rect 7252 -282 7300 -248
rect 7170 -314 7300 -282
rect 7170 -330 7200 -314
rect 7270 -330 7300 -314
rect 7370 -226 7400 -210
rect 7470 -226 7500 -210
rect 7370 -248 7500 -226
rect 7370 -282 7418 -248
rect 7452 -282 7500 -248
rect 7370 -314 7500 -282
rect 7370 -330 7400 -314
rect 7470 -330 7500 -314
rect 7570 -226 7600 -210
rect 7670 -226 7700 -210
rect 7570 -248 7700 -226
rect 7570 -282 7618 -248
rect 7652 -282 7700 -248
rect 7570 -314 7700 -282
rect 7570 -330 7600 -314
rect 7670 -330 7700 -314
rect 7770 -226 7800 -210
rect 7870 -226 7900 -210
rect 7770 -248 7900 -226
rect 7770 -282 7818 -248
rect 7852 -282 7900 -248
rect 7770 -314 7900 -282
rect 7770 -330 7800 -314
rect 7870 -330 7900 -314
rect 7970 -226 8000 -210
rect 8070 -226 8100 -210
rect 7970 -248 8100 -226
rect 7970 -282 8018 -248
rect 8052 -282 8100 -248
rect 7970 -314 8100 -282
rect 7970 -330 8000 -314
rect 8070 -330 8100 -314
rect 8170 -226 8200 -210
rect 8270 -226 8300 -210
rect 8170 -248 8300 -226
rect 8170 -282 8218 -248
rect 8252 -282 8300 -248
rect 8170 -314 8300 -282
rect 8170 -330 8200 -314
rect 8270 -330 8300 -314
rect 8370 -226 8400 -210
rect 8470 -226 8500 -210
rect 8370 -248 8500 -226
rect 8370 -282 8418 -248
rect 8452 -282 8500 -248
rect 8370 -314 8500 -282
rect 8370 -330 8400 -314
rect 8470 -330 8500 -314
rect 8570 -226 8600 -210
rect 8670 -226 8700 -210
rect 8570 -248 8700 -226
rect 8570 -282 8618 -248
rect 8652 -282 8700 -248
rect 8570 -314 8700 -282
rect 8570 -330 8600 -314
rect 8670 -330 8700 -314
rect 8770 -226 8800 -210
rect 8870 -226 8900 -210
rect 8770 -248 8900 -226
rect 8770 -282 8818 -248
rect 8852 -282 8900 -248
rect 8770 -314 8900 -282
rect 8770 -330 8800 -314
rect 8870 -330 8900 -314
rect 8970 -226 9000 -210
rect 9070 -226 9100 -210
rect 8970 -248 9100 -226
rect 8970 -282 9018 -248
rect 9052 -282 9100 -248
rect 8970 -314 9100 -282
rect 8970 -330 9000 -314
rect 9070 -330 9100 -314
rect 9170 -226 9200 -210
rect 9270 -226 9300 -210
rect 9170 -248 9300 -226
rect 9170 -282 9218 -248
rect 9252 -282 9300 -248
rect 9170 -314 9300 -282
rect 9170 -330 9200 -314
rect 9270 -330 9300 -314
rect 9370 -226 9400 -210
rect 9470 -226 9500 -210
rect 9370 -248 9500 -226
rect 9370 -282 9418 -248
rect 9452 -282 9500 -248
rect 9370 -314 9500 -282
rect 9370 -330 9400 -314
rect 9470 -330 9500 -314
rect 9570 -226 9600 -210
rect 9670 -226 9700 -210
rect 9570 -248 9700 -226
rect 9570 -282 9618 -248
rect 9652 -282 9700 -248
rect 9570 -314 9700 -282
rect 9570 -330 9600 -314
rect 9670 -330 9700 -314
rect 9770 -226 9800 -210
rect 9870 -226 9900 -210
rect 9770 -248 9900 -226
rect 9770 -282 9818 -248
rect 9852 -282 9900 -248
rect 9770 -314 9900 -282
rect 9770 -330 9800 -314
rect 9870 -330 9900 -314
rect 9970 -226 10000 -210
rect 10070 -226 10100 -210
rect 9970 -248 10100 -226
rect 9970 -282 10018 -248
rect 10052 -282 10100 -248
rect 9970 -314 10100 -282
rect 9970 -330 10000 -314
rect 10070 -330 10100 -314
rect 10170 -226 10200 -210
rect 10270 -226 10300 -210
rect 10170 -248 10300 -226
rect 10170 -282 10218 -248
rect 10252 -282 10300 -248
rect 10170 -314 10300 -282
rect 10170 -330 10200 -314
rect 10270 -330 10300 -314
rect 10370 -226 10400 -210
rect 10470 -226 10500 -210
rect 10370 -248 10500 -226
rect 10370 -282 10418 -248
rect 10452 -282 10500 -248
rect 10370 -314 10500 -282
rect 10370 -330 10400 -314
rect 10470 -330 10500 -314
rect 10570 -226 10600 -210
rect 10670 -226 10700 -210
rect 10570 -248 10700 -226
rect 10570 -282 10618 -248
rect 10652 -282 10700 -248
rect 10570 -314 10700 -282
rect 10570 -330 10600 -314
rect 10670 -330 10700 -314
rect 10770 -226 10800 -210
rect 10870 -226 10900 -210
rect 10770 -248 10900 -226
rect 10770 -282 10818 -248
rect 10852 -282 10900 -248
rect 10770 -314 10900 -282
rect 10770 -330 10800 -314
rect 10870 -330 10900 -314
rect 10970 -226 11000 -210
rect 11070 -226 11100 -210
rect 10970 -248 11100 -226
rect 10970 -282 11018 -248
rect 11052 -282 11100 -248
rect 10970 -314 11100 -282
rect 10970 -330 11000 -314
rect 11070 -330 11100 -314
rect 11170 -226 11200 -210
rect 11270 -226 11300 -210
rect 11170 -248 11300 -226
rect 11170 -282 11218 -248
rect 11252 -282 11300 -248
rect 11170 -314 11300 -282
rect 11170 -330 11200 -314
rect 11270 -330 11300 -314
rect 11370 -226 11400 -210
rect 11470 -226 11500 -210
rect 11370 -248 11500 -226
rect 11370 -282 11418 -248
rect 11452 -282 11500 -248
rect 11370 -314 11500 -282
rect 11370 -330 11400 -314
rect 11470 -330 11500 -314
rect 11570 -226 11600 -210
rect 11670 -226 11700 -210
rect 11570 -248 11700 -226
rect 11570 -282 11618 -248
rect 11652 -282 11700 -248
rect 11570 -314 11700 -282
rect 11570 -330 11600 -314
rect 11670 -330 11700 -314
rect 11770 -226 11800 -210
rect 11870 -226 11900 -210
rect 11770 -248 11900 -226
rect 11770 -282 11818 -248
rect 11852 -282 11900 -248
rect 11770 -314 11900 -282
rect 11770 -330 11800 -314
rect 11870 -330 11900 -314
rect 11970 -226 12000 -210
rect 12070 -226 12100 -210
rect 11970 -248 12100 -226
rect 11970 -282 12018 -248
rect 12052 -282 12100 -248
rect 11970 -314 12100 -282
rect 11970 -330 12000 -314
rect 12070 -330 12100 -314
rect 12170 -226 12200 -210
rect 12270 -226 12300 -210
rect 12170 -248 12300 -226
rect 12170 -282 12218 -248
rect 12252 -282 12300 -248
rect 12170 -314 12300 -282
rect 12170 -330 12200 -314
rect 12270 -330 12300 -314
rect 12370 -226 12400 -210
rect 12470 -226 12500 -210
rect 12370 -248 12500 -226
rect 12370 -282 12418 -248
rect 12452 -282 12500 -248
rect 12370 -314 12500 -282
rect 12370 -330 12400 -314
rect 12470 -330 12500 -314
rect 12570 -226 12600 -210
rect 12670 -226 12700 -210
rect 12570 -248 12700 -226
rect 12570 -282 12618 -248
rect 12652 -282 12700 -248
rect 12570 -314 12700 -282
rect 14514 -290 14540 -260
rect 14690 -290 14816 -260
rect 15116 -290 15142 -260
rect 15200 -290 15226 -260
rect 15526 -290 15652 -260
rect 15802 -290 15828 -260
rect 12570 -330 12600 -314
rect 12670 -330 12700 -314
rect 14706 -309 14800 -290
rect 14706 -343 14734 -309
rect 14768 -343 14800 -309
rect 14706 -360 14800 -343
rect 15542 -309 15636 -290
rect 15542 -343 15574 -309
rect 15608 -343 15636 -309
rect 15542 -360 15636 -343
rect 14514 -390 14540 -360
rect 14690 -390 14816 -360
rect 15116 -390 15142 -360
rect 15200 -390 15226 -360
rect 15526 -390 15652 -360
rect 15802 -390 15828 -360
rect 14514 -490 14540 -460
rect 14690 -490 14816 -460
rect 15116 -490 15142 -460
rect 15200 -490 15226 -460
rect 15526 -490 15652 -460
rect 15802 -490 15828 -460
rect -30 -524 0 -498
rect 70 -524 100 -498
rect 170 -524 200 -498
rect 270 -524 300 -498
rect 370 -524 400 -498
rect 470 -524 500 -498
rect 570 -524 600 -498
rect 670 -524 700 -498
rect 770 -524 800 -498
rect 870 -524 900 -498
rect 970 -524 1000 -498
rect 1070 -524 1100 -498
rect 1170 -524 1200 -498
rect 1270 -524 1300 -498
rect 1370 -524 1400 -498
rect 1470 -524 1500 -498
rect 1570 -524 1600 -498
rect 1670 -524 1700 -498
rect 1770 -524 1800 -498
rect 1870 -524 1900 -498
rect 1970 -524 2000 -498
rect 2070 -524 2100 -498
rect 2170 -524 2200 -498
rect 2270 -524 2300 -498
rect 2370 -524 2400 -498
rect 2470 -524 2500 -498
rect 2570 -524 2600 -498
rect 2670 -524 2700 -498
rect 2770 -524 2800 -498
rect 2870 -524 2900 -498
rect 2970 -524 3000 -498
rect 3070 -524 3100 -498
rect 3170 -524 3200 -498
rect 3270 -524 3300 -498
rect 3370 -524 3400 -498
rect 3470 -524 3500 -498
rect 3570 -524 3600 -498
rect 3670 -524 3700 -498
rect 3770 -524 3800 -498
rect 3870 -524 3900 -498
rect 3970 -524 4000 -498
rect 4070 -524 4100 -498
rect 4170 -524 4200 -498
rect 4270 -524 4300 -498
rect 4370 -524 4400 -498
rect 4470 -524 4500 -498
rect 4570 -524 4600 -498
rect 4670 -524 4700 -498
rect 4770 -524 4800 -498
rect 4870 -524 4900 -498
rect 4970 -524 5000 -498
rect 5070 -524 5100 -498
rect 5170 -524 5200 -498
rect 5270 -524 5300 -498
rect 5370 -524 5400 -498
rect 5470 -524 5500 -498
rect 5570 -524 5600 -498
rect 5670 -524 5700 -498
rect 5770 -524 5800 -498
rect 5870 -524 5900 -498
rect 5970 -524 6000 -498
rect 6070 -524 6100 -498
rect 6170 -524 6200 -498
rect 6270 -524 6300 -498
rect 6370 -524 6400 -498
rect 6470 -524 6500 -498
rect 6570 -524 6600 -498
rect 6670 -524 6700 -498
rect 6770 -524 6800 -498
rect 6870 -524 6900 -498
rect 6970 -524 7000 -498
rect 7070 -524 7100 -498
rect 7170 -524 7200 -498
rect 7270 -524 7300 -498
rect 7370 -524 7400 -498
rect 7470 -524 7500 -498
rect 7570 -524 7600 -498
rect 7670 -524 7700 -498
rect 7770 -524 7800 -498
rect 7870 -524 7900 -498
rect 7970 -524 8000 -498
rect 8070 -524 8100 -498
rect 8170 -524 8200 -498
rect 8270 -524 8300 -498
rect 8370 -524 8400 -498
rect 8470 -524 8500 -498
rect 8570 -524 8600 -498
rect 8670 -524 8700 -498
rect 8770 -524 8800 -498
rect 8870 -524 8900 -498
rect 8970 -524 9000 -498
rect 9070 -524 9100 -498
rect 9170 -524 9200 -498
rect 9270 -524 9300 -498
rect 9370 -524 9400 -498
rect 9470 -524 9500 -498
rect 9570 -524 9600 -498
rect 9670 -524 9700 -498
rect 9770 -524 9800 -498
rect 9870 -524 9900 -498
rect 9970 -524 10000 -498
rect 10070 -524 10100 -498
rect 10170 -524 10200 -498
rect 10270 -524 10300 -498
rect 10370 -524 10400 -498
rect 10470 -524 10500 -498
rect 10570 -524 10600 -498
rect 10670 -524 10700 -498
rect 10770 -524 10800 -498
rect 10870 -524 10900 -498
rect 10970 -524 11000 -498
rect 11070 -524 11100 -498
rect 11170 -524 11200 -498
rect 11270 -524 11300 -498
rect 11370 -524 11400 -498
rect 11470 -524 11500 -498
rect 11570 -524 11600 -498
rect 11670 -524 11700 -498
rect 11770 -524 11800 -498
rect 11870 -524 11900 -498
rect 11970 -524 12000 -498
rect 12070 -524 12100 -498
rect 12170 -524 12200 -498
rect 12270 -524 12300 -498
rect 12370 -524 12400 -498
rect 12470 -524 12500 -498
rect 12570 -524 12600 -498
rect 12670 -524 12700 -498
rect 14706 -509 14800 -490
rect 14706 -543 14734 -509
rect 14768 -543 14800 -509
rect 14706 -560 14800 -543
rect 15542 -509 15636 -490
rect 15542 -543 15574 -509
rect 15608 -543 15636 -509
rect 15542 -560 15636 -543
rect 15 -577 107 -567
rect 15 -611 44 -577
rect 78 -611 107 -577
rect 15 -658 107 -611
rect 163 -577 255 -567
rect 163 -611 192 -577
rect 226 -611 255 -577
rect 415 -577 507 -567
rect 163 -658 255 -611
rect 415 -611 444 -577
rect 478 -611 507 -577
rect 415 -658 507 -611
rect 563 -577 655 -567
rect 563 -611 592 -577
rect 626 -611 655 -577
rect 815 -577 907 -567
rect 563 -658 655 -611
rect 815 -611 844 -577
rect 878 -611 907 -577
rect 815 -658 907 -611
rect 963 -577 1055 -567
rect 963 -611 992 -577
rect 1026 -611 1055 -577
rect 1215 -577 1307 -567
rect 963 -658 1055 -611
rect 1215 -611 1244 -577
rect 1278 -611 1307 -577
rect 1215 -658 1307 -611
rect 1363 -577 1455 -567
rect 1363 -611 1392 -577
rect 1426 -611 1455 -577
rect 1615 -577 1707 -567
rect 1363 -658 1455 -611
rect 1615 -611 1644 -577
rect 1678 -611 1707 -577
rect 1615 -658 1707 -611
rect 1763 -577 1855 -567
rect 1763 -611 1792 -577
rect 1826 -611 1855 -577
rect 2015 -577 2107 -567
rect 1763 -658 1855 -611
rect 2015 -611 2044 -577
rect 2078 -611 2107 -577
rect 2015 -658 2107 -611
rect 2163 -577 2255 -567
rect 2163 -611 2192 -577
rect 2226 -611 2255 -577
rect 2415 -577 2507 -567
rect 2163 -658 2255 -611
rect 2415 -611 2444 -577
rect 2478 -611 2507 -577
rect 2415 -658 2507 -611
rect 2563 -577 2655 -567
rect 2563 -611 2592 -577
rect 2626 -611 2655 -577
rect 2815 -577 2907 -567
rect 2563 -658 2655 -611
rect 2815 -611 2844 -577
rect 2878 -611 2907 -577
rect 2815 -658 2907 -611
rect 2963 -577 3055 -567
rect 2963 -611 2992 -577
rect 3026 -611 3055 -577
rect 3215 -577 3307 -567
rect 2963 -658 3055 -611
rect 3215 -611 3244 -577
rect 3278 -611 3307 -577
rect 3215 -658 3307 -611
rect 3363 -577 3455 -567
rect 3363 -611 3392 -577
rect 3426 -611 3455 -577
rect 3615 -577 3707 -567
rect 3363 -658 3455 -611
rect 3615 -611 3644 -577
rect 3678 -611 3707 -577
rect 3615 -658 3707 -611
rect 3763 -577 3855 -567
rect 3763 -611 3792 -577
rect 3826 -611 3855 -577
rect 4015 -577 4107 -567
rect 3763 -658 3855 -611
rect 4015 -611 4044 -577
rect 4078 -611 4107 -577
rect 4015 -658 4107 -611
rect 4163 -577 4255 -567
rect 4163 -611 4192 -577
rect 4226 -611 4255 -577
rect 4415 -577 4507 -567
rect 4163 -658 4255 -611
rect 4415 -611 4444 -577
rect 4478 -611 4507 -577
rect 4415 -658 4507 -611
rect 4563 -577 4655 -567
rect 4563 -611 4592 -577
rect 4626 -611 4655 -577
rect 4815 -577 4907 -567
rect 4563 -658 4655 -611
rect 4815 -611 4844 -577
rect 4878 -611 4907 -577
rect 4815 -658 4907 -611
rect 4963 -577 5055 -567
rect 4963 -611 4992 -577
rect 5026 -611 5055 -577
rect 5215 -577 5307 -567
rect 4963 -658 5055 -611
rect 5215 -611 5244 -577
rect 5278 -611 5307 -577
rect 5215 -658 5307 -611
rect 5363 -577 5455 -567
rect 5363 -611 5392 -577
rect 5426 -611 5455 -577
rect 5615 -577 5707 -567
rect 5363 -658 5455 -611
rect 5615 -611 5644 -577
rect 5678 -611 5707 -577
rect 5615 -658 5707 -611
rect 5763 -577 5855 -567
rect 5763 -611 5792 -577
rect 5826 -611 5855 -577
rect 6015 -577 6107 -567
rect 5763 -658 5855 -611
rect 6015 -611 6044 -577
rect 6078 -611 6107 -577
rect 6015 -658 6107 -611
rect 6163 -577 6255 -567
rect 6163 -611 6192 -577
rect 6226 -611 6255 -577
rect 6415 -577 6507 -567
rect 6163 -658 6255 -611
rect 6415 -611 6444 -577
rect 6478 -611 6507 -577
rect 6415 -658 6507 -611
rect 6563 -577 6655 -567
rect 6563 -611 6592 -577
rect 6626 -611 6655 -577
rect 6815 -577 6907 -567
rect 6563 -658 6655 -611
rect 6815 -611 6844 -577
rect 6878 -611 6907 -577
rect 6815 -658 6907 -611
rect 6963 -577 7055 -567
rect 6963 -611 6992 -577
rect 7026 -611 7055 -577
rect 7215 -577 7307 -567
rect 6963 -658 7055 -611
rect 7215 -611 7244 -577
rect 7278 -611 7307 -577
rect 7215 -658 7307 -611
rect 7363 -577 7455 -567
rect 7363 -611 7392 -577
rect 7426 -611 7455 -577
rect 7615 -577 7707 -567
rect 7363 -658 7455 -611
rect 7615 -611 7644 -577
rect 7678 -611 7707 -577
rect 7615 -658 7707 -611
rect 7763 -577 7855 -567
rect 7763 -611 7792 -577
rect 7826 -611 7855 -577
rect 8015 -577 8107 -567
rect 7763 -658 7855 -611
rect 8015 -611 8044 -577
rect 8078 -611 8107 -577
rect 8015 -658 8107 -611
rect 8163 -577 8255 -567
rect 8163 -611 8192 -577
rect 8226 -611 8255 -577
rect 8415 -577 8507 -567
rect 8163 -658 8255 -611
rect 8415 -611 8444 -577
rect 8478 -611 8507 -577
rect 8415 -658 8507 -611
rect 8563 -577 8655 -567
rect 8563 -611 8592 -577
rect 8626 -611 8655 -577
rect 8815 -577 8907 -567
rect 8563 -658 8655 -611
rect 8815 -611 8844 -577
rect 8878 -611 8907 -577
rect 8815 -658 8907 -611
rect 8963 -577 9055 -567
rect 8963 -611 8992 -577
rect 9026 -611 9055 -577
rect 9215 -577 9307 -567
rect 8963 -658 9055 -611
rect 9215 -611 9244 -577
rect 9278 -611 9307 -577
rect 9215 -658 9307 -611
rect 9363 -577 9455 -567
rect 9363 -611 9392 -577
rect 9426 -611 9455 -577
rect 9615 -577 9707 -567
rect 9363 -658 9455 -611
rect 9615 -611 9644 -577
rect 9678 -611 9707 -577
rect 9615 -658 9707 -611
rect 9763 -577 9855 -567
rect 9763 -611 9792 -577
rect 9826 -611 9855 -577
rect 10015 -577 10107 -567
rect 9763 -658 9855 -611
rect 10015 -611 10044 -577
rect 10078 -611 10107 -577
rect 10015 -658 10107 -611
rect 10163 -577 10255 -567
rect 10163 -611 10192 -577
rect 10226 -611 10255 -577
rect 10415 -577 10507 -567
rect 10163 -658 10255 -611
rect 10415 -611 10444 -577
rect 10478 -611 10507 -577
rect 10415 -658 10507 -611
rect 10563 -577 10655 -567
rect 10563 -611 10592 -577
rect 10626 -611 10655 -577
rect 10815 -577 10907 -567
rect 10563 -658 10655 -611
rect 10815 -611 10844 -577
rect 10878 -611 10907 -577
rect 10815 -658 10907 -611
rect 10963 -577 11055 -567
rect 10963 -611 10992 -577
rect 11026 -611 11055 -577
rect 11215 -577 11307 -567
rect 10963 -658 11055 -611
rect 11215 -611 11244 -577
rect 11278 -611 11307 -577
rect 11215 -658 11307 -611
rect 11363 -577 11455 -567
rect 11363 -611 11392 -577
rect 11426 -611 11455 -577
rect 11615 -577 11707 -567
rect 11363 -658 11455 -611
rect 11615 -611 11644 -577
rect 11678 -611 11707 -577
rect 11615 -658 11707 -611
rect 11763 -577 11855 -567
rect 11763 -611 11792 -577
rect 11826 -611 11855 -577
rect 12015 -577 12107 -567
rect 11763 -658 11855 -611
rect 12015 -611 12044 -577
rect 12078 -611 12107 -577
rect 12015 -658 12107 -611
rect 12163 -577 12255 -567
rect 12163 -611 12192 -577
rect 12226 -611 12255 -577
rect 12415 -577 12507 -567
rect 12163 -658 12255 -611
rect 12415 -611 12444 -577
rect 12478 -611 12507 -577
rect 12415 -658 12507 -611
rect 12563 -577 12655 -567
rect 12563 -611 12592 -577
rect 12626 -611 12655 -577
rect 14514 -590 14540 -560
rect 14690 -590 14816 -560
rect 15116 -590 15142 -560
rect 15200 -590 15226 -560
rect 15526 -590 15652 -560
rect 15802 -590 15828 -560
rect 12563 -658 12655 -611
rect 14514 -690 14540 -660
rect 14690 -690 14816 -660
rect 15116 -690 15142 -660
rect 15200 -690 15226 -660
rect 15526 -690 15652 -660
rect 15802 -690 15828 -660
rect 15 -768 107 -742
rect 163 -768 255 -742
rect 415 -768 507 -742
rect 563 -768 655 -742
rect 815 -768 907 -742
rect 963 -768 1055 -742
rect 1215 -768 1307 -742
rect 1363 -768 1455 -742
rect 1615 -768 1707 -742
rect 1763 -768 1855 -742
rect 2015 -768 2107 -742
rect 2163 -768 2255 -742
rect 2415 -768 2507 -742
rect 2563 -768 2655 -742
rect 2815 -768 2907 -742
rect 2963 -768 3055 -742
rect 3215 -768 3307 -742
rect 3363 -768 3455 -742
rect 3615 -768 3707 -742
rect 3763 -768 3855 -742
rect 4015 -768 4107 -742
rect 4163 -768 4255 -742
rect 4415 -768 4507 -742
rect 4563 -768 4655 -742
rect 4815 -768 4907 -742
rect 4963 -768 5055 -742
rect 5215 -768 5307 -742
rect 5363 -768 5455 -742
rect 5615 -768 5707 -742
rect 5763 -768 5855 -742
rect 6015 -768 6107 -742
rect 6163 -768 6255 -742
rect 6415 -768 6507 -742
rect 6563 -768 6655 -742
rect 6815 -768 6907 -742
rect 6963 -768 7055 -742
rect 7215 -768 7307 -742
rect 7363 -768 7455 -742
rect 7615 -768 7707 -742
rect 7763 -768 7855 -742
rect 8015 -768 8107 -742
rect 8163 -768 8255 -742
rect 8415 -768 8507 -742
rect 8563 -768 8655 -742
rect 8815 -768 8907 -742
rect 8963 -768 9055 -742
rect 9215 -768 9307 -742
rect 9363 -768 9455 -742
rect 9615 -768 9707 -742
rect 9763 -768 9855 -742
rect 10015 -768 10107 -742
rect 10163 -768 10255 -742
rect 10415 -768 10507 -742
rect 10563 -768 10655 -742
rect 10815 -768 10907 -742
rect 10963 -768 11055 -742
rect 11215 -768 11307 -742
rect 11363 -768 11455 -742
rect 11615 -768 11707 -742
rect 11763 -768 11855 -742
rect 12015 -768 12107 -742
rect 12163 -768 12255 -742
rect 12415 -768 12507 -742
rect 12563 -768 12655 -742
rect 14706 -709 14800 -690
rect 14706 -743 14734 -709
rect 14768 -743 14800 -709
rect 14706 -760 14800 -743
rect 15542 -709 15636 -690
rect 15542 -743 15574 -709
rect 15608 -743 15636 -709
rect 15542 -760 15636 -743
rect 14514 -790 14540 -760
rect 14690 -790 14816 -760
rect 15116 -790 15142 -760
rect 15200 -790 15226 -760
rect 15526 -790 15652 -760
rect 15802 -790 15828 -760
rect -98 -908 -32 -898
rect -98 -910 -82 -908
rect -106 -940 -82 -910
rect -98 -942 -82 -940
rect -48 -910 -32 -908
rect 702 -908 768 -898
rect 702 -910 718 -908
rect -48 -940 -10 -910
rect 108 -940 162 -910
rect 280 -940 390 -910
rect 508 -940 562 -910
rect 680 -940 718 -910
rect -48 -942 -32 -940
rect -98 -952 -32 -942
rect -98 -1008 -32 -998
rect -98 -1010 -82 -1008
rect -106 -1040 -82 -1010
rect -98 -1042 -82 -1040
rect -48 -1010 -32 -1008
rect 702 -942 718 -940
rect 752 -910 768 -908
rect 1502 -908 1568 -898
rect 1502 -910 1518 -908
rect 752 -940 790 -910
rect 908 -940 962 -910
rect 1080 -940 1190 -910
rect 1308 -940 1362 -910
rect 1480 -940 1518 -910
rect 752 -942 768 -940
rect 702 -952 768 -942
rect 702 -1008 768 -998
rect 702 -1010 718 -1008
rect -48 -1040 -10 -1010
rect 108 -1040 162 -1010
rect 280 -1040 390 -1010
rect 508 -1040 562 -1010
rect 680 -1040 718 -1010
rect -48 -1042 -32 -1040
rect -98 -1052 -32 -1042
rect -98 -1108 -32 -1098
rect -98 -1110 -82 -1108
rect -106 -1140 -82 -1110
rect -98 -1142 -82 -1140
rect -48 -1110 -32 -1108
rect 702 -1042 718 -1040
rect 752 -1010 768 -1008
rect 1502 -942 1518 -940
rect 1552 -910 1568 -908
rect 2302 -908 2368 -898
rect 2302 -910 2318 -908
rect 1552 -940 1590 -910
rect 1708 -940 1762 -910
rect 1880 -940 1990 -910
rect 2108 -940 2162 -910
rect 2280 -940 2318 -910
rect 1552 -942 1568 -940
rect 1502 -952 1568 -942
rect 1502 -1008 1568 -998
rect 1502 -1010 1518 -1008
rect 752 -1040 790 -1010
rect 908 -1040 962 -1010
rect 1080 -1040 1190 -1010
rect 1308 -1040 1362 -1010
rect 1480 -1040 1518 -1010
rect 752 -1042 768 -1040
rect 702 -1052 768 -1042
rect 702 -1108 768 -1098
rect 702 -1110 718 -1108
rect -48 -1140 -10 -1110
rect 108 -1140 162 -1110
rect 280 -1140 390 -1110
rect 508 -1140 562 -1110
rect 680 -1140 718 -1110
rect -48 -1142 -32 -1140
rect -98 -1152 -32 -1142
rect -98 -1208 -32 -1198
rect -98 -1210 -82 -1208
rect -106 -1240 -82 -1210
rect -98 -1242 -82 -1240
rect -48 -1210 -32 -1208
rect 702 -1142 718 -1140
rect 752 -1110 768 -1108
rect 1502 -1042 1518 -1040
rect 1552 -1010 1568 -1008
rect 2302 -942 2318 -940
rect 2352 -910 2368 -908
rect 3102 -908 3168 -898
rect 3102 -910 3118 -908
rect 2352 -940 2390 -910
rect 2508 -940 2562 -910
rect 2680 -940 2790 -910
rect 2908 -940 2962 -910
rect 3080 -940 3118 -910
rect 2352 -942 2368 -940
rect 2302 -952 2368 -942
rect 2302 -1008 2368 -998
rect 2302 -1010 2318 -1008
rect 1552 -1040 1590 -1010
rect 1708 -1040 1762 -1010
rect 1880 -1040 1990 -1010
rect 2108 -1040 2162 -1010
rect 2280 -1040 2318 -1010
rect 1552 -1042 1568 -1040
rect 1502 -1052 1568 -1042
rect 1502 -1108 1568 -1098
rect 1502 -1110 1518 -1108
rect 752 -1140 790 -1110
rect 908 -1140 962 -1110
rect 1080 -1140 1190 -1110
rect 1308 -1140 1362 -1110
rect 1480 -1140 1518 -1110
rect 752 -1142 768 -1140
rect 702 -1152 768 -1142
rect 702 -1208 768 -1198
rect 702 -1210 718 -1208
rect -48 -1240 -10 -1210
rect 108 -1240 162 -1210
rect 280 -1240 390 -1210
rect 508 -1240 562 -1210
rect 680 -1240 718 -1210
rect -48 -1242 -32 -1240
rect -98 -1252 -32 -1242
rect -98 -1308 -32 -1298
rect -98 -1310 -82 -1308
rect -106 -1340 -82 -1310
rect -98 -1342 -82 -1340
rect -48 -1310 -32 -1308
rect 702 -1242 718 -1240
rect 752 -1210 768 -1208
rect 1502 -1142 1518 -1140
rect 1552 -1110 1568 -1108
rect 2302 -1042 2318 -1040
rect 2352 -1010 2368 -1008
rect 3102 -942 3118 -940
rect 3152 -910 3168 -908
rect 3902 -908 3968 -898
rect 3902 -910 3918 -908
rect 3152 -940 3190 -910
rect 3308 -940 3362 -910
rect 3480 -940 3590 -910
rect 3708 -940 3762 -910
rect 3880 -940 3918 -910
rect 3152 -942 3168 -940
rect 3102 -952 3168 -942
rect 3102 -1008 3168 -998
rect 3102 -1010 3118 -1008
rect 2352 -1040 2390 -1010
rect 2508 -1040 2562 -1010
rect 2680 -1040 2790 -1010
rect 2908 -1040 2962 -1010
rect 3080 -1040 3118 -1010
rect 2352 -1042 2368 -1040
rect 2302 -1052 2368 -1042
rect 2302 -1108 2368 -1098
rect 2302 -1110 2318 -1108
rect 1552 -1140 1590 -1110
rect 1708 -1140 1762 -1110
rect 1880 -1140 1990 -1110
rect 2108 -1140 2162 -1110
rect 2280 -1140 2318 -1110
rect 1552 -1142 1568 -1140
rect 1502 -1152 1568 -1142
rect 1502 -1208 1568 -1198
rect 1502 -1210 1518 -1208
rect 752 -1240 790 -1210
rect 908 -1240 962 -1210
rect 1080 -1240 1190 -1210
rect 1308 -1240 1362 -1210
rect 1480 -1240 1518 -1210
rect 752 -1242 768 -1240
rect 702 -1252 768 -1242
rect 702 -1308 768 -1298
rect 702 -1310 718 -1308
rect -48 -1340 -10 -1310
rect 108 -1340 162 -1310
rect 280 -1340 390 -1310
rect 508 -1340 562 -1310
rect 680 -1340 718 -1310
rect -48 -1342 -32 -1340
rect -98 -1352 -32 -1342
rect -98 -1408 -32 -1398
rect -98 -1410 -82 -1408
rect -106 -1440 -82 -1410
rect -98 -1442 -82 -1440
rect -48 -1410 -32 -1408
rect 702 -1342 718 -1340
rect 752 -1310 768 -1308
rect 1502 -1242 1518 -1240
rect 1552 -1210 1568 -1208
rect 2302 -1142 2318 -1140
rect 2352 -1110 2368 -1108
rect 3102 -1042 3118 -1040
rect 3152 -1010 3168 -1008
rect 3902 -942 3918 -940
rect 3952 -910 3968 -908
rect 4702 -908 4768 -898
rect 4702 -910 4718 -908
rect 3952 -940 3990 -910
rect 4108 -940 4162 -910
rect 4280 -940 4390 -910
rect 4508 -940 4562 -910
rect 4680 -940 4718 -910
rect 3952 -942 3968 -940
rect 3902 -952 3968 -942
rect 3902 -1008 3968 -998
rect 3902 -1010 3918 -1008
rect 3152 -1040 3190 -1010
rect 3308 -1040 3362 -1010
rect 3480 -1040 3590 -1010
rect 3708 -1040 3762 -1010
rect 3880 -1040 3918 -1010
rect 3152 -1042 3168 -1040
rect 3102 -1052 3168 -1042
rect 3102 -1108 3168 -1098
rect 3102 -1110 3118 -1108
rect 2352 -1140 2390 -1110
rect 2508 -1140 2562 -1110
rect 2680 -1140 2790 -1110
rect 2908 -1140 2962 -1110
rect 3080 -1140 3118 -1110
rect 2352 -1142 2368 -1140
rect 2302 -1152 2368 -1142
rect 2302 -1208 2368 -1198
rect 2302 -1210 2318 -1208
rect 1552 -1240 1590 -1210
rect 1708 -1240 1762 -1210
rect 1880 -1240 1990 -1210
rect 2108 -1240 2162 -1210
rect 2280 -1240 2318 -1210
rect 1552 -1242 1568 -1240
rect 1502 -1252 1568 -1242
rect 1502 -1308 1568 -1298
rect 1502 -1310 1518 -1308
rect 752 -1340 790 -1310
rect 908 -1340 962 -1310
rect 1080 -1340 1190 -1310
rect 1308 -1340 1362 -1310
rect 1480 -1340 1518 -1310
rect 752 -1342 768 -1340
rect 702 -1352 768 -1342
rect 702 -1408 768 -1398
rect 702 -1410 718 -1408
rect -48 -1440 -10 -1410
rect 108 -1440 162 -1410
rect 280 -1440 390 -1410
rect 508 -1440 562 -1410
rect 680 -1440 718 -1410
rect -48 -1442 -32 -1440
rect -98 -1452 -32 -1442
rect -98 -1508 -32 -1498
rect -98 -1510 -82 -1508
rect -106 -1540 -82 -1510
rect -98 -1542 -82 -1540
rect -48 -1510 -32 -1508
rect 702 -1442 718 -1440
rect 752 -1410 768 -1408
rect 1502 -1342 1518 -1340
rect 1552 -1310 1568 -1308
rect 2302 -1242 2318 -1240
rect 2352 -1210 2368 -1208
rect 3102 -1142 3118 -1140
rect 3152 -1110 3168 -1108
rect 3902 -1042 3918 -1040
rect 3952 -1010 3968 -1008
rect 4702 -942 4718 -940
rect 4752 -910 4768 -908
rect 5502 -908 5568 -898
rect 5502 -910 5518 -908
rect 4752 -940 4790 -910
rect 4908 -940 4962 -910
rect 5080 -940 5190 -910
rect 5308 -940 5362 -910
rect 5480 -940 5518 -910
rect 4752 -942 4768 -940
rect 4702 -952 4768 -942
rect 4702 -1008 4768 -998
rect 4702 -1010 4718 -1008
rect 3952 -1040 3990 -1010
rect 4108 -1040 4162 -1010
rect 4280 -1040 4390 -1010
rect 4508 -1040 4562 -1010
rect 4680 -1040 4718 -1010
rect 3952 -1042 3968 -1040
rect 3902 -1052 3968 -1042
rect 3902 -1108 3968 -1098
rect 3902 -1110 3918 -1108
rect 3152 -1140 3190 -1110
rect 3308 -1140 3362 -1110
rect 3480 -1140 3590 -1110
rect 3708 -1140 3762 -1110
rect 3880 -1140 3918 -1110
rect 3152 -1142 3168 -1140
rect 3102 -1152 3168 -1142
rect 3102 -1208 3168 -1198
rect 3102 -1210 3118 -1208
rect 2352 -1240 2390 -1210
rect 2508 -1240 2562 -1210
rect 2680 -1240 2790 -1210
rect 2908 -1240 2962 -1210
rect 3080 -1240 3118 -1210
rect 2352 -1242 2368 -1240
rect 2302 -1252 2368 -1242
rect 2302 -1308 2368 -1298
rect 2302 -1310 2318 -1308
rect 1552 -1340 1590 -1310
rect 1708 -1340 1762 -1310
rect 1880 -1340 1990 -1310
rect 2108 -1340 2162 -1310
rect 2280 -1340 2318 -1310
rect 1552 -1342 1568 -1340
rect 1502 -1352 1568 -1342
rect 1502 -1408 1568 -1398
rect 1502 -1410 1518 -1408
rect 752 -1440 790 -1410
rect 908 -1440 962 -1410
rect 1080 -1440 1190 -1410
rect 1308 -1440 1362 -1410
rect 1480 -1440 1518 -1410
rect 752 -1442 768 -1440
rect 702 -1452 768 -1442
rect 702 -1508 768 -1498
rect 702 -1510 718 -1508
rect -48 -1540 -10 -1510
rect 108 -1540 162 -1510
rect 280 -1540 390 -1510
rect 508 -1540 562 -1510
rect 680 -1540 718 -1510
rect -48 -1542 -32 -1540
rect -98 -1552 -32 -1542
rect -98 -1608 -32 -1598
rect -98 -1610 -82 -1608
rect -106 -1640 -82 -1610
rect -98 -1642 -82 -1640
rect -48 -1610 -32 -1608
rect 702 -1542 718 -1540
rect 752 -1510 768 -1508
rect 1502 -1442 1518 -1440
rect 1552 -1410 1568 -1408
rect 2302 -1342 2318 -1340
rect 2352 -1310 2368 -1308
rect 3102 -1242 3118 -1240
rect 3152 -1210 3168 -1208
rect 3902 -1142 3918 -1140
rect 3952 -1110 3968 -1108
rect 4702 -1042 4718 -1040
rect 4752 -1010 4768 -1008
rect 5502 -942 5518 -940
rect 5552 -910 5568 -908
rect 6302 -908 6368 -898
rect 6302 -910 6318 -908
rect 5552 -940 5590 -910
rect 5708 -940 5762 -910
rect 5880 -940 5990 -910
rect 6108 -940 6162 -910
rect 6280 -940 6318 -910
rect 5552 -942 5568 -940
rect 5502 -952 5568 -942
rect 5502 -1008 5568 -998
rect 5502 -1010 5518 -1008
rect 4752 -1040 4790 -1010
rect 4908 -1040 4962 -1010
rect 5080 -1040 5190 -1010
rect 5308 -1040 5362 -1010
rect 5480 -1040 5518 -1010
rect 4752 -1042 4768 -1040
rect 4702 -1052 4768 -1042
rect 4702 -1108 4768 -1098
rect 4702 -1110 4718 -1108
rect 3952 -1140 3990 -1110
rect 4108 -1140 4162 -1110
rect 4280 -1140 4390 -1110
rect 4508 -1140 4562 -1110
rect 4680 -1140 4718 -1110
rect 3952 -1142 3968 -1140
rect 3902 -1152 3968 -1142
rect 3902 -1208 3968 -1198
rect 3902 -1210 3918 -1208
rect 3152 -1240 3190 -1210
rect 3308 -1240 3362 -1210
rect 3480 -1240 3590 -1210
rect 3708 -1240 3762 -1210
rect 3880 -1240 3918 -1210
rect 3152 -1242 3168 -1240
rect 3102 -1252 3168 -1242
rect 3102 -1308 3168 -1298
rect 3102 -1310 3118 -1308
rect 2352 -1340 2390 -1310
rect 2508 -1340 2562 -1310
rect 2680 -1340 2790 -1310
rect 2908 -1340 2962 -1310
rect 3080 -1340 3118 -1310
rect 2352 -1342 2368 -1340
rect 2302 -1352 2368 -1342
rect 2302 -1408 2368 -1398
rect 2302 -1410 2318 -1408
rect 1552 -1440 1590 -1410
rect 1708 -1440 1762 -1410
rect 1880 -1440 1990 -1410
rect 2108 -1440 2162 -1410
rect 2280 -1440 2318 -1410
rect 1552 -1442 1568 -1440
rect 1502 -1452 1568 -1442
rect 1502 -1508 1568 -1498
rect 1502 -1510 1518 -1508
rect 752 -1540 790 -1510
rect 908 -1540 962 -1510
rect 1080 -1540 1190 -1510
rect 1308 -1540 1362 -1510
rect 1480 -1540 1518 -1510
rect 752 -1542 768 -1540
rect 702 -1552 768 -1542
rect 702 -1608 768 -1598
rect 702 -1610 718 -1608
rect -48 -1640 -10 -1610
rect 108 -1640 162 -1610
rect 280 -1640 390 -1610
rect 508 -1640 562 -1610
rect 680 -1640 718 -1610
rect -48 -1642 -32 -1640
rect -98 -1652 -32 -1642
rect -98 -1708 -32 -1698
rect -98 -1710 -82 -1708
rect -106 -1740 -82 -1710
rect -98 -1742 -82 -1740
rect -48 -1710 -32 -1708
rect 702 -1642 718 -1640
rect 752 -1610 768 -1608
rect 1502 -1542 1518 -1540
rect 1552 -1510 1568 -1508
rect 2302 -1442 2318 -1440
rect 2352 -1410 2368 -1408
rect 3102 -1342 3118 -1340
rect 3152 -1310 3168 -1308
rect 3902 -1242 3918 -1240
rect 3952 -1210 3968 -1208
rect 4702 -1142 4718 -1140
rect 4752 -1110 4768 -1108
rect 5502 -1042 5518 -1040
rect 5552 -1010 5568 -1008
rect 6302 -942 6318 -940
rect 6352 -910 6368 -908
rect 7102 -908 7168 -898
rect 7102 -910 7118 -908
rect 6352 -940 6390 -910
rect 6508 -940 6562 -910
rect 6680 -940 6790 -910
rect 6908 -940 6962 -910
rect 7080 -940 7118 -910
rect 6352 -942 6368 -940
rect 6302 -952 6368 -942
rect 6302 -1008 6368 -998
rect 6302 -1010 6318 -1008
rect 5552 -1040 5590 -1010
rect 5708 -1040 5762 -1010
rect 5880 -1040 5990 -1010
rect 6108 -1040 6162 -1010
rect 6280 -1040 6318 -1010
rect 5552 -1042 5568 -1040
rect 5502 -1052 5568 -1042
rect 5502 -1108 5568 -1098
rect 5502 -1110 5518 -1108
rect 4752 -1140 4790 -1110
rect 4908 -1140 4962 -1110
rect 5080 -1140 5190 -1110
rect 5308 -1140 5362 -1110
rect 5480 -1140 5518 -1110
rect 4752 -1142 4768 -1140
rect 4702 -1152 4768 -1142
rect 4702 -1208 4768 -1198
rect 4702 -1210 4718 -1208
rect 3952 -1240 3990 -1210
rect 4108 -1240 4162 -1210
rect 4280 -1240 4390 -1210
rect 4508 -1240 4562 -1210
rect 4680 -1240 4718 -1210
rect 3952 -1242 3968 -1240
rect 3902 -1252 3968 -1242
rect 3902 -1308 3968 -1298
rect 3902 -1310 3918 -1308
rect 3152 -1340 3190 -1310
rect 3308 -1340 3362 -1310
rect 3480 -1340 3590 -1310
rect 3708 -1340 3762 -1310
rect 3880 -1340 3918 -1310
rect 3152 -1342 3168 -1340
rect 3102 -1352 3168 -1342
rect 3102 -1408 3168 -1398
rect 3102 -1410 3118 -1408
rect 2352 -1440 2390 -1410
rect 2508 -1440 2562 -1410
rect 2680 -1440 2790 -1410
rect 2908 -1440 2962 -1410
rect 3080 -1440 3118 -1410
rect 2352 -1442 2368 -1440
rect 2302 -1452 2368 -1442
rect 2302 -1508 2368 -1498
rect 2302 -1510 2318 -1508
rect 1552 -1540 1590 -1510
rect 1708 -1540 1762 -1510
rect 1880 -1540 1990 -1510
rect 2108 -1540 2162 -1510
rect 2280 -1540 2318 -1510
rect 1552 -1542 1568 -1540
rect 1502 -1552 1568 -1542
rect 1502 -1608 1568 -1598
rect 1502 -1610 1518 -1608
rect 752 -1640 790 -1610
rect 908 -1640 962 -1610
rect 1080 -1640 1190 -1610
rect 1308 -1640 1362 -1610
rect 1480 -1640 1518 -1610
rect 752 -1642 768 -1640
rect 702 -1652 768 -1642
rect 702 -1708 768 -1698
rect 702 -1710 718 -1708
rect -48 -1740 -10 -1710
rect 108 -1740 162 -1710
rect 280 -1740 390 -1710
rect 508 -1740 562 -1710
rect 680 -1740 718 -1710
rect -48 -1742 -32 -1740
rect -98 -1752 -32 -1742
rect -98 -1808 -32 -1798
rect -98 -1810 -82 -1808
rect -106 -1840 -82 -1810
rect -98 -1842 -82 -1840
rect -48 -1810 -32 -1808
rect 702 -1742 718 -1740
rect 752 -1710 768 -1708
rect 1502 -1642 1518 -1640
rect 1552 -1610 1568 -1608
rect 2302 -1542 2318 -1540
rect 2352 -1510 2368 -1508
rect 3102 -1442 3118 -1440
rect 3152 -1410 3168 -1408
rect 3902 -1342 3918 -1340
rect 3952 -1310 3968 -1308
rect 4702 -1242 4718 -1240
rect 4752 -1210 4768 -1208
rect 5502 -1142 5518 -1140
rect 5552 -1110 5568 -1108
rect 6302 -1042 6318 -1040
rect 6352 -1010 6368 -1008
rect 7102 -942 7118 -940
rect 7152 -910 7168 -908
rect 7902 -908 7968 -898
rect 7902 -910 7918 -908
rect 7152 -940 7190 -910
rect 7308 -940 7362 -910
rect 7480 -940 7590 -910
rect 7708 -940 7762 -910
rect 7880 -940 7918 -910
rect 7152 -942 7168 -940
rect 7102 -952 7168 -942
rect 7102 -1008 7168 -998
rect 7102 -1010 7118 -1008
rect 6352 -1040 6390 -1010
rect 6508 -1040 6562 -1010
rect 6680 -1040 6790 -1010
rect 6908 -1040 6962 -1010
rect 7080 -1040 7118 -1010
rect 6352 -1042 6368 -1040
rect 6302 -1052 6368 -1042
rect 6302 -1108 6368 -1098
rect 6302 -1110 6318 -1108
rect 5552 -1140 5590 -1110
rect 5708 -1140 5762 -1110
rect 5880 -1140 5990 -1110
rect 6108 -1140 6162 -1110
rect 6280 -1140 6318 -1110
rect 5552 -1142 5568 -1140
rect 5502 -1152 5568 -1142
rect 5502 -1208 5568 -1198
rect 5502 -1210 5518 -1208
rect 4752 -1240 4790 -1210
rect 4908 -1240 4962 -1210
rect 5080 -1240 5190 -1210
rect 5308 -1240 5362 -1210
rect 5480 -1240 5518 -1210
rect 4752 -1242 4768 -1240
rect 4702 -1252 4768 -1242
rect 4702 -1308 4768 -1298
rect 4702 -1310 4718 -1308
rect 3952 -1340 3990 -1310
rect 4108 -1340 4162 -1310
rect 4280 -1340 4390 -1310
rect 4508 -1340 4562 -1310
rect 4680 -1340 4718 -1310
rect 3952 -1342 3968 -1340
rect 3902 -1352 3968 -1342
rect 3902 -1408 3968 -1398
rect 3902 -1410 3918 -1408
rect 3152 -1440 3190 -1410
rect 3308 -1440 3362 -1410
rect 3480 -1440 3590 -1410
rect 3708 -1440 3762 -1410
rect 3880 -1440 3918 -1410
rect 3152 -1442 3168 -1440
rect 3102 -1452 3168 -1442
rect 3102 -1508 3168 -1498
rect 3102 -1510 3118 -1508
rect 2352 -1540 2390 -1510
rect 2508 -1540 2562 -1510
rect 2680 -1540 2790 -1510
rect 2908 -1540 2962 -1510
rect 3080 -1540 3118 -1510
rect 2352 -1542 2368 -1540
rect 2302 -1552 2368 -1542
rect 2302 -1608 2368 -1598
rect 2302 -1610 2318 -1608
rect 1552 -1640 1590 -1610
rect 1708 -1640 1762 -1610
rect 1880 -1640 1990 -1610
rect 2108 -1640 2162 -1610
rect 2280 -1640 2318 -1610
rect 1552 -1642 1568 -1640
rect 1502 -1652 1568 -1642
rect 1502 -1708 1568 -1698
rect 1502 -1710 1518 -1708
rect 752 -1740 790 -1710
rect 908 -1740 962 -1710
rect 1080 -1740 1190 -1710
rect 1308 -1740 1362 -1710
rect 1480 -1740 1518 -1710
rect 752 -1742 768 -1740
rect 702 -1752 768 -1742
rect 702 -1808 768 -1798
rect 702 -1810 718 -1808
rect -48 -1840 -10 -1810
rect 108 -1840 162 -1810
rect 280 -1840 390 -1810
rect 508 -1840 562 -1810
rect 680 -1840 718 -1810
rect -48 -1842 -32 -1840
rect -98 -1852 -32 -1842
rect -98 -1908 -32 -1898
rect -98 -1910 -82 -1908
rect -106 -1940 -82 -1910
rect -98 -1942 -82 -1940
rect -48 -1910 -32 -1908
rect 702 -1842 718 -1840
rect 752 -1810 768 -1808
rect 1502 -1742 1518 -1740
rect 1552 -1710 1568 -1708
rect 2302 -1642 2318 -1640
rect 2352 -1610 2368 -1608
rect 3102 -1542 3118 -1540
rect 3152 -1510 3168 -1508
rect 3902 -1442 3918 -1440
rect 3952 -1410 3968 -1408
rect 4702 -1342 4718 -1340
rect 4752 -1310 4768 -1308
rect 5502 -1242 5518 -1240
rect 5552 -1210 5568 -1208
rect 6302 -1142 6318 -1140
rect 6352 -1110 6368 -1108
rect 7102 -1042 7118 -1040
rect 7152 -1010 7168 -1008
rect 7902 -942 7918 -940
rect 7952 -910 7968 -908
rect 8702 -908 8768 -898
rect 8702 -910 8718 -908
rect 7952 -940 7990 -910
rect 8108 -940 8162 -910
rect 8280 -940 8390 -910
rect 8508 -940 8562 -910
rect 8680 -940 8718 -910
rect 7952 -942 7968 -940
rect 7902 -952 7968 -942
rect 7902 -1008 7968 -998
rect 7902 -1010 7918 -1008
rect 7152 -1040 7190 -1010
rect 7308 -1040 7362 -1010
rect 7480 -1040 7590 -1010
rect 7708 -1040 7762 -1010
rect 7880 -1040 7918 -1010
rect 7152 -1042 7168 -1040
rect 7102 -1052 7168 -1042
rect 7102 -1108 7168 -1098
rect 7102 -1110 7118 -1108
rect 6352 -1140 6390 -1110
rect 6508 -1140 6562 -1110
rect 6680 -1140 6790 -1110
rect 6908 -1140 6962 -1110
rect 7080 -1140 7118 -1110
rect 6352 -1142 6368 -1140
rect 6302 -1152 6368 -1142
rect 6302 -1208 6368 -1198
rect 6302 -1210 6318 -1208
rect 5552 -1240 5590 -1210
rect 5708 -1240 5762 -1210
rect 5880 -1240 5990 -1210
rect 6108 -1240 6162 -1210
rect 6280 -1240 6318 -1210
rect 5552 -1242 5568 -1240
rect 5502 -1252 5568 -1242
rect 5502 -1308 5568 -1298
rect 5502 -1310 5518 -1308
rect 4752 -1340 4790 -1310
rect 4908 -1340 4962 -1310
rect 5080 -1340 5190 -1310
rect 5308 -1340 5362 -1310
rect 5480 -1340 5518 -1310
rect 4752 -1342 4768 -1340
rect 4702 -1352 4768 -1342
rect 4702 -1408 4768 -1398
rect 4702 -1410 4718 -1408
rect 3952 -1440 3990 -1410
rect 4108 -1440 4162 -1410
rect 4280 -1440 4390 -1410
rect 4508 -1440 4562 -1410
rect 4680 -1440 4718 -1410
rect 3952 -1442 3968 -1440
rect 3902 -1452 3968 -1442
rect 3902 -1508 3968 -1498
rect 3902 -1510 3918 -1508
rect 3152 -1540 3190 -1510
rect 3308 -1540 3362 -1510
rect 3480 -1540 3590 -1510
rect 3708 -1540 3762 -1510
rect 3880 -1540 3918 -1510
rect 3152 -1542 3168 -1540
rect 3102 -1552 3168 -1542
rect 3102 -1608 3168 -1598
rect 3102 -1610 3118 -1608
rect 2352 -1640 2390 -1610
rect 2508 -1640 2562 -1610
rect 2680 -1640 2790 -1610
rect 2908 -1640 2962 -1610
rect 3080 -1640 3118 -1610
rect 2352 -1642 2368 -1640
rect 2302 -1652 2368 -1642
rect 2302 -1708 2368 -1698
rect 2302 -1710 2318 -1708
rect 1552 -1740 1590 -1710
rect 1708 -1740 1762 -1710
rect 1880 -1740 1990 -1710
rect 2108 -1740 2162 -1710
rect 2280 -1740 2318 -1710
rect 1552 -1742 1568 -1740
rect 1502 -1752 1568 -1742
rect 1502 -1808 1568 -1798
rect 1502 -1810 1518 -1808
rect 752 -1840 790 -1810
rect 908 -1840 962 -1810
rect 1080 -1840 1190 -1810
rect 1308 -1840 1362 -1810
rect 1480 -1840 1518 -1810
rect 752 -1842 768 -1840
rect 702 -1852 768 -1842
rect 702 -1908 768 -1898
rect 702 -1910 718 -1908
rect -48 -1940 -10 -1910
rect 108 -1940 162 -1910
rect 280 -1940 390 -1910
rect 508 -1940 562 -1910
rect 680 -1940 718 -1910
rect -48 -1942 -32 -1940
rect -98 -1952 -32 -1942
rect -98 -2008 -32 -1998
rect -98 -2010 -82 -2008
rect -106 -2040 -82 -2010
rect -98 -2042 -82 -2040
rect -48 -2010 -32 -2008
rect 702 -1942 718 -1940
rect 752 -1910 768 -1908
rect 1502 -1842 1518 -1840
rect 1552 -1810 1568 -1808
rect 2302 -1742 2318 -1740
rect 2352 -1710 2368 -1708
rect 3102 -1642 3118 -1640
rect 3152 -1610 3168 -1608
rect 3902 -1542 3918 -1540
rect 3952 -1510 3968 -1508
rect 4702 -1442 4718 -1440
rect 4752 -1410 4768 -1408
rect 5502 -1342 5518 -1340
rect 5552 -1310 5568 -1308
rect 6302 -1242 6318 -1240
rect 6352 -1210 6368 -1208
rect 7102 -1142 7118 -1140
rect 7152 -1110 7168 -1108
rect 7902 -1042 7918 -1040
rect 7952 -1010 7968 -1008
rect 8702 -942 8718 -940
rect 8752 -910 8768 -908
rect 9502 -908 9568 -898
rect 9502 -910 9518 -908
rect 8752 -940 8790 -910
rect 8908 -940 8962 -910
rect 9080 -940 9190 -910
rect 9308 -940 9362 -910
rect 9480 -940 9518 -910
rect 8752 -942 8768 -940
rect 8702 -952 8768 -942
rect 8702 -1008 8768 -998
rect 8702 -1010 8718 -1008
rect 7952 -1040 7990 -1010
rect 8108 -1040 8162 -1010
rect 8280 -1040 8390 -1010
rect 8508 -1040 8562 -1010
rect 8680 -1040 8718 -1010
rect 7952 -1042 7968 -1040
rect 7902 -1052 7968 -1042
rect 7902 -1108 7968 -1098
rect 7902 -1110 7918 -1108
rect 7152 -1140 7190 -1110
rect 7308 -1140 7362 -1110
rect 7480 -1140 7590 -1110
rect 7708 -1140 7762 -1110
rect 7880 -1140 7918 -1110
rect 7152 -1142 7168 -1140
rect 7102 -1152 7168 -1142
rect 7102 -1208 7168 -1198
rect 7102 -1210 7118 -1208
rect 6352 -1240 6390 -1210
rect 6508 -1240 6562 -1210
rect 6680 -1240 6790 -1210
rect 6908 -1240 6962 -1210
rect 7080 -1240 7118 -1210
rect 6352 -1242 6368 -1240
rect 6302 -1252 6368 -1242
rect 6302 -1308 6368 -1298
rect 6302 -1310 6318 -1308
rect 5552 -1340 5590 -1310
rect 5708 -1340 5762 -1310
rect 5880 -1340 5990 -1310
rect 6108 -1340 6162 -1310
rect 6280 -1340 6318 -1310
rect 5552 -1342 5568 -1340
rect 5502 -1352 5568 -1342
rect 5502 -1408 5568 -1398
rect 5502 -1410 5518 -1408
rect 4752 -1440 4790 -1410
rect 4908 -1440 4962 -1410
rect 5080 -1440 5190 -1410
rect 5308 -1440 5362 -1410
rect 5480 -1440 5518 -1410
rect 4752 -1442 4768 -1440
rect 4702 -1452 4768 -1442
rect 4702 -1508 4768 -1498
rect 4702 -1510 4718 -1508
rect 3952 -1540 3990 -1510
rect 4108 -1540 4162 -1510
rect 4280 -1540 4390 -1510
rect 4508 -1540 4562 -1510
rect 4680 -1540 4718 -1510
rect 3952 -1542 3968 -1540
rect 3902 -1552 3968 -1542
rect 3902 -1608 3968 -1598
rect 3902 -1610 3918 -1608
rect 3152 -1640 3190 -1610
rect 3308 -1640 3362 -1610
rect 3480 -1640 3590 -1610
rect 3708 -1640 3762 -1610
rect 3880 -1640 3918 -1610
rect 3152 -1642 3168 -1640
rect 3102 -1652 3168 -1642
rect 3102 -1708 3168 -1698
rect 3102 -1710 3118 -1708
rect 2352 -1740 2390 -1710
rect 2508 -1740 2562 -1710
rect 2680 -1740 2790 -1710
rect 2908 -1740 2962 -1710
rect 3080 -1740 3118 -1710
rect 2352 -1742 2368 -1740
rect 2302 -1752 2368 -1742
rect 2302 -1808 2368 -1798
rect 2302 -1810 2318 -1808
rect 1552 -1840 1590 -1810
rect 1708 -1840 1762 -1810
rect 1880 -1840 1990 -1810
rect 2108 -1840 2162 -1810
rect 2280 -1840 2318 -1810
rect 1552 -1842 1568 -1840
rect 1502 -1852 1568 -1842
rect 1502 -1908 1568 -1898
rect 1502 -1910 1518 -1908
rect 752 -1940 790 -1910
rect 908 -1940 962 -1910
rect 1080 -1940 1190 -1910
rect 1308 -1940 1362 -1910
rect 1480 -1940 1518 -1910
rect 752 -1942 768 -1940
rect 702 -1952 768 -1942
rect 702 -2008 768 -1998
rect 702 -2010 718 -2008
rect -48 -2040 -10 -2010
rect 108 -2040 162 -2010
rect 280 -2040 390 -2010
rect 508 -2040 562 -2010
rect 680 -2040 718 -2010
rect -48 -2042 -32 -2040
rect -98 -2052 -32 -2042
rect 702 -2042 718 -2040
rect 752 -2010 768 -2008
rect 1502 -1942 1518 -1940
rect 1552 -1910 1568 -1908
rect 2302 -1842 2318 -1840
rect 2352 -1810 2368 -1808
rect 3102 -1742 3118 -1740
rect 3152 -1710 3168 -1708
rect 3902 -1642 3918 -1640
rect 3952 -1610 3968 -1608
rect 4702 -1542 4718 -1540
rect 4752 -1510 4768 -1508
rect 5502 -1442 5518 -1440
rect 5552 -1410 5568 -1408
rect 6302 -1342 6318 -1340
rect 6352 -1310 6368 -1308
rect 7102 -1242 7118 -1240
rect 7152 -1210 7168 -1208
rect 7902 -1142 7918 -1140
rect 7952 -1110 7968 -1108
rect 8702 -1042 8718 -1040
rect 8752 -1010 8768 -1008
rect 9502 -942 9518 -940
rect 9552 -910 9568 -908
rect 10302 -908 10368 -898
rect 10302 -910 10318 -908
rect 9552 -940 9590 -910
rect 9708 -940 9762 -910
rect 9880 -940 9990 -910
rect 10108 -940 10162 -910
rect 10280 -940 10318 -910
rect 9552 -942 9568 -940
rect 9502 -952 9568 -942
rect 9502 -1008 9568 -998
rect 9502 -1010 9518 -1008
rect 8752 -1040 8790 -1010
rect 8908 -1040 8962 -1010
rect 9080 -1040 9190 -1010
rect 9308 -1040 9362 -1010
rect 9480 -1040 9518 -1010
rect 8752 -1042 8768 -1040
rect 8702 -1052 8768 -1042
rect 8702 -1108 8768 -1098
rect 8702 -1110 8718 -1108
rect 7952 -1140 7990 -1110
rect 8108 -1140 8162 -1110
rect 8280 -1140 8390 -1110
rect 8508 -1140 8562 -1110
rect 8680 -1140 8718 -1110
rect 7952 -1142 7968 -1140
rect 7902 -1152 7968 -1142
rect 7902 -1208 7968 -1198
rect 7902 -1210 7918 -1208
rect 7152 -1240 7190 -1210
rect 7308 -1240 7362 -1210
rect 7480 -1240 7590 -1210
rect 7708 -1240 7762 -1210
rect 7880 -1240 7918 -1210
rect 7152 -1242 7168 -1240
rect 7102 -1252 7168 -1242
rect 7102 -1308 7168 -1298
rect 7102 -1310 7118 -1308
rect 6352 -1340 6390 -1310
rect 6508 -1340 6562 -1310
rect 6680 -1340 6790 -1310
rect 6908 -1340 6962 -1310
rect 7080 -1340 7118 -1310
rect 6352 -1342 6368 -1340
rect 6302 -1352 6368 -1342
rect 6302 -1408 6368 -1398
rect 6302 -1410 6318 -1408
rect 5552 -1440 5590 -1410
rect 5708 -1440 5762 -1410
rect 5880 -1440 5990 -1410
rect 6108 -1440 6162 -1410
rect 6280 -1440 6318 -1410
rect 5552 -1442 5568 -1440
rect 5502 -1452 5568 -1442
rect 5502 -1508 5568 -1498
rect 5502 -1510 5518 -1508
rect 4752 -1540 4790 -1510
rect 4908 -1540 4962 -1510
rect 5080 -1540 5190 -1510
rect 5308 -1540 5362 -1510
rect 5480 -1540 5518 -1510
rect 4752 -1542 4768 -1540
rect 4702 -1552 4768 -1542
rect 4702 -1608 4768 -1598
rect 4702 -1610 4718 -1608
rect 3952 -1640 3990 -1610
rect 4108 -1640 4162 -1610
rect 4280 -1640 4390 -1610
rect 4508 -1640 4562 -1610
rect 4680 -1640 4718 -1610
rect 3952 -1642 3968 -1640
rect 3902 -1652 3968 -1642
rect 3902 -1708 3968 -1698
rect 3902 -1710 3918 -1708
rect 3152 -1740 3190 -1710
rect 3308 -1740 3362 -1710
rect 3480 -1740 3590 -1710
rect 3708 -1740 3762 -1710
rect 3880 -1740 3918 -1710
rect 3152 -1742 3168 -1740
rect 3102 -1752 3168 -1742
rect 3102 -1808 3168 -1798
rect 3102 -1810 3118 -1808
rect 2352 -1840 2390 -1810
rect 2508 -1840 2562 -1810
rect 2680 -1840 2790 -1810
rect 2908 -1840 2962 -1810
rect 3080 -1840 3118 -1810
rect 2352 -1842 2368 -1840
rect 2302 -1852 2368 -1842
rect 2302 -1908 2368 -1898
rect 2302 -1910 2318 -1908
rect 1552 -1940 1590 -1910
rect 1708 -1940 1762 -1910
rect 1880 -1940 1990 -1910
rect 2108 -1940 2162 -1910
rect 2280 -1940 2318 -1910
rect 1552 -1942 1568 -1940
rect 1502 -1952 1568 -1942
rect 1502 -2008 1568 -1998
rect 1502 -2010 1518 -2008
rect 752 -2040 790 -2010
rect 908 -2040 962 -2010
rect 1080 -2040 1190 -2010
rect 1308 -2040 1362 -2010
rect 1480 -2040 1518 -2010
rect 752 -2042 768 -2040
rect 702 -2052 768 -2042
rect 1502 -2042 1518 -2040
rect 1552 -2010 1568 -2008
rect 2302 -1942 2318 -1940
rect 2352 -1910 2368 -1908
rect 3102 -1842 3118 -1840
rect 3152 -1810 3168 -1808
rect 3902 -1742 3918 -1740
rect 3952 -1710 3968 -1708
rect 4702 -1642 4718 -1640
rect 4752 -1610 4768 -1608
rect 5502 -1542 5518 -1540
rect 5552 -1510 5568 -1508
rect 6302 -1442 6318 -1440
rect 6352 -1410 6368 -1408
rect 7102 -1342 7118 -1340
rect 7152 -1310 7168 -1308
rect 7902 -1242 7918 -1240
rect 7952 -1210 7968 -1208
rect 8702 -1142 8718 -1140
rect 8752 -1110 8768 -1108
rect 9502 -1042 9518 -1040
rect 9552 -1010 9568 -1008
rect 10302 -942 10318 -940
rect 10352 -910 10368 -908
rect 11102 -908 11168 -898
rect 11102 -910 11118 -908
rect 10352 -940 10390 -910
rect 10508 -940 10562 -910
rect 10680 -940 10790 -910
rect 10908 -940 10962 -910
rect 11080 -940 11118 -910
rect 10352 -942 10368 -940
rect 10302 -952 10368 -942
rect 10302 -1008 10368 -998
rect 10302 -1010 10318 -1008
rect 9552 -1040 9590 -1010
rect 9708 -1040 9762 -1010
rect 9880 -1040 9990 -1010
rect 10108 -1040 10162 -1010
rect 10280 -1040 10318 -1010
rect 9552 -1042 9568 -1040
rect 9502 -1052 9568 -1042
rect 9502 -1108 9568 -1098
rect 9502 -1110 9518 -1108
rect 8752 -1140 8790 -1110
rect 8908 -1140 8962 -1110
rect 9080 -1140 9190 -1110
rect 9308 -1140 9362 -1110
rect 9480 -1140 9518 -1110
rect 8752 -1142 8768 -1140
rect 8702 -1152 8768 -1142
rect 8702 -1208 8768 -1198
rect 8702 -1210 8718 -1208
rect 7952 -1240 7990 -1210
rect 8108 -1240 8162 -1210
rect 8280 -1240 8390 -1210
rect 8508 -1240 8562 -1210
rect 8680 -1240 8718 -1210
rect 7952 -1242 7968 -1240
rect 7902 -1252 7968 -1242
rect 7902 -1308 7968 -1298
rect 7902 -1310 7918 -1308
rect 7152 -1340 7190 -1310
rect 7308 -1340 7362 -1310
rect 7480 -1340 7590 -1310
rect 7708 -1340 7762 -1310
rect 7880 -1340 7918 -1310
rect 7152 -1342 7168 -1340
rect 7102 -1352 7168 -1342
rect 7102 -1408 7168 -1398
rect 7102 -1410 7118 -1408
rect 6352 -1440 6390 -1410
rect 6508 -1440 6562 -1410
rect 6680 -1440 6790 -1410
rect 6908 -1440 6962 -1410
rect 7080 -1440 7118 -1410
rect 6352 -1442 6368 -1440
rect 6302 -1452 6368 -1442
rect 6302 -1508 6368 -1498
rect 6302 -1510 6318 -1508
rect 5552 -1540 5590 -1510
rect 5708 -1540 5762 -1510
rect 5880 -1540 5990 -1510
rect 6108 -1540 6162 -1510
rect 6280 -1540 6318 -1510
rect 5552 -1542 5568 -1540
rect 5502 -1552 5568 -1542
rect 5502 -1608 5568 -1598
rect 5502 -1610 5518 -1608
rect 4752 -1640 4790 -1610
rect 4908 -1640 4962 -1610
rect 5080 -1640 5190 -1610
rect 5308 -1640 5362 -1610
rect 5480 -1640 5518 -1610
rect 4752 -1642 4768 -1640
rect 4702 -1652 4768 -1642
rect 4702 -1708 4768 -1698
rect 4702 -1710 4718 -1708
rect 3952 -1740 3990 -1710
rect 4108 -1740 4162 -1710
rect 4280 -1740 4390 -1710
rect 4508 -1740 4562 -1710
rect 4680 -1740 4718 -1710
rect 3952 -1742 3968 -1740
rect 3902 -1752 3968 -1742
rect 3902 -1808 3968 -1798
rect 3902 -1810 3918 -1808
rect 3152 -1840 3190 -1810
rect 3308 -1840 3362 -1810
rect 3480 -1840 3590 -1810
rect 3708 -1840 3762 -1810
rect 3880 -1840 3918 -1810
rect 3152 -1842 3168 -1840
rect 3102 -1852 3168 -1842
rect 3102 -1908 3168 -1898
rect 3102 -1910 3118 -1908
rect 2352 -1940 2390 -1910
rect 2508 -1940 2562 -1910
rect 2680 -1940 2790 -1910
rect 2908 -1940 2962 -1910
rect 3080 -1940 3118 -1910
rect 2352 -1942 2368 -1940
rect 2302 -1952 2368 -1942
rect 2302 -2008 2368 -1998
rect 2302 -2010 2318 -2008
rect 1552 -2040 1590 -2010
rect 1708 -2040 1762 -2010
rect 1880 -2040 1990 -2010
rect 2108 -2040 2162 -2010
rect 2280 -2040 2318 -2010
rect 1552 -2042 1568 -2040
rect 1502 -2052 1568 -2042
rect 2302 -2042 2318 -2040
rect 2352 -2010 2368 -2008
rect 3102 -1942 3118 -1940
rect 3152 -1910 3168 -1908
rect 3902 -1842 3918 -1840
rect 3952 -1810 3968 -1808
rect 4702 -1742 4718 -1740
rect 4752 -1710 4768 -1708
rect 5502 -1642 5518 -1640
rect 5552 -1610 5568 -1608
rect 6302 -1542 6318 -1540
rect 6352 -1510 6368 -1508
rect 7102 -1442 7118 -1440
rect 7152 -1410 7168 -1408
rect 7902 -1342 7918 -1340
rect 7952 -1310 7968 -1308
rect 8702 -1242 8718 -1240
rect 8752 -1210 8768 -1208
rect 9502 -1142 9518 -1140
rect 9552 -1110 9568 -1108
rect 10302 -1042 10318 -1040
rect 10352 -1010 10368 -1008
rect 11102 -942 11118 -940
rect 11152 -910 11168 -908
rect 11902 -908 11968 -898
rect 11902 -910 11918 -908
rect 11152 -940 11190 -910
rect 11308 -940 11362 -910
rect 11480 -940 11590 -910
rect 11708 -940 11762 -910
rect 11880 -940 11918 -910
rect 11152 -942 11168 -940
rect 11102 -952 11168 -942
rect 11102 -1008 11168 -998
rect 11102 -1010 11118 -1008
rect 10352 -1040 10390 -1010
rect 10508 -1040 10562 -1010
rect 10680 -1040 10790 -1010
rect 10908 -1040 10962 -1010
rect 11080 -1040 11118 -1010
rect 10352 -1042 10368 -1040
rect 10302 -1052 10368 -1042
rect 10302 -1108 10368 -1098
rect 10302 -1110 10318 -1108
rect 9552 -1140 9590 -1110
rect 9708 -1140 9762 -1110
rect 9880 -1140 9990 -1110
rect 10108 -1140 10162 -1110
rect 10280 -1140 10318 -1110
rect 9552 -1142 9568 -1140
rect 9502 -1152 9568 -1142
rect 9502 -1208 9568 -1198
rect 9502 -1210 9518 -1208
rect 8752 -1240 8790 -1210
rect 8908 -1240 8962 -1210
rect 9080 -1240 9190 -1210
rect 9308 -1240 9362 -1210
rect 9480 -1240 9518 -1210
rect 8752 -1242 8768 -1240
rect 8702 -1252 8768 -1242
rect 8702 -1308 8768 -1298
rect 8702 -1310 8718 -1308
rect 7952 -1340 7990 -1310
rect 8108 -1340 8162 -1310
rect 8280 -1340 8390 -1310
rect 8508 -1340 8562 -1310
rect 8680 -1340 8718 -1310
rect 7952 -1342 7968 -1340
rect 7902 -1352 7968 -1342
rect 7902 -1408 7968 -1398
rect 7902 -1410 7918 -1408
rect 7152 -1440 7190 -1410
rect 7308 -1440 7362 -1410
rect 7480 -1440 7590 -1410
rect 7708 -1440 7762 -1410
rect 7880 -1440 7918 -1410
rect 7152 -1442 7168 -1440
rect 7102 -1452 7168 -1442
rect 7102 -1508 7168 -1498
rect 7102 -1510 7118 -1508
rect 6352 -1540 6390 -1510
rect 6508 -1540 6562 -1510
rect 6680 -1540 6790 -1510
rect 6908 -1540 6962 -1510
rect 7080 -1540 7118 -1510
rect 6352 -1542 6368 -1540
rect 6302 -1552 6368 -1542
rect 6302 -1608 6368 -1598
rect 6302 -1610 6318 -1608
rect 5552 -1640 5590 -1610
rect 5708 -1640 5762 -1610
rect 5880 -1640 5990 -1610
rect 6108 -1640 6162 -1610
rect 6280 -1640 6318 -1610
rect 5552 -1642 5568 -1640
rect 5502 -1652 5568 -1642
rect 5502 -1708 5568 -1698
rect 5502 -1710 5518 -1708
rect 4752 -1740 4790 -1710
rect 4908 -1740 4962 -1710
rect 5080 -1740 5190 -1710
rect 5308 -1740 5362 -1710
rect 5480 -1740 5518 -1710
rect 4752 -1742 4768 -1740
rect 4702 -1752 4768 -1742
rect 4702 -1808 4768 -1798
rect 4702 -1810 4718 -1808
rect 3952 -1840 3990 -1810
rect 4108 -1840 4162 -1810
rect 4280 -1840 4390 -1810
rect 4508 -1840 4562 -1810
rect 4680 -1840 4718 -1810
rect 3952 -1842 3968 -1840
rect 3902 -1852 3968 -1842
rect 3902 -1908 3968 -1898
rect 3902 -1910 3918 -1908
rect 3152 -1940 3190 -1910
rect 3308 -1940 3362 -1910
rect 3480 -1940 3590 -1910
rect 3708 -1940 3762 -1910
rect 3880 -1940 3918 -1910
rect 3152 -1942 3168 -1940
rect 3102 -1952 3168 -1942
rect 3102 -2008 3168 -1998
rect 3102 -2010 3118 -2008
rect 2352 -2040 2390 -2010
rect 2508 -2040 2562 -2010
rect 2680 -2040 2790 -2010
rect 2908 -2040 2962 -2010
rect 3080 -2040 3118 -2010
rect 2352 -2042 2368 -2040
rect 2302 -2052 2368 -2042
rect 3102 -2042 3118 -2040
rect 3152 -2010 3168 -2008
rect 3902 -1942 3918 -1940
rect 3952 -1910 3968 -1908
rect 4702 -1842 4718 -1840
rect 4752 -1810 4768 -1808
rect 5502 -1742 5518 -1740
rect 5552 -1710 5568 -1708
rect 6302 -1642 6318 -1640
rect 6352 -1610 6368 -1608
rect 7102 -1542 7118 -1540
rect 7152 -1510 7168 -1508
rect 7902 -1442 7918 -1440
rect 7952 -1410 7968 -1408
rect 8702 -1342 8718 -1340
rect 8752 -1310 8768 -1308
rect 9502 -1242 9518 -1240
rect 9552 -1210 9568 -1208
rect 10302 -1142 10318 -1140
rect 10352 -1110 10368 -1108
rect 11102 -1042 11118 -1040
rect 11152 -1010 11168 -1008
rect 11902 -942 11918 -940
rect 11952 -910 11968 -908
rect 14514 -890 14540 -860
rect 14690 -890 14816 -860
rect 15116 -890 15142 -860
rect 15200 -890 15226 -860
rect 15526 -890 15652 -860
rect 15802 -890 15828 -860
rect 12702 -908 12768 -898
rect 12702 -910 12718 -908
rect 11952 -940 11990 -910
rect 12108 -940 12162 -910
rect 12280 -940 12390 -910
rect 12508 -940 12562 -910
rect 12680 -940 12718 -910
rect 11952 -942 11968 -940
rect 11902 -952 11968 -942
rect 11902 -1008 11968 -998
rect 11902 -1010 11918 -1008
rect 11152 -1040 11190 -1010
rect 11308 -1040 11362 -1010
rect 11480 -1040 11590 -1010
rect 11708 -1040 11762 -1010
rect 11880 -1040 11918 -1010
rect 11152 -1042 11168 -1040
rect 11102 -1052 11168 -1042
rect 11102 -1108 11168 -1098
rect 11102 -1110 11118 -1108
rect 10352 -1140 10390 -1110
rect 10508 -1140 10562 -1110
rect 10680 -1140 10790 -1110
rect 10908 -1140 10962 -1110
rect 11080 -1140 11118 -1110
rect 10352 -1142 10368 -1140
rect 10302 -1152 10368 -1142
rect 10302 -1208 10368 -1198
rect 10302 -1210 10318 -1208
rect 9552 -1240 9590 -1210
rect 9708 -1240 9762 -1210
rect 9880 -1240 9990 -1210
rect 10108 -1240 10162 -1210
rect 10280 -1240 10318 -1210
rect 9552 -1242 9568 -1240
rect 9502 -1252 9568 -1242
rect 9502 -1308 9568 -1298
rect 9502 -1310 9518 -1308
rect 8752 -1340 8790 -1310
rect 8908 -1340 8962 -1310
rect 9080 -1340 9190 -1310
rect 9308 -1340 9362 -1310
rect 9480 -1340 9518 -1310
rect 8752 -1342 8768 -1340
rect 8702 -1352 8768 -1342
rect 8702 -1408 8768 -1398
rect 8702 -1410 8718 -1408
rect 7952 -1440 7990 -1410
rect 8108 -1440 8162 -1410
rect 8280 -1440 8390 -1410
rect 8508 -1440 8562 -1410
rect 8680 -1440 8718 -1410
rect 7952 -1442 7968 -1440
rect 7902 -1452 7968 -1442
rect 7902 -1508 7968 -1498
rect 7902 -1510 7918 -1508
rect 7152 -1540 7190 -1510
rect 7308 -1540 7362 -1510
rect 7480 -1540 7590 -1510
rect 7708 -1540 7762 -1510
rect 7880 -1540 7918 -1510
rect 7152 -1542 7168 -1540
rect 7102 -1552 7168 -1542
rect 7102 -1608 7168 -1598
rect 7102 -1610 7118 -1608
rect 6352 -1640 6390 -1610
rect 6508 -1640 6562 -1610
rect 6680 -1640 6790 -1610
rect 6908 -1640 6962 -1610
rect 7080 -1640 7118 -1610
rect 6352 -1642 6368 -1640
rect 6302 -1652 6368 -1642
rect 6302 -1708 6368 -1698
rect 6302 -1710 6318 -1708
rect 5552 -1740 5590 -1710
rect 5708 -1740 5762 -1710
rect 5880 -1740 5990 -1710
rect 6108 -1740 6162 -1710
rect 6280 -1740 6318 -1710
rect 5552 -1742 5568 -1740
rect 5502 -1752 5568 -1742
rect 5502 -1808 5568 -1798
rect 5502 -1810 5518 -1808
rect 4752 -1840 4790 -1810
rect 4908 -1840 4962 -1810
rect 5080 -1840 5190 -1810
rect 5308 -1840 5362 -1810
rect 5480 -1840 5518 -1810
rect 4752 -1842 4768 -1840
rect 4702 -1852 4768 -1842
rect 4702 -1908 4768 -1898
rect 4702 -1910 4718 -1908
rect 3952 -1940 3990 -1910
rect 4108 -1940 4162 -1910
rect 4280 -1940 4390 -1910
rect 4508 -1940 4562 -1910
rect 4680 -1940 4718 -1910
rect 3952 -1942 3968 -1940
rect 3902 -1952 3968 -1942
rect 3902 -2008 3968 -1998
rect 3902 -2010 3918 -2008
rect 3152 -2040 3190 -2010
rect 3308 -2040 3362 -2010
rect 3480 -2040 3590 -2010
rect 3708 -2040 3762 -2010
rect 3880 -2040 3918 -2010
rect 3152 -2042 3168 -2040
rect 3102 -2052 3168 -2042
rect 3902 -2042 3918 -2040
rect 3952 -2010 3968 -2008
rect 4702 -1942 4718 -1940
rect 4752 -1910 4768 -1908
rect 5502 -1842 5518 -1840
rect 5552 -1810 5568 -1808
rect 6302 -1742 6318 -1740
rect 6352 -1710 6368 -1708
rect 7102 -1642 7118 -1640
rect 7152 -1610 7168 -1608
rect 7902 -1542 7918 -1540
rect 7952 -1510 7968 -1508
rect 8702 -1442 8718 -1440
rect 8752 -1410 8768 -1408
rect 9502 -1342 9518 -1340
rect 9552 -1310 9568 -1308
rect 10302 -1242 10318 -1240
rect 10352 -1210 10368 -1208
rect 11102 -1142 11118 -1140
rect 11152 -1110 11168 -1108
rect 11902 -1042 11918 -1040
rect 11952 -1010 11968 -1008
rect 12702 -942 12718 -940
rect 12752 -910 12768 -908
rect 12752 -940 12776 -910
rect 12752 -942 12768 -940
rect 12702 -952 12768 -942
rect 14706 -909 14800 -890
rect 14706 -943 14734 -909
rect 14768 -943 14800 -909
rect 14706 -960 14800 -943
rect 15542 -909 15636 -890
rect 15542 -943 15574 -909
rect 15608 -943 15636 -909
rect 15542 -960 15636 -943
rect 14514 -990 14540 -960
rect 14690 -990 14816 -960
rect 15116 -990 15142 -960
rect 15200 -990 15226 -960
rect 15526 -990 15652 -960
rect 15802 -990 15828 -960
rect 12702 -1008 12768 -998
rect 12702 -1010 12718 -1008
rect 11952 -1040 11990 -1010
rect 12108 -1040 12162 -1010
rect 12280 -1040 12390 -1010
rect 12508 -1040 12562 -1010
rect 12680 -1040 12718 -1010
rect 11952 -1042 11968 -1040
rect 11902 -1052 11968 -1042
rect 11902 -1108 11968 -1098
rect 11902 -1110 11918 -1108
rect 11152 -1140 11190 -1110
rect 11308 -1140 11362 -1110
rect 11480 -1140 11590 -1110
rect 11708 -1140 11762 -1110
rect 11880 -1140 11918 -1110
rect 11152 -1142 11168 -1140
rect 11102 -1152 11168 -1142
rect 11102 -1208 11168 -1198
rect 11102 -1210 11118 -1208
rect 10352 -1240 10390 -1210
rect 10508 -1240 10562 -1210
rect 10680 -1240 10790 -1210
rect 10908 -1240 10962 -1210
rect 11080 -1240 11118 -1210
rect 10352 -1242 10368 -1240
rect 10302 -1252 10368 -1242
rect 10302 -1308 10368 -1298
rect 10302 -1310 10318 -1308
rect 9552 -1340 9590 -1310
rect 9708 -1340 9762 -1310
rect 9880 -1340 9990 -1310
rect 10108 -1340 10162 -1310
rect 10280 -1340 10318 -1310
rect 9552 -1342 9568 -1340
rect 9502 -1352 9568 -1342
rect 9502 -1408 9568 -1398
rect 9502 -1410 9518 -1408
rect 8752 -1440 8790 -1410
rect 8908 -1440 8962 -1410
rect 9080 -1440 9190 -1410
rect 9308 -1440 9362 -1410
rect 9480 -1440 9518 -1410
rect 8752 -1442 8768 -1440
rect 8702 -1452 8768 -1442
rect 8702 -1508 8768 -1498
rect 8702 -1510 8718 -1508
rect 7952 -1540 7990 -1510
rect 8108 -1540 8162 -1510
rect 8280 -1540 8390 -1510
rect 8508 -1540 8562 -1510
rect 8680 -1540 8718 -1510
rect 7952 -1542 7968 -1540
rect 7902 -1552 7968 -1542
rect 7902 -1608 7968 -1598
rect 7902 -1610 7918 -1608
rect 7152 -1640 7190 -1610
rect 7308 -1640 7362 -1610
rect 7480 -1640 7590 -1610
rect 7708 -1640 7762 -1610
rect 7880 -1640 7918 -1610
rect 7152 -1642 7168 -1640
rect 7102 -1652 7168 -1642
rect 7102 -1708 7168 -1698
rect 7102 -1710 7118 -1708
rect 6352 -1740 6390 -1710
rect 6508 -1740 6562 -1710
rect 6680 -1740 6790 -1710
rect 6908 -1740 6962 -1710
rect 7080 -1740 7118 -1710
rect 6352 -1742 6368 -1740
rect 6302 -1752 6368 -1742
rect 6302 -1808 6368 -1798
rect 6302 -1810 6318 -1808
rect 5552 -1840 5590 -1810
rect 5708 -1840 5762 -1810
rect 5880 -1840 5990 -1810
rect 6108 -1840 6162 -1810
rect 6280 -1840 6318 -1810
rect 5552 -1842 5568 -1840
rect 5502 -1852 5568 -1842
rect 5502 -1908 5568 -1898
rect 5502 -1910 5518 -1908
rect 4752 -1940 4790 -1910
rect 4908 -1940 4962 -1910
rect 5080 -1940 5190 -1910
rect 5308 -1940 5362 -1910
rect 5480 -1940 5518 -1910
rect 4752 -1942 4768 -1940
rect 4702 -1952 4768 -1942
rect 4702 -2008 4768 -1998
rect 4702 -2010 4718 -2008
rect 3952 -2040 3990 -2010
rect 4108 -2040 4162 -2010
rect 4280 -2040 4390 -2010
rect 4508 -2040 4562 -2010
rect 4680 -2040 4718 -2010
rect 3952 -2042 3968 -2040
rect 3902 -2052 3968 -2042
rect 4702 -2042 4718 -2040
rect 4752 -2010 4768 -2008
rect 5502 -1942 5518 -1940
rect 5552 -1910 5568 -1908
rect 6302 -1842 6318 -1840
rect 6352 -1810 6368 -1808
rect 7102 -1742 7118 -1740
rect 7152 -1710 7168 -1708
rect 7902 -1642 7918 -1640
rect 7952 -1610 7968 -1608
rect 8702 -1542 8718 -1540
rect 8752 -1510 8768 -1508
rect 9502 -1442 9518 -1440
rect 9552 -1410 9568 -1408
rect 10302 -1342 10318 -1340
rect 10352 -1310 10368 -1308
rect 11102 -1242 11118 -1240
rect 11152 -1210 11168 -1208
rect 11902 -1142 11918 -1140
rect 11952 -1110 11968 -1108
rect 12702 -1042 12718 -1040
rect 12752 -1010 12768 -1008
rect 12752 -1040 12776 -1010
rect 12752 -1042 12768 -1040
rect 12702 -1052 12768 -1042
rect 14514 -1090 14540 -1060
rect 14690 -1090 14816 -1060
rect 15116 -1090 15142 -1060
rect 15200 -1090 15226 -1060
rect 15526 -1090 15652 -1060
rect 15802 -1090 15828 -1060
rect 12702 -1108 12768 -1098
rect 12702 -1110 12718 -1108
rect 11952 -1140 11990 -1110
rect 12108 -1140 12162 -1110
rect 12280 -1140 12390 -1110
rect 12508 -1140 12562 -1110
rect 12680 -1140 12718 -1110
rect 11952 -1142 11968 -1140
rect 11902 -1152 11968 -1142
rect 11902 -1208 11968 -1198
rect 11902 -1210 11918 -1208
rect 11152 -1240 11190 -1210
rect 11308 -1240 11362 -1210
rect 11480 -1240 11590 -1210
rect 11708 -1240 11762 -1210
rect 11880 -1240 11918 -1210
rect 11152 -1242 11168 -1240
rect 11102 -1252 11168 -1242
rect 11102 -1308 11168 -1298
rect 11102 -1310 11118 -1308
rect 10352 -1340 10390 -1310
rect 10508 -1340 10562 -1310
rect 10680 -1340 10790 -1310
rect 10908 -1340 10962 -1310
rect 11080 -1340 11118 -1310
rect 10352 -1342 10368 -1340
rect 10302 -1352 10368 -1342
rect 10302 -1408 10368 -1398
rect 10302 -1410 10318 -1408
rect 9552 -1440 9590 -1410
rect 9708 -1440 9762 -1410
rect 9880 -1440 9990 -1410
rect 10108 -1440 10162 -1410
rect 10280 -1440 10318 -1410
rect 9552 -1442 9568 -1440
rect 9502 -1452 9568 -1442
rect 9502 -1508 9568 -1498
rect 9502 -1510 9518 -1508
rect 8752 -1540 8790 -1510
rect 8908 -1540 8962 -1510
rect 9080 -1540 9190 -1510
rect 9308 -1540 9362 -1510
rect 9480 -1540 9518 -1510
rect 8752 -1542 8768 -1540
rect 8702 -1552 8768 -1542
rect 8702 -1608 8768 -1598
rect 8702 -1610 8718 -1608
rect 7952 -1640 7990 -1610
rect 8108 -1640 8162 -1610
rect 8280 -1640 8390 -1610
rect 8508 -1640 8562 -1610
rect 8680 -1640 8718 -1610
rect 7952 -1642 7968 -1640
rect 7902 -1652 7968 -1642
rect 7902 -1708 7968 -1698
rect 7902 -1710 7918 -1708
rect 7152 -1740 7190 -1710
rect 7308 -1740 7362 -1710
rect 7480 -1740 7590 -1710
rect 7708 -1740 7762 -1710
rect 7880 -1740 7918 -1710
rect 7152 -1742 7168 -1740
rect 7102 -1752 7168 -1742
rect 7102 -1808 7168 -1798
rect 7102 -1810 7118 -1808
rect 6352 -1840 6390 -1810
rect 6508 -1840 6562 -1810
rect 6680 -1840 6790 -1810
rect 6908 -1840 6962 -1810
rect 7080 -1840 7118 -1810
rect 6352 -1842 6368 -1840
rect 6302 -1852 6368 -1842
rect 6302 -1908 6368 -1898
rect 6302 -1910 6318 -1908
rect 5552 -1940 5590 -1910
rect 5708 -1940 5762 -1910
rect 5880 -1940 5990 -1910
rect 6108 -1940 6162 -1910
rect 6280 -1940 6318 -1910
rect 5552 -1942 5568 -1940
rect 5502 -1952 5568 -1942
rect 5502 -2008 5568 -1998
rect 5502 -2010 5518 -2008
rect 4752 -2040 4790 -2010
rect 4908 -2040 4962 -2010
rect 5080 -2040 5190 -2010
rect 5308 -2040 5362 -2010
rect 5480 -2040 5518 -2010
rect 4752 -2042 4768 -2040
rect 4702 -2052 4768 -2042
rect 5502 -2042 5518 -2040
rect 5552 -2010 5568 -2008
rect 6302 -1942 6318 -1940
rect 6352 -1910 6368 -1908
rect 7102 -1842 7118 -1840
rect 7152 -1810 7168 -1808
rect 7902 -1742 7918 -1740
rect 7952 -1710 7968 -1708
rect 8702 -1642 8718 -1640
rect 8752 -1610 8768 -1608
rect 9502 -1542 9518 -1540
rect 9552 -1510 9568 -1508
rect 10302 -1442 10318 -1440
rect 10352 -1410 10368 -1408
rect 11102 -1342 11118 -1340
rect 11152 -1310 11168 -1308
rect 11902 -1242 11918 -1240
rect 11952 -1210 11968 -1208
rect 12702 -1142 12718 -1140
rect 12752 -1110 12768 -1108
rect 12752 -1140 12776 -1110
rect 12752 -1142 12768 -1140
rect 12702 -1152 12768 -1142
rect 14706 -1109 14800 -1090
rect 14706 -1143 14734 -1109
rect 14768 -1143 14800 -1109
rect 14706 -1160 14800 -1143
rect 15542 -1109 15636 -1090
rect 15542 -1143 15574 -1109
rect 15608 -1143 15636 -1109
rect 15542 -1160 15636 -1143
rect 14514 -1190 14540 -1160
rect 14690 -1190 14816 -1160
rect 15116 -1190 15142 -1160
rect 15200 -1190 15226 -1160
rect 15526 -1190 15652 -1160
rect 15802 -1190 15828 -1160
rect 12702 -1208 12768 -1198
rect 12702 -1210 12718 -1208
rect 11952 -1240 11990 -1210
rect 12108 -1240 12162 -1210
rect 12280 -1240 12390 -1210
rect 12508 -1240 12562 -1210
rect 12680 -1240 12718 -1210
rect 11952 -1242 11968 -1240
rect 11902 -1252 11968 -1242
rect 11902 -1308 11968 -1298
rect 11902 -1310 11918 -1308
rect 11152 -1340 11190 -1310
rect 11308 -1340 11362 -1310
rect 11480 -1340 11590 -1310
rect 11708 -1340 11762 -1310
rect 11880 -1340 11918 -1310
rect 11152 -1342 11168 -1340
rect 11102 -1352 11168 -1342
rect 11102 -1408 11168 -1398
rect 11102 -1410 11118 -1408
rect 10352 -1440 10390 -1410
rect 10508 -1440 10562 -1410
rect 10680 -1440 10790 -1410
rect 10908 -1440 10962 -1410
rect 11080 -1440 11118 -1410
rect 10352 -1442 10368 -1440
rect 10302 -1452 10368 -1442
rect 10302 -1508 10368 -1498
rect 10302 -1510 10318 -1508
rect 9552 -1540 9590 -1510
rect 9708 -1540 9762 -1510
rect 9880 -1540 9990 -1510
rect 10108 -1540 10162 -1510
rect 10280 -1540 10318 -1510
rect 9552 -1542 9568 -1540
rect 9502 -1552 9568 -1542
rect 9502 -1608 9568 -1598
rect 9502 -1610 9518 -1608
rect 8752 -1640 8790 -1610
rect 8908 -1640 8962 -1610
rect 9080 -1640 9190 -1610
rect 9308 -1640 9362 -1610
rect 9480 -1640 9518 -1610
rect 8752 -1642 8768 -1640
rect 8702 -1652 8768 -1642
rect 8702 -1708 8768 -1698
rect 8702 -1710 8718 -1708
rect 7952 -1740 7990 -1710
rect 8108 -1740 8162 -1710
rect 8280 -1740 8390 -1710
rect 8508 -1740 8562 -1710
rect 8680 -1740 8718 -1710
rect 7952 -1742 7968 -1740
rect 7902 -1752 7968 -1742
rect 7902 -1808 7968 -1798
rect 7902 -1810 7918 -1808
rect 7152 -1840 7190 -1810
rect 7308 -1840 7362 -1810
rect 7480 -1840 7590 -1810
rect 7708 -1840 7762 -1810
rect 7880 -1840 7918 -1810
rect 7152 -1842 7168 -1840
rect 7102 -1852 7168 -1842
rect 7102 -1908 7168 -1898
rect 7102 -1910 7118 -1908
rect 6352 -1940 6390 -1910
rect 6508 -1940 6562 -1910
rect 6680 -1940 6790 -1910
rect 6908 -1940 6962 -1910
rect 7080 -1940 7118 -1910
rect 6352 -1942 6368 -1940
rect 6302 -1952 6368 -1942
rect 6302 -2008 6368 -1998
rect 6302 -2010 6318 -2008
rect 5552 -2040 5590 -2010
rect 5708 -2040 5762 -2010
rect 5880 -2040 5990 -2010
rect 6108 -2040 6162 -2010
rect 6280 -2040 6318 -2010
rect 5552 -2042 5568 -2040
rect 5502 -2052 5568 -2042
rect 6302 -2042 6318 -2040
rect 6352 -2010 6368 -2008
rect 7102 -1942 7118 -1940
rect 7152 -1910 7168 -1908
rect 7902 -1842 7918 -1840
rect 7952 -1810 7968 -1808
rect 8702 -1742 8718 -1740
rect 8752 -1710 8768 -1708
rect 9502 -1642 9518 -1640
rect 9552 -1610 9568 -1608
rect 10302 -1542 10318 -1540
rect 10352 -1510 10368 -1508
rect 11102 -1442 11118 -1440
rect 11152 -1410 11168 -1408
rect 11902 -1342 11918 -1340
rect 11952 -1310 11968 -1308
rect 12702 -1242 12718 -1240
rect 12752 -1210 12768 -1208
rect 12752 -1240 12776 -1210
rect 12752 -1242 12768 -1240
rect 12702 -1252 12768 -1242
rect 14514 -1290 14540 -1260
rect 14690 -1290 14816 -1260
rect 15116 -1290 15142 -1260
rect 15200 -1290 15226 -1260
rect 15526 -1290 15652 -1260
rect 15802 -1290 15828 -1260
rect 12702 -1308 12768 -1298
rect 12702 -1310 12718 -1308
rect 11952 -1340 11990 -1310
rect 12108 -1340 12162 -1310
rect 12280 -1340 12390 -1310
rect 12508 -1340 12562 -1310
rect 12680 -1340 12718 -1310
rect 11952 -1342 11968 -1340
rect 11902 -1352 11968 -1342
rect 11902 -1408 11968 -1398
rect 11902 -1410 11918 -1408
rect 11152 -1440 11190 -1410
rect 11308 -1440 11362 -1410
rect 11480 -1440 11590 -1410
rect 11708 -1440 11762 -1410
rect 11880 -1440 11918 -1410
rect 11152 -1442 11168 -1440
rect 11102 -1452 11168 -1442
rect 11102 -1508 11168 -1498
rect 11102 -1510 11118 -1508
rect 10352 -1540 10390 -1510
rect 10508 -1540 10562 -1510
rect 10680 -1540 10790 -1510
rect 10908 -1540 10962 -1510
rect 11080 -1540 11118 -1510
rect 10352 -1542 10368 -1540
rect 10302 -1552 10368 -1542
rect 10302 -1608 10368 -1598
rect 10302 -1610 10318 -1608
rect 9552 -1640 9590 -1610
rect 9708 -1640 9762 -1610
rect 9880 -1640 9990 -1610
rect 10108 -1640 10162 -1610
rect 10280 -1640 10318 -1610
rect 9552 -1642 9568 -1640
rect 9502 -1652 9568 -1642
rect 9502 -1708 9568 -1698
rect 9502 -1710 9518 -1708
rect 8752 -1740 8790 -1710
rect 8908 -1740 8962 -1710
rect 9080 -1740 9190 -1710
rect 9308 -1740 9362 -1710
rect 9480 -1740 9518 -1710
rect 8752 -1742 8768 -1740
rect 8702 -1752 8768 -1742
rect 8702 -1808 8768 -1798
rect 8702 -1810 8718 -1808
rect 7952 -1840 7990 -1810
rect 8108 -1840 8162 -1810
rect 8280 -1840 8390 -1810
rect 8508 -1840 8562 -1810
rect 8680 -1840 8718 -1810
rect 7952 -1842 7968 -1840
rect 7902 -1852 7968 -1842
rect 7902 -1908 7968 -1898
rect 7902 -1910 7918 -1908
rect 7152 -1940 7190 -1910
rect 7308 -1940 7362 -1910
rect 7480 -1940 7590 -1910
rect 7708 -1940 7762 -1910
rect 7880 -1940 7918 -1910
rect 7152 -1942 7168 -1940
rect 7102 -1952 7168 -1942
rect 7102 -2008 7168 -1998
rect 7102 -2010 7118 -2008
rect 6352 -2040 6390 -2010
rect 6508 -2040 6562 -2010
rect 6680 -2040 6790 -2010
rect 6908 -2040 6962 -2010
rect 7080 -2040 7118 -2010
rect 6352 -2042 6368 -2040
rect 6302 -2052 6368 -2042
rect 7102 -2042 7118 -2040
rect 7152 -2010 7168 -2008
rect 7902 -1942 7918 -1940
rect 7952 -1910 7968 -1908
rect 8702 -1842 8718 -1840
rect 8752 -1810 8768 -1808
rect 9502 -1742 9518 -1740
rect 9552 -1710 9568 -1708
rect 10302 -1642 10318 -1640
rect 10352 -1610 10368 -1608
rect 11102 -1542 11118 -1540
rect 11152 -1510 11168 -1508
rect 11902 -1442 11918 -1440
rect 11952 -1410 11968 -1408
rect 12702 -1342 12718 -1340
rect 12752 -1310 12768 -1308
rect 12752 -1340 12776 -1310
rect 12752 -1342 12768 -1340
rect 12702 -1352 12768 -1342
rect 14706 -1309 14800 -1290
rect 14706 -1343 14734 -1309
rect 14768 -1343 14800 -1309
rect 14706 -1360 14800 -1343
rect 15542 -1309 15636 -1290
rect 15542 -1343 15574 -1309
rect 15608 -1343 15636 -1309
rect 15542 -1360 15636 -1343
rect 14514 -1390 14540 -1360
rect 14690 -1390 14816 -1360
rect 15116 -1390 15142 -1360
rect 15200 -1390 15226 -1360
rect 15526 -1390 15652 -1360
rect 15802 -1390 15828 -1360
rect 12702 -1408 12768 -1398
rect 12702 -1410 12718 -1408
rect 11952 -1440 11990 -1410
rect 12108 -1440 12162 -1410
rect 12280 -1440 12390 -1410
rect 12508 -1440 12562 -1410
rect 12680 -1440 12718 -1410
rect 11952 -1442 11968 -1440
rect 11902 -1452 11968 -1442
rect 11902 -1508 11968 -1498
rect 11902 -1510 11918 -1508
rect 11152 -1540 11190 -1510
rect 11308 -1540 11362 -1510
rect 11480 -1540 11590 -1510
rect 11708 -1540 11762 -1510
rect 11880 -1540 11918 -1510
rect 11152 -1542 11168 -1540
rect 11102 -1552 11168 -1542
rect 11102 -1608 11168 -1598
rect 11102 -1610 11118 -1608
rect 10352 -1640 10390 -1610
rect 10508 -1640 10562 -1610
rect 10680 -1640 10790 -1610
rect 10908 -1640 10962 -1610
rect 11080 -1640 11118 -1610
rect 10352 -1642 10368 -1640
rect 10302 -1652 10368 -1642
rect 10302 -1708 10368 -1698
rect 10302 -1710 10318 -1708
rect 9552 -1740 9590 -1710
rect 9708 -1740 9762 -1710
rect 9880 -1740 9990 -1710
rect 10108 -1740 10162 -1710
rect 10280 -1740 10318 -1710
rect 9552 -1742 9568 -1740
rect 9502 -1752 9568 -1742
rect 9502 -1808 9568 -1798
rect 9502 -1810 9518 -1808
rect 8752 -1840 8790 -1810
rect 8908 -1840 8962 -1810
rect 9080 -1840 9190 -1810
rect 9308 -1840 9362 -1810
rect 9480 -1840 9518 -1810
rect 8752 -1842 8768 -1840
rect 8702 -1852 8768 -1842
rect 8702 -1908 8768 -1898
rect 8702 -1910 8718 -1908
rect 7952 -1940 7990 -1910
rect 8108 -1940 8162 -1910
rect 8280 -1940 8390 -1910
rect 8508 -1940 8562 -1910
rect 8680 -1940 8718 -1910
rect 7952 -1942 7968 -1940
rect 7902 -1952 7968 -1942
rect 7902 -2008 7968 -1998
rect 7902 -2010 7918 -2008
rect 7152 -2040 7190 -2010
rect 7308 -2040 7362 -2010
rect 7480 -2040 7590 -2010
rect 7708 -2040 7762 -2010
rect 7880 -2040 7918 -2010
rect 7152 -2042 7168 -2040
rect 7102 -2052 7168 -2042
rect 7902 -2042 7918 -2040
rect 7952 -2010 7968 -2008
rect 8702 -1942 8718 -1940
rect 8752 -1910 8768 -1908
rect 9502 -1842 9518 -1840
rect 9552 -1810 9568 -1808
rect 10302 -1742 10318 -1740
rect 10352 -1710 10368 -1708
rect 11102 -1642 11118 -1640
rect 11152 -1610 11168 -1608
rect 11902 -1542 11918 -1540
rect 11952 -1510 11968 -1508
rect 12702 -1442 12718 -1440
rect 12752 -1410 12768 -1408
rect 12752 -1440 12776 -1410
rect 12752 -1442 12768 -1440
rect 12702 -1452 12768 -1442
rect 14514 -1490 14540 -1460
rect 14690 -1490 14816 -1460
rect 15116 -1490 15142 -1460
rect 15200 -1490 15226 -1460
rect 15526 -1490 15652 -1460
rect 15802 -1490 15828 -1460
rect 12702 -1508 12768 -1498
rect 12702 -1510 12718 -1508
rect 11952 -1540 11990 -1510
rect 12108 -1540 12162 -1510
rect 12280 -1540 12390 -1510
rect 12508 -1540 12562 -1510
rect 12680 -1540 12718 -1510
rect 11952 -1542 11968 -1540
rect 11902 -1552 11968 -1542
rect 11902 -1608 11968 -1598
rect 11902 -1610 11918 -1608
rect 11152 -1640 11190 -1610
rect 11308 -1640 11362 -1610
rect 11480 -1640 11590 -1610
rect 11708 -1640 11762 -1610
rect 11880 -1640 11918 -1610
rect 11152 -1642 11168 -1640
rect 11102 -1652 11168 -1642
rect 11102 -1708 11168 -1698
rect 11102 -1710 11118 -1708
rect 10352 -1740 10390 -1710
rect 10508 -1740 10562 -1710
rect 10680 -1740 10790 -1710
rect 10908 -1740 10962 -1710
rect 11080 -1740 11118 -1710
rect 10352 -1742 10368 -1740
rect 10302 -1752 10368 -1742
rect 10302 -1808 10368 -1798
rect 10302 -1810 10318 -1808
rect 9552 -1840 9590 -1810
rect 9708 -1840 9762 -1810
rect 9880 -1840 9990 -1810
rect 10108 -1840 10162 -1810
rect 10280 -1840 10318 -1810
rect 9552 -1842 9568 -1840
rect 9502 -1852 9568 -1842
rect 9502 -1908 9568 -1898
rect 9502 -1910 9518 -1908
rect 8752 -1940 8790 -1910
rect 8908 -1940 8962 -1910
rect 9080 -1940 9190 -1910
rect 9308 -1940 9362 -1910
rect 9480 -1940 9518 -1910
rect 8752 -1942 8768 -1940
rect 8702 -1952 8768 -1942
rect 8702 -2008 8768 -1998
rect 8702 -2010 8718 -2008
rect 7952 -2040 7990 -2010
rect 8108 -2040 8162 -2010
rect 8280 -2040 8390 -2010
rect 8508 -2040 8562 -2010
rect 8680 -2040 8718 -2010
rect 7952 -2042 7968 -2040
rect 7902 -2052 7968 -2042
rect 8702 -2042 8718 -2040
rect 8752 -2010 8768 -2008
rect 9502 -1942 9518 -1940
rect 9552 -1910 9568 -1908
rect 10302 -1842 10318 -1840
rect 10352 -1810 10368 -1808
rect 11102 -1742 11118 -1740
rect 11152 -1710 11168 -1708
rect 11902 -1642 11918 -1640
rect 11952 -1610 11968 -1608
rect 12702 -1542 12718 -1540
rect 12752 -1510 12768 -1508
rect 12752 -1540 12776 -1510
rect 12752 -1542 12768 -1540
rect 12702 -1552 12768 -1542
rect 14706 -1509 14800 -1490
rect 14706 -1543 14734 -1509
rect 14768 -1543 14800 -1509
rect 14706 -1560 14800 -1543
rect 15542 -1509 15636 -1490
rect 15542 -1543 15574 -1509
rect 15608 -1543 15636 -1509
rect 15542 -1560 15636 -1543
rect 14514 -1590 14540 -1560
rect 14690 -1590 14816 -1560
rect 15116 -1590 15142 -1560
rect 15200 -1590 15226 -1560
rect 15526 -1590 15652 -1560
rect 15802 -1590 15828 -1560
rect 12702 -1608 12768 -1598
rect 12702 -1610 12718 -1608
rect 11952 -1640 11990 -1610
rect 12108 -1640 12162 -1610
rect 12280 -1640 12390 -1610
rect 12508 -1640 12562 -1610
rect 12680 -1640 12718 -1610
rect 11952 -1642 11968 -1640
rect 11902 -1652 11968 -1642
rect 11902 -1708 11968 -1698
rect 11902 -1710 11918 -1708
rect 11152 -1740 11190 -1710
rect 11308 -1740 11362 -1710
rect 11480 -1740 11590 -1710
rect 11708 -1740 11762 -1710
rect 11880 -1740 11918 -1710
rect 11152 -1742 11168 -1740
rect 11102 -1752 11168 -1742
rect 11102 -1808 11168 -1798
rect 11102 -1810 11118 -1808
rect 10352 -1840 10390 -1810
rect 10508 -1840 10562 -1810
rect 10680 -1840 10790 -1810
rect 10908 -1840 10962 -1810
rect 11080 -1840 11118 -1810
rect 10352 -1842 10368 -1840
rect 10302 -1852 10368 -1842
rect 10302 -1908 10368 -1898
rect 10302 -1910 10318 -1908
rect 9552 -1940 9590 -1910
rect 9708 -1940 9762 -1910
rect 9880 -1940 9990 -1910
rect 10108 -1940 10162 -1910
rect 10280 -1940 10318 -1910
rect 9552 -1942 9568 -1940
rect 9502 -1952 9568 -1942
rect 9502 -2008 9568 -1998
rect 9502 -2010 9518 -2008
rect 8752 -2040 8790 -2010
rect 8908 -2040 8962 -2010
rect 9080 -2040 9190 -2010
rect 9308 -2040 9362 -2010
rect 9480 -2040 9518 -2010
rect 8752 -2042 8768 -2040
rect 8702 -2052 8768 -2042
rect 9502 -2042 9518 -2040
rect 9552 -2010 9568 -2008
rect 10302 -1942 10318 -1940
rect 10352 -1910 10368 -1908
rect 11102 -1842 11118 -1840
rect 11152 -1810 11168 -1808
rect 11902 -1742 11918 -1740
rect 11952 -1710 11968 -1708
rect 12702 -1642 12718 -1640
rect 12752 -1610 12768 -1608
rect 12752 -1640 12776 -1610
rect 12752 -1642 12768 -1640
rect 12702 -1652 12768 -1642
rect 14514 -1690 14540 -1660
rect 14690 -1690 14816 -1660
rect 15116 -1690 15142 -1660
rect 15200 -1690 15226 -1660
rect 15526 -1690 15652 -1660
rect 15802 -1690 15828 -1660
rect 12702 -1708 12768 -1698
rect 12702 -1710 12718 -1708
rect 11952 -1740 11990 -1710
rect 12108 -1740 12162 -1710
rect 12280 -1740 12390 -1710
rect 12508 -1740 12562 -1710
rect 12680 -1740 12718 -1710
rect 11952 -1742 11968 -1740
rect 11902 -1752 11968 -1742
rect 11902 -1808 11968 -1798
rect 11902 -1810 11918 -1808
rect 11152 -1840 11190 -1810
rect 11308 -1840 11362 -1810
rect 11480 -1840 11590 -1810
rect 11708 -1840 11762 -1810
rect 11880 -1840 11918 -1810
rect 11152 -1842 11168 -1840
rect 11102 -1852 11168 -1842
rect 11102 -1908 11168 -1898
rect 11102 -1910 11118 -1908
rect 10352 -1940 10390 -1910
rect 10508 -1940 10562 -1910
rect 10680 -1940 10790 -1910
rect 10908 -1940 10962 -1910
rect 11080 -1940 11118 -1910
rect 10352 -1942 10368 -1940
rect 10302 -1952 10368 -1942
rect 10302 -2008 10368 -1998
rect 10302 -2010 10318 -2008
rect 9552 -2040 9590 -2010
rect 9708 -2040 9762 -2010
rect 9880 -2040 9990 -2010
rect 10108 -2040 10162 -2010
rect 10280 -2040 10318 -2010
rect 9552 -2042 9568 -2040
rect 9502 -2052 9568 -2042
rect 10302 -2042 10318 -2040
rect 10352 -2010 10368 -2008
rect 11102 -1942 11118 -1940
rect 11152 -1910 11168 -1908
rect 11902 -1842 11918 -1840
rect 11952 -1810 11968 -1808
rect 12702 -1742 12718 -1740
rect 12752 -1710 12768 -1708
rect 12752 -1740 12776 -1710
rect 12752 -1742 12768 -1740
rect 12702 -1752 12768 -1742
rect 14706 -1709 14800 -1690
rect 14706 -1743 14734 -1709
rect 14768 -1743 14800 -1709
rect 14706 -1760 14800 -1743
rect 15542 -1709 15636 -1690
rect 15542 -1743 15574 -1709
rect 15608 -1743 15636 -1709
rect 15542 -1760 15636 -1743
rect 14514 -1790 14540 -1760
rect 14690 -1790 14816 -1760
rect 15116 -1790 15142 -1760
rect 15200 -1790 15226 -1760
rect 15526 -1790 15652 -1760
rect 15802 -1790 15828 -1760
rect 12702 -1808 12768 -1798
rect 12702 -1810 12718 -1808
rect 11952 -1840 11990 -1810
rect 12108 -1840 12162 -1810
rect 12280 -1840 12390 -1810
rect 12508 -1840 12562 -1810
rect 12680 -1840 12718 -1810
rect 11952 -1842 11968 -1840
rect 11902 -1852 11968 -1842
rect 11902 -1908 11968 -1898
rect 11902 -1910 11918 -1908
rect 11152 -1940 11190 -1910
rect 11308 -1940 11362 -1910
rect 11480 -1940 11590 -1910
rect 11708 -1940 11762 -1910
rect 11880 -1940 11918 -1910
rect 11152 -1942 11168 -1940
rect 11102 -1952 11168 -1942
rect 11102 -2008 11168 -1998
rect 11102 -2010 11118 -2008
rect 10352 -2040 10390 -2010
rect 10508 -2040 10562 -2010
rect 10680 -2040 10790 -2010
rect 10908 -2040 10962 -2010
rect 11080 -2040 11118 -2010
rect 10352 -2042 10368 -2040
rect 10302 -2052 10368 -2042
rect 11102 -2042 11118 -2040
rect 11152 -2010 11168 -2008
rect 11902 -1942 11918 -1940
rect 11952 -1910 11968 -1908
rect 12702 -1842 12718 -1840
rect 12752 -1810 12768 -1808
rect 12752 -1840 12776 -1810
rect 12752 -1842 12768 -1840
rect 12702 -1852 12768 -1842
rect 14514 -1890 14540 -1860
rect 14690 -1890 14816 -1860
rect 15116 -1890 15142 -1860
rect 15200 -1890 15226 -1860
rect 15526 -1890 15652 -1860
rect 15802 -1890 15828 -1860
rect 12702 -1908 12768 -1898
rect 12702 -1910 12718 -1908
rect 11952 -1940 11990 -1910
rect 12108 -1940 12162 -1910
rect 12280 -1940 12390 -1910
rect 12508 -1940 12562 -1910
rect 12680 -1940 12718 -1910
rect 11952 -1942 11968 -1940
rect 11902 -1952 11968 -1942
rect 11902 -2008 11968 -1998
rect 11902 -2010 11918 -2008
rect 11152 -2040 11190 -2010
rect 11308 -2040 11362 -2010
rect 11480 -2040 11590 -2010
rect 11708 -2040 11762 -2010
rect 11880 -2040 11918 -2010
rect 11152 -2042 11168 -2040
rect 11102 -2052 11168 -2042
rect 11902 -2042 11918 -2040
rect 11952 -2010 11968 -2008
rect 12702 -1942 12718 -1940
rect 12752 -1910 12768 -1908
rect 12752 -1940 12776 -1910
rect 12752 -1942 12768 -1940
rect 12702 -1952 12768 -1942
rect 14706 -1909 14800 -1890
rect 14706 -1943 14734 -1909
rect 14768 -1943 14800 -1909
rect 14706 -1960 14800 -1943
rect 15542 -1909 15636 -1890
rect 15542 -1943 15574 -1909
rect 15608 -1943 15636 -1909
rect 15542 -1960 15636 -1943
rect 14514 -1990 14540 -1960
rect 14690 -1990 14816 -1960
rect 15116 -1990 15142 -1960
rect 15200 -1990 15226 -1960
rect 15526 -1990 15652 -1960
rect 15802 -1990 15828 -1960
rect 12702 -2008 12768 -1998
rect 12702 -2010 12718 -2008
rect 11952 -2040 11990 -2010
rect 12108 -2040 12162 -2010
rect 12280 -2040 12390 -2010
rect 12508 -2040 12562 -2010
rect 12680 -2040 12718 -2010
rect 11952 -2042 11968 -2040
rect 11902 -2052 11968 -2042
rect 12702 -2042 12718 -2040
rect 12752 -2010 12768 -2008
rect 12752 -2040 12776 -2010
rect 12752 -2042 12768 -2040
rect 12702 -2052 12768 -2042
<< polycont >>
rect 118 4860 152 4894
rect 318 4876 352 4910
rect 518 4860 552 4894
rect 718 4876 752 4910
rect 918 4860 952 4894
rect 1118 4876 1152 4910
rect 1318 4860 1352 4894
rect 1518 4876 1552 4910
rect 1718 4860 1752 4894
rect 1918 4876 1952 4910
rect 2118 4860 2152 4894
rect 2318 4876 2352 4910
rect 2518 4860 2552 4894
rect 2718 4876 2752 4910
rect 2918 4860 2952 4894
rect 3118 4876 3152 4910
rect 3318 4860 3352 4894
rect 3518 4876 3552 4910
rect 3718 4860 3752 4894
rect 3918 4876 3952 4910
rect 4118 4860 4152 4894
rect 4318 4876 4352 4910
rect 4518 4860 4552 4894
rect 4718 4876 4752 4910
rect 4918 4860 4952 4894
rect 5118 4876 5152 4910
rect 5318 4860 5352 4894
rect 5518 4876 5552 4910
rect 5718 4860 5752 4894
rect 5918 4876 5952 4910
rect 6118 4860 6152 4894
rect 6318 4876 6352 4910
rect 6518 4860 6552 4894
rect 118 3650 152 3684
rect 318 3666 352 3700
rect 518 3650 552 3684
rect 718 3666 752 3700
rect 918 3650 952 3684
rect 1118 3666 1152 3700
rect 1318 3650 1352 3684
rect 1518 3666 1552 3700
rect 1718 3650 1752 3684
rect 1918 3666 1952 3700
rect 2118 3650 2152 3684
rect 2318 3666 2352 3700
rect 2518 3650 2552 3684
rect 2718 3666 2752 3700
rect 2918 3650 2952 3684
rect 3118 3666 3152 3700
rect 3318 3650 3352 3684
rect 3518 3666 3552 3700
rect 3718 3650 3752 3684
rect 3918 3666 3952 3700
rect 4118 3650 4152 3684
rect 4318 3666 4352 3700
rect 4518 3650 4552 3684
rect 4718 3666 4752 3700
rect 4918 3650 4952 3684
rect 5118 3666 5152 3700
rect 5318 3650 5352 3684
rect 6718 4876 6752 4910
rect 6918 4860 6952 4894
rect 7118 4876 7152 4910
rect 7318 4860 7352 4894
rect 7518 4876 7552 4910
rect 7718 4860 7752 4894
rect 7918 4876 7952 4910
rect 8118 4860 8152 4894
rect 8318 4876 8352 4910
rect 8518 4860 8552 4894
rect 8718 4876 8752 4910
rect 8918 4860 8952 4894
rect 9118 4876 9152 4910
rect 9318 4860 9352 4894
rect 9518 4876 9552 4910
rect 9718 4860 9752 4894
rect 9918 4876 9952 4910
rect 10118 4860 10152 4894
rect 10318 4876 10352 4910
rect 10518 4860 10552 4894
rect 10718 4876 10752 4910
rect 10918 4860 10952 4894
rect 11118 4876 11152 4910
rect 11318 4860 11352 4894
rect 11518 4876 11552 4910
rect 11718 4860 11752 4894
rect 11918 4876 11952 4910
rect 12118 4860 12152 4894
rect 12318 4876 12352 4910
rect 12518 4860 12552 4894
rect 12718 4876 12752 4910
rect 12968 4874 13002 4908
rect 13068 4874 13102 4908
rect 13278 4874 13312 4908
rect 13378 4874 13412 4908
rect 13478 4874 13512 4908
rect 13578 4874 13612 4908
rect 5518 3666 5552 3700
rect 5718 3650 5752 3684
rect 5918 3666 5952 3700
rect 6118 3650 6152 3684
rect 6318 3666 6352 3700
rect 6518 3650 6552 3684
rect 6718 3666 6752 3700
rect 6918 3650 6952 3684
rect 7118 3666 7152 3700
rect 7318 3650 7352 3684
rect 7518 3666 7552 3700
rect 7718 3650 7752 3684
rect 7918 3666 7952 3700
rect 8118 3650 8152 3684
rect 8318 3666 8352 3700
rect 8518 3650 8552 3684
rect 8718 3666 8752 3700
rect 8918 3650 8952 3684
rect 9118 3666 9152 3700
rect 9318 3650 9352 3684
rect 9518 3666 9552 3700
rect 9718 3650 9752 3684
rect 9918 3666 9952 3700
rect 10118 3650 10152 3684
rect 118 2440 152 2474
rect 318 2456 352 2490
rect 518 2440 552 2474
rect 718 2456 752 2490
rect 918 2440 952 2474
rect 1118 2456 1152 2490
rect 1318 2440 1352 2474
rect 1518 2456 1552 2490
rect 1718 2440 1752 2474
rect 1918 2456 1952 2490
rect 2118 2440 2152 2474
rect 2318 2456 2352 2490
rect 2518 2440 2552 2474
rect 2718 2456 2752 2490
rect 2918 2440 2952 2474
rect 3118 2456 3152 2490
rect 3318 2440 3352 2474
rect 3518 2456 3552 2490
rect 3718 2440 3752 2474
rect 3918 2456 3952 2490
rect 4118 2440 4152 2474
rect 4318 2456 4352 2490
rect 4518 2440 4552 2474
rect 4718 2456 4752 2490
rect 4918 2440 4952 2474
rect 5118 2456 5152 2490
rect 5318 2440 5352 2474
rect 5518 2456 5552 2490
rect 5718 2440 5752 2474
rect 5918 2456 5952 2490
rect 6118 2440 6152 2474
rect 6318 2456 6352 2490
rect 6518 2440 6552 2474
rect 6718 2456 6752 2490
rect 6918 2440 6952 2474
rect 118 1230 152 1264
rect 318 1246 352 1280
rect 518 1230 552 1264
rect 718 1246 752 1280
rect 918 1230 952 1264
rect 1118 1246 1152 1280
rect 1318 1230 1352 1264
rect 1518 1246 1552 1280
rect 1718 1230 1752 1264
rect 1918 1246 1952 1280
rect 2118 1230 2152 1264
rect 2318 1246 2352 1280
rect 2518 1230 2552 1264
rect 2718 1246 2752 1280
rect 2918 1230 2952 1264
rect 3118 1246 3152 1280
rect 3318 1230 3352 1264
rect 118 20 152 54
rect 318 36 352 70
rect 518 20 552 54
rect 718 36 752 70
rect 918 20 952 54
rect 1118 36 1152 70
rect 1318 20 1352 54
rect 1518 36 1552 70
rect 3518 1246 3552 1280
rect 3718 1230 3752 1264
rect 3918 1246 3952 1280
rect 4118 1230 4152 1264
rect 4318 1246 4352 1280
rect 4518 1230 4552 1264
rect 4718 1246 4752 1280
rect 4918 1230 4952 1264
rect 7118 2456 7152 2490
rect 7318 2440 7352 2474
rect 7518 2456 7552 2490
rect 7718 2440 7752 2474
rect 7918 2456 7952 2490
rect 8118 2440 8152 2474
rect 8318 2456 8352 2490
rect 8518 2440 8552 2474
rect 10318 3666 10352 3700
rect 10518 3650 10552 3684
rect 10718 3666 10752 3700
rect 10918 3650 10952 3684
rect 11118 3666 11152 3700
rect 11318 3650 11352 3684
rect 11518 3666 11552 3700
rect 11718 3650 11752 3684
rect 11918 3666 11952 3700
rect 12118 3650 12152 3684
rect 12318 3666 12352 3700
rect 12518 3650 12552 3684
rect 12718 3666 12752 3700
rect 12968 3664 13002 3698
rect 13068 3664 13102 3698
rect 13278 3664 13312 3698
rect 13378 3664 13412 3698
rect 13478 3664 13512 3698
rect 13578 3664 13612 3698
rect 8718 2456 8752 2490
rect 8918 2440 8952 2474
rect 9118 2456 9152 2490
rect 9318 2440 9352 2474
rect 9518 2456 9552 2490
rect 9718 2440 9752 2474
rect 9918 2456 9952 2490
rect 10118 2440 10152 2474
rect 10318 2456 10352 2490
rect 10518 2440 10552 2474
rect 10718 2456 10752 2490
rect 10918 2440 10952 2474
rect 11118 2456 11152 2490
rect 11318 2440 11352 2474
rect 11518 2456 11552 2490
rect 11718 2440 11752 2474
rect 11918 2456 11952 2490
rect 12118 2440 12152 2474
rect 12318 2456 12352 2490
rect 12518 2440 12552 2474
rect 5118 1246 5152 1280
rect 5318 1230 5352 1264
rect 5518 1246 5552 1280
rect 5718 1230 5752 1264
rect 5918 1246 5952 1280
rect 6118 1230 6152 1264
rect 6318 1246 6352 1280
rect 6518 1230 6552 1264
rect 6718 1246 6752 1280
rect 6918 1230 6952 1264
rect 7118 1246 7152 1280
rect 7318 1230 7352 1264
rect 7518 1246 7552 1280
rect 7718 1230 7752 1264
rect 7918 1246 7952 1280
rect 8118 1230 8152 1264
rect 8318 1246 8352 1280
rect 8518 1230 8552 1264
rect 8718 1246 8752 1280
rect 8918 1230 8952 1264
rect 9118 1246 9152 1280
rect 12718 2456 12752 2490
rect 12968 2454 13002 2488
rect 13068 2454 13102 2488
rect 13278 2454 13312 2488
rect 13378 2454 13412 2488
rect 13478 2454 13512 2488
rect 13578 2454 13612 2488
rect 9318 1230 9352 1264
rect 9518 1246 9552 1280
rect 9718 1230 9752 1264
rect 1718 20 1752 54
rect 9918 1246 9952 1280
rect 10118 1230 10152 1264
rect 10318 1246 10352 1280
rect 10518 1230 10552 1264
rect 10718 1246 10752 1280
rect 10918 1230 10952 1264
rect 11118 1246 11152 1280
rect 1918 36 1952 70
rect 2118 20 2152 54
rect 2318 36 2352 70
rect 2518 20 2552 54
rect 2718 36 2752 70
rect 2918 20 2952 54
rect 3118 36 3152 70
rect 3318 20 3352 54
rect 3518 36 3552 70
rect 3718 20 3752 54
rect 3918 36 3952 70
rect 4118 20 4152 54
rect 4318 36 4352 70
rect 4518 20 4552 54
rect 4718 36 4752 70
rect 4918 20 4952 54
rect 5118 36 5152 70
rect 5318 20 5352 54
rect 5518 36 5552 70
rect 5718 20 5752 54
rect 5918 36 5952 70
rect 6118 20 6152 54
rect 6318 36 6352 70
rect 6518 20 6552 54
rect 6718 36 6752 70
rect 6918 20 6952 54
rect 11318 1230 11352 1264
rect 11518 1246 11552 1280
rect 11718 1230 11752 1264
rect 11918 1246 11952 1280
rect 12118 1230 12152 1264
rect 12318 1246 12352 1280
rect 12518 1230 12552 1264
rect 12718 1246 12752 1280
rect 12968 1244 13002 1278
rect 13068 1244 13102 1278
rect 13278 1244 13312 1278
rect 13378 1244 13412 1278
rect 13478 1244 13512 1278
rect 13578 1244 13612 1278
rect 7118 36 7152 70
rect 7318 20 7352 54
rect 7518 36 7552 70
rect 7718 20 7752 54
rect 7918 36 7952 70
rect 8118 20 8152 54
rect 8318 36 8352 70
rect 8518 20 8552 54
rect 8718 36 8752 70
rect 8918 20 8952 54
rect 9118 36 9152 70
rect 9318 20 9352 54
rect 9518 36 9552 70
rect 9718 20 9752 54
rect 9918 36 9952 70
rect 10118 20 10152 54
rect 10318 36 10352 70
rect 10518 20 10552 54
rect 10718 36 10752 70
rect 10918 20 10952 54
rect 11118 36 11152 70
rect 11318 20 11352 54
rect 11518 36 11552 70
rect 11718 20 11752 54
rect 11918 36 11952 70
rect 12118 20 12152 54
rect 12318 36 12352 70
rect 12518 20 12552 54
rect 12718 36 12752 70
rect 12968 34 13002 68
rect 13068 34 13102 68
rect 13278 34 13312 68
rect 13378 34 13412 68
rect 13478 34 13512 68
rect 13578 34 13612 68
rect 18 -282 52 -248
rect 218 -282 252 -248
rect 418 -282 452 -248
rect 618 -282 652 -248
rect 818 -282 852 -248
rect 1018 -282 1052 -248
rect 1218 -282 1252 -248
rect 1418 -282 1452 -248
rect 1618 -282 1652 -248
rect 1818 -282 1852 -248
rect 2018 -282 2052 -248
rect 2218 -282 2252 -248
rect 2418 -282 2452 -248
rect 2618 -282 2652 -248
rect 2818 -282 2852 -248
rect 3018 -282 3052 -248
rect 3218 -282 3252 -248
rect 3418 -282 3452 -248
rect 3618 -282 3652 -248
rect 3818 -282 3852 -248
rect 4018 -282 4052 -248
rect 4218 -282 4252 -248
rect 4418 -282 4452 -248
rect 4618 -282 4652 -248
rect 4818 -282 4852 -248
rect 5018 -282 5052 -248
rect 5218 -282 5252 -248
rect 5418 -282 5452 -248
rect 5618 -282 5652 -248
rect 5818 -282 5852 -248
rect 6018 -282 6052 -248
rect 6218 -282 6252 -248
rect 6418 -282 6452 -248
rect 6618 -282 6652 -248
rect 6818 -282 6852 -248
rect 7018 -282 7052 -248
rect 7218 -282 7252 -248
rect 7418 -282 7452 -248
rect 7618 -282 7652 -248
rect 7818 -282 7852 -248
rect 8018 -282 8052 -248
rect 8218 -282 8252 -248
rect 8418 -282 8452 -248
rect 8618 -282 8652 -248
rect 8818 -282 8852 -248
rect 9018 -282 9052 -248
rect 9218 -282 9252 -248
rect 9418 -282 9452 -248
rect 9618 -282 9652 -248
rect 9818 -282 9852 -248
rect 10018 -282 10052 -248
rect 10218 -282 10252 -248
rect 10418 -282 10452 -248
rect 10618 -282 10652 -248
rect 10818 -282 10852 -248
rect 11018 -282 11052 -248
rect 11218 -282 11252 -248
rect 11418 -282 11452 -248
rect 11618 -282 11652 -248
rect 11818 -282 11852 -248
rect 12018 -282 12052 -248
rect 12218 -282 12252 -248
rect 12418 -282 12452 -248
rect 12618 -282 12652 -248
rect 14734 -343 14768 -309
rect 15574 -343 15608 -309
rect 14734 -543 14768 -509
rect 15574 -543 15608 -509
rect 44 -611 78 -577
rect 192 -611 226 -577
rect 444 -611 478 -577
rect 592 -611 626 -577
rect 844 -611 878 -577
rect 992 -611 1026 -577
rect 1244 -611 1278 -577
rect 1392 -611 1426 -577
rect 1644 -611 1678 -577
rect 1792 -611 1826 -577
rect 2044 -611 2078 -577
rect 2192 -611 2226 -577
rect 2444 -611 2478 -577
rect 2592 -611 2626 -577
rect 2844 -611 2878 -577
rect 2992 -611 3026 -577
rect 3244 -611 3278 -577
rect 3392 -611 3426 -577
rect 3644 -611 3678 -577
rect 3792 -611 3826 -577
rect 4044 -611 4078 -577
rect 4192 -611 4226 -577
rect 4444 -611 4478 -577
rect 4592 -611 4626 -577
rect 4844 -611 4878 -577
rect 4992 -611 5026 -577
rect 5244 -611 5278 -577
rect 5392 -611 5426 -577
rect 5644 -611 5678 -577
rect 5792 -611 5826 -577
rect 6044 -611 6078 -577
rect 6192 -611 6226 -577
rect 6444 -611 6478 -577
rect 6592 -611 6626 -577
rect 6844 -611 6878 -577
rect 6992 -611 7026 -577
rect 7244 -611 7278 -577
rect 7392 -611 7426 -577
rect 7644 -611 7678 -577
rect 7792 -611 7826 -577
rect 8044 -611 8078 -577
rect 8192 -611 8226 -577
rect 8444 -611 8478 -577
rect 8592 -611 8626 -577
rect 8844 -611 8878 -577
rect 8992 -611 9026 -577
rect 9244 -611 9278 -577
rect 9392 -611 9426 -577
rect 9644 -611 9678 -577
rect 9792 -611 9826 -577
rect 10044 -611 10078 -577
rect 10192 -611 10226 -577
rect 10444 -611 10478 -577
rect 10592 -611 10626 -577
rect 10844 -611 10878 -577
rect 10992 -611 11026 -577
rect 11244 -611 11278 -577
rect 11392 -611 11426 -577
rect 11644 -611 11678 -577
rect 11792 -611 11826 -577
rect 12044 -611 12078 -577
rect 12192 -611 12226 -577
rect 12444 -611 12478 -577
rect 12592 -611 12626 -577
rect 14734 -743 14768 -709
rect 15574 -743 15608 -709
rect -82 -942 -48 -908
rect -82 -1042 -48 -1008
rect 718 -942 752 -908
rect -82 -1142 -48 -1108
rect 718 -1042 752 -1008
rect 1518 -942 1552 -908
rect -82 -1242 -48 -1208
rect 718 -1142 752 -1108
rect 1518 -1042 1552 -1008
rect 2318 -942 2352 -908
rect -82 -1342 -48 -1308
rect 718 -1242 752 -1208
rect 1518 -1142 1552 -1108
rect 2318 -1042 2352 -1008
rect 3118 -942 3152 -908
rect -82 -1442 -48 -1408
rect 718 -1342 752 -1308
rect 1518 -1242 1552 -1208
rect 2318 -1142 2352 -1108
rect 3118 -1042 3152 -1008
rect 3918 -942 3952 -908
rect -82 -1542 -48 -1508
rect 718 -1442 752 -1408
rect 1518 -1342 1552 -1308
rect 2318 -1242 2352 -1208
rect 3118 -1142 3152 -1108
rect 3918 -1042 3952 -1008
rect 4718 -942 4752 -908
rect -82 -1642 -48 -1608
rect 718 -1542 752 -1508
rect 1518 -1442 1552 -1408
rect 2318 -1342 2352 -1308
rect 3118 -1242 3152 -1208
rect 3918 -1142 3952 -1108
rect 4718 -1042 4752 -1008
rect 5518 -942 5552 -908
rect -82 -1742 -48 -1708
rect 718 -1642 752 -1608
rect 1518 -1542 1552 -1508
rect 2318 -1442 2352 -1408
rect 3118 -1342 3152 -1308
rect 3918 -1242 3952 -1208
rect 4718 -1142 4752 -1108
rect 5518 -1042 5552 -1008
rect 6318 -942 6352 -908
rect -82 -1842 -48 -1808
rect 718 -1742 752 -1708
rect 1518 -1642 1552 -1608
rect 2318 -1542 2352 -1508
rect 3118 -1442 3152 -1408
rect 3918 -1342 3952 -1308
rect 4718 -1242 4752 -1208
rect 5518 -1142 5552 -1108
rect 6318 -1042 6352 -1008
rect 7118 -942 7152 -908
rect -82 -1942 -48 -1908
rect 718 -1842 752 -1808
rect 1518 -1742 1552 -1708
rect 2318 -1642 2352 -1608
rect 3118 -1542 3152 -1508
rect 3918 -1442 3952 -1408
rect 4718 -1342 4752 -1308
rect 5518 -1242 5552 -1208
rect 6318 -1142 6352 -1108
rect 7118 -1042 7152 -1008
rect 7918 -942 7952 -908
rect -82 -2042 -48 -2008
rect 718 -1942 752 -1908
rect 1518 -1842 1552 -1808
rect 2318 -1742 2352 -1708
rect 3118 -1642 3152 -1608
rect 3918 -1542 3952 -1508
rect 4718 -1442 4752 -1408
rect 5518 -1342 5552 -1308
rect 6318 -1242 6352 -1208
rect 7118 -1142 7152 -1108
rect 7918 -1042 7952 -1008
rect 8718 -942 8752 -908
rect 718 -2042 752 -2008
rect 1518 -1942 1552 -1908
rect 2318 -1842 2352 -1808
rect 3118 -1742 3152 -1708
rect 3918 -1642 3952 -1608
rect 4718 -1542 4752 -1508
rect 5518 -1442 5552 -1408
rect 6318 -1342 6352 -1308
rect 7118 -1242 7152 -1208
rect 7918 -1142 7952 -1108
rect 8718 -1042 8752 -1008
rect 9518 -942 9552 -908
rect 1518 -2042 1552 -2008
rect 2318 -1942 2352 -1908
rect 3118 -1842 3152 -1808
rect 3918 -1742 3952 -1708
rect 4718 -1642 4752 -1608
rect 5518 -1542 5552 -1508
rect 6318 -1442 6352 -1408
rect 7118 -1342 7152 -1308
rect 7918 -1242 7952 -1208
rect 8718 -1142 8752 -1108
rect 9518 -1042 9552 -1008
rect 10318 -942 10352 -908
rect 2318 -2042 2352 -2008
rect 3118 -1942 3152 -1908
rect 3918 -1842 3952 -1808
rect 4718 -1742 4752 -1708
rect 5518 -1642 5552 -1608
rect 6318 -1542 6352 -1508
rect 7118 -1442 7152 -1408
rect 7918 -1342 7952 -1308
rect 8718 -1242 8752 -1208
rect 9518 -1142 9552 -1108
rect 10318 -1042 10352 -1008
rect 11118 -942 11152 -908
rect 3118 -2042 3152 -2008
rect 3918 -1942 3952 -1908
rect 4718 -1842 4752 -1808
rect 5518 -1742 5552 -1708
rect 6318 -1642 6352 -1608
rect 7118 -1542 7152 -1508
rect 7918 -1442 7952 -1408
rect 8718 -1342 8752 -1308
rect 9518 -1242 9552 -1208
rect 10318 -1142 10352 -1108
rect 11118 -1042 11152 -1008
rect 11918 -942 11952 -908
rect 3918 -2042 3952 -2008
rect 4718 -1942 4752 -1908
rect 5518 -1842 5552 -1808
rect 6318 -1742 6352 -1708
rect 7118 -1642 7152 -1608
rect 7918 -1542 7952 -1508
rect 8718 -1442 8752 -1408
rect 9518 -1342 9552 -1308
rect 10318 -1242 10352 -1208
rect 11118 -1142 11152 -1108
rect 11918 -1042 11952 -1008
rect 12718 -942 12752 -908
rect 14734 -943 14768 -909
rect 15574 -943 15608 -909
rect 4718 -2042 4752 -2008
rect 5518 -1942 5552 -1908
rect 6318 -1842 6352 -1808
rect 7118 -1742 7152 -1708
rect 7918 -1642 7952 -1608
rect 8718 -1542 8752 -1508
rect 9518 -1442 9552 -1408
rect 10318 -1342 10352 -1308
rect 11118 -1242 11152 -1208
rect 11918 -1142 11952 -1108
rect 12718 -1042 12752 -1008
rect 5518 -2042 5552 -2008
rect 6318 -1942 6352 -1908
rect 7118 -1842 7152 -1808
rect 7918 -1742 7952 -1708
rect 8718 -1642 8752 -1608
rect 9518 -1542 9552 -1508
rect 10318 -1442 10352 -1408
rect 11118 -1342 11152 -1308
rect 11918 -1242 11952 -1208
rect 12718 -1142 12752 -1108
rect 14734 -1143 14768 -1109
rect 15574 -1143 15608 -1109
rect 6318 -2042 6352 -2008
rect 7118 -1942 7152 -1908
rect 7918 -1842 7952 -1808
rect 8718 -1742 8752 -1708
rect 9518 -1642 9552 -1608
rect 10318 -1542 10352 -1508
rect 11118 -1442 11152 -1408
rect 11918 -1342 11952 -1308
rect 12718 -1242 12752 -1208
rect 7118 -2042 7152 -2008
rect 7918 -1942 7952 -1908
rect 8718 -1842 8752 -1808
rect 9518 -1742 9552 -1708
rect 10318 -1642 10352 -1608
rect 11118 -1542 11152 -1508
rect 11918 -1442 11952 -1408
rect 12718 -1342 12752 -1308
rect 14734 -1343 14768 -1309
rect 15574 -1343 15608 -1309
rect 7918 -2042 7952 -2008
rect 8718 -1942 8752 -1908
rect 9518 -1842 9552 -1808
rect 10318 -1742 10352 -1708
rect 11118 -1642 11152 -1608
rect 11918 -1542 11952 -1508
rect 12718 -1442 12752 -1408
rect 8718 -2042 8752 -2008
rect 9518 -1942 9552 -1908
rect 10318 -1842 10352 -1808
rect 11118 -1742 11152 -1708
rect 11918 -1642 11952 -1608
rect 12718 -1542 12752 -1508
rect 14734 -1543 14768 -1509
rect 15574 -1543 15608 -1509
rect 9518 -2042 9552 -2008
rect 10318 -1942 10352 -1908
rect 11118 -1842 11152 -1808
rect 11918 -1742 11952 -1708
rect 12718 -1642 12752 -1608
rect 10318 -2042 10352 -2008
rect 11118 -1942 11152 -1908
rect 11918 -1842 11952 -1808
rect 12718 -1742 12752 -1708
rect 14734 -1743 14768 -1709
rect 15574 -1743 15608 -1709
rect 11118 -2042 11152 -2008
rect 11918 -1942 11952 -1908
rect 12718 -1842 12752 -1808
rect 11918 -2042 11952 -2008
rect 12718 -1942 12752 -1908
rect 14734 -1943 14768 -1909
rect 15574 -1943 15608 -1909
rect 12718 -2042 12752 -2008
<< locali >>
rect 106 5017 164 5043
rect 106 4983 118 5017
rect 152 4983 164 5017
rect 106 4957 164 4983
rect 306 5017 364 5043
rect 306 4983 318 5017
rect 352 4983 364 5017
rect 306 4957 364 4983
rect 506 5017 564 5043
rect 506 4983 518 5017
rect 552 4983 564 5017
rect 506 4957 564 4983
rect 706 5017 764 5043
rect 706 4983 718 5017
rect 752 4983 764 5017
rect 706 4957 764 4983
rect 906 5017 964 5043
rect 906 4983 918 5017
rect 952 4983 964 5017
rect 906 4957 964 4983
rect 1106 5017 1164 5043
rect 1106 4983 1118 5017
rect 1152 4983 1164 5017
rect 1106 4957 1164 4983
rect 1306 5017 1364 5043
rect 1306 4983 1318 5017
rect 1352 4983 1364 5017
rect 1306 4957 1364 4983
rect 1506 5017 1564 5043
rect 1506 4983 1518 5017
rect 1552 4983 1564 5017
rect 1506 4957 1564 4983
rect 1706 5017 1764 5043
rect 1706 4983 1718 5017
rect 1752 4983 1764 5017
rect 1706 4957 1764 4983
rect 1906 5017 1964 5043
rect 1906 4983 1918 5017
rect 1952 4983 1964 5017
rect 1906 4957 1964 4983
rect 2106 5017 2164 5043
rect 2106 4983 2118 5017
rect 2152 4983 2164 5017
rect 2106 4957 2164 4983
rect 2306 5017 2364 5043
rect 2306 4983 2318 5017
rect 2352 4983 2364 5017
rect 2306 4957 2364 4983
rect 2506 5017 2564 5043
rect 2506 4983 2518 5017
rect 2552 4983 2564 5017
rect 2506 4957 2564 4983
rect 2706 5017 2764 5043
rect 2706 4983 2718 5017
rect 2752 4983 2764 5017
rect 2706 4957 2764 4983
rect 2906 5017 2964 5043
rect 2906 4983 2918 5017
rect 2952 4983 2964 5017
rect 2906 4957 2964 4983
rect 3106 5017 3164 5043
rect 3106 4983 3118 5017
rect 3152 4983 3164 5017
rect 3106 4957 3164 4983
rect 3306 5017 3364 5043
rect 3306 4983 3318 5017
rect 3352 4983 3364 5017
rect 3306 4957 3364 4983
rect 3506 5017 3564 5043
rect 3506 4983 3518 5017
rect 3552 4983 3564 5017
rect 3506 4957 3564 4983
rect 3706 5017 3764 5043
rect 3706 4983 3718 5017
rect 3752 4983 3764 5017
rect 3706 4957 3764 4983
rect 3906 5017 3964 5043
rect 3906 4983 3918 5017
rect 3952 4983 3964 5017
rect 3906 4957 3964 4983
rect 4106 5017 4164 5043
rect 4106 4983 4118 5017
rect 4152 4983 4164 5017
rect 4106 4957 4164 4983
rect 4306 5017 4364 5043
rect 4306 4983 4318 5017
rect 4352 4983 4364 5017
rect 4306 4957 4364 4983
rect 4506 5017 4564 5043
rect 4506 4983 4518 5017
rect 4552 4983 4564 5017
rect 4506 4957 4564 4983
rect 4706 5017 4764 5043
rect 4706 4983 4718 5017
rect 4752 4983 4764 5017
rect 4706 4957 4764 4983
rect 4906 5017 4964 5043
rect 4906 4983 4918 5017
rect 4952 4983 4964 5017
rect 4906 4957 4964 4983
rect 5106 5017 5164 5043
rect 5106 4983 5118 5017
rect 5152 4983 5164 5017
rect 5106 4957 5164 4983
rect 5306 5017 5364 5043
rect 5306 4983 5318 5017
rect 5352 4983 5364 5017
rect 5306 4957 5364 4983
rect 5506 5017 5564 5043
rect 5506 4983 5518 5017
rect 5552 4983 5564 5017
rect 5506 4957 5564 4983
rect 5706 5017 5764 5043
rect 5706 4983 5718 5017
rect 5752 4983 5764 5017
rect 5706 4957 5764 4983
rect 5906 5017 5964 5043
rect 5906 4983 5918 5017
rect 5952 4983 5964 5017
rect 5906 4957 5964 4983
rect 6106 5017 6164 5043
rect 6106 4983 6118 5017
rect 6152 4983 6164 5017
rect 6106 4957 6164 4983
rect 6306 5017 6364 5043
rect 6306 4983 6318 5017
rect 6352 4983 6364 5017
rect 6306 4957 6364 4983
rect 6506 5017 6564 5043
rect 6506 4983 6518 5017
rect 6552 4983 6564 5017
rect 6506 4957 6564 4983
rect 6706 5017 6764 5043
rect 6706 4983 6718 5017
rect 6752 4983 6764 5017
rect 6706 4957 6764 4983
rect 6906 5017 6964 5043
rect 6906 4983 6918 5017
rect 6952 4983 6964 5017
rect 6906 4957 6964 4983
rect 7106 5017 7164 5043
rect 7106 4983 7118 5017
rect 7152 4983 7164 5017
rect 7106 4957 7164 4983
rect 7306 5017 7364 5043
rect 7306 4983 7318 5017
rect 7352 4983 7364 5017
rect 7306 4957 7364 4983
rect 7506 5017 7564 5043
rect 7506 4983 7518 5017
rect 7552 4983 7564 5017
rect 7506 4957 7564 4983
rect 7706 5017 7764 5043
rect 7706 4983 7718 5017
rect 7752 4983 7764 5017
rect 7706 4957 7764 4983
rect 7906 5017 7964 5043
rect 7906 4983 7918 5017
rect 7952 4983 7964 5017
rect 7906 4957 7964 4983
rect 8106 5017 8164 5043
rect 8106 4983 8118 5017
rect 8152 4983 8164 5017
rect 8106 4957 8164 4983
rect 8306 5017 8364 5043
rect 8306 4983 8318 5017
rect 8352 4983 8364 5017
rect 8306 4957 8364 4983
rect 8506 5017 8564 5043
rect 8506 4983 8518 5017
rect 8552 4983 8564 5017
rect 8506 4957 8564 4983
rect 8706 5017 8764 5043
rect 8706 4983 8718 5017
rect 8752 4983 8764 5017
rect 8706 4957 8764 4983
rect 8906 5017 8964 5043
rect 8906 4983 8918 5017
rect 8952 4983 8964 5017
rect 8906 4957 8964 4983
rect 9106 5017 9164 5043
rect 9106 4983 9118 5017
rect 9152 4983 9164 5017
rect 9106 4957 9164 4983
rect 9306 5017 9364 5043
rect 9306 4983 9318 5017
rect 9352 4983 9364 5017
rect 9306 4957 9364 4983
rect 9506 5017 9564 5043
rect 9506 4983 9518 5017
rect 9552 4983 9564 5017
rect 9506 4957 9564 4983
rect 9706 5017 9764 5043
rect 9706 4983 9718 5017
rect 9752 4983 9764 5017
rect 9706 4957 9764 4983
rect 9906 5017 9964 5043
rect 9906 4983 9918 5017
rect 9952 4983 9964 5017
rect 9906 4957 9964 4983
rect 10106 5017 10164 5043
rect 10106 4983 10118 5017
rect 10152 4983 10164 5017
rect 10106 4957 10164 4983
rect 10306 5017 10364 5043
rect 10306 4983 10318 5017
rect 10352 4983 10364 5017
rect 10306 4957 10364 4983
rect 10506 5017 10564 5043
rect 10506 4983 10518 5017
rect 10552 4983 10564 5017
rect 10506 4957 10564 4983
rect 10706 5017 10764 5043
rect 10706 4983 10718 5017
rect 10752 4983 10764 5017
rect 10706 4957 10764 4983
rect 10906 5017 10964 5043
rect 10906 4983 10918 5017
rect 10952 4983 10964 5017
rect 10906 4957 10964 4983
rect 11106 5017 11164 5043
rect 11106 4983 11118 5017
rect 11152 4983 11164 5017
rect 11106 4957 11164 4983
rect 11306 5017 11364 5043
rect 11306 4983 11318 5017
rect 11352 4983 11364 5017
rect 11306 4957 11364 4983
rect 11506 5017 11564 5043
rect 11506 4983 11518 5017
rect 11552 4983 11564 5017
rect 11506 4957 11564 4983
rect 11706 5017 11764 5043
rect 11706 4983 11718 5017
rect 11752 4983 11764 5017
rect 11706 4957 11764 4983
rect 11906 5017 11964 5043
rect 11906 4983 11918 5017
rect 11952 4983 11964 5017
rect 11906 4957 11964 4983
rect 12106 5017 12164 5043
rect 12106 4983 12118 5017
rect 12152 4983 12164 5017
rect 12106 4957 12164 4983
rect 12306 5017 12364 5043
rect 12306 4983 12318 5017
rect 12352 4983 12364 5017
rect 12306 4957 12364 4983
rect 12506 5017 12564 5043
rect 12506 4983 12518 5017
rect 12552 4983 12564 5017
rect 12506 4957 12564 4983
rect 12706 5017 12764 5043
rect 12706 4983 12718 5017
rect 12752 4983 12764 5017
rect 12706 4957 12764 4983
rect 8 4860 18 4894
rect 52 4860 118 4894
rect 152 4860 168 4894
rect 208 4876 218 4910
rect 252 4876 318 4910
rect 352 4876 368 4910
rect 408 4860 418 4894
rect 452 4860 518 4894
rect 552 4860 568 4894
rect 608 4876 618 4910
rect 652 4876 718 4910
rect 752 4876 768 4910
rect 808 4860 818 4894
rect 852 4860 918 4894
rect 952 4860 968 4894
rect 1008 4876 1018 4910
rect 1052 4876 1118 4910
rect 1152 4876 1168 4910
rect 1208 4860 1218 4894
rect 1252 4860 1318 4894
rect 1352 4860 1368 4894
rect 1408 4876 1418 4910
rect 1452 4876 1518 4910
rect 1552 4876 1568 4910
rect 1608 4860 1618 4894
rect 1652 4860 1718 4894
rect 1752 4860 1768 4894
rect 1808 4876 1818 4910
rect 1852 4876 1918 4910
rect 1952 4876 1968 4910
rect 2008 4860 2018 4894
rect 2052 4860 2118 4894
rect 2152 4860 2168 4894
rect 2208 4876 2218 4910
rect 2252 4876 2318 4910
rect 2352 4876 2368 4910
rect 2408 4860 2418 4894
rect 2452 4860 2518 4894
rect 2552 4860 2568 4894
rect 2608 4876 2618 4910
rect 2652 4876 2718 4910
rect 2752 4876 2768 4910
rect 2808 4860 2818 4894
rect 2852 4860 2918 4894
rect 2952 4860 2968 4894
rect 3008 4876 3018 4910
rect 3052 4876 3118 4910
rect 3152 4876 3168 4910
rect 3208 4860 3218 4894
rect 3252 4860 3318 4894
rect 3352 4860 3368 4894
rect 3408 4876 3418 4910
rect 3452 4876 3518 4910
rect 3552 4876 3568 4910
rect 3608 4860 3618 4894
rect 3652 4860 3718 4894
rect 3752 4860 3768 4894
rect 3808 4876 3818 4910
rect 3852 4876 3918 4910
rect 3952 4876 3968 4910
rect 4008 4860 4018 4894
rect 4052 4860 4118 4894
rect 4152 4860 4168 4894
rect 4208 4876 4218 4910
rect 4252 4876 4318 4910
rect 4352 4876 4368 4910
rect 4408 4860 4418 4894
rect 4452 4860 4518 4894
rect 4552 4860 4568 4894
rect 4608 4876 4618 4910
rect 4652 4876 4718 4910
rect 4752 4876 4768 4910
rect 4808 4860 4818 4894
rect 4852 4860 4918 4894
rect 4952 4860 4968 4894
rect 5008 4876 5018 4910
rect 5052 4876 5118 4910
rect 5152 4876 5168 4910
rect 5208 4860 5218 4894
rect 5252 4860 5318 4894
rect 5352 4860 5368 4894
rect 5408 4876 5418 4910
rect 5452 4876 5518 4910
rect 5552 4876 5568 4910
rect 5608 4860 5618 4894
rect 5652 4860 5718 4894
rect 5752 4860 5768 4894
rect 5808 4876 5818 4910
rect 5852 4876 5918 4910
rect 5952 4876 5968 4910
rect 6008 4860 6018 4894
rect 6052 4860 6118 4894
rect 6152 4860 6168 4894
rect 6208 4876 6218 4910
rect 6252 4876 6318 4910
rect 6352 4876 6368 4910
rect 6408 4860 6418 4894
rect 6452 4860 6518 4894
rect 6552 4860 6568 4894
rect 6608 4876 6618 4910
rect 6652 4876 6718 4910
rect 6752 4876 6768 4910
rect 6808 4860 6818 4894
rect 6852 4860 6918 4894
rect 6952 4860 6968 4894
rect 7008 4876 7018 4910
rect 7052 4876 7118 4910
rect 7152 4876 7168 4910
rect 7208 4860 7218 4894
rect 7252 4860 7318 4894
rect 7352 4860 7368 4894
rect 7408 4876 7418 4910
rect 7452 4876 7518 4910
rect 7552 4876 7568 4910
rect 7608 4860 7618 4894
rect 7652 4860 7718 4894
rect 7752 4860 7768 4894
rect 7808 4876 7818 4910
rect 7852 4876 7918 4910
rect 7952 4876 7968 4910
rect 8008 4860 8018 4894
rect 8052 4860 8118 4894
rect 8152 4860 8168 4894
rect 8208 4876 8218 4910
rect 8252 4876 8318 4910
rect 8352 4876 8368 4910
rect 8408 4860 8418 4894
rect 8452 4860 8518 4894
rect 8552 4860 8568 4894
rect 8608 4876 8618 4910
rect 8652 4876 8718 4910
rect 8752 4876 8768 4910
rect 8808 4860 8818 4894
rect 8852 4860 8918 4894
rect 8952 4860 8968 4894
rect 9008 4876 9018 4910
rect 9052 4876 9118 4910
rect 9152 4876 9168 4910
rect 9208 4860 9218 4894
rect 9252 4860 9318 4894
rect 9352 4860 9368 4894
rect 9408 4876 9418 4910
rect 9452 4876 9518 4910
rect 9552 4876 9568 4910
rect 9608 4860 9618 4894
rect 9652 4860 9718 4894
rect 9752 4860 9768 4894
rect 9808 4876 9818 4910
rect 9852 4876 9918 4910
rect 9952 4876 9968 4910
rect 10008 4860 10018 4894
rect 10052 4860 10118 4894
rect 10152 4860 10168 4894
rect 10208 4876 10218 4910
rect 10252 4876 10318 4910
rect 10352 4876 10368 4910
rect 10408 4860 10418 4894
rect 10452 4860 10518 4894
rect 10552 4860 10568 4894
rect 10608 4876 10618 4910
rect 10652 4876 10718 4910
rect 10752 4876 10768 4910
rect 10808 4860 10818 4894
rect 10852 4860 10918 4894
rect 10952 4860 10968 4894
rect 11008 4876 11018 4910
rect 11052 4876 11118 4910
rect 11152 4876 11168 4910
rect 11208 4860 11218 4894
rect 11252 4860 11318 4894
rect 11352 4860 11368 4894
rect 11408 4876 11418 4910
rect 11452 4876 11518 4910
rect 11552 4876 11568 4910
rect 11608 4860 11618 4894
rect 11652 4860 11718 4894
rect 11752 4860 11768 4894
rect 11808 4876 11818 4910
rect 11852 4876 11918 4910
rect 11952 4876 11968 4910
rect 12008 4860 12018 4894
rect 12052 4860 12118 4894
rect 12152 4860 12168 4894
rect 12208 4876 12218 4910
rect 12252 4876 12318 4910
rect 12352 4876 12368 4910
rect 12408 4860 12418 4894
rect 12452 4860 12518 4894
rect 12552 4860 12568 4894
rect 12608 4876 12618 4910
rect 12652 4876 12718 4910
rect 12752 4876 12768 4910
rect 12916 4891 12968 4908
rect 12950 4874 12968 4891
rect 13002 4874 13018 4908
rect 13052 4874 13068 4908
rect 13102 4879 13120 4908
rect 13102 4874 13154 4879
rect 13262 4874 13278 4908
rect 13312 4874 13328 4908
rect 13362 4874 13378 4908
rect 13412 4874 13428 4908
rect 13462 4874 13478 4908
rect 13512 4874 13528 4908
rect 13562 4874 13578 4908
rect 13612 4874 13628 4908
rect 6 4787 64 4813
rect 6 4753 18 4787
rect 58 4753 64 4787
rect 6 4727 64 4753
rect 106 4787 164 4813
rect 106 4753 118 4787
rect 152 4753 164 4787
rect 106 4727 164 4753
rect 206 4787 264 4813
rect 206 4753 218 4787
rect 252 4753 264 4787
rect 206 4727 264 4753
rect 306 4787 364 4813
rect 306 4753 312 4787
rect 352 4753 364 4787
rect 306 4727 364 4753
rect 406 4787 464 4813
rect 406 4753 418 4787
rect 458 4753 464 4787
rect 406 4727 464 4753
rect 506 4787 564 4813
rect 506 4753 518 4787
rect 552 4753 564 4787
rect 506 4727 564 4753
rect 606 4787 664 4813
rect 606 4753 618 4787
rect 652 4753 664 4787
rect 606 4727 664 4753
rect 706 4787 764 4813
rect 706 4753 718 4787
rect 752 4753 764 4787
rect 706 4727 764 4753
rect 806 4787 864 4813
rect 806 4753 818 4787
rect 852 4753 864 4787
rect 806 4727 864 4753
rect 906 4787 964 4813
rect 906 4753 918 4787
rect 952 4753 964 4787
rect 906 4727 964 4753
rect 1006 4787 1064 4813
rect 1006 4753 1018 4787
rect 1052 4753 1064 4787
rect 1006 4727 1064 4753
rect 1106 4787 1164 4813
rect 1106 4753 1112 4787
rect 1152 4753 1164 4787
rect 1106 4727 1164 4753
rect 1206 4787 1264 4813
rect 1206 4753 1218 4787
rect 1258 4753 1264 4787
rect 1206 4727 1264 4753
rect 1306 4787 1364 4813
rect 1306 4753 1318 4787
rect 1352 4753 1364 4787
rect 1306 4727 1364 4753
rect 1406 4787 1464 4813
rect 1406 4753 1418 4787
rect 1452 4753 1464 4787
rect 1406 4727 1464 4753
rect 1506 4787 1564 4813
rect 1506 4753 1518 4787
rect 1552 4753 1564 4787
rect 1506 4727 1564 4753
rect 1606 4787 1664 4813
rect 1606 4753 1618 4787
rect 1652 4753 1664 4787
rect 1606 4727 1664 4753
rect 1706 4787 1764 4813
rect 1706 4753 1718 4787
rect 1752 4753 1764 4787
rect 1706 4727 1764 4753
rect 1806 4787 1864 4813
rect 1806 4753 1818 4787
rect 1852 4753 1864 4787
rect 1806 4727 1864 4753
rect 1906 4787 1964 4813
rect 1906 4753 1918 4787
rect 1952 4753 1964 4787
rect 1906 4727 1964 4753
rect 2006 4787 2064 4813
rect 2006 4753 2018 4787
rect 2052 4753 2064 4787
rect 2006 4727 2064 4753
rect 2106 4787 2164 4813
rect 2106 4753 2118 4787
rect 2152 4753 2164 4787
rect 2106 4727 2164 4753
rect 2206 4787 2264 4813
rect 2206 4753 2218 4787
rect 2252 4753 2264 4787
rect 2206 4727 2264 4753
rect 2306 4787 2364 4813
rect 2306 4753 2312 4787
rect 2352 4753 2364 4787
rect 2306 4727 2364 4753
rect 2406 4787 2464 4813
rect 2406 4753 2418 4787
rect 2458 4753 2464 4787
rect 2406 4727 2464 4753
rect 2506 4787 2564 4813
rect 2506 4753 2518 4787
rect 2552 4753 2564 4787
rect 2506 4727 2564 4753
rect 2606 4787 2664 4813
rect 2606 4753 2618 4787
rect 2652 4753 2664 4787
rect 2606 4727 2664 4753
rect 2706 4787 2764 4813
rect 2706 4753 2718 4787
rect 2752 4753 2764 4787
rect 2706 4727 2764 4753
rect 2806 4787 2864 4813
rect 2806 4753 2818 4787
rect 2852 4753 2864 4787
rect 2806 4727 2864 4753
rect 2906 4787 2964 4813
rect 2906 4753 2918 4787
rect 2952 4753 2964 4787
rect 2906 4727 2964 4753
rect 3006 4787 3064 4813
rect 3006 4753 3018 4787
rect 3052 4753 3064 4787
rect 3006 4727 3064 4753
rect 3106 4787 3164 4813
rect 3106 4753 3112 4787
rect 3152 4753 3164 4787
rect 3106 4727 3164 4753
rect 3206 4787 3264 4813
rect 3206 4753 3218 4787
rect 3258 4753 3264 4787
rect 3206 4727 3264 4753
rect 3306 4787 3364 4813
rect 3306 4753 3318 4787
rect 3352 4753 3364 4787
rect 3306 4727 3364 4753
rect 3406 4787 3464 4813
rect 3406 4753 3412 4787
rect 3452 4753 3464 4787
rect 3406 4727 3464 4753
rect 3506 4787 3564 4813
rect 3506 4753 3518 4787
rect 3558 4753 3564 4787
rect 3506 4727 3564 4753
rect 3606 4787 3664 4813
rect 3606 4753 3618 4787
rect 3652 4753 3664 4787
rect 3606 4727 3664 4753
rect 3706 4787 3764 4813
rect 3706 4753 3718 4787
rect 3752 4753 3764 4787
rect 3706 4727 3764 4753
rect 3806 4787 3864 4813
rect 3806 4753 3818 4787
rect 3852 4753 3864 4787
rect 3806 4727 3864 4753
rect 3906 4787 3964 4813
rect 3906 4753 3918 4787
rect 3952 4753 3964 4787
rect 3906 4727 3964 4753
rect 4006 4787 4064 4813
rect 4006 4753 4018 4787
rect 4052 4753 4064 4787
rect 4006 4727 4064 4753
rect 4106 4787 4164 4813
rect 4106 4753 4118 4787
rect 4152 4753 4164 4787
rect 4106 4727 4164 4753
rect 4206 4787 4264 4813
rect 4206 4753 4212 4787
rect 4252 4753 4264 4787
rect 4206 4727 4264 4753
rect 4306 4787 4364 4813
rect 4306 4753 4318 4787
rect 4358 4753 4364 4787
rect 4306 4727 4364 4753
rect 4406 4787 4464 4813
rect 4406 4753 4418 4787
rect 4452 4753 4464 4787
rect 4406 4727 4464 4753
rect 4506 4787 4564 4813
rect 4506 4753 4518 4787
rect 4552 4753 4564 4787
rect 4506 4727 4564 4753
rect 4606 4787 4664 4813
rect 4606 4753 4618 4787
rect 4652 4753 4664 4787
rect 4606 4727 4664 4753
rect 4706 4787 4764 4813
rect 4706 4753 4718 4787
rect 4752 4753 4764 4787
rect 4706 4727 4764 4753
rect 4806 4787 4864 4813
rect 4806 4753 4818 4787
rect 4852 4753 4864 4787
rect 4806 4727 4864 4753
rect 4906 4787 4964 4813
rect 4906 4753 4918 4787
rect 4952 4753 4964 4787
rect 4906 4727 4964 4753
rect 5006 4787 5064 4813
rect 5006 4753 5018 4787
rect 5052 4753 5064 4787
rect 5006 4727 5064 4753
rect 5106 4787 5164 4813
rect 5106 4753 5118 4787
rect 5152 4753 5164 4787
rect 5106 4727 5164 4753
rect 5206 4787 5264 4813
rect 5206 4753 5218 4787
rect 5252 4753 5264 4787
rect 5206 4727 5264 4753
rect 5306 4787 5364 4813
rect 5306 4753 5318 4787
rect 5352 4753 5364 4787
rect 5306 4727 5364 4753
rect 5406 4787 5464 4813
rect 5406 4753 5418 4787
rect 5452 4753 5464 4787
rect 5406 4727 5464 4753
rect 5506 4787 5564 4813
rect 5506 4753 5518 4787
rect 5552 4753 5564 4787
rect 5506 4727 5564 4753
rect 5606 4787 5664 4813
rect 5606 4753 5618 4787
rect 5652 4753 5664 4787
rect 5606 4727 5664 4753
rect 5706 4787 5764 4813
rect 5706 4753 5718 4787
rect 5752 4753 5764 4787
rect 5706 4727 5764 4753
rect 5806 4787 5864 4813
rect 5806 4753 5818 4787
rect 5852 4753 5864 4787
rect 5806 4727 5864 4753
rect 5906 4787 5964 4813
rect 5906 4753 5918 4787
rect 5952 4753 5964 4787
rect 5906 4727 5964 4753
rect 6006 4787 6064 4813
rect 6006 4753 6018 4787
rect 6052 4753 6064 4787
rect 6006 4727 6064 4753
rect 6106 4787 6164 4813
rect 6106 4753 6118 4787
rect 6152 4753 6164 4787
rect 6106 4727 6164 4753
rect 6206 4787 6264 4813
rect 6206 4753 6218 4787
rect 6252 4753 6264 4787
rect 6206 4727 6264 4753
rect 6306 4787 6364 4813
rect 6306 4753 6318 4787
rect 6352 4753 6364 4787
rect 6306 4727 6364 4753
rect 6406 4787 6464 4813
rect 6406 4753 6412 4787
rect 6452 4753 6464 4787
rect 6406 4727 6464 4753
rect 6506 4787 6564 4813
rect 6506 4753 6518 4787
rect 6558 4753 6564 4787
rect 6506 4727 6564 4753
rect 6606 4787 6664 4813
rect 6606 4753 6618 4787
rect 6652 4753 6664 4787
rect 6606 4727 6664 4753
rect 6706 4787 6764 4813
rect 6706 4753 6718 4787
rect 6752 4753 6764 4787
rect 6706 4727 6764 4753
rect 6806 4787 6864 4813
rect 6806 4753 6818 4787
rect 6852 4753 6864 4787
rect 6806 4727 6864 4753
rect 6906 4787 6964 4813
rect 6906 4753 6918 4787
rect 6952 4753 6964 4787
rect 6906 4727 6964 4753
rect 7006 4787 7064 4813
rect 7006 4753 7018 4787
rect 7052 4753 7064 4787
rect 7006 4727 7064 4753
rect 7106 4787 7164 4813
rect 7106 4753 7118 4787
rect 7152 4753 7164 4787
rect 7106 4727 7164 4753
rect 7206 4787 7264 4813
rect 7206 4753 7218 4787
rect 7252 4753 7264 4787
rect 7206 4727 7264 4753
rect 7306 4787 7364 4813
rect 7306 4753 7318 4787
rect 7352 4753 7364 4787
rect 7306 4727 7364 4753
rect 7406 4787 7464 4813
rect 7406 4753 7418 4787
rect 7452 4753 7464 4787
rect 7406 4727 7464 4753
rect 7506 4787 7564 4813
rect 7506 4753 7518 4787
rect 7552 4753 7564 4787
rect 7506 4727 7564 4753
rect 7606 4787 7664 4813
rect 7606 4753 7618 4787
rect 7652 4753 7664 4787
rect 7606 4727 7664 4753
rect 7706 4787 7764 4813
rect 7706 4753 7718 4787
rect 7752 4753 7764 4787
rect 7706 4727 7764 4753
rect 7806 4787 7864 4813
rect 7806 4753 7818 4787
rect 7852 4753 7864 4787
rect 7806 4727 7864 4753
rect 7906 4787 7964 4813
rect 7906 4753 7918 4787
rect 7952 4753 7964 4787
rect 7906 4727 7964 4753
rect 8006 4787 8064 4813
rect 8006 4753 8018 4787
rect 8052 4753 8064 4787
rect 8006 4727 8064 4753
rect 8106 4787 8164 4813
rect 8106 4753 8118 4787
rect 8152 4753 8164 4787
rect 8106 4727 8164 4753
rect 8206 4787 8264 4813
rect 8206 4753 8218 4787
rect 8252 4753 8264 4787
rect 8206 4727 8264 4753
rect 8306 4787 8364 4813
rect 8306 4753 8318 4787
rect 8352 4753 8364 4787
rect 8306 4727 8364 4753
rect 8406 4787 8464 4813
rect 8406 4753 8418 4787
rect 8452 4753 8464 4787
rect 8406 4727 8464 4753
rect 8506 4787 8564 4813
rect 8506 4753 8518 4787
rect 8552 4753 8564 4787
rect 8506 4727 8564 4753
rect 8606 4787 8664 4813
rect 8606 4753 8618 4787
rect 8652 4753 8664 4787
rect 8606 4727 8664 4753
rect 8706 4787 8764 4813
rect 8706 4753 8718 4787
rect 8752 4753 8764 4787
rect 8706 4727 8764 4753
rect 8806 4787 8864 4813
rect 8806 4753 8818 4787
rect 8852 4753 8864 4787
rect 8806 4727 8864 4753
rect 8906 4787 8964 4813
rect 8906 4753 8918 4787
rect 8952 4753 8964 4787
rect 8906 4727 8964 4753
rect 9006 4787 9064 4813
rect 9006 4753 9018 4787
rect 9052 4753 9064 4787
rect 9006 4727 9064 4753
rect 9106 4787 9164 4813
rect 9106 4753 9118 4787
rect 9152 4753 9164 4787
rect 9106 4727 9164 4753
rect 9206 4787 9264 4813
rect 9206 4753 9218 4787
rect 9252 4753 9264 4787
rect 9206 4727 9264 4753
rect 9306 4787 9364 4813
rect 9306 4753 9318 4787
rect 9352 4753 9364 4787
rect 9306 4727 9364 4753
rect 9406 4787 9464 4813
rect 9406 4753 9418 4787
rect 9452 4753 9464 4787
rect 9406 4727 9464 4753
rect 9506 4787 9564 4813
rect 9506 4753 9518 4787
rect 9552 4753 9564 4787
rect 9506 4727 9564 4753
rect 9606 4787 9664 4813
rect 9606 4753 9618 4787
rect 9652 4753 9664 4787
rect 9606 4727 9664 4753
rect 9706 4787 9764 4813
rect 9706 4753 9718 4787
rect 9752 4753 9764 4787
rect 9706 4727 9764 4753
rect 9806 4787 9864 4813
rect 9806 4753 9812 4787
rect 9852 4753 9864 4787
rect 9806 4727 9864 4753
rect 9906 4787 9964 4813
rect 9906 4753 9918 4787
rect 9958 4753 9964 4787
rect 9906 4727 9964 4753
rect 10006 4787 10064 4813
rect 10006 4753 10018 4787
rect 10052 4753 10064 4787
rect 10006 4727 10064 4753
rect 10106 4787 10164 4813
rect 10106 4753 10118 4787
rect 10152 4753 10164 4787
rect 10106 4727 10164 4753
rect 10206 4787 10264 4813
rect 10206 4753 10218 4787
rect 10252 4753 10264 4787
rect 10206 4727 10264 4753
rect 10306 4787 10364 4813
rect 10306 4753 10318 4787
rect 10352 4753 10364 4787
rect 10306 4727 10364 4753
rect 10406 4787 10464 4813
rect 10406 4753 10418 4787
rect 10452 4753 10464 4787
rect 10406 4727 10464 4753
rect 10506 4787 10564 4813
rect 10506 4753 10518 4787
rect 10552 4753 10564 4787
rect 10506 4727 10564 4753
rect 10606 4787 10664 4813
rect 10606 4753 10618 4787
rect 10652 4753 10664 4787
rect 10606 4727 10664 4753
rect 10706 4787 10764 4813
rect 10706 4753 10712 4787
rect 10752 4753 10764 4787
rect 10706 4727 10764 4753
rect 10806 4787 10864 4813
rect 10806 4753 10818 4787
rect 10858 4753 10864 4787
rect 10806 4727 10864 4753
rect 10906 4787 10964 4813
rect 10906 4753 10918 4787
rect 10952 4753 10964 4787
rect 10906 4727 10964 4753
rect 11006 4787 11064 4813
rect 11006 4753 11018 4787
rect 11052 4753 11064 4787
rect 11006 4727 11064 4753
rect 11106 4787 11164 4813
rect 11106 4753 11118 4787
rect 11152 4753 11164 4787
rect 11106 4727 11164 4753
rect 11206 4787 11264 4813
rect 11206 4753 11218 4787
rect 11252 4753 11264 4787
rect 11206 4727 11264 4753
rect 11306 4787 11364 4813
rect 11306 4753 11318 4787
rect 11352 4753 11364 4787
rect 11306 4727 11364 4753
rect 11406 4787 11464 4813
rect 11406 4753 11418 4787
rect 11452 4753 11464 4787
rect 11406 4727 11464 4753
rect 11506 4787 11564 4813
rect 11506 4753 11518 4787
rect 11552 4753 11564 4787
rect 11506 4727 11564 4753
rect 11606 4787 11664 4813
rect 11606 4753 11612 4787
rect 11652 4753 11664 4787
rect 11606 4727 11664 4753
rect 11706 4787 11764 4813
rect 11706 4753 11718 4787
rect 11758 4753 11764 4787
rect 11706 4727 11764 4753
rect 11806 4787 11864 4813
rect 11806 4753 11818 4787
rect 11852 4753 11864 4787
rect 11806 4727 11864 4753
rect 11906 4787 11964 4813
rect 11906 4753 11918 4787
rect 11952 4753 11964 4787
rect 11906 4727 11964 4753
rect 12006 4787 12064 4813
rect 12006 4753 12018 4787
rect 12052 4753 12064 4787
rect 12006 4727 12064 4753
rect 12106 4787 12164 4813
rect 12106 4753 12118 4787
rect 12152 4753 12164 4787
rect 12106 4727 12164 4753
rect 12206 4787 12264 4813
rect 12206 4753 12218 4787
rect 12252 4753 12264 4787
rect 12206 4727 12264 4753
rect 12306 4787 12364 4813
rect 12306 4753 12318 4787
rect 12352 4753 12364 4787
rect 12306 4727 12364 4753
rect 12406 4787 12464 4813
rect 12406 4753 12412 4787
rect 12452 4753 12464 4787
rect 12406 4727 12464 4753
rect 12506 4787 12564 4813
rect 12506 4753 12518 4787
rect 12558 4753 12564 4787
rect 12506 4727 12564 4753
rect 12606 4787 12664 4813
rect 12606 4753 12618 4787
rect 12652 4753 12664 4787
rect 12606 4727 12664 4753
rect 12706 4787 12764 4813
rect 12706 4753 12718 4787
rect 12752 4753 12764 4787
rect 12706 4727 12764 4753
rect 12806 4787 12864 4813
rect 13018 4806 13262 4840
rect 12806 4753 12812 4787
rect 12852 4753 12864 4787
rect 12908 4768 12916 4802
rect 12958 4768 12974 4802
rect 13018 4787 13052 4806
rect 12806 4727 12864 4753
rect 13228 4803 13262 4806
rect 13228 4787 13362 4803
rect 13018 4737 13052 4753
rect 13096 4738 13112 4772
rect 13154 4738 13162 4772
rect 13262 4753 13328 4787
rect 13228 4737 13362 4753
rect 13428 4787 13562 4803
rect 13462 4753 13528 4787
rect 13428 4737 13562 4753
rect 13628 4787 13662 4803
rect 13628 4737 13662 4753
rect 6 4647 64 4673
rect 6 4613 18 4647
rect 52 4613 64 4647
rect 6 4587 64 4613
rect 106 4647 164 4673
rect 106 4613 118 4647
rect 152 4613 164 4647
rect 106 4587 164 4613
rect 206 4647 264 4673
rect 206 4613 218 4647
rect 252 4613 264 4647
rect 206 4587 264 4613
rect 306 4647 364 4673
rect 306 4613 318 4647
rect 352 4613 364 4647
rect 306 4587 364 4613
rect 406 4647 464 4673
rect 406 4613 418 4647
rect 452 4613 464 4647
rect 406 4587 464 4613
rect 506 4647 564 4673
rect 506 4613 518 4647
rect 552 4613 564 4647
rect 506 4587 564 4613
rect 606 4647 664 4673
rect 606 4613 618 4647
rect 652 4613 664 4647
rect 606 4587 664 4613
rect 706 4647 764 4673
rect 706 4613 718 4647
rect 752 4613 764 4647
rect 706 4587 764 4613
rect 806 4647 864 4673
rect 806 4613 818 4647
rect 852 4613 864 4647
rect 806 4587 864 4613
rect 906 4647 964 4673
rect 906 4613 918 4647
rect 952 4613 964 4647
rect 906 4587 964 4613
rect 1006 4647 1064 4673
rect 1006 4613 1018 4647
rect 1052 4613 1064 4647
rect 1006 4587 1064 4613
rect 1106 4647 1164 4673
rect 1106 4613 1112 4647
rect 1152 4613 1164 4647
rect 1106 4587 1164 4613
rect 1206 4647 1264 4673
rect 1206 4613 1218 4647
rect 1258 4613 1264 4647
rect 1206 4587 1264 4613
rect 1306 4647 1364 4673
rect 1306 4613 1318 4647
rect 1352 4613 1364 4647
rect 1306 4587 1364 4613
rect 1406 4647 1464 4673
rect 1406 4613 1418 4647
rect 1452 4613 1464 4647
rect 1406 4587 1464 4613
rect 1506 4647 1564 4673
rect 1506 4613 1518 4647
rect 1552 4613 1564 4647
rect 1506 4587 1564 4613
rect 1606 4647 1664 4673
rect 1606 4613 1618 4647
rect 1652 4613 1664 4647
rect 1606 4587 1664 4613
rect 1706 4647 1764 4673
rect 1706 4613 1718 4647
rect 1752 4613 1764 4647
rect 1706 4587 1764 4613
rect 1806 4647 1864 4673
rect 1806 4613 1818 4647
rect 1852 4613 1864 4647
rect 1806 4587 1864 4613
rect 1906 4647 1964 4673
rect 1906 4613 1918 4647
rect 1952 4613 1964 4647
rect 1906 4587 1964 4613
rect 2006 4647 2064 4673
rect 2006 4613 2018 4647
rect 2052 4613 2064 4647
rect 2006 4587 2064 4613
rect 2106 4647 2164 4673
rect 2106 4613 2118 4647
rect 2152 4613 2164 4647
rect 2106 4587 2164 4613
rect 2206 4647 2264 4673
rect 2206 4613 2218 4647
rect 2252 4613 2264 4647
rect 2206 4587 2264 4613
rect 2306 4647 2364 4673
rect 2306 4613 2318 4647
rect 2352 4613 2364 4647
rect 2306 4587 2364 4613
rect 2406 4647 2464 4673
rect 2406 4613 2418 4647
rect 2452 4613 2464 4647
rect 2406 4587 2464 4613
rect 2506 4647 2564 4673
rect 2506 4613 2518 4647
rect 2552 4613 2564 4647
rect 2506 4587 2564 4613
rect 2606 4647 2664 4673
rect 2606 4613 2618 4647
rect 2652 4613 2664 4647
rect 2606 4587 2664 4613
rect 2706 4647 2764 4673
rect 2706 4613 2718 4647
rect 2752 4613 2764 4647
rect 2706 4587 2764 4613
rect 2806 4647 2864 4673
rect 2806 4613 2818 4647
rect 2852 4613 2864 4647
rect 2806 4587 2864 4613
rect 2906 4647 2964 4673
rect 2906 4613 2912 4647
rect 2952 4613 2964 4647
rect 2906 4587 2964 4613
rect 3006 4647 3064 4673
rect 3006 4613 3018 4647
rect 3058 4613 3064 4647
rect 3006 4587 3064 4613
rect 3106 4647 3164 4673
rect 3106 4613 3118 4647
rect 3152 4613 3164 4647
rect 3106 4587 3164 4613
rect 3206 4647 3264 4673
rect 3206 4613 3218 4647
rect 3252 4613 3264 4647
rect 3206 4587 3264 4613
rect 3306 4647 3364 4673
rect 3306 4613 3318 4647
rect 3352 4613 3364 4647
rect 3306 4587 3364 4613
rect 3406 4647 3464 4673
rect 3406 4613 3418 4647
rect 3452 4613 3464 4647
rect 3406 4587 3464 4613
rect 3506 4647 3564 4673
rect 3506 4613 3518 4647
rect 3552 4613 3564 4647
rect 3506 4587 3564 4613
rect 3606 4647 3664 4673
rect 3606 4613 3612 4647
rect 3652 4613 3664 4647
rect 3606 4587 3664 4613
rect 3706 4647 3764 4673
rect 3706 4613 3718 4647
rect 3758 4613 3764 4647
rect 3706 4587 3764 4613
rect 3806 4647 3864 4673
rect 3806 4613 3818 4647
rect 3852 4613 3864 4647
rect 3806 4587 3864 4613
rect 3906 4647 3964 4673
rect 3906 4613 3918 4647
rect 3952 4613 3964 4647
rect 3906 4587 3964 4613
rect 4006 4647 4064 4673
rect 4006 4613 4018 4647
rect 4052 4613 4064 4647
rect 4006 4587 4064 4613
rect 4106 4647 4164 4673
rect 4106 4613 4118 4647
rect 4152 4613 4164 4647
rect 4106 4587 4164 4613
rect 4206 4647 4264 4673
rect 4206 4613 4218 4647
rect 4252 4613 4264 4647
rect 4206 4587 4264 4613
rect 4306 4647 4364 4673
rect 4306 4613 4318 4647
rect 4352 4613 4364 4647
rect 4306 4587 4364 4613
rect 4406 4647 4464 4673
rect 4406 4613 4418 4647
rect 4452 4613 4464 4647
rect 4406 4587 4464 4613
rect 4506 4647 4564 4673
rect 4506 4613 4518 4647
rect 4552 4613 4564 4647
rect 4506 4587 4564 4613
rect 4606 4647 4664 4673
rect 4606 4613 4618 4647
rect 4652 4613 4664 4647
rect 4606 4587 4664 4613
rect 4706 4647 4764 4673
rect 4706 4613 4712 4647
rect 4752 4613 4764 4647
rect 4706 4587 4764 4613
rect 4806 4647 4864 4673
rect 4806 4613 4818 4647
rect 4858 4613 4864 4647
rect 4806 4587 4864 4613
rect 4906 4647 4964 4673
rect 4906 4613 4918 4647
rect 4952 4613 4964 4647
rect 4906 4587 4964 4613
rect 5006 4647 5064 4673
rect 5006 4613 5012 4647
rect 5052 4613 5064 4647
rect 5006 4587 5064 4613
rect 5106 4647 5164 4673
rect 5106 4613 5118 4647
rect 5158 4613 5164 4647
rect 5106 4587 5164 4613
rect 5206 4647 5264 4673
rect 5206 4613 5218 4647
rect 5252 4613 5264 4647
rect 5206 4587 5264 4613
rect 5306 4647 5364 4673
rect 5306 4613 5318 4647
rect 5352 4613 5364 4647
rect 5306 4587 5364 4613
rect 5406 4647 5464 4673
rect 5406 4613 5418 4647
rect 5452 4613 5464 4647
rect 5406 4587 5464 4613
rect 5506 4647 5564 4673
rect 5506 4613 5518 4647
rect 5552 4613 5564 4647
rect 5506 4587 5564 4613
rect 5606 4647 5664 4673
rect 5606 4613 5618 4647
rect 5652 4613 5664 4647
rect 5606 4587 5664 4613
rect 5706 4647 5764 4673
rect 5706 4613 5718 4647
rect 5752 4613 5764 4647
rect 5706 4587 5764 4613
rect 5806 4647 5864 4673
rect 5806 4613 5812 4647
rect 5852 4613 5864 4647
rect 5806 4587 5864 4613
rect 5906 4647 5964 4673
rect 5906 4613 5918 4647
rect 5958 4613 5964 4647
rect 5906 4587 5964 4613
rect 6006 4647 6064 4673
rect 6006 4613 6018 4647
rect 6052 4613 6064 4647
rect 6006 4587 6064 4613
rect 6106 4647 6164 4673
rect 6106 4613 6118 4647
rect 6152 4613 6164 4647
rect 6106 4587 6164 4613
rect 6206 4647 6264 4673
rect 6206 4613 6218 4647
rect 6252 4613 6264 4647
rect 6206 4587 6264 4613
rect 6306 4647 6364 4673
rect 6306 4613 6318 4647
rect 6352 4613 6364 4647
rect 6306 4587 6364 4613
rect 6406 4647 6464 4673
rect 6406 4613 6412 4647
rect 6452 4613 6464 4647
rect 6406 4587 6464 4613
rect 6506 4647 6564 4673
rect 6506 4613 6518 4647
rect 6558 4613 6564 4647
rect 6506 4587 6564 4613
rect 6606 4647 6664 4673
rect 6606 4613 6618 4647
rect 6652 4613 6664 4647
rect 6606 4587 6664 4613
rect 6706 4647 6764 4673
rect 6706 4613 6718 4647
rect 6752 4613 6764 4647
rect 6706 4587 6764 4613
rect 6806 4647 6864 4673
rect 6806 4613 6818 4647
rect 6852 4613 6864 4647
rect 6806 4587 6864 4613
rect 6906 4647 6964 4673
rect 6906 4613 6918 4647
rect 6952 4613 6964 4647
rect 6906 4587 6964 4613
rect 7006 4647 7064 4673
rect 7006 4613 7018 4647
rect 7052 4613 7064 4647
rect 7006 4587 7064 4613
rect 7106 4647 7164 4673
rect 7106 4613 7118 4647
rect 7152 4613 7164 4647
rect 7106 4587 7164 4613
rect 7206 4647 7264 4673
rect 7206 4613 7218 4647
rect 7252 4613 7264 4647
rect 7206 4587 7264 4613
rect 7306 4647 7364 4673
rect 7306 4613 7318 4647
rect 7352 4613 7364 4647
rect 7306 4587 7364 4613
rect 7406 4647 7464 4673
rect 7406 4613 7418 4647
rect 7452 4613 7464 4647
rect 7406 4587 7464 4613
rect 7506 4647 7564 4673
rect 7506 4613 7518 4647
rect 7552 4613 7564 4647
rect 7506 4587 7564 4613
rect 7606 4647 7664 4673
rect 7606 4613 7618 4647
rect 7652 4613 7664 4647
rect 7606 4587 7664 4613
rect 7706 4647 7764 4673
rect 7706 4613 7718 4647
rect 7752 4613 7764 4647
rect 7706 4587 7764 4613
rect 7806 4647 7864 4673
rect 7806 4613 7818 4647
rect 7852 4613 7864 4647
rect 7806 4587 7864 4613
rect 7906 4647 7964 4673
rect 7906 4613 7918 4647
rect 7952 4613 7964 4647
rect 7906 4587 7964 4613
rect 8006 4647 8064 4673
rect 8006 4613 8018 4647
rect 8052 4613 8064 4647
rect 8006 4587 8064 4613
rect 8106 4647 8164 4673
rect 8106 4613 8118 4647
rect 8152 4613 8164 4647
rect 8106 4587 8164 4613
rect 8206 4647 8264 4673
rect 8206 4613 8218 4647
rect 8252 4613 8264 4647
rect 8206 4587 8264 4613
rect 8306 4647 8364 4673
rect 8306 4613 8318 4647
rect 8352 4613 8364 4647
rect 8306 4587 8364 4613
rect 8406 4647 8464 4673
rect 8406 4613 8418 4647
rect 8452 4613 8464 4647
rect 8406 4587 8464 4613
rect 8506 4647 8564 4673
rect 8506 4613 8518 4647
rect 8552 4613 8564 4647
rect 8506 4587 8564 4613
rect 8606 4647 8664 4673
rect 8606 4613 8618 4647
rect 8652 4613 8664 4647
rect 8606 4587 8664 4613
rect 8706 4647 8764 4673
rect 8706 4613 8712 4647
rect 8752 4613 8764 4647
rect 8706 4587 8764 4613
rect 8806 4647 8864 4673
rect 8806 4613 8818 4647
rect 8858 4613 8864 4647
rect 8806 4587 8864 4613
rect 8906 4647 8964 4673
rect 8906 4613 8918 4647
rect 8952 4613 8964 4647
rect 8906 4587 8964 4613
rect 9006 4647 9064 4673
rect 9006 4613 9018 4647
rect 9052 4613 9064 4647
rect 9006 4587 9064 4613
rect 9106 4647 9164 4673
rect 9106 4613 9118 4647
rect 9152 4613 9164 4647
rect 9106 4587 9164 4613
rect 9206 4647 9264 4673
rect 9206 4613 9218 4647
rect 9252 4613 9264 4647
rect 9206 4587 9264 4613
rect 9306 4647 9364 4673
rect 9306 4613 9318 4647
rect 9352 4613 9364 4647
rect 9306 4587 9364 4613
rect 9406 4647 9464 4673
rect 9406 4613 9418 4647
rect 9452 4613 9464 4647
rect 9406 4587 9464 4613
rect 9506 4647 9564 4673
rect 9506 4613 9518 4647
rect 9552 4613 9564 4647
rect 9506 4587 9564 4613
rect 9606 4647 9664 4673
rect 9606 4613 9618 4647
rect 9652 4613 9664 4647
rect 9606 4587 9664 4613
rect 9706 4647 9764 4673
rect 9706 4613 9718 4647
rect 9752 4613 9764 4647
rect 9706 4587 9764 4613
rect 9806 4647 9864 4673
rect 9806 4613 9818 4647
rect 9852 4613 9864 4647
rect 9806 4587 9864 4613
rect 9906 4647 9964 4673
rect 9906 4613 9918 4647
rect 9952 4613 9964 4647
rect 9906 4587 9964 4613
rect 10006 4647 10064 4673
rect 10006 4613 10018 4647
rect 10052 4613 10064 4647
rect 10006 4587 10064 4613
rect 10106 4647 10164 4673
rect 10106 4613 10118 4647
rect 10152 4613 10164 4647
rect 10106 4587 10164 4613
rect 10206 4647 10264 4673
rect 10206 4613 10218 4647
rect 10252 4613 10264 4647
rect 10206 4587 10264 4613
rect 10306 4647 10364 4673
rect 10306 4613 10318 4647
rect 10352 4613 10364 4647
rect 10306 4587 10364 4613
rect 10406 4647 10464 4673
rect 10406 4613 10418 4647
rect 10452 4613 10464 4647
rect 10406 4587 10464 4613
rect 10506 4647 10564 4673
rect 10506 4613 10518 4647
rect 10552 4613 10564 4647
rect 10506 4587 10564 4613
rect 10606 4647 10664 4673
rect 10606 4613 10618 4647
rect 10652 4613 10664 4647
rect 10606 4587 10664 4613
rect 10706 4647 10764 4673
rect 10706 4613 10718 4647
rect 10752 4613 10764 4647
rect 10706 4587 10764 4613
rect 10806 4647 10864 4673
rect 10806 4613 10818 4647
rect 10852 4613 10864 4647
rect 10806 4587 10864 4613
rect 10906 4647 10964 4673
rect 10906 4613 10918 4647
rect 10952 4613 10964 4647
rect 10906 4587 10964 4613
rect 11006 4647 11064 4673
rect 11006 4613 11018 4647
rect 11052 4613 11064 4647
rect 11006 4587 11064 4613
rect 11106 4647 11164 4673
rect 11106 4613 11118 4647
rect 11152 4613 11164 4647
rect 11106 4587 11164 4613
rect 11206 4647 11264 4673
rect 11206 4613 11218 4647
rect 11252 4613 11264 4647
rect 11206 4587 11264 4613
rect 11306 4647 11364 4673
rect 11306 4613 11318 4647
rect 11352 4613 11364 4647
rect 11306 4587 11364 4613
rect 11406 4647 11464 4673
rect 11406 4613 11418 4647
rect 11452 4613 11464 4647
rect 11406 4587 11464 4613
rect 11506 4647 11564 4673
rect 11506 4613 11518 4647
rect 11552 4613 11564 4647
rect 11506 4587 11564 4613
rect 11606 4647 11664 4673
rect 11606 4613 11618 4647
rect 11652 4613 11664 4647
rect 11606 4587 11664 4613
rect 11706 4647 11764 4673
rect 11706 4613 11718 4647
rect 11752 4613 11764 4647
rect 11706 4587 11764 4613
rect 11806 4647 11864 4673
rect 11806 4613 11818 4647
rect 11852 4613 11864 4647
rect 11806 4587 11864 4613
rect 11906 4647 11964 4673
rect 11906 4613 11918 4647
rect 11952 4613 11964 4647
rect 11906 4587 11964 4613
rect 12006 4647 12064 4673
rect 12006 4613 12018 4647
rect 12052 4613 12064 4647
rect 12006 4587 12064 4613
rect 12106 4647 12164 4673
rect 12106 4613 12118 4647
rect 12152 4613 12164 4647
rect 12106 4587 12164 4613
rect 12206 4647 12264 4673
rect 12206 4613 12218 4647
rect 12252 4613 12264 4647
rect 12206 4587 12264 4613
rect 12306 4647 12364 4673
rect 12306 4613 12318 4647
rect 12352 4613 12364 4647
rect 12306 4587 12364 4613
rect 12406 4647 12464 4673
rect 12406 4613 12418 4647
rect 12452 4613 12464 4647
rect 12406 4587 12464 4613
rect 12506 4647 12564 4673
rect 12506 4613 12518 4647
rect 12552 4613 12564 4647
rect 12506 4587 12564 4613
rect 12606 4647 12664 4673
rect 12606 4613 12612 4647
rect 12652 4613 12664 4647
rect 12606 4587 12664 4613
rect 12706 4647 12764 4673
rect 12706 4613 12718 4647
rect 12758 4613 12764 4647
rect 12706 4587 12764 4613
rect 12806 4647 12864 4673
rect 13018 4666 13262 4700
rect 12806 4613 12812 4647
rect 12852 4613 12864 4647
rect 12908 4628 12916 4662
rect 12958 4628 12974 4662
rect 13018 4647 13052 4666
rect 12806 4587 12864 4613
rect 13228 4647 13262 4666
rect 13018 4597 13052 4613
rect 13096 4598 13112 4632
rect 13154 4598 13162 4632
rect 13228 4597 13262 4613
rect 13328 4647 13562 4663
rect 13362 4613 13428 4647
rect 13462 4613 13528 4647
rect 13328 4597 13562 4613
rect 13628 4647 13662 4663
rect 13628 4597 13662 4613
rect 6 4507 64 4533
rect 6 4473 18 4507
rect 52 4473 64 4507
rect 6 4447 64 4473
rect 106 4507 164 4533
rect 106 4473 118 4507
rect 152 4473 164 4507
rect 106 4447 164 4473
rect 206 4507 264 4533
rect 206 4473 218 4507
rect 252 4473 264 4507
rect 206 4447 264 4473
rect 306 4507 364 4533
rect 306 4473 312 4507
rect 352 4473 364 4507
rect 306 4447 364 4473
rect 406 4507 464 4533
rect 406 4473 418 4507
rect 458 4473 464 4507
rect 406 4447 464 4473
rect 506 4507 564 4533
rect 506 4473 518 4507
rect 552 4473 564 4507
rect 506 4447 564 4473
rect 606 4507 664 4533
rect 606 4473 618 4507
rect 652 4473 664 4507
rect 606 4447 664 4473
rect 706 4507 764 4533
rect 706 4473 718 4507
rect 752 4473 764 4507
rect 706 4447 764 4473
rect 806 4507 864 4533
rect 806 4473 818 4507
rect 852 4473 864 4507
rect 806 4447 864 4473
rect 906 4507 964 4533
rect 906 4473 918 4507
rect 952 4473 964 4507
rect 906 4447 964 4473
rect 1006 4507 1064 4533
rect 1006 4473 1018 4507
rect 1052 4473 1064 4507
rect 1006 4447 1064 4473
rect 1106 4507 1164 4533
rect 1106 4473 1118 4507
rect 1152 4473 1164 4507
rect 1106 4447 1164 4473
rect 1206 4507 1264 4533
rect 1206 4473 1218 4507
rect 1252 4473 1264 4507
rect 1206 4447 1264 4473
rect 1306 4507 1364 4533
rect 1306 4473 1318 4507
rect 1352 4473 1364 4507
rect 1306 4447 1364 4473
rect 1406 4507 1464 4533
rect 1406 4473 1418 4507
rect 1452 4473 1464 4507
rect 1406 4447 1464 4473
rect 1506 4507 1564 4533
rect 1506 4473 1518 4507
rect 1552 4473 1564 4507
rect 1506 4447 1564 4473
rect 1606 4507 1664 4533
rect 1606 4473 1612 4507
rect 1652 4473 1664 4507
rect 1606 4447 1664 4473
rect 1706 4507 1764 4533
rect 1706 4473 1718 4507
rect 1758 4473 1764 4507
rect 1706 4447 1764 4473
rect 1806 4507 1864 4533
rect 1806 4473 1812 4507
rect 1852 4473 1864 4507
rect 1806 4447 1864 4473
rect 1906 4507 1964 4533
rect 1906 4473 1918 4507
rect 1958 4473 1964 4507
rect 1906 4447 1964 4473
rect 2006 4507 2064 4533
rect 2006 4473 2018 4507
rect 2052 4473 2064 4507
rect 2006 4447 2064 4473
rect 2106 4507 2164 4533
rect 2106 4473 2118 4507
rect 2152 4473 2164 4507
rect 2106 4447 2164 4473
rect 2206 4507 2264 4533
rect 2206 4473 2218 4507
rect 2252 4473 2264 4507
rect 2206 4447 2264 4473
rect 2306 4507 2364 4533
rect 2306 4473 2312 4507
rect 2352 4473 2364 4507
rect 2306 4447 2364 4473
rect 2406 4507 2464 4533
rect 2406 4473 2418 4507
rect 2458 4473 2464 4507
rect 2406 4447 2464 4473
rect 2506 4507 2564 4533
rect 2506 4473 2518 4507
rect 2552 4473 2564 4507
rect 2506 4447 2564 4473
rect 2606 4507 2664 4533
rect 2606 4473 2612 4507
rect 2652 4473 2664 4507
rect 2606 4447 2664 4473
rect 2706 4507 2764 4533
rect 2706 4473 2718 4507
rect 2758 4473 2764 4507
rect 2706 4447 2764 4473
rect 2806 4507 2864 4533
rect 2806 4473 2812 4507
rect 2852 4473 2864 4507
rect 2806 4447 2864 4473
rect 2906 4507 2964 4533
rect 2906 4473 2918 4507
rect 2958 4473 2964 4507
rect 2906 4447 2964 4473
rect 3006 4507 3064 4533
rect 3006 4473 3018 4507
rect 3052 4473 3064 4507
rect 3006 4447 3064 4473
rect 3106 4507 3164 4533
rect 3106 4473 3118 4507
rect 3152 4473 3164 4507
rect 3106 4447 3164 4473
rect 3206 4507 3264 4533
rect 3206 4473 3218 4507
rect 3252 4473 3264 4507
rect 3206 4447 3264 4473
rect 3306 4507 3364 4533
rect 3306 4473 3318 4507
rect 3352 4473 3364 4507
rect 3306 4447 3364 4473
rect 3406 4507 3464 4533
rect 3406 4473 3418 4507
rect 3452 4473 3464 4507
rect 3406 4447 3464 4473
rect 3506 4507 3564 4533
rect 3506 4473 3518 4507
rect 3552 4473 3564 4507
rect 3506 4447 3564 4473
rect 3606 4507 3664 4533
rect 3606 4473 3618 4507
rect 3652 4473 3664 4507
rect 3606 4447 3664 4473
rect 3706 4507 3764 4533
rect 3706 4473 3712 4507
rect 3752 4473 3764 4507
rect 3706 4447 3764 4473
rect 3806 4507 3864 4533
rect 3806 4473 3818 4507
rect 3858 4473 3864 4507
rect 3806 4447 3864 4473
rect 3906 4507 3964 4533
rect 3906 4473 3918 4507
rect 3952 4473 3964 4507
rect 3906 4447 3964 4473
rect 4006 4507 4064 4533
rect 4006 4473 4018 4507
rect 4052 4473 4064 4507
rect 4006 4447 4064 4473
rect 4106 4507 4164 4533
rect 4106 4473 4118 4507
rect 4152 4473 4164 4507
rect 4106 4447 4164 4473
rect 4206 4507 4264 4533
rect 4206 4473 4218 4507
rect 4252 4473 4264 4507
rect 4206 4447 4264 4473
rect 4306 4507 4364 4533
rect 4306 4473 4318 4507
rect 4352 4473 4364 4507
rect 4306 4447 4364 4473
rect 4406 4507 4464 4533
rect 4406 4473 4418 4507
rect 4452 4473 4464 4507
rect 4406 4447 4464 4473
rect 4506 4507 4564 4533
rect 4506 4473 4518 4507
rect 4552 4473 4564 4507
rect 4506 4447 4564 4473
rect 4606 4507 4664 4533
rect 4606 4473 4618 4507
rect 4652 4473 4664 4507
rect 4606 4447 4664 4473
rect 4706 4507 4764 4533
rect 4706 4473 4718 4507
rect 4752 4473 4764 4507
rect 4706 4447 4764 4473
rect 4806 4507 4864 4533
rect 4806 4473 4818 4507
rect 4852 4473 4864 4507
rect 4806 4447 4864 4473
rect 4906 4507 4964 4533
rect 4906 4473 4918 4507
rect 4952 4473 4964 4507
rect 4906 4447 4964 4473
rect 5006 4507 5064 4533
rect 5006 4473 5012 4507
rect 5052 4473 5064 4507
rect 5006 4447 5064 4473
rect 5106 4507 5164 4533
rect 5106 4473 5118 4507
rect 5158 4473 5164 4507
rect 5106 4447 5164 4473
rect 5206 4507 5264 4533
rect 5206 4473 5218 4507
rect 5252 4473 5264 4507
rect 5206 4447 5264 4473
rect 5306 4507 5364 4533
rect 5306 4473 5312 4507
rect 5352 4473 5364 4507
rect 5306 4447 5364 4473
rect 5406 4507 5464 4533
rect 5406 4473 5418 4507
rect 5458 4473 5464 4507
rect 5406 4447 5464 4473
rect 5506 4507 5564 4533
rect 5506 4473 5518 4507
rect 5552 4473 5564 4507
rect 5506 4447 5564 4473
rect 5606 4507 5664 4533
rect 5606 4473 5618 4507
rect 5652 4473 5664 4507
rect 5606 4447 5664 4473
rect 5706 4507 5764 4533
rect 5706 4473 5718 4507
rect 5752 4473 5764 4507
rect 5706 4447 5764 4473
rect 5806 4507 5864 4533
rect 5806 4473 5818 4507
rect 5852 4473 5864 4507
rect 5806 4447 5864 4473
rect 5906 4507 5964 4533
rect 5906 4473 5918 4507
rect 5952 4473 5964 4507
rect 5906 4447 5964 4473
rect 6006 4507 6064 4533
rect 6006 4473 6012 4507
rect 6052 4473 6064 4507
rect 6006 4447 6064 4473
rect 6106 4507 6164 4533
rect 6106 4473 6118 4507
rect 6158 4473 6164 4507
rect 6106 4447 6164 4473
rect 6206 4507 6264 4533
rect 6206 4473 6218 4507
rect 6252 4473 6264 4507
rect 6206 4447 6264 4473
rect 6306 4507 6364 4533
rect 6306 4473 6318 4507
rect 6352 4473 6364 4507
rect 6306 4447 6364 4473
rect 6406 4507 6464 4533
rect 6406 4473 6418 4507
rect 6452 4473 6464 4507
rect 6406 4447 6464 4473
rect 6506 4507 6564 4533
rect 6506 4473 6518 4507
rect 6552 4473 6564 4507
rect 6506 4447 6564 4473
rect 6606 4507 6664 4533
rect 6606 4473 6618 4507
rect 6652 4473 6664 4507
rect 6606 4447 6664 4473
rect 6706 4507 6764 4533
rect 6706 4473 6718 4507
rect 6752 4473 6764 4507
rect 6706 4447 6764 4473
rect 6806 4507 6864 4533
rect 6806 4473 6818 4507
rect 6852 4473 6864 4507
rect 6806 4447 6864 4473
rect 6906 4507 6964 4533
rect 6906 4473 6918 4507
rect 6952 4473 6964 4507
rect 6906 4447 6964 4473
rect 7006 4507 7064 4533
rect 7006 4473 7018 4507
rect 7052 4473 7064 4507
rect 7006 4447 7064 4473
rect 7106 4507 7164 4533
rect 7106 4473 7118 4507
rect 7152 4473 7164 4507
rect 7106 4447 7164 4473
rect 7206 4507 7264 4533
rect 7206 4473 7218 4507
rect 7252 4473 7264 4507
rect 7206 4447 7264 4473
rect 7306 4507 7364 4533
rect 7306 4473 7318 4507
rect 7352 4473 7364 4507
rect 7306 4447 7364 4473
rect 7406 4507 7464 4533
rect 7406 4473 7418 4507
rect 7452 4473 7464 4507
rect 7406 4447 7464 4473
rect 7506 4507 7564 4533
rect 7506 4473 7518 4507
rect 7552 4473 7564 4507
rect 7506 4447 7564 4473
rect 7606 4507 7664 4533
rect 7606 4473 7618 4507
rect 7652 4473 7664 4507
rect 7606 4447 7664 4473
rect 7706 4507 7764 4533
rect 7706 4473 7718 4507
rect 7752 4473 7764 4507
rect 7706 4447 7764 4473
rect 7806 4507 7864 4533
rect 7806 4473 7818 4507
rect 7852 4473 7864 4507
rect 7806 4447 7864 4473
rect 7906 4507 7964 4533
rect 7906 4473 7918 4507
rect 7952 4473 7964 4507
rect 7906 4447 7964 4473
rect 8006 4507 8064 4533
rect 8006 4473 8012 4507
rect 8052 4473 8064 4507
rect 8006 4447 8064 4473
rect 8106 4507 8164 4533
rect 8106 4473 8118 4507
rect 8158 4473 8164 4507
rect 8106 4447 8164 4473
rect 8206 4507 8264 4533
rect 8206 4473 8218 4507
rect 8252 4473 8264 4507
rect 8206 4447 8264 4473
rect 8306 4507 8364 4533
rect 8306 4473 8312 4507
rect 8352 4473 8364 4507
rect 8306 4447 8364 4473
rect 8406 4507 8464 4533
rect 8406 4473 8418 4507
rect 8458 4473 8464 4507
rect 8406 4447 8464 4473
rect 8506 4507 8564 4533
rect 8506 4473 8518 4507
rect 8552 4473 8564 4507
rect 8506 4447 8564 4473
rect 8606 4507 8664 4533
rect 8606 4473 8618 4507
rect 8652 4473 8664 4507
rect 8606 4447 8664 4473
rect 8706 4507 8764 4533
rect 8706 4473 8718 4507
rect 8752 4473 8764 4507
rect 8706 4447 8764 4473
rect 8806 4507 8864 4533
rect 8806 4473 8812 4507
rect 8852 4473 8864 4507
rect 8806 4447 8864 4473
rect 8906 4507 8964 4533
rect 8906 4473 8918 4507
rect 8958 4473 8964 4507
rect 8906 4447 8964 4473
rect 9006 4507 9064 4533
rect 9006 4473 9012 4507
rect 9052 4473 9064 4507
rect 9006 4447 9064 4473
rect 9106 4507 9164 4533
rect 9106 4473 9118 4507
rect 9158 4473 9164 4507
rect 9106 4447 9164 4473
rect 9206 4507 9264 4533
rect 9206 4473 9218 4507
rect 9252 4473 9264 4507
rect 9206 4447 9264 4473
rect 9306 4507 9364 4533
rect 9306 4473 9312 4507
rect 9352 4473 9364 4507
rect 9306 4447 9364 4473
rect 9406 4507 9464 4533
rect 9406 4473 9418 4507
rect 9458 4473 9464 4507
rect 9406 4447 9464 4473
rect 9506 4507 9564 4533
rect 9506 4473 9518 4507
rect 9552 4473 9564 4507
rect 9506 4447 9564 4473
rect 9606 4507 9664 4533
rect 9606 4473 9612 4507
rect 9652 4473 9664 4507
rect 9606 4447 9664 4473
rect 9706 4507 9764 4533
rect 9706 4473 9718 4507
rect 9758 4473 9764 4507
rect 9706 4447 9764 4473
rect 9806 4507 9864 4533
rect 9806 4473 9818 4507
rect 9852 4473 9864 4507
rect 9806 4447 9864 4473
rect 9906 4507 9964 4533
rect 9906 4473 9912 4507
rect 9952 4473 9964 4507
rect 9906 4447 9964 4473
rect 10006 4507 10064 4533
rect 10006 4473 10018 4507
rect 10058 4473 10064 4507
rect 10006 4447 10064 4473
rect 10106 4507 10164 4533
rect 10106 4473 10118 4507
rect 10152 4473 10164 4507
rect 10106 4447 10164 4473
rect 10206 4507 10264 4533
rect 10206 4473 10212 4507
rect 10252 4473 10264 4507
rect 10206 4447 10264 4473
rect 10306 4507 10364 4533
rect 10306 4473 10318 4507
rect 10358 4473 10364 4507
rect 10306 4447 10364 4473
rect 10406 4507 10464 4533
rect 10406 4473 10418 4507
rect 10452 4473 10464 4507
rect 10406 4447 10464 4473
rect 10506 4507 10564 4533
rect 10506 4473 10512 4507
rect 10552 4473 10564 4507
rect 10506 4447 10564 4473
rect 10606 4507 10664 4533
rect 10606 4473 10618 4507
rect 10658 4473 10664 4507
rect 10606 4447 10664 4473
rect 10706 4507 10764 4533
rect 10706 4473 10712 4507
rect 10752 4473 10764 4507
rect 10706 4447 10764 4473
rect 10806 4507 10864 4533
rect 10806 4473 10818 4507
rect 10858 4473 10864 4507
rect 10806 4447 10864 4473
rect 10906 4507 10964 4533
rect 10906 4473 10912 4507
rect 10952 4473 10964 4507
rect 10906 4447 10964 4473
rect 11006 4507 11064 4533
rect 11006 4473 11018 4507
rect 11058 4473 11064 4507
rect 11006 4447 11064 4473
rect 11106 4507 11164 4533
rect 11106 4473 11118 4507
rect 11152 4473 11164 4507
rect 11106 4447 11164 4473
rect 11206 4507 11264 4533
rect 11206 4473 11212 4507
rect 11252 4473 11264 4507
rect 11206 4447 11264 4473
rect 11306 4507 11364 4533
rect 11306 4473 11318 4507
rect 11358 4473 11364 4507
rect 11306 4447 11364 4473
rect 11406 4507 11464 4533
rect 11406 4473 11418 4507
rect 11452 4473 11464 4507
rect 11406 4447 11464 4473
rect 11506 4507 11564 4533
rect 11506 4473 11518 4507
rect 11552 4473 11564 4507
rect 11506 4447 11564 4473
rect 11606 4507 11664 4533
rect 11606 4473 11618 4507
rect 11652 4473 11664 4507
rect 11606 4447 11664 4473
rect 11706 4507 11764 4533
rect 11706 4473 11718 4507
rect 11752 4473 11764 4507
rect 11706 4447 11764 4473
rect 11806 4507 11864 4533
rect 11806 4473 11818 4507
rect 11852 4473 11864 4507
rect 11806 4447 11864 4473
rect 11906 4507 11964 4533
rect 11906 4473 11918 4507
rect 11952 4473 11964 4507
rect 11906 4447 11964 4473
rect 12006 4507 12064 4533
rect 12006 4473 12018 4507
rect 12052 4473 12064 4507
rect 12006 4447 12064 4473
rect 12106 4507 12164 4533
rect 12106 4473 12118 4507
rect 12152 4473 12164 4507
rect 12106 4447 12164 4473
rect 12206 4507 12264 4533
rect 12206 4473 12218 4507
rect 12252 4473 12264 4507
rect 12206 4447 12264 4473
rect 12306 4507 12364 4533
rect 12306 4473 12318 4507
rect 12352 4473 12364 4507
rect 12306 4447 12364 4473
rect 12406 4507 12464 4533
rect 12406 4473 12412 4507
rect 12452 4473 12464 4507
rect 12406 4447 12464 4473
rect 12506 4507 12564 4533
rect 12506 4473 12518 4507
rect 12558 4473 12564 4507
rect 12506 4447 12564 4473
rect 12606 4507 12664 4533
rect 12606 4473 12618 4507
rect 12652 4473 12664 4507
rect 12606 4447 12664 4473
rect 12706 4507 12764 4533
rect 12706 4473 12718 4507
rect 12752 4473 12764 4507
rect 12706 4447 12764 4473
rect 12806 4507 12864 4533
rect 13018 4526 13262 4560
rect 12806 4473 12812 4507
rect 12852 4473 12864 4507
rect 12908 4488 12916 4522
rect 12958 4488 12974 4522
rect 13018 4507 13052 4526
rect 12806 4447 12864 4473
rect 13228 4523 13262 4526
rect 13228 4507 13362 4523
rect 13018 4457 13052 4473
rect 13096 4458 13112 4492
rect 13154 4458 13162 4492
rect 13262 4473 13328 4507
rect 13228 4457 13362 4473
rect 13428 4507 13462 4523
rect 13428 4457 13462 4473
rect 13528 4507 13662 4523
rect 13562 4473 13628 4507
rect 13528 4457 13662 4473
rect 6 4367 64 4393
rect 6 4333 18 4367
rect 58 4333 64 4367
rect 6 4307 64 4333
rect 106 4367 164 4393
rect 106 4333 118 4367
rect 152 4333 164 4367
rect 106 4307 164 4333
rect 206 4367 264 4393
rect 206 4333 218 4367
rect 252 4333 264 4367
rect 206 4307 264 4333
rect 306 4367 364 4393
rect 306 4333 318 4367
rect 352 4333 364 4367
rect 306 4307 364 4333
rect 406 4367 464 4393
rect 406 4333 418 4367
rect 452 4333 464 4367
rect 406 4307 464 4333
rect 506 4367 564 4393
rect 506 4333 518 4367
rect 552 4333 564 4367
rect 506 4307 564 4333
rect 606 4367 664 4393
rect 606 4333 618 4367
rect 652 4333 664 4367
rect 606 4307 664 4333
rect 706 4367 764 4393
rect 706 4333 718 4367
rect 752 4333 764 4367
rect 706 4307 764 4333
rect 806 4367 864 4393
rect 806 4333 818 4367
rect 852 4333 864 4367
rect 806 4307 864 4333
rect 906 4367 964 4393
rect 906 4333 918 4367
rect 952 4333 964 4367
rect 906 4307 964 4333
rect 1006 4367 1064 4393
rect 1006 4333 1018 4367
rect 1052 4333 1064 4367
rect 1006 4307 1064 4333
rect 1106 4367 1164 4393
rect 1106 4333 1118 4367
rect 1152 4333 1164 4367
rect 1106 4307 1164 4333
rect 1206 4367 1264 4393
rect 1206 4333 1212 4367
rect 1252 4333 1264 4367
rect 1206 4307 1264 4333
rect 1306 4367 1364 4393
rect 1306 4333 1318 4367
rect 1358 4333 1364 4367
rect 1306 4307 1364 4333
rect 1406 4367 1464 4393
rect 1406 4333 1418 4367
rect 1452 4333 1464 4367
rect 1406 4307 1464 4333
rect 1506 4367 1564 4393
rect 1506 4333 1518 4367
rect 1552 4333 1564 4367
rect 1506 4307 1564 4333
rect 1606 4367 1664 4393
rect 1606 4333 1618 4367
rect 1652 4333 1664 4367
rect 1606 4307 1664 4333
rect 1706 4367 1764 4393
rect 1706 4333 1718 4367
rect 1752 4333 1764 4367
rect 1706 4307 1764 4333
rect 1806 4367 1864 4393
rect 1806 4333 1818 4367
rect 1852 4333 1864 4367
rect 1806 4307 1864 4333
rect 1906 4367 1964 4393
rect 1906 4333 1912 4367
rect 1952 4333 1964 4367
rect 1906 4307 1964 4333
rect 2006 4367 2064 4393
rect 2006 4333 2018 4367
rect 2058 4333 2064 4367
rect 2006 4307 2064 4333
rect 2106 4367 2164 4393
rect 2106 4333 2118 4367
rect 2152 4333 2164 4367
rect 2106 4307 2164 4333
rect 2206 4367 2264 4393
rect 2206 4333 2218 4367
rect 2252 4333 2264 4367
rect 2206 4307 2264 4333
rect 2306 4367 2364 4393
rect 2306 4333 2318 4367
rect 2352 4333 2364 4367
rect 2306 4307 2364 4333
rect 2406 4367 2464 4393
rect 2406 4333 2418 4367
rect 2452 4333 2464 4367
rect 2406 4307 2464 4333
rect 2506 4367 2564 4393
rect 2506 4333 2518 4367
rect 2552 4333 2564 4367
rect 2506 4307 2564 4333
rect 2606 4367 2664 4393
rect 2606 4333 2618 4367
rect 2652 4333 2664 4367
rect 2606 4307 2664 4333
rect 2706 4367 2764 4393
rect 2706 4333 2718 4367
rect 2752 4333 2764 4367
rect 2706 4307 2764 4333
rect 2806 4367 2864 4393
rect 2806 4333 2818 4367
rect 2852 4333 2864 4367
rect 2806 4307 2864 4333
rect 2906 4367 2964 4393
rect 2906 4333 2918 4367
rect 2952 4333 2964 4367
rect 2906 4307 2964 4333
rect 3006 4367 3064 4393
rect 3006 4333 3018 4367
rect 3052 4333 3064 4367
rect 3006 4307 3064 4333
rect 3106 4367 3164 4393
rect 3106 4333 3118 4367
rect 3152 4333 3164 4367
rect 3106 4307 3164 4333
rect 3206 4367 3264 4393
rect 3206 4333 3218 4367
rect 3252 4333 3264 4367
rect 3206 4307 3264 4333
rect 3306 4367 3364 4393
rect 3306 4333 3318 4367
rect 3352 4333 3364 4367
rect 3306 4307 3364 4333
rect 3406 4367 3464 4393
rect 3406 4333 3418 4367
rect 3452 4333 3464 4367
rect 3406 4307 3464 4333
rect 3506 4367 3564 4393
rect 3506 4333 3518 4367
rect 3552 4333 3564 4367
rect 3506 4307 3564 4333
rect 3606 4367 3664 4393
rect 3606 4333 3618 4367
rect 3652 4333 3664 4367
rect 3606 4307 3664 4333
rect 3706 4367 3764 4393
rect 3706 4333 3712 4367
rect 3752 4333 3764 4367
rect 3706 4307 3764 4333
rect 3806 4367 3864 4393
rect 3806 4333 3818 4367
rect 3858 4333 3864 4367
rect 3806 4307 3864 4333
rect 3906 4367 3964 4393
rect 3906 4333 3918 4367
rect 3952 4333 3964 4367
rect 3906 4307 3964 4333
rect 4006 4367 4064 4393
rect 4006 4333 4018 4367
rect 4052 4333 4064 4367
rect 4006 4307 4064 4333
rect 4106 4367 4164 4393
rect 4106 4333 4118 4367
rect 4152 4333 4164 4367
rect 4106 4307 4164 4333
rect 4206 4367 4264 4393
rect 4206 4333 4218 4367
rect 4252 4333 4264 4367
rect 4206 4307 4264 4333
rect 4306 4367 4364 4393
rect 4306 4333 4318 4367
rect 4352 4333 4364 4367
rect 4306 4307 4364 4333
rect 4406 4367 4464 4393
rect 4406 4333 4418 4367
rect 4452 4333 4464 4367
rect 4406 4307 4464 4333
rect 4506 4367 4564 4393
rect 4506 4333 4518 4367
rect 4552 4333 4564 4367
rect 4506 4307 4564 4333
rect 4606 4367 4664 4393
rect 4606 4333 4618 4367
rect 4652 4333 4664 4367
rect 4606 4307 4664 4333
rect 4706 4367 4764 4393
rect 4706 4333 4718 4367
rect 4752 4333 4764 4367
rect 4706 4307 4764 4333
rect 4806 4367 4864 4393
rect 4806 4333 4818 4367
rect 4852 4333 4864 4367
rect 4806 4307 4864 4333
rect 4906 4367 4964 4393
rect 4906 4333 4918 4367
rect 4952 4333 4964 4367
rect 4906 4307 4964 4333
rect 5006 4367 5064 4393
rect 5006 4333 5018 4367
rect 5052 4333 5064 4367
rect 5006 4307 5064 4333
rect 5106 4367 5164 4393
rect 5106 4333 5118 4367
rect 5152 4333 5164 4367
rect 5106 4307 5164 4333
rect 5206 4367 5264 4393
rect 5206 4333 5218 4367
rect 5252 4333 5264 4367
rect 5206 4307 5264 4333
rect 5306 4367 5364 4393
rect 5306 4333 5318 4367
rect 5352 4333 5364 4367
rect 5306 4307 5364 4333
rect 5406 4367 5464 4393
rect 5406 4333 5418 4367
rect 5452 4333 5464 4367
rect 5406 4307 5464 4333
rect 5506 4367 5564 4393
rect 5506 4333 5518 4367
rect 5552 4333 5564 4367
rect 5506 4307 5564 4333
rect 5606 4367 5664 4393
rect 5606 4333 5618 4367
rect 5652 4333 5664 4367
rect 5606 4307 5664 4333
rect 5706 4367 5764 4393
rect 5706 4333 5718 4367
rect 5752 4333 5764 4367
rect 5706 4307 5764 4333
rect 5806 4367 5864 4393
rect 5806 4333 5818 4367
rect 5852 4333 5864 4367
rect 5806 4307 5864 4333
rect 5906 4367 5964 4393
rect 5906 4333 5918 4367
rect 5952 4333 5964 4367
rect 5906 4307 5964 4333
rect 6006 4367 6064 4393
rect 6006 4333 6012 4367
rect 6052 4333 6064 4367
rect 6006 4307 6064 4333
rect 6106 4367 6164 4393
rect 6106 4333 6118 4367
rect 6158 4333 6164 4367
rect 6106 4307 6164 4333
rect 6206 4367 6264 4393
rect 6206 4333 6218 4367
rect 6252 4333 6264 4367
rect 6206 4307 6264 4333
rect 6306 4367 6364 4393
rect 6306 4333 6318 4367
rect 6352 4333 6364 4367
rect 6306 4307 6364 4333
rect 6406 4367 6464 4393
rect 6406 4333 6418 4367
rect 6452 4333 6464 4367
rect 6406 4307 6464 4333
rect 6506 4367 6564 4393
rect 6506 4333 6518 4367
rect 6552 4333 6564 4367
rect 6506 4307 6564 4333
rect 6606 4367 6664 4393
rect 6606 4333 6612 4367
rect 6652 4333 6664 4367
rect 6606 4307 6664 4333
rect 6706 4367 6764 4393
rect 6706 4333 6718 4367
rect 6758 4333 6764 4367
rect 6706 4307 6764 4333
rect 6806 4367 6864 4393
rect 6806 4333 6818 4367
rect 6852 4333 6864 4367
rect 6806 4307 6864 4333
rect 6906 4367 6964 4393
rect 6906 4333 6918 4367
rect 6952 4333 6964 4367
rect 6906 4307 6964 4333
rect 7006 4367 7064 4393
rect 7006 4333 7018 4367
rect 7052 4333 7064 4367
rect 7006 4307 7064 4333
rect 7106 4367 7164 4393
rect 7106 4333 7118 4367
rect 7152 4333 7164 4367
rect 7106 4307 7164 4333
rect 7206 4367 7264 4393
rect 7206 4333 7218 4367
rect 7252 4333 7264 4367
rect 7206 4307 7264 4333
rect 7306 4367 7364 4393
rect 7306 4333 7312 4367
rect 7352 4333 7364 4367
rect 7306 4307 7364 4333
rect 7406 4367 7464 4393
rect 7406 4333 7418 4367
rect 7458 4333 7464 4367
rect 7406 4307 7464 4333
rect 7506 4367 7564 4393
rect 7506 4333 7518 4367
rect 7552 4333 7564 4367
rect 7506 4307 7564 4333
rect 7606 4367 7664 4393
rect 7606 4333 7618 4367
rect 7652 4333 7664 4367
rect 7606 4307 7664 4333
rect 7706 4367 7764 4393
rect 7706 4333 7718 4367
rect 7752 4333 7764 4367
rect 7706 4307 7764 4333
rect 7806 4367 7864 4393
rect 7806 4333 7818 4367
rect 7852 4333 7864 4367
rect 7806 4307 7864 4333
rect 7906 4367 7964 4393
rect 7906 4333 7918 4367
rect 7952 4333 7964 4367
rect 7906 4307 7964 4333
rect 8006 4367 8064 4393
rect 8006 4333 8018 4367
rect 8052 4333 8064 4367
rect 8006 4307 8064 4333
rect 8106 4367 8164 4393
rect 8106 4333 8118 4367
rect 8152 4333 8164 4367
rect 8106 4307 8164 4333
rect 8206 4367 8264 4393
rect 8206 4333 8218 4367
rect 8252 4333 8264 4367
rect 8206 4307 8264 4333
rect 8306 4367 8364 4393
rect 8306 4333 8318 4367
rect 8352 4333 8364 4367
rect 8306 4307 8364 4333
rect 8406 4367 8464 4393
rect 8406 4333 8418 4367
rect 8452 4333 8464 4367
rect 8406 4307 8464 4333
rect 8506 4367 8564 4393
rect 8506 4333 8518 4367
rect 8552 4333 8564 4367
rect 8506 4307 8564 4333
rect 8606 4367 8664 4393
rect 8606 4333 8618 4367
rect 8652 4333 8664 4367
rect 8606 4307 8664 4333
rect 8706 4367 8764 4393
rect 8706 4333 8718 4367
rect 8752 4333 8764 4367
rect 8706 4307 8764 4333
rect 8806 4367 8864 4393
rect 8806 4333 8818 4367
rect 8852 4333 8864 4367
rect 8806 4307 8864 4333
rect 8906 4367 8964 4393
rect 8906 4333 8918 4367
rect 8952 4333 8964 4367
rect 8906 4307 8964 4333
rect 9006 4367 9064 4393
rect 9006 4333 9018 4367
rect 9052 4333 9064 4367
rect 9006 4307 9064 4333
rect 9106 4367 9164 4393
rect 9106 4333 9118 4367
rect 9152 4333 9164 4367
rect 9106 4307 9164 4333
rect 9206 4367 9264 4393
rect 9206 4333 9218 4367
rect 9252 4333 9264 4367
rect 9206 4307 9264 4333
rect 9306 4367 9364 4393
rect 9306 4333 9318 4367
rect 9352 4333 9364 4367
rect 9306 4307 9364 4333
rect 9406 4367 9464 4393
rect 9406 4333 9418 4367
rect 9452 4333 9464 4367
rect 9406 4307 9464 4333
rect 9506 4367 9564 4393
rect 9506 4333 9518 4367
rect 9552 4333 9564 4367
rect 9506 4307 9564 4333
rect 9606 4367 9664 4393
rect 9606 4333 9618 4367
rect 9652 4333 9664 4367
rect 9606 4307 9664 4333
rect 9706 4367 9764 4393
rect 9706 4333 9718 4367
rect 9752 4333 9764 4367
rect 9706 4307 9764 4333
rect 9806 4367 9864 4393
rect 9806 4333 9818 4367
rect 9852 4333 9864 4367
rect 9806 4307 9864 4333
rect 9906 4367 9964 4393
rect 9906 4333 9918 4367
rect 9952 4333 9964 4367
rect 9906 4307 9964 4333
rect 10006 4367 10064 4393
rect 10006 4333 10018 4367
rect 10052 4333 10064 4367
rect 10006 4307 10064 4333
rect 10106 4367 10164 4393
rect 10106 4333 10118 4367
rect 10152 4333 10164 4367
rect 10106 4307 10164 4333
rect 10206 4367 10264 4393
rect 10206 4333 10218 4367
rect 10252 4333 10264 4367
rect 10206 4307 10264 4333
rect 10306 4367 10364 4393
rect 10306 4333 10318 4367
rect 10352 4333 10364 4367
rect 10306 4307 10364 4333
rect 10406 4367 10464 4393
rect 10406 4333 10418 4367
rect 10452 4333 10464 4367
rect 10406 4307 10464 4333
rect 10506 4367 10564 4393
rect 10506 4333 10518 4367
rect 10552 4333 10564 4367
rect 10506 4307 10564 4333
rect 10606 4367 10664 4393
rect 10606 4333 10618 4367
rect 10652 4333 10664 4367
rect 10606 4307 10664 4333
rect 10706 4367 10764 4393
rect 10706 4333 10718 4367
rect 10752 4333 10764 4367
rect 10706 4307 10764 4333
rect 10806 4367 10864 4393
rect 10806 4333 10812 4367
rect 10852 4333 10864 4367
rect 10806 4307 10864 4333
rect 10906 4367 10964 4393
rect 10906 4333 10918 4367
rect 10958 4333 10964 4367
rect 10906 4307 10964 4333
rect 11006 4367 11064 4393
rect 11006 4333 11018 4367
rect 11052 4333 11064 4367
rect 11006 4307 11064 4333
rect 11106 4367 11164 4393
rect 11106 4333 11112 4367
rect 11152 4333 11164 4367
rect 11106 4307 11164 4333
rect 11206 4367 11264 4393
rect 11206 4333 11218 4367
rect 11258 4333 11264 4367
rect 11206 4307 11264 4333
rect 11306 4367 11364 4393
rect 11306 4333 11318 4367
rect 11352 4333 11364 4367
rect 11306 4307 11364 4333
rect 11406 4367 11464 4393
rect 11406 4333 11418 4367
rect 11452 4333 11464 4367
rect 11406 4307 11464 4333
rect 11506 4367 11564 4393
rect 11506 4333 11518 4367
rect 11552 4333 11564 4367
rect 11506 4307 11564 4333
rect 11606 4367 11664 4393
rect 11606 4333 11618 4367
rect 11652 4333 11664 4367
rect 11606 4307 11664 4333
rect 11706 4367 11764 4393
rect 11706 4333 11718 4367
rect 11752 4333 11764 4367
rect 11706 4307 11764 4333
rect 11806 4367 11864 4393
rect 11806 4333 11818 4367
rect 11852 4333 11864 4367
rect 11806 4307 11864 4333
rect 11906 4367 11964 4393
rect 11906 4333 11912 4367
rect 11952 4333 11964 4367
rect 11906 4307 11964 4333
rect 12006 4367 12064 4393
rect 12006 4333 12018 4367
rect 12058 4333 12064 4367
rect 12006 4307 12064 4333
rect 12106 4367 12164 4393
rect 12106 4333 12118 4367
rect 12152 4333 12164 4367
rect 12106 4307 12164 4333
rect 12206 4367 12264 4393
rect 12206 4333 12218 4367
rect 12252 4333 12264 4367
rect 12206 4307 12264 4333
rect 12306 4367 12364 4393
rect 12306 4333 12318 4367
rect 12352 4333 12364 4367
rect 12306 4307 12364 4333
rect 12406 4367 12464 4393
rect 12406 4333 12418 4367
rect 12452 4333 12464 4367
rect 12406 4307 12464 4333
rect 12506 4367 12564 4393
rect 12506 4333 12518 4367
rect 12552 4333 12564 4367
rect 12506 4307 12564 4333
rect 12606 4367 12664 4393
rect 12606 4333 12618 4367
rect 12652 4333 12664 4367
rect 12606 4307 12664 4333
rect 12706 4367 12764 4393
rect 12706 4333 12718 4367
rect 12752 4333 12764 4367
rect 12706 4307 12764 4333
rect 12806 4367 12864 4393
rect 13018 4386 13262 4420
rect 12806 4333 12812 4367
rect 12852 4333 12864 4367
rect 12908 4348 12916 4382
rect 12958 4348 12974 4382
rect 13018 4367 13052 4386
rect 12806 4307 12864 4333
rect 13228 4367 13262 4386
rect 13018 4317 13052 4333
rect 13096 4318 13112 4352
rect 13154 4318 13162 4352
rect 13228 4317 13262 4333
rect 13328 4367 13462 4383
rect 13362 4333 13428 4367
rect 13328 4317 13462 4333
rect 13528 4367 13662 4383
rect 13562 4333 13628 4367
rect 13528 4317 13662 4333
rect 6 4227 64 4253
rect 6 4193 18 4227
rect 52 4193 64 4227
rect 6 4167 64 4193
rect 106 4227 164 4253
rect 106 4193 118 4227
rect 152 4193 164 4227
rect 106 4167 164 4193
rect 206 4227 264 4253
rect 206 4193 218 4227
rect 252 4193 264 4227
rect 206 4167 264 4193
rect 306 4227 364 4253
rect 306 4193 318 4227
rect 352 4193 364 4227
rect 306 4167 364 4193
rect 406 4227 464 4253
rect 406 4193 418 4227
rect 452 4193 464 4227
rect 406 4167 464 4193
rect 506 4227 564 4253
rect 506 4193 512 4227
rect 552 4193 564 4227
rect 506 4167 564 4193
rect 606 4227 664 4253
rect 606 4193 618 4227
rect 658 4193 664 4227
rect 606 4167 664 4193
rect 706 4227 764 4253
rect 706 4193 718 4227
rect 752 4193 764 4227
rect 706 4167 764 4193
rect 806 4227 864 4253
rect 806 4193 818 4227
rect 852 4193 864 4227
rect 806 4167 864 4193
rect 906 4227 964 4253
rect 906 4193 918 4227
rect 952 4193 964 4227
rect 906 4167 964 4193
rect 1006 4227 1064 4253
rect 1006 4193 1018 4227
rect 1052 4193 1064 4227
rect 1006 4167 1064 4193
rect 1106 4227 1164 4253
rect 1106 4193 1112 4227
rect 1152 4193 1164 4227
rect 1106 4167 1164 4193
rect 1206 4227 1264 4253
rect 1206 4193 1218 4227
rect 1258 4193 1264 4227
rect 1206 4167 1264 4193
rect 1306 4227 1364 4253
rect 1306 4193 1318 4227
rect 1352 4193 1364 4227
rect 1306 4167 1364 4193
rect 1406 4227 1464 4253
rect 1406 4193 1418 4227
rect 1452 4193 1464 4227
rect 1406 4167 1464 4193
rect 1506 4227 1564 4253
rect 1506 4193 1518 4227
rect 1552 4193 1564 4227
rect 1506 4167 1564 4193
rect 1606 4227 1664 4253
rect 1606 4193 1618 4227
rect 1652 4193 1664 4227
rect 1606 4167 1664 4193
rect 1706 4227 1764 4253
rect 1706 4193 1718 4227
rect 1752 4193 1764 4227
rect 1706 4167 1764 4193
rect 1806 4227 1864 4253
rect 1806 4193 1818 4227
rect 1852 4193 1864 4227
rect 1806 4167 1864 4193
rect 1906 4227 1964 4253
rect 1906 4193 1912 4227
rect 1952 4193 1964 4227
rect 1906 4167 1964 4193
rect 2006 4227 2064 4253
rect 2006 4193 2018 4227
rect 2058 4193 2064 4227
rect 2006 4167 2064 4193
rect 2106 4227 2164 4253
rect 2106 4193 2118 4227
rect 2152 4193 2164 4227
rect 2106 4167 2164 4193
rect 2206 4227 2264 4253
rect 2206 4193 2218 4227
rect 2252 4193 2264 4227
rect 2206 4167 2264 4193
rect 2306 4227 2364 4253
rect 2306 4193 2318 4227
rect 2352 4193 2364 4227
rect 2306 4167 2364 4193
rect 2406 4227 2464 4253
rect 2406 4193 2418 4227
rect 2452 4193 2464 4227
rect 2406 4167 2464 4193
rect 2506 4227 2564 4253
rect 2506 4193 2518 4227
rect 2552 4193 2564 4227
rect 2506 4167 2564 4193
rect 2606 4227 2664 4253
rect 2606 4193 2618 4227
rect 2652 4193 2664 4227
rect 2606 4167 2664 4193
rect 2706 4227 2764 4253
rect 2706 4193 2718 4227
rect 2752 4193 2764 4227
rect 2706 4167 2764 4193
rect 2806 4227 2864 4253
rect 2806 4193 2818 4227
rect 2852 4193 2864 4227
rect 2806 4167 2864 4193
rect 2906 4227 2964 4253
rect 2906 4193 2918 4227
rect 2952 4193 2964 4227
rect 2906 4167 2964 4193
rect 3006 4227 3064 4253
rect 3006 4193 3018 4227
rect 3052 4193 3064 4227
rect 3006 4167 3064 4193
rect 3106 4227 3164 4253
rect 3106 4193 3118 4227
rect 3152 4193 3164 4227
rect 3106 4167 3164 4193
rect 3206 4227 3264 4253
rect 3206 4193 3218 4227
rect 3252 4193 3264 4227
rect 3206 4167 3264 4193
rect 3306 4227 3364 4253
rect 3306 4193 3318 4227
rect 3352 4193 3364 4227
rect 3306 4167 3364 4193
rect 3406 4227 3464 4253
rect 3406 4193 3418 4227
rect 3452 4193 3464 4227
rect 3406 4167 3464 4193
rect 3506 4227 3564 4253
rect 3506 4193 3518 4227
rect 3552 4193 3564 4227
rect 3506 4167 3564 4193
rect 3606 4227 3664 4253
rect 3606 4193 3618 4227
rect 3652 4193 3664 4227
rect 3606 4167 3664 4193
rect 3706 4227 3764 4253
rect 3706 4193 3718 4227
rect 3752 4193 3764 4227
rect 3706 4167 3764 4193
rect 3806 4227 3864 4253
rect 3806 4193 3818 4227
rect 3852 4193 3864 4227
rect 3806 4167 3864 4193
rect 3906 4227 3964 4253
rect 3906 4193 3918 4227
rect 3952 4193 3964 4227
rect 3906 4167 3964 4193
rect 4006 4227 4064 4253
rect 4006 4193 4012 4227
rect 4052 4193 4064 4227
rect 4006 4167 4064 4193
rect 4106 4227 4164 4253
rect 4106 4193 4118 4227
rect 4158 4193 4164 4227
rect 4106 4167 4164 4193
rect 4206 4227 4264 4253
rect 4206 4193 4212 4227
rect 4252 4193 4264 4227
rect 4206 4167 4264 4193
rect 4306 4227 4364 4253
rect 4306 4193 4318 4227
rect 4358 4193 4364 4227
rect 4306 4167 4364 4193
rect 4406 4227 4464 4253
rect 4406 4193 4412 4227
rect 4452 4193 4464 4227
rect 4406 4167 4464 4193
rect 4506 4227 4564 4253
rect 4506 4193 4518 4227
rect 4558 4193 4564 4227
rect 4506 4167 4564 4193
rect 4606 4227 4664 4253
rect 4606 4193 4612 4227
rect 4652 4193 4664 4227
rect 4606 4167 4664 4193
rect 4706 4227 4764 4253
rect 4706 4193 4718 4227
rect 4758 4193 4764 4227
rect 4706 4167 4764 4193
rect 4806 4227 4864 4253
rect 4806 4193 4812 4227
rect 4852 4193 4864 4227
rect 4806 4167 4864 4193
rect 4906 4227 4964 4253
rect 4906 4193 4918 4227
rect 4958 4193 4964 4227
rect 4906 4167 4964 4193
rect 5006 4227 5064 4253
rect 5006 4193 5018 4227
rect 5052 4193 5064 4227
rect 5006 4167 5064 4193
rect 5106 4227 5164 4253
rect 5106 4193 5118 4227
rect 5152 4193 5164 4227
rect 5106 4167 5164 4193
rect 5206 4227 5264 4253
rect 5206 4193 5218 4227
rect 5252 4193 5264 4227
rect 5206 4167 5264 4193
rect 5306 4227 5364 4253
rect 5306 4193 5318 4227
rect 5352 4193 5364 4227
rect 5306 4167 5364 4193
rect 5406 4227 5464 4253
rect 5406 4193 5418 4227
rect 5452 4193 5464 4227
rect 5406 4167 5464 4193
rect 5506 4227 5564 4253
rect 5506 4193 5512 4227
rect 5552 4193 5564 4227
rect 5506 4167 5564 4193
rect 5606 4227 5664 4253
rect 5606 4193 5618 4227
rect 5658 4193 5664 4227
rect 5606 4167 5664 4193
rect 5706 4227 5764 4253
rect 5706 4193 5718 4227
rect 5752 4193 5764 4227
rect 5706 4167 5764 4193
rect 5806 4227 5864 4253
rect 5806 4193 5818 4227
rect 5852 4193 5864 4227
rect 5806 4167 5864 4193
rect 5906 4227 5964 4253
rect 5906 4193 5918 4227
rect 5952 4193 5964 4227
rect 5906 4167 5964 4193
rect 6006 4227 6064 4253
rect 6006 4193 6012 4227
rect 6052 4193 6064 4227
rect 6006 4167 6064 4193
rect 6106 4227 6164 4253
rect 6106 4193 6118 4227
rect 6158 4193 6164 4227
rect 6106 4167 6164 4193
rect 6206 4227 6264 4253
rect 6206 4193 6212 4227
rect 6252 4193 6264 4227
rect 6206 4167 6264 4193
rect 6306 4227 6364 4253
rect 6306 4193 6318 4227
rect 6358 4193 6364 4227
rect 6306 4167 6364 4193
rect 6406 4227 6464 4253
rect 6406 4193 6412 4227
rect 6452 4193 6464 4227
rect 6406 4167 6464 4193
rect 6506 4227 6564 4253
rect 6506 4193 6518 4227
rect 6558 4193 6564 4227
rect 6506 4167 6564 4193
rect 6606 4227 6664 4253
rect 6606 4193 6612 4227
rect 6652 4193 6664 4227
rect 6606 4167 6664 4193
rect 6706 4227 6764 4253
rect 6706 4193 6718 4227
rect 6758 4193 6764 4227
rect 6706 4167 6764 4193
rect 6806 4227 6864 4253
rect 6806 4193 6818 4227
rect 6852 4193 6864 4227
rect 6806 4167 6864 4193
rect 6906 4227 6964 4253
rect 6906 4193 6918 4227
rect 6952 4193 6964 4227
rect 6906 4167 6964 4193
rect 7006 4227 7064 4253
rect 7006 4193 7018 4227
rect 7052 4193 7064 4227
rect 7006 4167 7064 4193
rect 7106 4227 7164 4253
rect 7106 4193 7112 4227
rect 7152 4193 7164 4227
rect 7106 4167 7164 4193
rect 7206 4227 7264 4253
rect 7206 4193 7218 4227
rect 7258 4193 7264 4227
rect 7206 4167 7264 4193
rect 7306 4227 7364 4253
rect 7306 4193 7318 4227
rect 7352 4193 7364 4227
rect 7306 4167 7364 4193
rect 7406 4227 7464 4253
rect 7406 4193 7418 4227
rect 7452 4193 7464 4227
rect 7406 4167 7464 4193
rect 7506 4227 7564 4253
rect 7506 4193 7518 4227
rect 7552 4193 7564 4227
rect 7506 4167 7564 4193
rect 7606 4227 7664 4253
rect 7606 4193 7618 4227
rect 7652 4193 7664 4227
rect 7606 4167 7664 4193
rect 7706 4227 7764 4253
rect 7706 4193 7718 4227
rect 7752 4193 7764 4227
rect 7706 4167 7764 4193
rect 7806 4227 7864 4253
rect 7806 4193 7818 4227
rect 7852 4193 7864 4227
rect 7806 4167 7864 4193
rect 7906 4227 7964 4253
rect 7906 4193 7918 4227
rect 7952 4193 7964 4227
rect 7906 4167 7964 4193
rect 8006 4227 8064 4253
rect 8006 4193 8018 4227
rect 8052 4193 8064 4227
rect 8006 4167 8064 4193
rect 8106 4227 8164 4253
rect 8106 4193 8112 4227
rect 8152 4193 8164 4227
rect 8106 4167 8164 4193
rect 8206 4227 8264 4253
rect 8206 4193 8218 4227
rect 8258 4193 8264 4227
rect 8206 4167 8264 4193
rect 8306 4227 8364 4253
rect 8306 4193 8312 4227
rect 8352 4193 8364 4227
rect 8306 4167 8364 4193
rect 8406 4227 8464 4253
rect 8406 4193 8418 4227
rect 8458 4193 8464 4227
rect 8406 4167 8464 4193
rect 8506 4227 8564 4253
rect 8506 4193 8512 4227
rect 8552 4193 8564 4227
rect 8506 4167 8564 4193
rect 8606 4227 8664 4253
rect 8606 4193 8618 4227
rect 8658 4193 8664 4227
rect 8606 4167 8664 4193
rect 8706 4227 8764 4253
rect 8706 4193 8712 4227
rect 8752 4193 8764 4227
rect 8706 4167 8764 4193
rect 8806 4227 8864 4253
rect 8806 4193 8818 4227
rect 8858 4193 8864 4227
rect 8806 4167 8864 4193
rect 8906 4227 8964 4253
rect 8906 4193 8912 4227
rect 8952 4193 8964 4227
rect 8906 4167 8964 4193
rect 9006 4227 9064 4253
rect 9006 4193 9018 4227
rect 9058 4193 9064 4227
rect 9006 4167 9064 4193
rect 9106 4227 9164 4253
rect 9106 4193 9118 4227
rect 9152 4193 9164 4227
rect 9106 4167 9164 4193
rect 9206 4227 9264 4253
rect 9206 4193 9218 4227
rect 9252 4193 9264 4227
rect 9206 4167 9264 4193
rect 9306 4227 9364 4253
rect 9306 4193 9312 4227
rect 9352 4193 9364 4227
rect 9306 4167 9364 4193
rect 9406 4227 9464 4253
rect 9406 4193 9418 4227
rect 9458 4193 9464 4227
rect 9406 4167 9464 4193
rect 9506 4227 9564 4253
rect 9506 4193 9512 4227
rect 9552 4193 9564 4227
rect 9506 4167 9564 4193
rect 9606 4227 9664 4253
rect 9606 4193 9618 4227
rect 9658 4193 9664 4227
rect 9606 4167 9664 4193
rect 9706 4227 9764 4253
rect 9706 4193 9712 4227
rect 9752 4193 9764 4227
rect 9706 4167 9764 4193
rect 9806 4227 9864 4253
rect 9806 4193 9818 4227
rect 9858 4193 9864 4227
rect 9806 4167 9864 4193
rect 9906 4227 9964 4253
rect 9906 4193 9918 4227
rect 9952 4193 9964 4227
rect 9906 4167 9964 4193
rect 10006 4227 10064 4253
rect 10006 4193 10012 4227
rect 10052 4193 10064 4227
rect 10006 4167 10064 4193
rect 10106 4227 10164 4253
rect 10106 4193 10118 4227
rect 10158 4193 10164 4227
rect 10106 4167 10164 4193
rect 10206 4227 10264 4253
rect 10206 4193 10218 4227
rect 10252 4193 10264 4227
rect 10206 4167 10264 4193
rect 10306 4227 10364 4253
rect 10306 4193 10318 4227
rect 10352 4193 10364 4227
rect 10306 4167 10364 4193
rect 10406 4227 10464 4253
rect 10406 4193 10418 4227
rect 10452 4193 10464 4227
rect 10406 4167 10464 4193
rect 10506 4227 10564 4253
rect 10506 4193 10518 4227
rect 10552 4193 10564 4227
rect 10506 4167 10564 4193
rect 10606 4227 10664 4253
rect 10606 4193 10618 4227
rect 10652 4193 10664 4227
rect 10606 4167 10664 4193
rect 10706 4227 10764 4253
rect 10706 4193 10718 4227
rect 10752 4193 10764 4227
rect 10706 4167 10764 4193
rect 10806 4227 10864 4253
rect 10806 4193 10818 4227
rect 10852 4193 10864 4227
rect 10806 4167 10864 4193
rect 10906 4227 10964 4253
rect 10906 4193 10912 4227
rect 10952 4193 10964 4227
rect 10906 4167 10964 4193
rect 11006 4227 11064 4253
rect 11006 4193 11018 4227
rect 11058 4193 11064 4227
rect 11006 4167 11064 4193
rect 11106 4227 11164 4253
rect 11106 4193 11118 4227
rect 11152 4193 11164 4227
rect 11106 4167 11164 4193
rect 11206 4227 11264 4253
rect 11206 4193 11218 4227
rect 11252 4193 11264 4227
rect 11206 4167 11264 4193
rect 11306 4227 11364 4253
rect 11306 4193 11312 4227
rect 11352 4193 11364 4227
rect 11306 4167 11364 4193
rect 11406 4227 11464 4253
rect 11406 4193 11418 4227
rect 11458 4193 11464 4227
rect 11406 4167 11464 4193
rect 11506 4227 11564 4253
rect 11506 4193 11512 4227
rect 11552 4193 11564 4227
rect 11506 4167 11564 4193
rect 11606 4227 11664 4253
rect 11606 4193 11618 4227
rect 11658 4193 11664 4227
rect 11606 4167 11664 4193
rect 11706 4227 11764 4253
rect 11706 4193 11718 4227
rect 11752 4193 11764 4227
rect 11706 4167 11764 4193
rect 11806 4227 11864 4253
rect 11806 4193 11818 4227
rect 11852 4193 11864 4227
rect 11806 4167 11864 4193
rect 11906 4227 11964 4253
rect 11906 4193 11918 4227
rect 11952 4193 11964 4227
rect 11906 4167 11964 4193
rect 12006 4227 12064 4253
rect 12006 4193 12018 4227
rect 12052 4193 12064 4227
rect 12006 4167 12064 4193
rect 12106 4227 12164 4253
rect 12106 4193 12118 4227
rect 12152 4193 12164 4227
rect 12106 4167 12164 4193
rect 12206 4227 12264 4253
rect 12206 4193 12218 4227
rect 12252 4193 12264 4227
rect 12206 4167 12264 4193
rect 12306 4227 12364 4253
rect 12306 4193 12318 4227
rect 12352 4193 12364 4227
rect 12306 4167 12364 4193
rect 12406 4227 12464 4253
rect 12406 4193 12418 4227
rect 12452 4193 12464 4227
rect 12406 4167 12464 4193
rect 12506 4227 12564 4253
rect 12506 4193 12518 4227
rect 12552 4193 12564 4227
rect 12506 4167 12564 4193
rect 12606 4227 12664 4253
rect 12606 4193 12618 4227
rect 12652 4193 12664 4227
rect 12606 4167 12664 4193
rect 12706 4227 12764 4253
rect 12706 4193 12718 4227
rect 12752 4193 12764 4227
rect 12706 4167 12764 4193
rect 12806 4227 12864 4253
rect 13018 4246 13262 4280
rect 12806 4193 12818 4227
rect 12852 4193 12864 4227
rect 12908 4208 12916 4242
rect 12958 4208 12974 4242
rect 13018 4227 13052 4246
rect 12806 4167 12864 4193
rect 13228 4243 13262 4246
rect 13228 4227 13362 4243
rect 13018 4177 13052 4193
rect 13096 4178 13112 4212
rect 13154 4178 13162 4212
rect 13262 4193 13328 4227
rect 13228 4177 13362 4193
rect 13428 4227 13562 4243
rect 13462 4193 13528 4227
rect 13428 4177 13562 4193
rect 13628 4227 13662 4243
rect 13628 4177 13662 4193
rect 6 4087 64 4113
rect 6 4053 18 4087
rect 58 4053 64 4087
rect 6 4027 64 4053
rect 106 4087 164 4113
rect 106 4053 118 4087
rect 152 4053 164 4087
rect 106 4027 164 4053
rect 206 4087 264 4113
rect 206 4053 212 4087
rect 252 4053 264 4087
rect 206 4027 264 4053
rect 306 4087 364 4113
rect 306 4053 318 4087
rect 358 4053 364 4087
rect 306 4027 364 4053
rect 406 4087 464 4113
rect 406 4053 412 4087
rect 452 4053 464 4087
rect 406 4027 464 4053
rect 506 4087 564 4113
rect 506 4053 518 4087
rect 558 4053 564 4087
rect 506 4027 564 4053
rect 606 4087 664 4113
rect 606 4053 618 4087
rect 652 4053 664 4087
rect 606 4027 664 4053
rect 706 4087 764 4113
rect 706 4053 718 4087
rect 752 4053 764 4087
rect 706 4027 764 4053
rect 806 4087 864 4113
rect 806 4053 818 4087
rect 852 4053 864 4087
rect 806 4027 864 4053
rect 906 4087 964 4113
rect 906 4053 918 4087
rect 952 4053 964 4087
rect 906 4027 964 4053
rect 1006 4087 1064 4113
rect 1006 4053 1018 4087
rect 1052 4053 1064 4087
rect 1006 4027 1064 4053
rect 1106 4087 1164 4113
rect 1106 4053 1118 4087
rect 1152 4053 1164 4087
rect 1106 4027 1164 4053
rect 1206 4087 1264 4113
rect 1206 4053 1218 4087
rect 1252 4053 1264 4087
rect 1206 4027 1264 4053
rect 1306 4087 1364 4113
rect 1306 4053 1312 4087
rect 1352 4053 1364 4087
rect 1306 4027 1364 4053
rect 1406 4087 1464 4113
rect 1406 4053 1418 4087
rect 1458 4053 1464 4087
rect 1406 4027 1464 4053
rect 1506 4087 1564 4113
rect 1506 4053 1518 4087
rect 1552 4053 1564 4087
rect 1506 4027 1564 4053
rect 1606 4087 1664 4113
rect 1606 4053 1612 4087
rect 1652 4053 1664 4087
rect 1606 4027 1664 4053
rect 1706 4087 1764 4113
rect 1706 4053 1718 4087
rect 1758 4053 1764 4087
rect 1706 4027 1764 4053
rect 1806 4087 1864 4113
rect 1806 4053 1818 4087
rect 1852 4053 1864 4087
rect 1806 4027 1864 4053
rect 1906 4087 1964 4113
rect 1906 4053 1918 4087
rect 1952 4053 1964 4087
rect 1906 4027 1964 4053
rect 2006 4087 2064 4113
rect 2006 4053 2018 4087
rect 2052 4053 2064 4087
rect 2006 4027 2064 4053
rect 2106 4087 2164 4113
rect 2106 4053 2118 4087
rect 2152 4053 2164 4087
rect 2106 4027 2164 4053
rect 2206 4087 2264 4113
rect 2206 4053 2212 4087
rect 2252 4053 2264 4087
rect 2206 4027 2264 4053
rect 2306 4087 2364 4113
rect 2306 4053 2318 4087
rect 2358 4053 2364 4087
rect 2306 4027 2364 4053
rect 2406 4087 2464 4113
rect 2406 4053 2418 4087
rect 2452 4053 2464 4087
rect 2406 4027 2464 4053
rect 2506 4087 2564 4113
rect 2506 4053 2518 4087
rect 2552 4053 2564 4087
rect 2506 4027 2564 4053
rect 2606 4087 2664 4113
rect 2606 4053 2612 4087
rect 2652 4053 2664 4087
rect 2606 4027 2664 4053
rect 2706 4087 2764 4113
rect 2706 4053 2718 4087
rect 2758 4053 2764 4087
rect 2706 4027 2764 4053
rect 2806 4087 2864 4113
rect 2806 4053 2818 4087
rect 2852 4053 2864 4087
rect 2806 4027 2864 4053
rect 2906 4087 2964 4113
rect 2906 4053 2912 4087
rect 2952 4053 2964 4087
rect 2906 4027 2964 4053
rect 3006 4087 3064 4113
rect 3006 4053 3018 4087
rect 3058 4053 3064 4087
rect 3006 4027 3064 4053
rect 3106 4087 3164 4113
rect 3106 4053 3118 4087
rect 3152 4053 3164 4087
rect 3106 4027 3164 4053
rect 3206 4087 3264 4113
rect 3206 4053 3212 4087
rect 3252 4053 3264 4087
rect 3206 4027 3264 4053
rect 3306 4087 3364 4113
rect 3306 4053 3318 4087
rect 3358 4053 3364 4087
rect 3306 4027 3364 4053
rect 3406 4087 3464 4113
rect 3406 4053 3418 4087
rect 3452 4053 3464 4087
rect 3406 4027 3464 4053
rect 3506 4087 3564 4113
rect 3506 4053 3518 4087
rect 3552 4053 3564 4087
rect 3506 4027 3564 4053
rect 3606 4087 3664 4113
rect 3606 4053 3618 4087
rect 3652 4053 3664 4087
rect 3606 4027 3664 4053
rect 3706 4087 3764 4113
rect 3706 4053 3718 4087
rect 3752 4053 3764 4087
rect 3706 4027 3764 4053
rect 3806 4087 3864 4113
rect 3806 4053 3818 4087
rect 3852 4053 3864 4087
rect 3806 4027 3864 4053
rect 3906 4087 3964 4113
rect 3906 4053 3918 4087
rect 3952 4053 3964 4087
rect 3906 4027 3964 4053
rect 4006 4087 4064 4113
rect 4006 4053 4018 4087
rect 4052 4053 4064 4087
rect 4006 4027 4064 4053
rect 4106 4087 4164 4113
rect 4106 4053 4112 4087
rect 4152 4053 4164 4087
rect 4106 4027 4164 4053
rect 4206 4087 4264 4113
rect 4206 4053 4218 4087
rect 4258 4053 4264 4087
rect 4206 4027 4264 4053
rect 4306 4087 4364 4113
rect 4306 4053 4312 4087
rect 4352 4053 4364 4087
rect 4306 4027 4364 4053
rect 4406 4087 4464 4113
rect 4406 4053 4418 4087
rect 4458 4053 4464 4087
rect 4406 4027 4464 4053
rect 4506 4087 4564 4113
rect 4506 4053 4512 4087
rect 4552 4053 4564 4087
rect 4506 4027 4564 4053
rect 4606 4087 4664 4113
rect 4606 4053 4618 4087
rect 4658 4053 4664 4087
rect 4606 4027 4664 4053
rect 4706 4087 4764 4113
rect 4706 4053 4712 4087
rect 4752 4053 4764 4087
rect 4706 4027 4764 4053
rect 4806 4087 4864 4113
rect 4806 4053 4818 4087
rect 4858 4053 4864 4087
rect 4806 4027 4864 4053
rect 4906 4087 4964 4113
rect 4906 4053 4912 4087
rect 4952 4053 4964 4087
rect 4906 4027 4964 4053
rect 5006 4087 5064 4113
rect 5006 4053 5018 4087
rect 5058 4053 5064 4087
rect 5006 4027 5064 4053
rect 5106 4087 5164 4113
rect 5106 4053 5118 4087
rect 5152 4053 5164 4087
rect 5106 4027 5164 4053
rect 5206 4087 5264 4113
rect 5206 4053 5212 4087
rect 5252 4053 5264 4087
rect 5206 4027 5264 4053
rect 5306 4087 5364 4113
rect 5306 4053 5318 4087
rect 5358 4053 5364 4087
rect 5306 4027 5364 4053
rect 5406 4087 5464 4113
rect 5406 4053 5418 4087
rect 5452 4053 5464 4087
rect 5406 4027 5464 4053
rect 5506 4087 5564 4113
rect 5506 4053 5518 4087
rect 5552 4053 5564 4087
rect 5506 4027 5564 4053
rect 5606 4087 5664 4113
rect 5606 4053 5612 4087
rect 5652 4053 5664 4087
rect 5606 4027 5664 4053
rect 5706 4087 5764 4113
rect 5706 4053 5718 4087
rect 5758 4053 5764 4087
rect 5706 4027 5764 4053
rect 5806 4087 5864 4113
rect 5806 4053 5818 4087
rect 5852 4053 5864 4087
rect 5806 4027 5864 4053
rect 5906 4087 5964 4113
rect 5906 4053 5918 4087
rect 5952 4053 5964 4087
rect 5906 4027 5964 4053
rect 6006 4087 6064 4113
rect 6006 4053 6018 4087
rect 6052 4053 6064 4087
rect 6006 4027 6064 4053
rect 6106 4087 6164 4113
rect 6106 4053 6118 4087
rect 6152 4053 6164 4087
rect 6106 4027 6164 4053
rect 6206 4087 6264 4113
rect 6206 4053 6218 4087
rect 6252 4053 6264 4087
rect 6206 4027 6264 4053
rect 6306 4087 6364 4113
rect 6306 4053 6318 4087
rect 6352 4053 6364 4087
rect 6306 4027 6364 4053
rect 6406 4087 6464 4113
rect 6406 4053 6418 4087
rect 6452 4053 6464 4087
rect 6406 4027 6464 4053
rect 6506 4087 6564 4113
rect 6506 4053 6518 4087
rect 6552 4053 6564 4087
rect 6506 4027 6564 4053
rect 6606 4087 6664 4113
rect 6606 4053 6618 4087
rect 6652 4053 6664 4087
rect 6606 4027 6664 4053
rect 6706 4087 6764 4113
rect 6706 4053 6718 4087
rect 6752 4053 6764 4087
rect 6706 4027 6764 4053
rect 6806 4087 6864 4113
rect 6806 4053 6818 4087
rect 6852 4053 6864 4087
rect 6806 4027 6864 4053
rect 6906 4087 6964 4113
rect 6906 4053 6918 4087
rect 6952 4053 6964 4087
rect 6906 4027 6964 4053
rect 7006 4087 7064 4113
rect 7006 4053 7018 4087
rect 7052 4053 7064 4087
rect 7006 4027 7064 4053
rect 7106 4087 7164 4113
rect 7106 4053 7118 4087
rect 7152 4053 7164 4087
rect 7106 4027 7164 4053
rect 7206 4087 7264 4113
rect 7206 4053 7218 4087
rect 7252 4053 7264 4087
rect 7206 4027 7264 4053
rect 7306 4087 7364 4113
rect 7306 4053 7312 4087
rect 7352 4053 7364 4087
rect 7306 4027 7364 4053
rect 7406 4087 7464 4113
rect 7406 4053 7418 4087
rect 7458 4053 7464 4087
rect 7406 4027 7464 4053
rect 7506 4087 7564 4113
rect 7506 4053 7518 4087
rect 7552 4053 7564 4087
rect 7506 4027 7564 4053
rect 7606 4087 7664 4113
rect 7606 4053 7612 4087
rect 7652 4053 7664 4087
rect 7606 4027 7664 4053
rect 7706 4087 7764 4113
rect 7706 4053 7718 4087
rect 7758 4053 7764 4087
rect 7706 4027 7764 4053
rect 7806 4087 7864 4113
rect 7806 4053 7812 4087
rect 7852 4053 7864 4087
rect 7806 4027 7864 4053
rect 7906 4087 7964 4113
rect 7906 4053 7918 4087
rect 7958 4053 7964 4087
rect 7906 4027 7964 4053
rect 8006 4087 8064 4113
rect 8006 4053 8018 4087
rect 8052 4053 8064 4087
rect 8006 4027 8064 4053
rect 8106 4087 8164 4113
rect 8106 4053 8118 4087
rect 8152 4053 8164 4087
rect 8106 4027 8164 4053
rect 8206 4087 8264 4113
rect 8206 4053 8218 4087
rect 8252 4053 8264 4087
rect 8206 4027 8264 4053
rect 8306 4087 8364 4113
rect 8306 4053 8318 4087
rect 8352 4053 8364 4087
rect 8306 4027 8364 4053
rect 8406 4087 8464 4113
rect 8406 4053 8418 4087
rect 8452 4053 8464 4087
rect 8406 4027 8464 4053
rect 8506 4087 8564 4113
rect 8506 4053 8518 4087
rect 8552 4053 8564 4087
rect 8506 4027 8564 4053
rect 8606 4087 8664 4113
rect 8606 4053 8618 4087
rect 8652 4053 8664 4087
rect 8606 4027 8664 4053
rect 8706 4087 8764 4113
rect 8706 4053 8712 4087
rect 8752 4053 8764 4087
rect 8706 4027 8764 4053
rect 8806 4087 8864 4113
rect 8806 4053 8818 4087
rect 8858 4053 8864 4087
rect 8806 4027 8864 4053
rect 8906 4087 8964 4113
rect 8906 4053 8912 4087
rect 8952 4053 8964 4087
rect 8906 4027 8964 4053
rect 9006 4087 9064 4113
rect 9006 4053 9018 4087
rect 9058 4053 9064 4087
rect 9006 4027 9064 4053
rect 9106 4087 9164 4113
rect 9106 4053 9118 4087
rect 9152 4053 9164 4087
rect 9106 4027 9164 4053
rect 9206 4087 9264 4113
rect 9206 4053 9218 4087
rect 9252 4053 9264 4087
rect 9206 4027 9264 4053
rect 9306 4087 9364 4113
rect 9306 4053 9318 4087
rect 9352 4053 9364 4087
rect 9306 4027 9364 4053
rect 9406 4087 9464 4113
rect 9406 4053 9418 4087
rect 9452 4053 9464 4087
rect 9406 4027 9464 4053
rect 9506 4087 9564 4113
rect 9506 4053 9512 4087
rect 9552 4053 9564 4087
rect 9506 4027 9564 4053
rect 9606 4087 9664 4113
rect 9606 4053 9618 4087
rect 9658 4053 9664 4087
rect 9606 4027 9664 4053
rect 9706 4087 9764 4113
rect 9706 4053 9718 4087
rect 9752 4053 9764 4087
rect 9706 4027 9764 4053
rect 9806 4087 9864 4113
rect 9806 4053 9818 4087
rect 9852 4053 9864 4087
rect 9806 4027 9864 4053
rect 9906 4087 9964 4113
rect 9906 4053 9918 4087
rect 9952 4053 9964 4087
rect 9906 4027 9964 4053
rect 10006 4087 10064 4113
rect 10006 4053 10018 4087
rect 10052 4053 10064 4087
rect 10006 4027 10064 4053
rect 10106 4087 10164 4113
rect 10106 4053 10118 4087
rect 10152 4053 10164 4087
rect 10106 4027 10164 4053
rect 10206 4087 10264 4113
rect 10206 4053 10218 4087
rect 10252 4053 10264 4087
rect 10206 4027 10264 4053
rect 10306 4087 10364 4113
rect 10306 4053 10318 4087
rect 10352 4053 10364 4087
rect 10306 4027 10364 4053
rect 10406 4087 10464 4113
rect 10406 4053 10418 4087
rect 10452 4053 10464 4087
rect 10406 4027 10464 4053
rect 10506 4087 10564 4113
rect 10506 4053 10518 4087
rect 10552 4053 10564 4087
rect 10506 4027 10564 4053
rect 10606 4087 10664 4113
rect 10606 4053 10612 4087
rect 10652 4053 10664 4087
rect 10606 4027 10664 4053
rect 10706 4087 10764 4113
rect 10706 4053 10718 4087
rect 10758 4053 10764 4087
rect 10706 4027 10764 4053
rect 10806 4087 10864 4113
rect 10806 4053 10812 4087
rect 10852 4053 10864 4087
rect 10806 4027 10864 4053
rect 10906 4087 10964 4113
rect 10906 4053 10918 4087
rect 10958 4053 10964 4087
rect 10906 4027 10964 4053
rect 11006 4087 11064 4113
rect 11006 4053 11018 4087
rect 11052 4053 11064 4087
rect 11006 4027 11064 4053
rect 11106 4087 11164 4113
rect 11106 4053 11118 4087
rect 11152 4053 11164 4087
rect 11106 4027 11164 4053
rect 11206 4087 11264 4113
rect 11206 4053 11218 4087
rect 11252 4053 11264 4087
rect 11206 4027 11264 4053
rect 11306 4087 11364 4113
rect 11306 4053 11312 4087
rect 11352 4053 11364 4087
rect 11306 4027 11364 4053
rect 11406 4087 11464 4113
rect 11406 4053 11418 4087
rect 11458 4053 11464 4087
rect 11406 4027 11464 4053
rect 11506 4087 11564 4113
rect 11506 4053 11512 4087
rect 11552 4053 11564 4087
rect 11506 4027 11564 4053
rect 11606 4087 11664 4113
rect 11606 4053 11618 4087
rect 11658 4053 11664 4087
rect 11606 4027 11664 4053
rect 11706 4087 11764 4113
rect 11706 4053 11718 4087
rect 11752 4053 11764 4087
rect 11706 4027 11764 4053
rect 11806 4087 11864 4113
rect 11806 4053 11812 4087
rect 11852 4053 11864 4087
rect 11806 4027 11864 4053
rect 11906 4087 11964 4113
rect 11906 4053 11918 4087
rect 11958 4053 11964 4087
rect 11906 4027 11964 4053
rect 12006 4087 12064 4113
rect 12006 4053 12018 4087
rect 12052 4053 12064 4087
rect 12006 4027 12064 4053
rect 12106 4087 12164 4113
rect 12106 4053 12118 4087
rect 12152 4053 12164 4087
rect 12106 4027 12164 4053
rect 12206 4087 12264 4113
rect 12206 4053 12218 4087
rect 12252 4053 12264 4087
rect 12206 4027 12264 4053
rect 12306 4087 12364 4113
rect 12306 4053 12318 4087
rect 12352 4053 12364 4087
rect 12306 4027 12364 4053
rect 12406 4087 12464 4113
rect 12406 4053 12418 4087
rect 12452 4053 12464 4087
rect 12406 4027 12464 4053
rect 12506 4087 12564 4113
rect 12506 4053 12518 4087
rect 12552 4053 12564 4087
rect 12506 4027 12564 4053
rect 12606 4087 12664 4113
rect 12606 4053 12612 4087
rect 12652 4053 12664 4087
rect 12606 4027 12664 4053
rect 12706 4087 12764 4113
rect 12706 4053 12718 4087
rect 12758 4053 12764 4087
rect 12706 4027 12764 4053
rect 12806 4087 12864 4113
rect 13018 4106 13262 4140
rect 12806 4053 12812 4087
rect 12852 4053 12864 4087
rect 12908 4068 12916 4102
rect 12958 4068 12974 4102
rect 13018 4087 13052 4106
rect 12806 4027 12864 4053
rect 13228 4087 13262 4106
rect 13018 4037 13052 4053
rect 13096 4038 13112 4072
rect 13154 4038 13162 4072
rect 13228 4037 13262 4053
rect 13328 4087 13562 4103
rect 13362 4053 13428 4087
rect 13462 4053 13528 4087
rect 13328 4037 13562 4053
rect 13628 4087 13662 4103
rect 13628 4037 13662 4053
rect 6 3947 64 3973
rect 6 3913 18 3947
rect 58 3913 64 3947
rect 6 3887 64 3913
rect 106 3947 164 3973
rect 106 3913 118 3947
rect 152 3913 164 3947
rect 106 3887 164 3913
rect 206 3947 264 3973
rect 206 3913 218 3947
rect 252 3913 264 3947
rect 206 3887 264 3913
rect 306 3947 364 3973
rect 306 3913 318 3947
rect 352 3913 364 3947
rect 306 3887 364 3913
rect 406 3947 464 3973
rect 406 3913 418 3947
rect 452 3913 464 3947
rect 406 3887 464 3913
rect 506 3947 564 3973
rect 506 3913 518 3947
rect 552 3913 564 3947
rect 506 3887 564 3913
rect 606 3947 664 3973
rect 606 3913 618 3947
rect 652 3913 664 3947
rect 606 3887 664 3913
rect 706 3947 764 3973
rect 706 3913 718 3947
rect 752 3913 764 3947
rect 706 3887 764 3913
rect 806 3947 864 3973
rect 806 3913 818 3947
rect 852 3913 864 3947
rect 806 3887 864 3913
rect 906 3947 964 3973
rect 906 3913 918 3947
rect 952 3913 964 3947
rect 906 3887 964 3913
rect 1006 3947 1064 3973
rect 1006 3913 1018 3947
rect 1052 3913 1064 3947
rect 1006 3887 1064 3913
rect 1106 3947 1164 3973
rect 1106 3913 1118 3947
rect 1152 3913 1164 3947
rect 1106 3887 1164 3913
rect 1206 3947 1264 3973
rect 1206 3913 1218 3947
rect 1252 3913 1264 3947
rect 1206 3887 1264 3913
rect 1306 3947 1364 3973
rect 1306 3913 1318 3947
rect 1352 3913 1364 3947
rect 1306 3887 1364 3913
rect 1406 3947 1464 3973
rect 1406 3913 1418 3947
rect 1452 3913 1464 3947
rect 1406 3887 1464 3913
rect 1506 3947 1564 3973
rect 1506 3913 1518 3947
rect 1552 3913 1564 3947
rect 1506 3887 1564 3913
rect 1606 3947 1664 3973
rect 1606 3913 1618 3947
rect 1652 3913 1664 3947
rect 1606 3887 1664 3913
rect 1706 3947 1764 3973
rect 1706 3913 1718 3947
rect 1752 3913 1764 3947
rect 1706 3887 1764 3913
rect 1806 3947 1864 3973
rect 1806 3913 1818 3947
rect 1852 3913 1864 3947
rect 1806 3887 1864 3913
rect 1906 3947 1964 3973
rect 1906 3913 1912 3947
rect 1952 3913 1964 3947
rect 1906 3887 1964 3913
rect 2006 3947 2064 3973
rect 2006 3913 2018 3947
rect 2058 3913 2064 3947
rect 2006 3887 2064 3913
rect 2106 3947 2164 3973
rect 2106 3913 2118 3947
rect 2152 3913 2164 3947
rect 2106 3887 2164 3913
rect 2206 3947 2264 3973
rect 2206 3913 2218 3947
rect 2252 3913 2264 3947
rect 2206 3887 2264 3913
rect 2306 3947 2364 3973
rect 2306 3913 2318 3947
rect 2352 3913 2364 3947
rect 2306 3887 2364 3913
rect 2406 3947 2464 3973
rect 2406 3913 2418 3947
rect 2452 3913 2464 3947
rect 2406 3887 2464 3913
rect 2506 3947 2564 3973
rect 2506 3913 2518 3947
rect 2552 3913 2564 3947
rect 2506 3887 2564 3913
rect 2606 3947 2664 3973
rect 2606 3913 2618 3947
rect 2652 3913 2664 3947
rect 2606 3887 2664 3913
rect 2706 3947 2764 3973
rect 2706 3913 2718 3947
rect 2752 3913 2764 3947
rect 2706 3887 2764 3913
rect 2806 3947 2864 3973
rect 2806 3913 2818 3947
rect 2852 3913 2864 3947
rect 2806 3887 2864 3913
rect 2906 3947 2964 3973
rect 2906 3913 2918 3947
rect 2952 3913 2964 3947
rect 2906 3887 2964 3913
rect 3006 3947 3064 3973
rect 3006 3913 3018 3947
rect 3052 3913 3064 3947
rect 3006 3887 3064 3913
rect 3106 3947 3164 3973
rect 3106 3913 3118 3947
rect 3152 3913 3164 3947
rect 3106 3887 3164 3913
rect 3206 3947 3264 3973
rect 3206 3913 3218 3947
rect 3252 3913 3264 3947
rect 3206 3887 3264 3913
rect 3306 3947 3364 3973
rect 3306 3913 3318 3947
rect 3352 3913 3364 3947
rect 3306 3887 3364 3913
rect 3406 3947 3464 3973
rect 3406 3913 3418 3947
rect 3452 3913 3464 3947
rect 3406 3887 3464 3913
rect 3506 3947 3564 3973
rect 3506 3913 3518 3947
rect 3552 3913 3564 3947
rect 3506 3887 3564 3913
rect 3606 3947 3664 3973
rect 3606 3913 3618 3947
rect 3652 3913 3664 3947
rect 3606 3887 3664 3913
rect 3706 3947 3764 3973
rect 3706 3913 3718 3947
rect 3752 3913 3764 3947
rect 3706 3887 3764 3913
rect 3806 3947 3864 3973
rect 3806 3913 3818 3947
rect 3852 3913 3864 3947
rect 3806 3887 3864 3913
rect 3906 3947 3964 3973
rect 3906 3913 3912 3947
rect 3952 3913 3964 3947
rect 3906 3887 3964 3913
rect 4006 3947 4064 3973
rect 4006 3913 4018 3947
rect 4058 3913 4064 3947
rect 4006 3887 4064 3913
rect 4106 3947 4164 3973
rect 4106 3913 4112 3947
rect 4152 3913 4164 3947
rect 4106 3887 4164 3913
rect 4206 3947 4264 3973
rect 4206 3913 4218 3947
rect 4258 3913 4264 3947
rect 4206 3887 4264 3913
rect 4306 3947 4364 3973
rect 4306 3913 4318 3947
rect 4352 3913 4364 3947
rect 4306 3887 4364 3913
rect 4406 3947 4464 3973
rect 4406 3913 4418 3947
rect 4452 3913 4464 3947
rect 4406 3887 4464 3913
rect 4506 3947 4564 3973
rect 4506 3913 4518 3947
rect 4552 3913 4564 3947
rect 4506 3887 4564 3913
rect 4606 3947 4664 3973
rect 4606 3913 4618 3947
rect 4652 3913 4664 3947
rect 4606 3887 4664 3913
rect 4706 3947 4764 3973
rect 4706 3913 4718 3947
rect 4752 3913 4764 3947
rect 4706 3887 4764 3913
rect 4806 3947 4864 3973
rect 4806 3913 4818 3947
rect 4852 3913 4864 3947
rect 4806 3887 4864 3913
rect 4906 3947 4964 3973
rect 4906 3913 4918 3947
rect 4952 3913 4964 3947
rect 4906 3887 4964 3913
rect 5006 3947 5064 3973
rect 5006 3913 5012 3947
rect 5052 3913 5064 3947
rect 5006 3887 5064 3913
rect 5106 3947 5164 3973
rect 5106 3913 5118 3947
rect 5158 3913 5164 3947
rect 5106 3887 5164 3913
rect 5206 3947 5264 3973
rect 5206 3913 5212 3947
rect 5252 3913 5264 3947
rect 5206 3887 5264 3913
rect 5306 3947 5364 3973
rect 5306 3913 5318 3947
rect 5358 3913 5364 3947
rect 5306 3887 5364 3913
rect 5406 3947 5464 3973
rect 5406 3913 5418 3947
rect 5452 3913 5464 3947
rect 5406 3887 5464 3913
rect 5506 3947 5564 3973
rect 5506 3913 5512 3947
rect 5552 3913 5564 3947
rect 5506 3887 5564 3913
rect 5606 3947 5664 3973
rect 5606 3913 5618 3947
rect 5658 3913 5664 3947
rect 5606 3887 5664 3913
rect 5706 3947 5764 3973
rect 5706 3913 5718 3947
rect 5752 3913 5764 3947
rect 5706 3887 5764 3913
rect 5806 3947 5864 3973
rect 5806 3913 5818 3947
rect 5852 3913 5864 3947
rect 5806 3887 5864 3913
rect 5906 3947 5964 3973
rect 5906 3913 5912 3947
rect 5952 3913 5964 3947
rect 5906 3887 5964 3913
rect 6006 3947 6064 3973
rect 6006 3913 6018 3947
rect 6058 3913 6064 3947
rect 6006 3887 6064 3913
rect 6106 3947 6164 3973
rect 6106 3913 6118 3947
rect 6152 3913 6164 3947
rect 6106 3887 6164 3913
rect 6206 3947 6264 3973
rect 6206 3913 6218 3947
rect 6252 3913 6264 3947
rect 6206 3887 6264 3913
rect 6306 3947 6364 3973
rect 6306 3913 6318 3947
rect 6352 3913 6364 3947
rect 6306 3887 6364 3913
rect 6406 3947 6464 3973
rect 6406 3913 6418 3947
rect 6452 3913 6464 3947
rect 6406 3887 6464 3913
rect 6506 3947 6564 3973
rect 6506 3913 6518 3947
rect 6552 3913 6564 3947
rect 6506 3887 6564 3913
rect 6606 3947 6664 3973
rect 6606 3913 6618 3947
rect 6652 3913 6664 3947
rect 6606 3887 6664 3913
rect 6706 3947 6764 3973
rect 6706 3913 6718 3947
rect 6752 3913 6764 3947
rect 6706 3887 6764 3913
rect 6806 3947 6864 3973
rect 6806 3913 6818 3947
rect 6852 3913 6864 3947
rect 6806 3887 6864 3913
rect 6906 3947 6964 3973
rect 6906 3913 6912 3947
rect 6952 3913 6964 3947
rect 6906 3887 6964 3913
rect 7006 3947 7064 3973
rect 7006 3913 7018 3947
rect 7058 3913 7064 3947
rect 7006 3887 7064 3913
rect 7106 3947 7164 3973
rect 7106 3913 7112 3947
rect 7152 3913 7164 3947
rect 7106 3887 7164 3913
rect 7206 3947 7264 3973
rect 7206 3913 7218 3947
rect 7258 3913 7264 3947
rect 7206 3887 7264 3913
rect 7306 3947 7364 3973
rect 7306 3913 7318 3947
rect 7352 3913 7364 3947
rect 7306 3887 7364 3913
rect 7406 3947 7464 3973
rect 7406 3913 7418 3947
rect 7452 3913 7464 3947
rect 7406 3887 7464 3913
rect 7506 3947 7564 3973
rect 7506 3913 7518 3947
rect 7552 3913 7564 3947
rect 7506 3887 7564 3913
rect 7606 3947 7664 3973
rect 7606 3913 7618 3947
rect 7652 3913 7664 3947
rect 7606 3887 7664 3913
rect 7706 3947 7764 3973
rect 7706 3913 7718 3947
rect 7752 3913 7764 3947
rect 7706 3887 7764 3913
rect 7806 3947 7864 3973
rect 7806 3913 7818 3947
rect 7852 3913 7864 3947
rect 7806 3887 7864 3913
rect 7906 3947 7964 3973
rect 7906 3913 7918 3947
rect 7952 3913 7964 3947
rect 7906 3887 7964 3913
rect 8006 3947 8064 3973
rect 8006 3913 8018 3947
rect 8052 3913 8064 3947
rect 8006 3887 8064 3913
rect 8106 3947 8164 3973
rect 8106 3913 8118 3947
rect 8152 3913 8164 3947
rect 8106 3887 8164 3913
rect 8206 3947 8264 3973
rect 8206 3913 8218 3947
rect 8252 3913 8264 3947
rect 8206 3887 8264 3913
rect 8306 3947 8364 3973
rect 8306 3913 8318 3947
rect 8352 3913 8364 3947
rect 8306 3887 8364 3913
rect 8406 3947 8464 3973
rect 8406 3913 8418 3947
rect 8452 3913 8464 3947
rect 8406 3887 8464 3913
rect 8506 3947 8564 3973
rect 8506 3913 8518 3947
rect 8552 3913 8564 3947
rect 8506 3887 8564 3913
rect 8606 3947 8664 3973
rect 8606 3913 8618 3947
rect 8652 3913 8664 3947
rect 8606 3887 8664 3913
rect 8706 3947 8764 3973
rect 8706 3913 8712 3947
rect 8752 3913 8764 3947
rect 8706 3887 8764 3913
rect 8806 3947 8864 3973
rect 8806 3913 8818 3947
rect 8858 3913 8864 3947
rect 8806 3887 8864 3913
rect 8906 3947 8964 3973
rect 8906 3913 8918 3947
rect 8952 3913 8964 3947
rect 8906 3887 8964 3913
rect 9006 3947 9064 3973
rect 9006 3913 9018 3947
rect 9052 3913 9064 3947
rect 9006 3887 9064 3913
rect 9106 3947 9164 3973
rect 9106 3913 9118 3947
rect 9152 3913 9164 3947
rect 9106 3887 9164 3913
rect 9206 3947 9264 3973
rect 9206 3913 9218 3947
rect 9252 3913 9264 3947
rect 9206 3887 9264 3913
rect 9306 3947 9364 3973
rect 9306 3913 9318 3947
rect 9352 3913 9364 3947
rect 9306 3887 9364 3913
rect 9406 3947 9464 3973
rect 9406 3913 9418 3947
rect 9452 3913 9464 3947
rect 9406 3887 9464 3913
rect 9506 3947 9564 3973
rect 9506 3913 9512 3947
rect 9552 3913 9564 3947
rect 9506 3887 9564 3913
rect 9606 3947 9664 3973
rect 9606 3913 9618 3947
rect 9658 3913 9664 3947
rect 9606 3887 9664 3913
rect 9706 3947 9764 3973
rect 9706 3913 9718 3947
rect 9752 3913 9764 3947
rect 9706 3887 9764 3913
rect 9806 3947 9864 3973
rect 9806 3913 9818 3947
rect 9852 3913 9864 3947
rect 9806 3887 9864 3913
rect 9906 3947 9964 3973
rect 9906 3913 9918 3947
rect 9952 3913 9964 3947
rect 9906 3887 9964 3913
rect 10006 3947 10064 3973
rect 10006 3913 10018 3947
rect 10052 3913 10064 3947
rect 10006 3887 10064 3913
rect 10106 3947 10164 3973
rect 10106 3913 10118 3947
rect 10152 3913 10164 3947
rect 10106 3887 10164 3913
rect 10206 3947 10264 3973
rect 10206 3913 10218 3947
rect 10252 3913 10264 3947
rect 10206 3887 10264 3913
rect 10306 3947 10364 3973
rect 10306 3913 10318 3947
rect 10352 3913 10364 3947
rect 10306 3887 10364 3913
rect 10406 3947 10464 3973
rect 10406 3913 10418 3947
rect 10452 3913 10464 3947
rect 10406 3887 10464 3913
rect 10506 3947 10564 3973
rect 10506 3913 10518 3947
rect 10552 3913 10564 3947
rect 10506 3887 10564 3913
rect 10606 3947 10664 3973
rect 10606 3913 10618 3947
rect 10652 3913 10664 3947
rect 10606 3887 10664 3913
rect 10706 3947 10764 3973
rect 10706 3913 10718 3947
rect 10752 3913 10764 3947
rect 10706 3887 10764 3913
rect 10806 3947 10864 3973
rect 10806 3913 10818 3947
rect 10852 3913 10864 3947
rect 10806 3887 10864 3913
rect 10906 3947 10964 3973
rect 10906 3913 10918 3947
rect 10952 3913 10964 3947
rect 10906 3887 10964 3913
rect 11006 3947 11064 3973
rect 11006 3913 11012 3947
rect 11052 3913 11064 3947
rect 11006 3887 11064 3913
rect 11106 3947 11164 3973
rect 11106 3913 11118 3947
rect 11158 3913 11164 3947
rect 11106 3887 11164 3913
rect 11206 3947 11264 3973
rect 11206 3913 11218 3947
rect 11252 3913 11264 3947
rect 11206 3887 11264 3913
rect 11306 3947 11364 3973
rect 11306 3913 11318 3947
rect 11352 3913 11364 3947
rect 11306 3887 11364 3913
rect 11406 3947 11464 3973
rect 11406 3913 11418 3947
rect 11452 3913 11464 3947
rect 11406 3887 11464 3913
rect 11506 3947 11564 3973
rect 11506 3913 11518 3947
rect 11552 3913 11564 3947
rect 11506 3887 11564 3913
rect 11606 3947 11664 3973
rect 11606 3913 11618 3947
rect 11652 3913 11664 3947
rect 11606 3887 11664 3913
rect 11706 3947 11764 3973
rect 11706 3913 11718 3947
rect 11752 3913 11764 3947
rect 11706 3887 11764 3913
rect 11806 3947 11864 3973
rect 11806 3913 11818 3947
rect 11852 3913 11864 3947
rect 11806 3887 11864 3913
rect 11906 3947 11964 3973
rect 11906 3913 11918 3947
rect 11952 3913 11964 3947
rect 11906 3887 11964 3913
rect 12006 3947 12064 3973
rect 12006 3913 12018 3947
rect 12052 3913 12064 3947
rect 12006 3887 12064 3913
rect 12106 3947 12164 3973
rect 12106 3913 12118 3947
rect 12152 3913 12164 3947
rect 12106 3887 12164 3913
rect 12206 3947 12264 3973
rect 12206 3913 12218 3947
rect 12252 3913 12264 3947
rect 12206 3887 12264 3913
rect 12306 3947 12364 3973
rect 12306 3913 12318 3947
rect 12352 3913 12364 3947
rect 12306 3887 12364 3913
rect 12406 3947 12464 3973
rect 12406 3913 12418 3947
rect 12452 3913 12464 3947
rect 12406 3887 12464 3913
rect 12506 3947 12564 3973
rect 12506 3913 12518 3947
rect 12552 3913 12564 3947
rect 12506 3887 12564 3913
rect 12606 3947 12664 3973
rect 12606 3913 12618 3947
rect 12652 3913 12664 3947
rect 12606 3887 12664 3913
rect 12706 3947 12764 3973
rect 12706 3913 12718 3947
rect 12752 3913 12764 3947
rect 12706 3887 12764 3913
rect 12806 3947 12864 3973
rect 13018 3966 13262 4000
rect 12806 3913 12812 3947
rect 12852 3913 12864 3947
rect 12908 3928 12916 3962
rect 12958 3928 12974 3962
rect 13018 3947 13052 3966
rect 12806 3887 12864 3913
rect 13228 3963 13262 3966
rect 13228 3947 13362 3963
rect 13018 3897 13052 3913
rect 13096 3898 13112 3932
rect 13154 3898 13162 3932
rect 13262 3913 13328 3947
rect 13228 3897 13362 3913
rect 13428 3947 13462 3963
rect 13428 3897 13462 3913
rect 13528 3947 13662 3963
rect 13562 3913 13628 3947
rect 13528 3897 13662 3913
rect 6 3807 64 3833
rect 6 3773 18 3807
rect 58 3773 64 3807
rect 6 3747 64 3773
rect 106 3807 164 3833
rect 106 3773 118 3807
rect 152 3773 164 3807
rect 106 3747 164 3773
rect 206 3807 264 3833
rect 206 3773 218 3807
rect 252 3773 264 3807
rect 206 3747 264 3773
rect 306 3807 364 3833
rect 306 3773 318 3807
rect 352 3773 364 3807
rect 306 3747 364 3773
rect 406 3807 464 3833
rect 406 3773 418 3807
rect 452 3773 464 3807
rect 406 3747 464 3773
rect 506 3807 564 3833
rect 506 3773 518 3807
rect 552 3773 564 3807
rect 506 3747 564 3773
rect 606 3807 664 3833
rect 606 3773 618 3807
rect 652 3773 664 3807
rect 606 3747 664 3773
rect 706 3807 764 3833
rect 706 3773 718 3807
rect 752 3773 764 3807
rect 706 3747 764 3773
rect 806 3807 864 3833
rect 806 3773 818 3807
rect 852 3773 864 3807
rect 806 3747 864 3773
rect 906 3807 964 3833
rect 906 3773 918 3807
rect 952 3773 964 3807
rect 906 3747 964 3773
rect 1006 3807 1064 3833
rect 1006 3773 1018 3807
rect 1052 3773 1064 3807
rect 1006 3747 1064 3773
rect 1106 3807 1164 3833
rect 1106 3773 1118 3807
rect 1152 3773 1164 3807
rect 1106 3747 1164 3773
rect 1206 3807 1264 3833
rect 1206 3773 1218 3807
rect 1252 3773 1264 3807
rect 1206 3747 1264 3773
rect 1306 3807 1364 3833
rect 1306 3773 1318 3807
rect 1352 3773 1364 3807
rect 1306 3747 1364 3773
rect 1406 3807 1464 3833
rect 1406 3773 1418 3807
rect 1452 3773 1464 3807
rect 1406 3747 1464 3773
rect 1506 3807 1564 3833
rect 1506 3773 1518 3807
rect 1552 3773 1564 3807
rect 1506 3747 1564 3773
rect 1606 3807 1664 3833
rect 1606 3773 1618 3807
rect 1652 3773 1664 3807
rect 1606 3747 1664 3773
rect 1706 3807 1764 3833
rect 1706 3773 1718 3807
rect 1752 3773 1764 3807
rect 1706 3747 1764 3773
rect 1806 3807 1864 3833
rect 1806 3773 1818 3807
rect 1852 3773 1864 3807
rect 1806 3747 1864 3773
rect 1906 3807 1964 3833
rect 1906 3773 1918 3807
rect 1952 3773 1964 3807
rect 1906 3747 1964 3773
rect 2006 3807 2064 3833
rect 2006 3773 2018 3807
rect 2052 3773 2064 3807
rect 2006 3747 2064 3773
rect 2106 3807 2164 3833
rect 2106 3773 2112 3807
rect 2152 3773 2164 3807
rect 2106 3747 2164 3773
rect 2206 3807 2264 3833
rect 2206 3773 2218 3807
rect 2258 3773 2264 3807
rect 2206 3747 2264 3773
rect 2306 3807 2364 3833
rect 2306 3773 2318 3807
rect 2352 3773 2364 3807
rect 2306 3747 2364 3773
rect 2406 3807 2464 3833
rect 2406 3773 2418 3807
rect 2452 3773 2464 3807
rect 2406 3747 2464 3773
rect 2506 3807 2564 3833
rect 2506 3773 2512 3807
rect 2552 3773 2564 3807
rect 2506 3747 2564 3773
rect 2606 3807 2664 3833
rect 2606 3773 2618 3807
rect 2658 3773 2664 3807
rect 2606 3747 2664 3773
rect 2706 3807 2764 3833
rect 2706 3773 2712 3807
rect 2752 3773 2764 3807
rect 2706 3747 2764 3773
rect 2806 3807 2864 3833
rect 2806 3773 2818 3807
rect 2858 3773 2864 3807
rect 2806 3747 2864 3773
rect 2906 3807 2964 3833
rect 2906 3773 2918 3807
rect 2952 3773 2964 3807
rect 2906 3747 2964 3773
rect 3006 3807 3064 3833
rect 3006 3773 3018 3807
rect 3052 3773 3064 3807
rect 3006 3747 3064 3773
rect 3106 3807 3164 3833
rect 3106 3773 3112 3807
rect 3152 3773 3164 3807
rect 3106 3747 3164 3773
rect 3206 3807 3264 3833
rect 3206 3773 3218 3807
rect 3258 3773 3264 3807
rect 3206 3747 3264 3773
rect 3306 3807 3364 3833
rect 3306 3773 3318 3807
rect 3352 3773 3364 3807
rect 3306 3747 3364 3773
rect 3406 3807 3464 3833
rect 3406 3773 3418 3807
rect 3452 3773 3464 3807
rect 3406 3747 3464 3773
rect 3506 3807 3564 3833
rect 3506 3773 3518 3807
rect 3552 3773 3564 3807
rect 3506 3747 3564 3773
rect 3606 3807 3664 3833
rect 3606 3773 3618 3807
rect 3652 3773 3664 3807
rect 3606 3747 3664 3773
rect 3706 3807 3764 3833
rect 3706 3773 3718 3807
rect 3752 3773 3764 3807
rect 3706 3747 3764 3773
rect 3806 3807 3864 3833
rect 3806 3773 3818 3807
rect 3852 3773 3864 3807
rect 3806 3747 3864 3773
rect 3906 3807 3964 3833
rect 3906 3773 3918 3807
rect 3952 3773 3964 3807
rect 3906 3747 3964 3773
rect 4006 3807 4064 3833
rect 4006 3773 4018 3807
rect 4052 3773 4064 3807
rect 4006 3747 4064 3773
rect 4106 3807 4164 3833
rect 4106 3773 4118 3807
rect 4152 3773 4164 3807
rect 4106 3747 4164 3773
rect 4206 3807 4264 3833
rect 4206 3773 4218 3807
rect 4252 3773 4264 3807
rect 4206 3747 4264 3773
rect 4306 3807 4364 3833
rect 4306 3773 4318 3807
rect 4352 3773 4364 3807
rect 4306 3747 4364 3773
rect 4406 3807 4464 3833
rect 4406 3773 4418 3807
rect 4452 3773 4464 3807
rect 4406 3747 4464 3773
rect 4506 3807 4564 3833
rect 4506 3773 4512 3807
rect 4552 3773 4564 3807
rect 4506 3747 4564 3773
rect 4606 3807 4664 3833
rect 4606 3773 4618 3807
rect 4658 3773 4664 3807
rect 4606 3747 4664 3773
rect 4706 3807 4764 3833
rect 4706 3773 4718 3807
rect 4752 3773 4764 3807
rect 4706 3747 4764 3773
rect 4806 3807 4864 3833
rect 4806 3773 4818 3807
rect 4852 3773 4864 3807
rect 4806 3747 4864 3773
rect 4906 3807 4964 3833
rect 4906 3773 4918 3807
rect 4952 3773 4964 3807
rect 4906 3747 4964 3773
rect 5006 3807 5064 3833
rect 5006 3773 5018 3807
rect 5052 3773 5064 3807
rect 5006 3747 5064 3773
rect 5106 3807 5164 3833
rect 5106 3773 5118 3807
rect 5152 3773 5164 3807
rect 5106 3747 5164 3773
rect 5206 3807 5264 3833
rect 5206 3773 5218 3807
rect 5252 3773 5264 3807
rect 5206 3747 5264 3773
rect 5306 3807 5364 3833
rect 5306 3773 5318 3807
rect 5352 3773 5364 3807
rect 5306 3747 5364 3773
rect 5406 3807 5464 3833
rect 5406 3773 5412 3807
rect 5452 3773 5464 3807
rect 5406 3747 5464 3773
rect 5506 3807 5564 3833
rect 5506 3773 5518 3807
rect 5558 3773 5564 3807
rect 5506 3747 5564 3773
rect 5606 3807 5664 3833
rect 5606 3773 5618 3807
rect 5652 3773 5664 3807
rect 5606 3747 5664 3773
rect 5706 3807 5764 3833
rect 5706 3773 5718 3807
rect 5752 3773 5764 3807
rect 5706 3747 5764 3773
rect 5806 3807 5864 3833
rect 5806 3773 5818 3807
rect 5852 3773 5864 3807
rect 5806 3747 5864 3773
rect 5906 3807 5964 3833
rect 5906 3773 5912 3807
rect 5952 3773 5964 3807
rect 5906 3747 5964 3773
rect 6006 3807 6064 3833
rect 6006 3773 6018 3807
rect 6058 3773 6064 3807
rect 6006 3747 6064 3773
rect 6106 3807 6164 3833
rect 6106 3773 6118 3807
rect 6152 3773 6164 3807
rect 6106 3747 6164 3773
rect 6206 3807 6264 3833
rect 6206 3773 6218 3807
rect 6252 3773 6264 3807
rect 6206 3747 6264 3773
rect 6306 3807 6364 3833
rect 6306 3773 6318 3807
rect 6352 3773 6364 3807
rect 6306 3747 6364 3773
rect 6406 3807 6464 3833
rect 6406 3773 6418 3807
rect 6452 3773 6464 3807
rect 6406 3747 6464 3773
rect 6506 3807 6564 3833
rect 6506 3773 6518 3807
rect 6552 3773 6564 3807
rect 6506 3747 6564 3773
rect 6606 3807 6664 3833
rect 6606 3773 6618 3807
rect 6652 3773 6664 3807
rect 6606 3747 6664 3773
rect 6706 3807 6764 3833
rect 6706 3773 6718 3807
rect 6752 3773 6764 3807
rect 6706 3747 6764 3773
rect 6806 3807 6864 3833
rect 6806 3773 6818 3807
rect 6852 3773 6864 3807
rect 6806 3747 6864 3773
rect 6906 3807 6964 3833
rect 6906 3773 6918 3807
rect 6952 3773 6964 3807
rect 6906 3747 6964 3773
rect 7006 3807 7064 3833
rect 7006 3773 7018 3807
rect 7052 3773 7064 3807
rect 7006 3747 7064 3773
rect 7106 3807 7164 3833
rect 7106 3773 7118 3807
rect 7152 3773 7164 3807
rect 7106 3747 7164 3773
rect 7206 3807 7264 3833
rect 7206 3773 7218 3807
rect 7252 3773 7264 3807
rect 7206 3747 7264 3773
rect 7306 3807 7364 3833
rect 7306 3773 7318 3807
rect 7352 3773 7364 3807
rect 7306 3747 7364 3773
rect 7406 3807 7464 3833
rect 7406 3773 7418 3807
rect 7452 3773 7464 3807
rect 7406 3747 7464 3773
rect 7506 3807 7564 3833
rect 7506 3773 7518 3807
rect 7552 3773 7564 3807
rect 7506 3747 7564 3773
rect 7606 3807 7664 3833
rect 7606 3773 7612 3807
rect 7652 3773 7664 3807
rect 7606 3747 7664 3773
rect 7706 3807 7764 3833
rect 7706 3773 7718 3807
rect 7758 3773 7764 3807
rect 7706 3747 7764 3773
rect 7806 3807 7864 3833
rect 7806 3773 7818 3807
rect 7852 3773 7864 3807
rect 7806 3747 7864 3773
rect 7906 3807 7964 3833
rect 7906 3773 7918 3807
rect 7952 3773 7964 3807
rect 7906 3747 7964 3773
rect 8006 3807 8064 3833
rect 8006 3773 8018 3807
rect 8052 3773 8064 3807
rect 8006 3747 8064 3773
rect 8106 3807 8164 3833
rect 8106 3773 8118 3807
rect 8152 3773 8164 3807
rect 8106 3747 8164 3773
rect 8206 3807 8264 3833
rect 8206 3773 8218 3807
rect 8252 3773 8264 3807
rect 8206 3747 8264 3773
rect 8306 3807 8364 3833
rect 8306 3773 8318 3807
rect 8352 3773 8364 3807
rect 8306 3747 8364 3773
rect 8406 3807 8464 3833
rect 8406 3773 8418 3807
rect 8452 3773 8464 3807
rect 8406 3747 8464 3773
rect 8506 3807 8564 3833
rect 8506 3773 8518 3807
rect 8552 3773 8564 3807
rect 8506 3747 8564 3773
rect 8606 3807 8664 3833
rect 8606 3773 8618 3807
rect 8652 3773 8664 3807
rect 8606 3747 8664 3773
rect 8706 3807 8764 3833
rect 8706 3773 8718 3807
rect 8752 3773 8764 3807
rect 8706 3747 8764 3773
rect 8806 3807 8864 3833
rect 8806 3773 8818 3807
rect 8852 3773 8864 3807
rect 8806 3747 8864 3773
rect 8906 3807 8964 3833
rect 8906 3773 8918 3807
rect 8952 3773 8964 3807
rect 8906 3747 8964 3773
rect 9006 3807 9064 3833
rect 9006 3773 9018 3807
rect 9052 3773 9064 3807
rect 9006 3747 9064 3773
rect 9106 3807 9164 3833
rect 9106 3773 9118 3807
rect 9152 3773 9164 3807
rect 9106 3747 9164 3773
rect 9206 3807 9264 3833
rect 9206 3773 9218 3807
rect 9252 3773 9264 3807
rect 9206 3747 9264 3773
rect 9306 3807 9364 3833
rect 9306 3773 9318 3807
rect 9352 3773 9364 3807
rect 9306 3747 9364 3773
rect 9406 3807 9464 3833
rect 9406 3773 9412 3807
rect 9452 3773 9464 3807
rect 9406 3747 9464 3773
rect 9506 3807 9564 3833
rect 9506 3773 9518 3807
rect 9558 3773 9564 3807
rect 9506 3747 9564 3773
rect 9606 3807 9664 3833
rect 9606 3773 9618 3807
rect 9652 3773 9664 3807
rect 9606 3747 9664 3773
rect 9706 3807 9764 3833
rect 9706 3773 9718 3807
rect 9752 3773 9764 3807
rect 9706 3747 9764 3773
rect 9806 3807 9864 3833
rect 9806 3773 9818 3807
rect 9852 3773 9864 3807
rect 9806 3747 9864 3773
rect 9906 3807 9964 3833
rect 9906 3773 9918 3807
rect 9952 3773 9964 3807
rect 9906 3747 9964 3773
rect 10006 3807 10064 3833
rect 10006 3773 10012 3807
rect 10052 3773 10064 3807
rect 10006 3747 10064 3773
rect 10106 3807 10164 3833
rect 10106 3773 10118 3807
rect 10158 3773 10164 3807
rect 10106 3747 10164 3773
rect 10206 3807 10264 3833
rect 10206 3773 10218 3807
rect 10252 3773 10264 3807
rect 10206 3747 10264 3773
rect 10306 3807 10364 3833
rect 10306 3773 10318 3807
rect 10352 3773 10364 3807
rect 10306 3747 10364 3773
rect 10406 3807 10464 3833
rect 10406 3773 10418 3807
rect 10452 3773 10464 3807
rect 10406 3747 10464 3773
rect 10506 3807 10564 3833
rect 10506 3773 10518 3807
rect 10552 3773 10564 3807
rect 10506 3747 10564 3773
rect 10606 3807 10664 3833
rect 10606 3773 10618 3807
rect 10652 3773 10664 3807
rect 10606 3747 10664 3773
rect 10706 3807 10764 3833
rect 10706 3773 10718 3807
rect 10752 3773 10764 3807
rect 10706 3747 10764 3773
rect 10806 3807 10864 3833
rect 10806 3773 10818 3807
rect 10852 3773 10864 3807
rect 10806 3747 10864 3773
rect 10906 3807 10964 3833
rect 10906 3773 10918 3807
rect 10952 3773 10964 3807
rect 10906 3747 10964 3773
rect 11006 3807 11064 3833
rect 11006 3773 11018 3807
rect 11052 3773 11064 3807
rect 11006 3747 11064 3773
rect 11106 3807 11164 3833
rect 11106 3773 11112 3807
rect 11152 3773 11164 3807
rect 11106 3747 11164 3773
rect 11206 3807 11264 3833
rect 11206 3773 11218 3807
rect 11258 3773 11264 3807
rect 11206 3747 11264 3773
rect 11306 3807 11364 3833
rect 11306 3773 11318 3807
rect 11352 3773 11364 3807
rect 11306 3747 11364 3773
rect 11406 3807 11464 3833
rect 11406 3773 11418 3807
rect 11452 3773 11464 3807
rect 11406 3747 11464 3773
rect 11506 3807 11564 3833
rect 11506 3773 11512 3807
rect 11552 3773 11564 3807
rect 11506 3747 11564 3773
rect 11606 3807 11664 3833
rect 11606 3773 11618 3807
rect 11658 3773 11664 3807
rect 11606 3747 11664 3773
rect 11706 3807 11764 3833
rect 11706 3773 11718 3807
rect 11752 3773 11764 3807
rect 11706 3747 11764 3773
rect 11806 3807 11864 3833
rect 11806 3773 11818 3807
rect 11852 3773 11864 3807
rect 11806 3747 11864 3773
rect 11906 3807 11964 3833
rect 11906 3773 11918 3807
rect 11952 3773 11964 3807
rect 11906 3747 11964 3773
rect 12006 3807 12064 3833
rect 12006 3773 12018 3807
rect 12052 3773 12064 3807
rect 12006 3747 12064 3773
rect 12106 3807 12164 3833
rect 12106 3773 12112 3807
rect 12152 3773 12164 3807
rect 12106 3747 12164 3773
rect 12206 3807 12264 3833
rect 12206 3773 12218 3807
rect 12258 3773 12264 3807
rect 12206 3747 12264 3773
rect 12306 3807 12364 3833
rect 12306 3773 12318 3807
rect 12352 3773 12364 3807
rect 12306 3747 12364 3773
rect 12406 3807 12464 3833
rect 12406 3773 12418 3807
rect 12452 3773 12464 3807
rect 12406 3747 12464 3773
rect 12506 3807 12564 3833
rect 12506 3773 12518 3807
rect 12552 3773 12564 3807
rect 12506 3747 12564 3773
rect 12606 3807 12664 3833
rect 12606 3773 12618 3807
rect 12652 3773 12664 3807
rect 12606 3747 12664 3773
rect 12706 3807 12764 3833
rect 12706 3773 12718 3807
rect 12752 3773 12764 3807
rect 12706 3747 12764 3773
rect 12806 3807 12864 3833
rect 13018 3826 13262 3860
rect 12806 3773 12818 3807
rect 12852 3773 12864 3807
rect 12908 3788 12916 3822
rect 12958 3788 12974 3822
rect 13018 3807 13052 3826
rect 12806 3747 12864 3773
rect 13228 3807 13262 3826
rect 13018 3757 13052 3773
rect 13096 3758 13112 3792
rect 13154 3758 13162 3792
rect 13228 3757 13262 3773
rect 13328 3807 13462 3823
rect 13362 3773 13428 3807
rect 13328 3757 13462 3773
rect 13528 3807 13662 3823
rect 13562 3773 13628 3807
rect 13528 3757 13662 3773
rect 8 3650 18 3684
rect 52 3650 118 3684
rect 152 3650 168 3684
rect 208 3666 218 3700
rect 252 3666 318 3700
rect 352 3666 368 3700
rect 408 3650 418 3684
rect 452 3650 518 3684
rect 552 3650 568 3684
rect 608 3666 618 3700
rect 652 3666 718 3700
rect 752 3666 768 3700
rect 808 3650 818 3684
rect 852 3650 918 3684
rect 952 3650 968 3684
rect 1008 3666 1018 3700
rect 1052 3666 1118 3700
rect 1152 3666 1168 3700
rect 1208 3650 1218 3684
rect 1252 3650 1318 3684
rect 1352 3650 1368 3684
rect 1408 3666 1418 3700
rect 1452 3666 1518 3700
rect 1552 3666 1568 3700
rect 1608 3650 1618 3684
rect 1652 3650 1718 3684
rect 1752 3650 1768 3684
rect 1808 3666 1818 3700
rect 1852 3666 1918 3700
rect 1952 3666 1968 3700
rect 2008 3650 2018 3684
rect 2052 3650 2118 3684
rect 2152 3650 2168 3684
rect 2208 3666 2218 3700
rect 2252 3666 2318 3700
rect 2352 3666 2368 3700
rect 2408 3650 2418 3684
rect 2452 3650 2518 3684
rect 2552 3650 2568 3684
rect 2608 3666 2618 3700
rect 2652 3666 2718 3700
rect 2752 3666 2768 3700
rect 2808 3650 2818 3684
rect 2852 3650 2918 3684
rect 2952 3650 2968 3684
rect 3008 3666 3018 3700
rect 3052 3666 3118 3700
rect 3152 3666 3168 3700
rect 3208 3650 3218 3684
rect 3252 3650 3318 3684
rect 3352 3650 3368 3684
rect 3408 3666 3418 3700
rect 3452 3666 3518 3700
rect 3552 3666 3568 3700
rect 3608 3650 3618 3684
rect 3652 3650 3718 3684
rect 3752 3650 3768 3684
rect 3808 3666 3818 3700
rect 3852 3666 3918 3700
rect 3952 3666 3968 3700
rect 4008 3650 4018 3684
rect 4052 3650 4118 3684
rect 4152 3650 4168 3684
rect 4208 3666 4218 3700
rect 4252 3666 4318 3700
rect 4352 3666 4368 3700
rect 4408 3650 4418 3684
rect 4452 3650 4518 3684
rect 4552 3650 4568 3684
rect 4608 3666 4618 3700
rect 4652 3666 4718 3700
rect 4752 3666 4768 3700
rect 4808 3650 4818 3684
rect 4852 3650 4918 3684
rect 4952 3650 4968 3684
rect 5008 3666 5018 3700
rect 5052 3666 5118 3700
rect 5152 3666 5168 3700
rect 5208 3650 5218 3684
rect 5252 3650 5318 3684
rect 5352 3650 5368 3684
rect 5408 3666 5418 3700
rect 5452 3666 5518 3700
rect 5552 3666 5568 3700
rect 5608 3650 5618 3684
rect 5652 3650 5718 3684
rect 5752 3650 5768 3684
rect 5808 3666 5818 3700
rect 5852 3666 5918 3700
rect 5952 3666 5968 3700
rect 6008 3650 6018 3684
rect 6052 3650 6118 3684
rect 6152 3650 6168 3684
rect 6208 3666 6218 3700
rect 6252 3666 6318 3700
rect 6352 3666 6368 3700
rect 6408 3650 6418 3684
rect 6452 3650 6518 3684
rect 6552 3650 6568 3684
rect 6608 3666 6618 3700
rect 6652 3666 6718 3700
rect 6752 3666 6768 3700
rect 6808 3650 6818 3684
rect 6852 3650 6918 3684
rect 6952 3650 6968 3684
rect 7008 3666 7018 3700
rect 7052 3666 7118 3700
rect 7152 3666 7168 3700
rect 7208 3650 7218 3684
rect 7252 3650 7318 3684
rect 7352 3650 7368 3684
rect 7408 3666 7418 3700
rect 7452 3666 7518 3700
rect 7552 3666 7568 3700
rect 7608 3650 7618 3684
rect 7652 3650 7718 3684
rect 7752 3650 7768 3684
rect 7808 3666 7818 3700
rect 7852 3666 7918 3700
rect 7952 3666 7968 3700
rect 8008 3650 8018 3684
rect 8052 3650 8118 3684
rect 8152 3650 8168 3684
rect 8208 3666 8218 3700
rect 8252 3666 8318 3700
rect 8352 3666 8368 3700
rect 8408 3650 8418 3684
rect 8452 3650 8518 3684
rect 8552 3650 8568 3684
rect 8608 3666 8618 3700
rect 8652 3666 8718 3700
rect 8752 3666 8768 3700
rect 8808 3650 8818 3684
rect 8852 3650 8918 3684
rect 8952 3650 8968 3684
rect 9008 3666 9018 3700
rect 9052 3666 9118 3700
rect 9152 3666 9168 3700
rect 9208 3650 9218 3684
rect 9252 3650 9318 3684
rect 9352 3650 9368 3684
rect 9408 3666 9418 3700
rect 9452 3666 9518 3700
rect 9552 3666 9568 3700
rect 9608 3650 9618 3684
rect 9652 3650 9718 3684
rect 9752 3650 9768 3684
rect 9808 3666 9818 3700
rect 9852 3666 9918 3700
rect 9952 3666 9968 3700
rect 10008 3650 10018 3684
rect 10052 3650 10118 3684
rect 10152 3650 10168 3684
rect 10208 3666 10218 3700
rect 10252 3666 10318 3700
rect 10352 3666 10368 3700
rect 10408 3650 10418 3684
rect 10452 3650 10518 3684
rect 10552 3650 10568 3684
rect 10608 3666 10618 3700
rect 10652 3666 10718 3700
rect 10752 3666 10768 3700
rect 10808 3650 10818 3684
rect 10852 3650 10918 3684
rect 10952 3650 10968 3684
rect 11008 3666 11018 3700
rect 11052 3666 11118 3700
rect 11152 3666 11168 3700
rect 11208 3650 11218 3684
rect 11252 3650 11318 3684
rect 11352 3650 11368 3684
rect 11408 3666 11418 3700
rect 11452 3666 11518 3700
rect 11552 3666 11568 3700
rect 11608 3650 11618 3684
rect 11652 3650 11718 3684
rect 11752 3650 11768 3684
rect 11808 3666 11818 3700
rect 11852 3666 11918 3700
rect 11952 3666 11968 3700
rect 12008 3650 12018 3684
rect 12052 3650 12118 3684
rect 12152 3650 12168 3684
rect 12208 3666 12218 3700
rect 12252 3666 12318 3700
rect 12352 3666 12368 3700
rect 12408 3650 12418 3684
rect 12452 3650 12518 3684
rect 12552 3650 12568 3684
rect 12608 3666 12618 3700
rect 12652 3666 12718 3700
rect 12752 3666 12768 3700
rect 12916 3681 12968 3698
rect 12950 3664 12968 3681
rect 13002 3664 13018 3698
rect 13052 3664 13068 3698
rect 13102 3669 13120 3698
rect 13102 3664 13154 3669
rect 13262 3664 13278 3698
rect 13312 3664 13328 3698
rect 13362 3664 13378 3698
rect 13412 3664 13428 3698
rect 13462 3664 13478 3698
rect 13512 3664 13528 3698
rect 13562 3664 13578 3698
rect 13612 3664 13628 3698
rect 6 3577 64 3603
rect 6 3543 18 3577
rect 52 3543 64 3577
rect 6 3517 64 3543
rect 106 3577 164 3603
rect 106 3543 118 3577
rect 152 3543 164 3577
rect 106 3517 164 3543
rect 206 3577 264 3603
rect 206 3543 218 3577
rect 252 3543 264 3577
rect 206 3517 264 3543
rect 306 3577 364 3603
rect 306 3543 318 3577
rect 352 3543 364 3577
rect 306 3517 364 3543
rect 406 3577 464 3603
rect 406 3543 418 3577
rect 452 3543 464 3577
rect 406 3517 464 3543
rect 506 3577 564 3603
rect 506 3543 518 3577
rect 552 3543 564 3577
rect 506 3517 564 3543
rect 606 3577 664 3603
rect 606 3543 618 3577
rect 652 3543 664 3577
rect 606 3517 664 3543
rect 706 3577 764 3603
rect 706 3543 718 3577
rect 752 3543 764 3577
rect 706 3517 764 3543
rect 806 3577 864 3603
rect 806 3543 812 3577
rect 852 3543 864 3577
rect 806 3517 864 3543
rect 906 3577 964 3603
rect 906 3543 918 3577
rect 958 3543 964 3577
rect 906 3517 964 3543
rect 1006 3577 1064 3603
rect 1006 3543 1012 3577
rect 1052 3543 1064 3577
rect 1006 3517 1064 3543
rect 1106 3577 1164 3603
rect 1106 3543 1118 3577
rect 1158 3543 1164 3577
rect 1106 3517 1164 3543
rect 1206 3577 1264 3603
rect 1206 3543 1218 3577
rect 1252 3543 1264 3577
rect 1206 3517 1264 3543
rect 1306 3577 1364 3603
rect 1306 3543 1318 3577
rect 1352 3543 1364 3577
rect 1306 3517 1364 3543
rect 1406 3577 1464 3603
rect 1406 3543 1418 3577
rect 1452 3543 1464 3577
rect 1406 3517 1464 3543
rect 1506 3577 1564 3603
rect 1506 3543 1518 3577
rect 1552 3543 1564 3577
rect 1506 3517 1564 3543
rect 1606 3577 1664 3603
rect 1606 3543 1618 3577
rect 1652 3543 1664 3577
rect 1606 3517 1664 3543
rect 1706 3577 1764 3603
rect 1706 3543 1718 3577
rect 1752 3543 1764 3577
rect 1706 3517 1764 3543
rect 1806 3577 1864 3603
rect 1806 3543 1818 3577
rect 1852 3543 1864 3577
rect 1806 3517 1864 3543
rect 1906 3577 1964 3603
rect 1906 3543 1918 3577
rect 1952 3543 1964 3577
rect 1906 3517 1964 3543
rect 2006 3577 2064 3603
rect 2006 3543 2018 3577
rect 2052 3543 2064 3577
rect 2006 3517 2064 3543
rect 2106 3577 2164 3603
rect 2106 3543 2118 3577
rect 2152 3543 2164 3577
rect 2106 3517 2164 3543
rect 2206 3577 2264 3603
rect 2206 3543 2218 3577
rect 2252 3543 2264 3577
rect 2206 3517 2264 3543
rect 2306 3577 2364 3603
rect 2306 3543 2318 3577
rect 2352 3543 2364 3577
rect 2306 3517 2364 3543
rect 2406 3577 2464 3603
rect 2406 3543 2418 3577
rect 2452 3543 2464 3577
rect 2406 3517 2464 3543
rect 2506 3577 2564 3603
rect 2506 3543 2512 3577
rect 2552 3543 2564 3577
rect 2506 3517 2564 3543
rect 2606 3577 2664 3603
rect 2606 3543 2618 3577
rect 2658 3543 2664 3577
rect 2606 3517 2664 3543
rect 2706 3577 2764 3603
rect 2706 3543 2718 3577
rect 2752 3543 2764 3577
rect 2706 3517 2764 3543
rect 2806 3577 2864 3603
rect 2806 3543 2818 3577
rect 2852 3543 2864 3577
rect 2806 3517 2864 3543
rect 2906 3577 2964 3603
rect 2906 3543 2918 3577
rect 2952 3543 2964 3577
rect 2906 3517 2964 3543
rect 3006 3577 3064 3603
rect 3006 3543 3018 3577
rect 3052 3543 3064 3577
rect 3006 3517 3064 3543
rect 3106 3577 3164 3603
rect 3106 3543 3112 3577
rect 3152 3543 3164 3577
rect 3106 3517 3164 3543
rect 3206 3577 3264 3603
rect 3206 3543 3218 3577
rect 3258 3543 3264 3577
rect 3206 3517 3264 3543
rect 3306 3577 3364 3603
rect 3306 3543 3318 3577
rect 3352 3543 3364 3577
rect 3306 3517 3364 3543
rect 3406 3577 3464 3603
rect 3406 3543 3418 3577
rect 3452 3543 3464 3577
rect 3406 3517 3464 3543
rect 3506 3577 3564 3603
rect 3506 3543 3518 3577
rect 3552 3543 3564 3577
rect 3506 3517 3564 3543
rect 3606 3577 3664 3603
rect 3606 3543 3618 3577
rect 3652 3543 3664 3577
rect 3606 3517 3664 3543
rect 3706 3577 3764 3603
rect 3706 3543 3718 3577
rect 3752 3543 3764 3577
rect 3706 3517 3764 3543
rect 3806 3577 3864 3603
rect 3806 3543 3818 3577
rect 3852 3543 3864 3577
rect 3806 3517 3864 3543
rect 3906 3577 3964 3603
rect 3906 3543 3918 3577
rect 3952 3543 3964 3577
rect 3906 3517 3964 3543
rect 4006 3577 4064 3603
rect 4006 3543 4018 3577
rect 4052 3543 4064 3577
rect 4006 3517 4064 3543
rect 4106 3577 4164 3603
rect 4106 3543 4118 3577
rect 4152 3543 4164 3577
rect 4106 3517 4164 3543
rect 4206 3577 4264 3603
rect 4206 3543 4218 3577
rect 4252 3543 4264 3577
rect 4206 3517 4264 3543
rect 4306 3577 4364 3603
rect 4306 3543 4318 3577
rect 4352 3543 4364 3577
rect 4306 3517 4364 3543
rect 4406 3577 4464 3603
rect 4406 3543 4412 3577
rect 4452 3543 4464 3577
rect 4406 3517 4464 3543
rect 4506 3577 4564 3603
rect 4506 3543 4518 3577
rect 4558 3543 4564 3577
rect 4506 3517 4564 3543
rect 4606 3577 4664 3603
rect 4606 3543 4618 3577
rect 4652 3543 4664 3577
rect 4606 3517 4664 3543
rect 4706 3577 4764 3603
rect 4706 3543 4718 3577
rect 4752 3543 4764 3577
rect 4706 3517 4764 3543
rect 4806 3577 4864 3603
rect 4806 3543 4818 3577
rect 4852 3543 4864 3577
rect 4806 3517 4864 3543
rect 4906 3577 4964 3603
rect 4906 3543 4918 3577
rect 4952 3543 4964 3577
rect 4906 3517 4964 3543
rect 5006 3577 5064 3603
rect 5006 3543 5018 3577
rect 5052 3543 5064 3577
rect 5006 3517 5064 3543
rect 5106 3577 5164 3603
rect 5106 3543 5118 3577
rect 5152 3543 5164 3577
rect 5106 3517 5164 3543
rect 5206 3577 5264 3603
rect 5206 3543 5218 3577
rect 5252 3543 5264 3577
rect 5206 3517 5264 3543
rect 5306 3577 5364 3603
rect 5306 3543 5318 3577
rect 5352 3543 5364 3577
rect 5306 3517 5364 3543
rect 5406 3577 5464 3603
rect 5406 3543 5418 3577
rect 5452 3543 5464 3577
rect 5406 3517 5464 3543
rect 5506 3577 5564 3603
rect 5506 3543 5518 3577
rect 5552 3543 5564 3577
rect 5506 3517 5564 3543
rect 5606 3577 5664 3603
rect 5606 3543 5618 3577
rect 5652 3543 5664 3577
rect 5606 3517 5664 3543
rect 5706 3577 5764 3603
rect 5706 3543 5712 3577
rect 5752 3543 5764 3577
rect 5706 3517 5764 3543
rect 5806 3577 5864 3603
rect 5806 3543 5818 3577
rect 5858 3543 5864 3577
rect 5806 3517 5864 3543
rect 5906 3577 5964 3603
rect 5906 3543 5918 3577
rect 5952 3543 5964 3577
rect 5906 3517 5964 3543
rect 6006 3577 6064 3603
rect 6006 3543 6018 3577
rect 6052 3543 6064 3577
rect 6006 3517 6064 3543
rect 6106 3577 6164 3603
rect 6106 3543 6118 3577
rect 6152 3543 6164 3577
rect 6106 3517 6164 3543
rect 6206 3577 6264 3603
rect 6206 3543 6218 3577
rect 6252 3543 6264 3577
rect 6206 3517 6264 3543
rect 6306 3577 6364 3603
rect 6306 3543 6318 3577
rect 6352 3543 6364 3577
rect 6306 3517 6364 3543
rect 6406 3577 6464 3603
rect 6406 3543 6418 3577
rect 6452 3543 6464 3577
rect 6406 3517 6464 3543
rect 6506 3577 6564 3603
rect 6506 3543 6518 3577
rect 6552 3543 6564 3577
rect 6506 3517 6564 3543
rect 6606 3577 6664 3603
rect 6606 3543 6618 3577
rect 6652 3543 6664 3577
rect 6606 3517 6664 3543
rect 6706 3577 6764 3603
rect 6706 3543 6718 3577
rect 6752 3543 6764 3577
rect 6706 3517 6764 3543
rect 6806 3577 6864 3603
rect 6806 3543 6818 3577
rect 6852 3543 6864 3577
rect 6806 3517 6864 3543
rect 6906 3577 6964 3603
rect 6906 3543 6918 3577
rect 6952 3543 6964 3577
rect 6906 3517 6964 3543
rect 7006 3577 7064 3603
rect 7006 3543 7018 3577
rect 7052 3543 7064 3577
rect 7006 3517 7064 3543
rect 7106 3577 7164 3603
rect 7106 3543 7118 3577
rect 7152 3543 7164 3577
rect 7106 3517 7164 3543
rect 7206 3577 7264 3603
rect 7206 3543 7218 3577
rect 7252 3543 7264 3577
rect 7206 3517 7264 3543
rect 7306 3577 7364 3603
rect 7306 3543 7318 3577
rect 7352 3543 7364 3577
rect 7306 3517 7364 3543
rect 7406 3577 7464 3603
rect 7406 3543 7418 3577
rect 7452 3543 7464 3577
rect 7406 3517 7464 3543
rect 7506 3577 7564 3603
rect 7506 3543 7518 3577
rect 7552 3543 7564 3577
rect 7506 3517 7564 3543
rect 7606 3577 7664 3603
rect 7606 3543 7618 3577
rect 7652 3543 7664 3577
rect 7606 3517 7664 3543
rect 7706 3577 7764 3603
rect 7706 3543 7718 3577
rect 7752 3543 7764 3577
rect 7706 3517 7764 3543
rect 7806 3577 7864 3603
rect 7806 3543 7818 3577
rect 7852 3543 7864 3577
rect 7806 3517 7864 3543
rect 7906 3577 7964 3603
rect 7906 3543 7918 3577
rect 7952 3543 7964 3577
rect 7906 3517 7964 3543
rect 8006 3577 8064 3603
rect 8006 3543 8018 3577
rect 8052 3543 8064 3577
rect 8006 3517 8064 3543
rect 8106 3577 8164 3603
rect 8106 3543 8118 3577
rect 8152 3543 8164 3577
rect 8106 3517 8164 3543
rect 8206 3577 8264 3603
rect 8206 3543 8218 3577
rect 8252 3543 8264 3577
rect 8206 3517 8264 3543
rect 8306 3577 8364 3603
rect 8306 3543 8318 3577
rect 8352 3543 8364 3577
rect 8306 3517 8364 3543
rect 8406 3577 8464 3603
rect 8406 3543 8418 3577
rect 8452 3543 8464 3577
rect 8406 3517 8464 3543
rect 8506 3577 8564 3603
rect 8506 3543 8518 3577
rect 8552 3543 8564 3577
rect 8506 3517 8564 3543
rect 8606 3577 8664 3603
rect 8606 3543 8618 3577
rect 8652 3543 8664 3577
rect 8606 3517 8664 3543
rect 8706 3577 8764 3603
rect 8706 3543 8718 3577
rect 8752 3543 8764 3577
rect 8706 3517 8764 3543
rect 8806 3577 8864 3603
rect 8806 3543 8818 3577
rect 8852 3543 8864 3577
rect 8806 3517 8864 3543
rect 8906 3577 8964 3603
rect 8906 3543 8912 3577
rect 8952 3543 8964 3577
rect 8906 3517 8964 3543
rect 9006 3577 9064 3603
rect 9006 3543 9018 3577
rect 9058 3543 9064 3577
rect 9006 3517 9064 3543
rect 9106 3577 9164 3603
rect 9106 3543 9112 3577
rect 9152 3543 9164 3577
rect 9106 3517 9164 3543
rect 9206 3577 9264 3603
rect 9206 3543 9218 3577
rect 9258 3543 9264 3577
rect 9206 3517 9264 3543
rect 9306 3577 9364 3603
rect 9306 3543 9312 3577
rect 9352 3543 9364 3577
rect 9306 3517 9364 3543
rect 9406 3577 9464 3603
rect 9406 3543 9418 3577
rect 9458 3543 9464 3577
rect 9406 3517 9464 3543
rect 9506 3577 9564 3603
rect 9506 3543 9518 3577
rect 9552 3543 9564 3577
rect 9506 3517 9564 3543
rect 9606 3577 9664 3603
rect 9606 3543 9618 3577
rect 9652 3543 9664 3577
rect 9606 3517 9664 3543
rect 9706 3577 9764 3603
rect 9706 3543 9718 3577
rect 9752 3543 9764 3577
rect 9706 3517 9764 3543
rect 9806 3577 9864 3603
rect 9806 3543 9818 3577
rect 9852 3543 9864 3577
rect 9806 3517 9864 3543
rect 9906 3577 9964 3603
rect 9906 3543 9918 3577
rect 9952 3543 9964 3577
rect 9906 3517 9964 3543
rect 10006 3577 10064 3603
rect 10006 3543 10012 3577
rect 10052 3543 10064 3577
rect 10006 3517 10064 3543
rect 10106 3577 10164 3603
rect 10106 3543 10118 3577
rect 10158 3543 10164 3577
rect 10106 3517 10164 3543
rect 10206 3577 10264 3603
rect 10206 3543 10218 3577
rect 10252 3543 10264 3577
rect 10206 3517 10264 3543
rect 10306 3577 10364 3603
rect 10306 3543 10318 3577
rect 10352 3543 10364 3577
rect 10306 3517 10364 3543
rect 10406 3577 10464 3603
rect 10406 3543 10418 3577
rect 10452 3543 10464 3577
rect 10406 3517 10464 3543
rect 10506 3577 10564 3603
rect 10506 3543 10518 3577
rect 10552 3543 10564 3577
rect 10506 3517 10564 3543
rect 10606 3577 10664 3603
rect 10606 3543 10612 3577
rect 10652 3543 10664 3577
rect 10606 3517 10664 3543
rect 10706 3577 10764 3603
rect 10706 3543 10718 3577
rect 10758 3543 10764 3577
rect 10706 3517 10764 3543
rect 10806 3577 10864 3603
rect 10806 3543 10818 3577
rect 10852 3543 10864 3577
rect 10806 3517 10864 3543
rect 10906 3577 10964 3603
rect 10906 3543 10918 3577
rect 10952 3543 10964 3577
rect 10906 3517 10964 3543
rect 11006 3577 11064 3603
rect 11006 3543 11018 3577
rect 11052 3543 11064 3577
rect 11006 3517 11064 3543
rect 11106 3577 11164 3603
rect 11106 3543 11118 3577
rect 11152 3543 11164 3577
rect 11106 3517 11164 3543
rect 11206 3577 11264 3603
rect 11206 3543 11218 3577
rect 11252 3543 11264 3577
rect 11206 3517 11264 3543
rect 11306 3577 11364 3603
rect 11306 3543 11318 3577
rect 11352 3543 11364 3577
rect 11306 3517 11364 3543
rect 11406 3577 11464 3603
rect 11406 3543 11412 3577
rect 11452 3543 11464 3577
rect 11406 3517 11464 3543
rect 11506 3577 11564 3603
rect 11506 3543 11518 3577
rect 11558 3543 11564 3577
rect 11506 3517 11564 3543
rect 11606 3577 11664 3603
rect 11606 3543 11618 3577
rect 11652 3543 11664 3577
rect 11606 3517 11664 3543
rect 11706 3577 11764 3603
rect 11706 3543 11718 3577
rect 11752 3543 11764 3577
rect 11706 3517 11764 3543
rect 11806 3577 11864 3603
rect 11806 3543 11818 3577
rect 11852 3543 11864 3577
rect 11806 3517 11864 3543
rect 11906 3577 11964 3603
rect 11906 3543 11918 3577
rect 11952 3543 11964 3577
rect 11906 3517 11964 3543
rect 12006 3577 12064 3603
rect 12006 3543 12018 3577
rect 12052 3543 12064 3577
rect 12006 3517 12064 3543
rect 12106 3577 12164 3603
rect 12106 3543 12118 3577
rect 12152 3543 12164 3577
rect 12106 3517 12164 3543
rect 12206 3577 12264 3603
rect 12206 3543 12218 3577
rect 12252 3543 12264 3577
rect 12206 3517 12264 3543
rect 12306 3577 12364 3603
rect 12306 3543 12318 3577
rect 12352 3543 12364 3577
rect 12306 3517 12364 3543
rect 12406 3577 12464 3603
rect 12406 3543 12418 3577
rect 12452 3543 12464 3577
rect 12406 3517 12464 3543
rect 12506 3577 12564 3603
rect 12506 3543 12518 3577
rect 12552 3543 12564 3577
rect 12506 3517 12564 3543
rect 12606 3577 12664 3603
rect 12606 3543 12618 3577
rect 12652 3543 12664 3577
rect 12606 3517 12664 3543
rect 12706 3577 12764 3603
rect 12706 3543 12718 3577
rect 12752 3543 12764 3577
rect 12706 3517 12764 3543
rect 12806 3577 12864 3603
rect 13018 3596 13262 3630
rect 12806 3543 12818 3577
rect 12852 3543 12864 3577
rect 12908 3558 12916 3592
rect 12958 3558 12974 3592
rect 13018 3577 13052 3596
rect 12806 3517 12864 3543
rect 13228 3593 13262 3596
rect 13228 3577 13362 3593
rect 13018 3527 13052 3543
rect 13096 3528 13112 3562
rect 13154 3528 13162 3562
rect 13262 3543 13328 3577
rect 13228 3527 13362 3543
rect 13428 3577 13562 3593
rect 13462 3543 13528 3577
rect 13428 3527 13562 3543
rect 13628 3577 13662 3593
rect 13628 3527 13662 3543
rect 6 3437 64 3463
rect 6 3403 18 3437
rect 58 3403 64 3437
rect 6 3377 64 3403
rect 106 3437 164 3463
rect 106 3403 118 3437
rect 152 3403 164 3437
rect 106 3377 164 3403
rect 206 3437 264 3463
rect 206 3403 218 3437
rect 252 3403 264 3437
rect 206 3377 264 3403
rect 306 3437 364 3463
rect 306 3403 312 3437
rect 352 3403 364 3437
rect 306 3377 364 3403
rect 406 3437 464 3463
rect 406 3403 418 3437
rect 458 3403 464 3437
rect 406 3377 464 3403
rect 506 3437 564 3463
rect 506 3403 512 3437
rect 552 3403 564 3437
rect 506 3377 564 3403
rect 606 3437 664 3463
rect 606 3403 618 3437
rect 658 3403 664 3437
rect 606 3377 664 3403
rect 706 3437 764 3463
rect 706 3403 712 3437
rect 752 3403 764 3437
rect 706 3377 764 3403
rect 806 3437 864 3463
rect 806 3403 818 3437
rect 858 3403 864 3437
rect 806 3377 864 3403
rect 906 3437 964 3463
rect 906 3403 912 3437
rect 952 3403 964 3437
rect 906 3377 964 3403
rect 1006 3437 1064 3463
rect 1006 3403 1018 3437
rect 1058 3403 1064 3437
rect 1006 3377 1064 3403
rect 1106 3437 1164 3463
rect 1106 3403 1118 3437
rect 1152 3403 1164 3437
rect 1106 3377 1164 3403
rect 1206 3437 1264 3463
rect 1206 3403 1218 3437
rect 1252 3403 1264 3437
rect 1206 3377 1264 3403
rect 1306 3437 1364 3463
rect 1306 3403 1318 3437
rect 1352 3403 1364 3437
rect 1306 3377 1364 3403
rect 1406 3437 1464 3463
rect 1406 3403 1418 3437
rect 1452 3403 1464 3437
rect 1406 3377 1464 3403
rect 1506 3437 1564 3463
rect 1506 3403 1518 3437
rect 1552 3403 1564 3437
rect 1506 3377 1564 3403
rect 1606 3437 1664 3463
rect 1606 3403 1618 3437
rect 1652 3403 1664 3437
rect 1606 3377 1664 3403
rect 1706 3437 1764 3463
rect 1706 3403 1718 3437
rect 1752 3403 1764 3437
rect 1706 3377 1764 3403
rect 1806 3437 1864 3463
rect 1806 3403 1818 3437
rect 1852 3403 1864 3437
rect 1806 3377 1864 3403
rect 1906 3437 1964 3463
rect 1906 3403 1918 3437
rect 1952 3403 1964 3437
rect 1906 3377 1964 3403
rect 2006 3437 2064 3463
rect 2006 3403 2018 3437
rect 2052 3403 2064 3437
rect 2006 3377 2064 3403
rect 2106 3437 2164 3463
rect 2106 3403 2118 3437
rect 2152 3403 2164 3437
rect 2106 3377 2164 3403
rect 2206 3437 2264 3463
rect 2206 3403 2218 3437
rect 2252 3403 2264 3437
rect 2206 3377 2264 3403
rect 2306 3437 2364 3463
rect 2306 3403 2318 3437
rect 2352 3403 2364 3437
rect 2306 3377 2364 3403
rect 2406 3437 2464 3463
rect 2406 3403 2418 3437
rect 2452 3403 2464 3437
rect 2406 3377 2464 3403
rect 2506 3437 2564 3463
rect 2506 3403 2518 3437
rect 2552 3403 2564 3437
rect 2506 3377 2564 3403
rect 2606 3437 2664 3463
rect 2606 3403 2618 3437
rect 2652 3403 2664 3437
rect 2606 3377 2664 3403
rect 2706 3437 2764 3463
rect 2706 3403 2718 3437
rect 2752 3403 2764 3437
rect 2706 3377 2764 3403
rect 2806 3437 2864 3463
rect 2806 3403 2818 3437
rect 2852 3403 2864 3437
rect 2806 3377 2864 3403
rect 2906 3437 2964 3463
rect 2906 3403 2918 3437
rect 2952 3403 2964 3437
rect 2906 3377 2964 3403
rect 3006 3437 3064 3463
rect 3006 3403 3018 3437
rect 3052 3403 3064 3437
rect 3006 3377 3064 3403
rect 3106 3437 3164 3463
rect 3106 3403 3118 3437
rect 3152 3403 3164 3437
rect 3106 3377 3164 3403
rect 3206 3437 3264 3463
rect 3206 3403 3218 3437
rect 3252 3403 3264 3437
rect 3206 3377 3264 3403
rect 3306 3437 3364 3463
rect 3306 3403 3318 3437
rect 3352 3403 3364 3437
rect 3306 3377 3364 3403
rect 3406 3437 3464 3463
rect 3406 3403 3418 3437
rect 3452 3403 3464 3437
rect 3406 3377 3464 3403
rect 3506 3437 3564 3463
rect 3506 3403 3518 3437
rect 3552 3403 3564 3437
rect 3506 3377 3564 3403
rect 3606 3437 3664 3463
rect 3606 3403 3618 3437
rect 3652 3403 3664 3437
rect 3606 3377 3664 3403
rect 3706 3437 3764 3463
rect 3706 3403 3718 3437
rect 3752 3403 3764 3437
rect 3706 3377 3764 3403
rect 3806 3437 3864 3463
rect 3806 3403 3812 3437
rect 3852 3403 3864 3437
rect 3806 3377 3864 3403
rect 3906 3437 3964 3463
rect 3906 3403 3918 3437
rect 3958 3403 3964 3437
rect 3906 3377 3964 3403
rect 4006 3437 4064 3463
rect 4006 3403 4018 3437
rect 4052 3403 4064 3437
rect 4006 3377 4064 3403
rect 4106 3437 4164 3463
rect 4106 3403 4118 3437
rect 4152 3403 4164 3437
rect 4106 3377 4164 3403
rect 4206 3437 4264 3463
rect 4206 3403 4218 3437
rect 4252 3403 4264 3437
rect 4206 3377 4264 3403
rect 4306 3437 4364 3463
rect 4306 3403 4318 3437
rect 4352 3403 4364 3437
rect 4306 3377 4364 3403
rect 4406 3437 4464 3463
rect 4406 3403 4412 3437
rect 4452 3403 4464 3437
rect 4406 3377 4464 3403
rect 4506 3437 4564 3463
rect 4506 3403 4518 3437
rect 4558 3403 4564 3437
rect 4506 3377 4564 3403
rect 4606 3437 4664 3463
rect 4606 3403 4618 3437
rect 4652 3403 4664 3437
rect 4606 3377 4664 3403
rect 4706 3437 4764 3463
rect 4706 3403 4718 3437
rect 4752 3403 4764 3437
rect 4706 3377 4764 3403
rect 4806 3437 4864 3463
rect 4806 3403 4812 3437
rect 4852 3403 4864 3437
rect 4806 3377 4864 3403
rect 4906 3437 4964 3463
rect 4906 3403 4918 3437
rect 4958 3403 4964 3437
rect 4906 3377 4964 3403
rect 5006 3437 5064 3463
rect 5006 3403 5012 3437
rect 5052 3403 5064 3437
rect 5006 3377 5064 3403
rect 5106 3437 5164 3463
rect 5106 3403 5118 3437
rect 5158 3403 5164 3437
rect 5106 3377 5164 3403
rect 5206 3437 5264 3463
rect 5206 3403 5218 3437
rect 5252 3403 5264 3437
rect 5206 3377 5264 3403
rect 5306 3437 5364 3463
rect 5306 3403 5318 3437
rect 5352 3403 5364 3437
rect 5306 3377 5364 3403
rect 5406 3437 5464 3463
rect 5406 3403 5418 3437
rect 5452 3403 5464 3437
rect 5406 3377 5464 3403
rect 5506 3437 5564 3463
rect 5506 3403 5518 3437
rect 5552 3403 5564 3437
rect 5506 3377 5564 3403
rect 5606 3437 5664 3463
rect 5606 3403 5618 3437
rect 5652 3403 5664 3437
rect 5606 3377 5664 3403
rect 5706 3437 5764 3463
rect 5706 3403 5718 3437
rect 5752 3403 5764 3437
rect 5706 3377 5764 3403
rect 5806 3437 5864 3463
rect 5806 3403 5818 3437
rect 5852 3403 5864 3437
rect 5806 3377 5864 3403
rect 5906 3437 5964 3463
rect 5906 3403 5918 3437
rect 5952 3403 5964 3437
rect 5906 3377 5964 3403
rect 6006 3437 6064 3463
rect 6006 3403 6012 3437
rect 6052 3403 6064 3437
rect 6006 3377 6064 3403
rect 6106 3437 6164 3463
rect 6106 3403 6118 3437
rect 6158 3403 6164 3437
rect 6106 3377 6164 3403
rect 6206 3437 6264 3463
rect 6206 3403 6218 3437
rect 6252 3403 6264 3437
rect 6206 3377 6264 3403
rect 6306 3437 6364 3463
rect 6306 3403 6318 3437
rect 6352 3403 6364 3437
rect 6306 3377 6364 3403
rect 6406 3437 6464 3463
rect 6406 3403 6412 3437
rect 6452 3403 6464 3437
rect 6406 3377 6464 3403
rect 6506 3437 6564 3463
rect 6506 3403 6518 3437
rect 6558 3403 6564 3437
rect 6506 3377 6564 3403
rect 6606 3437 6664 3463
rect 6606 3403 6618 3437
rect 6652 3403 6664 3437
rect 6606 3377 6664 3403
rect 6706 3437 6764 3463
rect 6706 3403 6712 3437
rect 6752 3403 6764 3437
rect 6706 3377 6764 3403
rect 6806 3437 6864 3463
rect 6806 3403 6818 3437
rect 6858 3403 6864 3437
rect 6806 3377 6864 3403
rect 6906 3437 6964 3463
rect 6906 3403 6918 3437
rect 6952 3403 6964 3437
rect 6906 3377 6964 3403
rect 7006 3437 7064 3463
rect 7006 3403 7018 3437
rect 7052 3403 7064 3437
rect 7006 3377 7064 3403
rect 7106 3437 7164 3463
rect 7106 3403 7118 3437
rect 7152 3403 7164 3437
rect 7106 3377 7164 3403
rect 7206 3437 7264 3463
rect 7206 3403 7218 3437
rect 7252 3403 7264 3437
rect 7206 3377 7264 3403
rect 7306 3437 7364 3463
rect 7306 3403 7318 3437
rect 7352 3403 7364 3437
rect 7306 3377 7364 3403
rect 7406 3437 7464 3463
rect 7406 3403 7418 3437
rect 7452 3403 7464 3437
rect 7406 3377 7464 3403
rect 7506 3437 7564 3463
rect 7506 3403 7518 3437
rect 7552 3403 7564 3437
rect 7506 3377 7564 3403
rect 7606 3437 7664 3463
rect 7606 3403 7618 3437
rect 7652 3403 7664 3437
rect 7606 3377 7664 3403
rect 7706 3437 7764 3463
rect 7706 3403 7718 3437
rect 7752 3403 7764 3437
rect 7706 3377 7764 3403
rect 7806 3437 7864 3463
rect 7806 3403 7818 3437
rect 7852 3403 7864 3437
rect 7806 3377 7864 3403
rect 7906 3437 7964 3463
rect 7906 3403 7918 3437
rect 7952 3403 7964 3437
rect 7906 3377 7964 3403
rect 8006 3437 8064 3463
rect 8006 3403 8018 3437
rect 8052 3403 8064 3437
rect 8006 3377 8064 3403
rect 8106 3437 8164 3463
rect 8106 3403 8118 3437
rect 8152 3403 8164 3437
rect 8106 3377 8164 3403
rect 8206 3437 8264 3463
rect 8206 3403 8218 3437
rect 8252 3403 8264 3437
rect 8206 3377 8264 3403
rect 8306 3437 8364 3463
rect 8306 3403 8318 3437
rect 8352 3403 8364 3437
rect 8306 3377 8364 3403
rect 8406 3437 8464 3463
rect 8406 3403 8418 3437
rect 8452 3403 8464 3437
rect 8406 3377 8464 3403
rect 8506 3437 8564 3463
rect 8506 3403 8518 3437
rect 8552 3403 8564 3437
rect 8506 3377 8564 3403
rect 8606 3437 8664 3463
rect 8606 3403 8618 3437
rect 8652 3403 8664 3437
rect 8606 3377 8664 3403
rect 8706 3437 8764 3463
rect 8706 3403 8718 3437
rect 8752 3403 8764 3437
rect 8706 3377 8764 3403
rect 8806 3437 8864 3463
rect 8806 3403 8818 3437
rect 8852 3403 8864 3437
rect 8806 3377 8864 3403
rect 8906 3437 8964 3463
rect 8906 3403 8918 3437
rect 8952 3403 8964 3437
rect 8906 3377 8964 3403
rect 9006 3437 9064 3463
rect 9006 3403 9018 3437
rect 9052 3403 9064 3437
rect 9006 3377 9064 3403
rect 9106 3437 9164 3463
rect 9106 3403 9118 3437
rect 9152 3403 9164 3437
rect 9106 3377 9164 3403
rect 9206 3437 9264 3463
rect 9206 3403 9218 3437
rect 9252 3403 9264 3437
rect 9206 3377 9264 3403
rect 9306 3437 9364 3463
rect 9306 3403 9318 3437
rect 9352 3403 9364 3437
rect 9306 3377 9364 3403
rect 9406 3437 9464 3463
rect 9406 3403 9412 3437
rect 9452 3403 9464 3437
rect 9406 3377 9464 3403
rect 9506 3437 9564 3463
rect 9506 3403 9518 3437
rect 9558 3403 9564 3437
rect 9506 3377 9564 3403
rect 9606 3437 9664 3463
rect 9606 3403 9618 3437
rect 9652 3403 9664 3437
rect 9606 3377 9664 3403
rect 9706 3437 9764 3463
rect 9706 3403 9712 3437
rect 9752 3403 9764 3437
rect 9706 3377 9764 3403
rect 9806 3437 9864 3463
rect 9806 3403 9818 3437
rect 9858 3403 9864 3437
rect 9806 3377 9864 3403
rect 9906 3437 9964 3463
rect 9906 3403 9918 3437
rect 9952 3403 9964 3437
rect 9906 3377 9964 3403
rect 10006 3437 10064 3463
rect 10006 3403 10018 3437
rect 10052 3403 10064 3437
rect 10006 3377 10064 3403
rect 10106 3437 10164 3463
rect 10106 3403 10118 3437
rect 10152 3403 10164 3437
rect 10106 3377 10164 3403
rect 10206 3437 10264 3463
rect 10206 3403 10218 3437
rect 10252 3403 10264 3437
rect 10206 3377 10264 3403
rect 10306 3437 10364 3463
rect 10306 3403 10318 3437
rect 10352 3403 10364 3437
rect 10306 3377 10364 3403
rect 10406 3437 10464 3463
rect 10406 3403 10418 3437
rect 10452 3403 10464 3437
rect 10406 3377 10464 3403
rect 10506 3437 10564 3463
rect 10506 3403 10518 3437
rect 10552 3403 10564 3437
rect 10506 3377 10564 3403
rect 10606 3437 10664 3463
rect 10606 3403 10618 3437
rect 10652 3403 10664 3437
rect 10606 3377 10664 3403
rect 10706 3437 10764 3463
rect 10706 3403 10718 3437
rect 10752 3403 10764 3437
rect 10706 3377 10764 3403
rect 10806 3437 10864 3463
rect 10806 3403 10818 3437
rect 10852 3403 10864 3437
rect 10806 3377 10864 3403
rect 10906 3437 10964 3463
rect 10906 3403 10918 3437
rect 10952 3403 10964 3437
rect 10906 3377 10964 3403
rect 11006 3437 11064 3463
rect 11006 3403 11018 3437
rect 11052 3403 11064 3437
rect 11006 3377 11064 3403
rect 11106 3437 11164 3463
rect 11106 3403 11118 3437
rect 11152 3403 11164 3437
rect 11106 3377 11164 3403
rect 11206 3437 11264 3463
rect 11206 3403 11218 3437
rect 11252 3403 11264 3437
rect 11206 3377 11264 3403
rect 11306 3437 11364 3463
rect 11306 3403 11318 3437
rect 11352 3403 11364 3437
rect 11306 3377 11364 3403
rect 11406 3437 11464 3463
rect 11406 3403 11412 3437
rect 11452 3403 11464 3437
rect 11406 3377 11464 3403
rect 11506 3437 11564 3463
rect 11506 3403 11518 3437
rect 11558 3403 11564 3437
rect 11506 3377 11564 3403
rect 11606 3437 11664 3463
rect 11606 3403 11618 3437
rect 11652 3403 11664 3437
rect 11606 3377 11664 3403
rect 11706 3437 11764 3463
rect 11706 3403 11718 3437
rect 11752 3403 11764 3437
rect 11706 3377 11764 3403
rect 11806 3437 11864 3463
rect 11806 3403 11818 3437
rect 11852 3403 11864 3437
rect 11806 3377 11864 3403
rect 11906 3437 11964 3463
rect 11906 3403 11918 3437
rect 11952 3403 11964 3437
rect 11906 3377 11964 3403
rect 12006 3437 12064 3463
rect 12006 3403 12018 3437
rect 12052 3403 12064 3437
rect 12006 3377 12064 3403
rect 12106 3437 12164 3463
rect 12106 3403 12112 3437
rect 12152 3403 12164 3437
rect 12106 3377 12164 3403
rect 12206 3437 12264 3463
rect 12206 3403 12218 3437
rect 12258 3403 12264 3437
rect 12206 3377 12264 3403
rect 12306 3437 12364 3463
rect 12306 3403 12318 3437
rect 12352 3403 12364 3437
rect 12306 3377 12364 3403
rect 12406 3437 12464 3463
rect 12406 3403 12418 3437
rect 12452 3403 12464 3437
rect 12406 3377 12464 3403
rect 12506 3437 12564 3463
rect 12506 3403 12518 3437
rect 12552 3403 12564 3437
rect 12506 3377 12564 3403
rect 12606 3437 12664 3463
rect 12606 3403 12618 3437
rect 12652 3403 12664 3437
rect 12606 3377 12664 3403
rect 12706 3437 12764 3463
rect 12706 3403 12718 3437
rect 12752 3403 12764 3437
rect 12706 3377 12764 3403
rect 12806 3437 12864 3463
rect 13018 3456 13262 3490
rect 12806 3403 12812 3437
rect 12852 3403 12864 3437
rect 12908 3418 12916 3452
rect 12958 3418 12974 3452
rect 13018 3437 13052 3456
rect 12806 3377 12864 3403
rect 13228 3437 13262 3456
rect 13018 3387 13052 3403
rect 13096 3388 13112 3422
rect 13154 3388 13162 3422
rect 13228 3387 13262 3403
rect 13328 3437 13562 3453
rect 13362 3403 13428 3437
rect 13462 3403 13528 3437
rect 13328 3387 13562 3403
rect 13628 3437 13662 3453
rect 13628 3387 13662 3403
rect 6 3297 64 3323
rect 6 3263 18 3297
rect 52 3263 64 3297
rect 6 3237 64 3263
rect 106 3297 164 3323
rect 106 3263 118 3297
rect 152 3263 164 3297
rect 106 3237 164 3263
rect 206 3297 264 3323
rect 206 3263 218 3297
rect 252 3263 264 3297
rect 206 3237 264 3263
rect 306 3297 364 3323
rect 306 3263 318 3297
rect 352 3263 364 3297
rect 306 3237 364 3263
rect 406 3297 464 3323
rect 406 3263 418 3297
rect 452 3263 464 3297
rect 406 3237 464 3263
rect 506 3297 564 3323
rect 506 3263 518 3297
rect 552 3263 564 3297
rect 506 3237 564 3263
rect 606 3297 664 3323
rect 606 3263 618 3297
rect 652 3263 664 3297
rect 606 3237 664 3263
rect 706 3297 764 3323
rect 706 3263 712 3297
rect 752 3263 764 3297
rect 706 3237 764 3263
rect 806 3297 864 3323
rect 806 3263 818 3297
rect 858 3263 864 3297
rect 806 3237 864 3263
rect 906 3297 964 3323
rect 906 3263 912 3297
rect 952 3263 964 3297
rect 906 3237 964 3263
rect 1006 3297 1064 3323
rect 1006 3263 1018 3297
rect 1058 3263 1064 3297
rect 1006 3237 1064 3263
rect 1106 3297 1164 3323
rect 1106 3263 1118 3297
rect 1152 3263 1164 3297
rect 1106 3237 1164 3263
rect 1206 3297 1264 3323
rect 1206 3263 1218 3297
rect 1252 3263 1264 3297
rect 1206 3237 1264 3263
rect 1306 3297 1364 3323
rect 1306 3263 1318 3297
rect 1352 3263 1364 3297
rect 1306 3237 1364 3263
rect 1406 3297 1464 3323
rect 1406 3263 1418 3297
rect 1452 3263 1464 3297
rect 1406 3237 1464 3263
rect 1506 3297 1564 3323
rect 1506 3263 1518 3297
rect 1552 3263 1564 3297
rect 1506 3237 1564 3263
rect 1606 3297 1664 3323
rect 1606 3263 1618 3297
rect 1652 3263 1664 3297
rect 1606 3237 1664 3263
rect 1706 3297 1764 3323
rect 1706 3263 1718 3297
rect 1752 3263 1764 3297
rect 1706 3237 1764 3263
rect 1806 3297 1864 3323
rect 1806 3263 1818 3297
rect 1852 3263 1864 3297
rect 1806 3237 1864 3263
rect 1906 3297 1964 3323
rect 1906 3263 1918 3297
rect 1952 3263 1964 3297
rect 1906 3237 1964 3263
rect 2006 3297 2064 3323
rect 2006 3263 2018 3297
rect 2052 3263 2064 3297
rect 2006 3237 2064 3263
rect 2106 3297 2164 3323
rect 2106 3263 2118 3297
rect 2152 3263 2164 3297
rect 2106 3237 2164 3263
rect 2206 3297 2264 3323
rect 2206 3263 2218 3297
rect 2252 3263 2264 3297
rect 2206 3237 2264 3263
rect 2306 3297 2364 3323
rect 2306 3263 2318 3297
rect 2352 3263 2364 3297
rect 2306 3237 2364 3263
rect 2406 3297 2464 3323
rect 2406 3263 2418 3297
rect 2452 3263 2464 3297
rect 2406 3237 2464 3263
rect 2506 3297 2564 3323
rect 2506 3263 2518 3297
rect 2552 3263 2564 3297
rect 2506 3237 2564 3263
rect 2606 3297 2664 3323
rect 2606 3263 2618 3297
rect 2652 3263 2664 3297
rect 2606 3237 2664 3263
rect 2706 3297 2764 3323
rect 2706 3263 2712 3297
rect 2752 3263 2764 3297
rect 2706 3237 2764 3263
rect 2806 3297 2864 3323
rect 2806 3263 2818 3297
rect 2858 3263 2864 3297
rect 2806 3237 2864 3263
rect 2906 3297 2964 3323
rect 2906 3263 2918 3297
rect 2952 3263 2964 3297
rect 2906 3237 2964 3263
rect 3006 3297 3064 3323
rect 3006 3263 3018 3297
rect 3052 3263 3064 3297
rect 3006 3237 3064 3263
rect 3106 3297 3164 3323
rect 3106 3263 3118 3297
rect 3152 3263 3164 3297
rect 3106 3237 3164 3263
rect 3206 3297 3264 3323
rect 3206 3263 3212 3297
rect 3252 3263 3264 3297
rect 3206 3237 3264 3263
rect 3306 3297 3364 3323
rect 3306 3263 3318 3297
rect 3358 3263 3364 3297
rect 3306 3237 3364 3263
rect 3406 3297 3464 3323
rect 3406 3263 3412 3297
rect 3452 3263 3464 3297
rect 3406 3237 3464 3263
rect 3506 3297 3564 3323
rect 3506 3263 3518 3297
rect 3558 3263 3564 3297
rect 3506 3237 3564 3263
rect 3606 3297 3664 3323
rect 3606 3263 3618 3297
rect 3652 3263 3664 3297
rect 3606 3237 3664 3263
rect 3706 3297 3764 3323
rect 3706 3263 3718 3297
rect 3752 3263 3764 3297
rect 3706 3237 3764 3263
rect 3806 3297 3864 3323
rect 3806 3263 3818 3297
rect 3852 3263 3864 3297
rect 3806 3237 3864 3263
rect 3906 3297 3964 3323
rect 3906 3263 3918 3297
rect 3952 3263 3964 3297
rect 3906 3237 3964 3263
rect 4006 3297 4064 3323
rect 4006 3263 4018 3297
rect 4052 3263 4064 3297
rect 4006 3237 4064 3263
rect 4106 3297 4164 3323
rect 4106 3263 4118 3297
rect 4152 3263 4164 3297
rect 4106 3237 4164 3263
rect 4206 3297 4264 3323
rect 4206 3263 4218 3297
rect 4252 3263 4264 3297
rect 4206 3237 4264 3263
rect 4306 3297 4364 3323
rect 4306 3263 4318 3297
rect 4352 3263 4364 3297
rect 4306 3237 4364 3263
rect 4406 3297 4464 3323
rect 4406 3263 4418 3297
rect 4452 3263 4464 3297
rect 4406 3237 4464 3263
rect 4506 3297 4564 3323
rect 4506 3263 4518 3297
rect 4552 3263 4564 3297
rect 4506 3237 4564 3263
rect 4606 3297 4664 3323
rect 4606 3263 4618 3297
rect 4652 3263 4664 3297
rect 4606 3237 4664 3263
rect 4706 3297 4764 3323
rect 4706 3263 4718 3297
rect 4752 3263 4764 3297
rect 4706 3237 4764 3263
rect 4806 3297 4864 3323
rect 4806 3263 4818 3297
rect 4852 3263 4864 3297
rect 4806 3237 4864 3263
rect 4906 3297 4964 3323
rect 4906 3263 4918 3297
rect 4952 3263 4964 3297
rect 4906 3237 4964 3263
rect 5006 3297 5064 3323
rect 5006 3263 5018 3297
rect 5052 3263 5064 3297
rect 5006 3237 5064 3263
rect 5106 3297 5164 3323
rect 5106 3263 5118 3297
rect 5152 3263 5164 3297
rect 5106 3237 5164 3263
rect 5206 3297 5264 3323
rect 5206 3263 5218 3297
rect 5252 3263 5264 3297
rect 5206 3237 5264 3263
rect 5306 3297 5364 3323
rect 5306 3263 5318 3297
rect 5352 3263 5364 3297
rect 5306 3237 5364 3263
rect 5406 3297 5464 3323
rect 5406 3263 5418 3297
rect 5452 3263 5464 3297
rect 5406 3237 5464 3263
rect 5506 3297 5564 3323
rect 5506 3263 5518 3297
rect 5552 3263 5564 3297
rect 5506 3237 5564 3263
rect 5606 3297 5664 3323
rect 5606 3263 5618 3297
rect 5652 3263 5664 3297
rect 5606 3237 5664 3263
rect 5706 3297 5764 3323
rect 5706 3263 5718 3297
rect 5752 3263 5764 3297
rect 5706 3237 5764 3263
rect 5806 3297 5864 3323
rect 5806 3263 5818 3297
rect 5852 3263 5864 3297
rect 5806 3237 5864 3263
rect 5906 3297 5964 3323
rect 5906 3263 5918 3297
rect 5952 3263 5964 3297
rect 5906 3237 5964 3263
rect 6006 3297 6064 3323
rect 6006 3263 6018 3297
rect 6052 3263 6064 3297
rect 6006 3237 6064 3263
rect 6106 3297 6164 3323
rect 6106 3263 6118 3297
rect 6152 3263 6164 3297
rect 6106 3237 6164 3263
rect 6206 3297 6264 3323
rect 6206 3263 6218 3297
rect 6252 3263 6264 3297
rect 6206 3237 6264 3263
rect 6306 3297 6364 3323
rect 6306 3263 6318 3297
rect 6352 3263 6364 3297
rect 6306 3237 6364 3263
rect 6406 3297 6464 3323
rect 6406 3263 6418 3297
rect 6452 3263 6464 3297
rect 6406 3237 6464 3263
rect 6506 3297 6564 3323
rect 6506 3263 6518 3297
rect 6552 3263 6564 3297
rect 6506 3237 6564 3263
rect 6606 3297 6664 3323
rect 6606 3263 6618 3297
rect 6652 3263 6664 3297
rect 6606 3237 6664 3263
rect 6706 3297 6764 3323
rect 6706 3263 6718 3297
rect 6752 3263 6764 3297
rect 6706 3237 6764 3263
rect 6806 3297 6864 3323
rect 6806 3263 6818 3297
rect 6852 3263 6864 3297
rect 6806 3237 6864 3263
rect 6906 3297 6964 3323
rect 6906 3263 6918 3297
rect 6952 3263 6964 3297
rect 6906 3237 6964 3263
rect 7006 3297 7064 3323
rect 7006 3263 7018 3297
rect 7052 3263 7064 3297
rect 7006 3237 7064 3263
rect 7106 3297 7164 3323
rect 7106 3263 7118 3297
rect 7152 3263 7164 3297
rect 7106 3237 7164 3263
rect 7206 3297 7264 3323
rect 7206 3263 7218 3297
rect 7252 3263 7264 3297
rect 7206 3237 7264 3263
rect 7306 3297 7364 3323
rect 7306 3263 7312 3297
rect 7352 3263 7364 3297
rect 7306 3237 7364 3263
rect 7406 3297 7464 3323
rect 7406 3263 7418 3297
rect 7458 3263 7464 3297
rect 7406 3237 7464 3263
rect 7506 3297 7564 3323
rect 7506 3263 7518 3297
rect 7552 3263 7564 3297
rect 7506 3237 7564 3263
rect 7606 3297 7664 3323
rect 7606 3263 7618 3297
rect 7652 3263 7664 3297
rect 7606 3237 7664 3263
rect 7706 3297 7764 3323
rect 7706 3263 7718 3297
rect 7752 3263 7764 3297
rect 7706 3237 7764 3263
rect 7806 3297 7864 3323
rect 7806 3263 7818 3297
rect 7852 3263 7864 3297
rect 7806 3237 7864 3263
rect 7906 3297 7964 3323
rect 7906 3263 7918 3297
rect 7952 3263 7964 3297
rect 7906 3237 7964 3263
rect 8006 3297 8064 3323
rect 8006 3263 8018 3297
rect 8052 3263 8064 3297
rect 8006 3237 8064 3263
rect 8106 3297 8164 3323
rect 8106 3263 8118 3297
rect 8152 3263 8164 3297
rect 8106 3237 8164 3263
rect 8206 3297 8264 3323
rect 8206 3263 8218 3297
rect 8252 3263 8264 3297
rect 8206 3237 8264 3263
rect 8306 3297 8364 3323
rect 8306 3263 8318 3297
rect 8352 3263 8364 3297
rect 8306 3237 8364 3263
rect 8406 3297 8464 3323
rect 8406 3263 8418 3297
rect 8452 3263 8464 3297
rect 8406 3237 8464 3263
rect 8506 3297 8564 3323
rect 8506 3263 8518 3297
rect 8552 3263 8564 3297
rect 8506 3237 8564 3263
rect 8606 3297 8664 3323
rect 8606 3263 8618 3297
rect 8652 3263 8664 3297
rect 8606 3237 8664 3263
rect 8706 3297 8764 3323
rect 8706 3263 8718 3297
rect 8752 3263 8764 3297
rect 8706 3237 8764 3263
rect 8806 3297 8864 3323
rect 8806 3263 8818 3297
rect 8852 3263 8864 3297
rect 8806 3237 8864 3263
rect 8906 3297 8964 3323
rect 8906 3263 8918 3297
rect 8952 3263 8964 3297
rect 8906 3237 8964 3263
rect 9006 3297 9064 3323
rect 9006 3263 9018 3297
rect 9052 3263 9064 3297
rect 9006 3237 9064 3263
rect 9106 3297 9164 3323
rect 9106 3263 9118 3297
rect 9152 3263 9164 3297
rect 9106 3237 9164 3263
rect 9206 3297 9264 3323
rect 9206 3263 9218 3297
rect 9252 3263 9264 3297
rect 9206 3237 9264 3263
rect 9306 3297 9364 3323
rect 9306 3263 9318 3297
rect 9352 3263 9364 3297
rect 9306 3237 9364 3263
rect 9406 3297 9464 3323
rect 9406 3263 9418 3297
rect 9452 3263 9464 3297
rect 9406 3237 9464 3263
rect 9506 3297 9564 3323
rect 9506 3263 9512 3297
rect 9552 3263 9564 3297
rect 9506 3237 9564 3263
rect 9606 3297 9664 3323
rect 9606 3263 9618 3297
rect 9658 3263 9664 3297
rect 9606 3237 9664 3263
rect 9706 3297 9764 3323
rect 9706 3263 9718 3297
rect 9752 3263 9764 3297
rect 9706 3237 9764 3263
rect 9806 3297 9864 3323
rect 9806 3263 9818 3297
rect 9852 3263 9864 3297
rect 9806 3237 9864 3263
rect 9906 3297 9964 3323
rect 9906 3263 9918 3297
rect 9952 3263 9964 3297
rect 9906 3237 9964 3263
rect 10006 3297 10064 3323
rect 10006 3263 10018 3297
rect 10052 3263 10064 3297
rect 10006 3237 10064 3263
rect 10106 3297 10164 3323
rect 10106 3263 10118 3297
rect 10152 3263 10164 3297
rect 10106 3237 10164 3263
rect 10206 3297 10264 3323
rect 10206 3263 10218 3297
rect 10252 3263 10264 3297
rect 10206 3237 10264 3263
rect 10306 3297 10364 3323
rect 10306 3263 10312 3297
rect 10352 3263 10364 3297
rect 10306 3237 10364 3263
rect 10406 3297 10464 3323
rect 10406 3263 10418 3297
rect 10458 3263 10464 3297
rect 10406 3237 10464 3263
rect 10506 3297 10564 3323
rect 10506 3263 10512 3297
rect 10552 3263 10564 3297
rect 10506 3237 10564 3263
rect 10606 3297 10664 3323
rect 10606 3263 10618 3297
rect 10658 3263 10664 3297
rect 10606 3237 10664 3263
rect 10706 3297 10764 3323
rect 10706 3263 10718 3297
rect 10752 3263 10764 3297
rect 10706 3237 10764 3263
rect 10806 3297 10864 3323
rect 10806 3263 10818 3297
rect 10852 3263 10864 3297
rect 10806 3237 10864 3263
rect 10906 3297 10964 3323
rect 10906 3263 10918 3297
rect 10952 3263 10964 3297
rect 10906 3237 10964 3263
rect 11006 3297 11064 3323
rect 11006 3263 11018 3297
rect 11052 3263 11064 3297
rect 11006 3237 11064 3263
rect 11106 3297 11164 3323
rect 11106 3263 11118 3297
rect 11152 3263 11164 3297
rect 11106 3237 11164 3263
rect 11206 3297 11264 3323
rect 11206 3263 11218 3297
rect 11252 3263 11264 3297
rect 11206 3237 11264 3263
rect 11306 3297 11364 3323
rect 11306 3263 11318 3297
rect 11352 3263 11364 3297
rect 11306 3237 11364 3263
rect 11406 3297 11464 3323
rect 11406 3263 11418 3297
rect 11452 3263 11464 3297
rect 11406 3237 11464 3263
rect 11506 3297 11564 3323
rect 11506 3263 11518 3297
rect 11552 3263 11564 3297
rect 11506 3237 11564 3263
rect 11606 3297 11664 3323
rect 11606 3263 11618 3297
rect 11652 3263 11664 3297
rect 11606 3237 11664 3263
rect 11706 3297 11764 3323
rect 11706 3263 11718 3297
rect 11752 3263 11764 3297
rect 11706 3237 11764 3263
rect 11806 3297 11864 3323
rect 11806 3263 11818 3297
rect 11852 3263 11864 3297
rect 11806 3237 11864 3263
rect 11906 3297 11964 3323
rect 11906 3263 11918 3297
rect 11952 3263 11964 3297
rect 11906 3237 11964 3263
rect 12006 3297 12064 3323
rect 12006 3263 12018 3297
rect 12052 3263 12064 3297
rect 12006 3237 12064 3263
rect 12106 3297 12164 3323
rect 12106 3263 12118 3297
rect 12152 3263 12164 3297
rect 12106 3237 12164 3263
rect 12206 3297 12264 3323
rect 12206 3263 12218 3297
rect 12252 3263 12264 3297
rect 12206 3237 12264 3263
rect 12306 3297 12364 3323
rect 12306 3263 12318 3297
rect 12352 3263 12364 3297
rect 12306 3237 12364 3263
rect 12406 3297 12464 3323
rect 12406 3263 12412 3297
rect 12452 3263 12464 3297
rect 12406 3237 12464 3263
rect 12506 3297 12564 3323
rect 12506 3263 12518 3297
rect 12558 3263 12564 3297
rect 12506 3237 12564 3263
rect 12606 3297 12664 3323
rect 12606 3263 12618 3297
rect 12652 3263 12664 3297
rect 12606 3237 12664 3263
rect 12706 3297 12764 3323
rect 12706 3263 12718 3297
rect 12752 3263 12764 3297
rect 12706 3237 12764 3263
rect 12806 3297 12864 3323
rect 13018 3316 13262 3350
rect 12806 3263 12818 3297
rect 12852 3263 12864 3297
rect 12908 3278 12916 3312
rect 12958 3278 12974 3312
rect 13018 3297 13052 3316
rect 12806 3237 12864 3263
rect 13228 3313 13262 3316
rect 13228 3297 13362 3313
rect 13018 3247 13052 3263
rect 13096 3248 13112 3282
rect 13154 3248 13162 3282
rect 13262 3263 13328 3297
rect 13228 3247 13362 3263
rect 13428 3297 13462 3313
rect 13428 3247 13462 3263
rect 13528 3297 13662 3313
rect 13562 3263 13628 3297
rect 13528 3247 13662 3263
rect 6 3157 64 3183
rect 6 3123 18 3157
rect 58 3123 64 3157
rect 6 3097 64 3123
rect 106 3157 164 3183
rect 106 3123 112 3157
rect 152 3123 164 3157
rect 106 3097 164 3123
rect 206 3157 264 3183
rect 206 3123 218 3157
rect 258 3123 264 3157
rect 206 3097 264 3123
rect 306 3157 364 3183
rect 306 3123 318 3157
rect 352 3123 364 3157
rect 306 3097 364 3123
rect 406 3157 464 3183
rect 406 3123 418 3157
rect 452 3123 464 3157
rect 406 3097 464 3123
rect 506 3157 564 3183
rect 506 3123 518 3157
rect 552 3123 564 3157
rect 506 3097 564 3123
rect 606 3157 664 3183
rect 606 3123 618 3157
rect 652 3123 664 3157
rect 606 3097 664 3123
rect 706 3157 764 3183
rect 706 3123 718 3157
rect 752 3123 764 3157
rect 706 3097 764 3123
rect 806 3157 864 3183
rect 806 3123 818 3157
rect 852 3123 864 3157
rect 806 3097 864 3123
rect 906 3157 964 3183
rect 906 3123 918 3157
rect 952 3123 964 3157
rect 906 3097 964 3123
rect 1006 3157 1064 3183
rect 1006 3123 1018 3157
rect 1052 3123 1064 3157
rect 1006 3097 1064 3123
rect 1106 3157 1164 3183
rect 1106 3123 1118 3157
rect 1152 3123 1164 3157
rect 1106 3097 1164 3123
rect 1206 3157 1264 3183
rect 1206 3123 1218 3157
rect 1252 3123 1264 3157
rect 1206 3097 1264 3123
rect 1306 3157 1364 3183
rect 1306 3123 1312 3157
rect 1352 3123 1364 3157
rect 1306 3097 1364 3123
rect 1406 3157 1464 3183
rect 1406 3123 1418 3157
rect 1458 3123 1464 3157
rect 1406 3097 1464 3123
rect 1506 3157 1564 3183
rect 1506 3123 1518 3157
rect 1552 3123 1564 3157
rect 1506 3097 1564 3123
rect 1606 3157 1664 3183
rect 1606 3123 1618 3157
rect 1652 3123 1664 3157
rect 1606 3097 1664 3123
rect 1706 3157 1764 3183
rect 1706 3123 1718 3157
rect 1752 3123 1764 3157
rect 1706 3097 1764 3123
rect 1806 3157 1864 3183
rect 1806 3123 1818 3157
rect 1852 3123 1864 3157
rect 1806 3097 1864 3123
rect 1906 3157 1964 3183
rect 1906 3123 1918 3157
rect 1952 3123 1964 3157
rect 1906 3097 1964 3123
rect 2006 3157 2064 3183
rect 2006 3123 2018 3157
rect 2052 3123 2064 3157
rect 2006 3097 2064 3123
rect 2106 3157 2164 3183
rect 2106 3123 2118 3157
rect 2152 3123 2164 3157
rect 2106 3097 2164 3123
rect 2206 3157 2264 3183
rect 2206 3123 2218 3157
rect 2252 3123 2264 3157
rect 2206 3097 2264 3123
rect 2306 3157 2364 3183
rect 2306 3123 2318 3157
rect 2352 3123 2364 3157
rect 2306 3097 2364 3123
rect 2406 3157 2464 3183
rect 2406 3123 2418 3157
rect 2452 3123 2464 3157
rect 2406 3097 2464 3123
rect 2506 3157 2564 3183
rect 2506 3123 2512 3157
rect 2552 3123 2564 3157
rect 2506 3097 2564 3123
rect 2606 3157 2664 3183
rect 2606 3123 2618 3157
rect 2658 3123 2664 3157
rect 2606 3097 2664 3123
rect 2706 3157 2764 3183
rect 2706 3123 2718 3157
rect 2752 3123 2764 3157
rect 2706 3097 2764 3123
rect 2806 3157 2864 3183
rect 2806 3123 2818 3157
rect 2852 3123 2864 3157
rect 2806 3097 2864 3123
rect 2906 3157 2964 3183
rect 2906 3123 2918 3157
rect 2952 3123 2964 3157
rect 2906 3097 2964 3123
rect 3006 3157 3064 3183
rect 3006 3123 3018 3157
rect 3052 3123 3064 3157
rect 3006 3097 3064 3123
rect 3106 3157 3164 3183
rect 3106 3123 3118 3157
rect 3152 3123 3164 3157
rect 3106 3097 3164 3123
rect 3206 3157 3264 3183
rect 3206 3123 3212 3157
rect 3252 3123 3264 3157
rect 3206 3097 3264 3123
rect 3306 3157 3364 3183
rect 3306 3123 3318 3157
rect 3358 3123 3364 3157
rect 3306 3097 3364 3123
rect 3406 3157 3464 3183
rect 3406 3123 3418 3157
rect 3452 3123 3464 3157
rect 3406 3097 3464 3123
rect 3506 3157 3564 3183
rect 3506 3123 3518 3157
rect 3552 3123 3564 3157
rect 3506 3097 3564 3123
rect 3606 3157 3664 3183
rect 3606 3123 3612 3157
rect 3652 3123 3664 3157
rect 3606 3097 3664 3123
rect 3706 3157 3764 3183
rect 3706 3123 3718 3157
rect 3758 3123 3764 3157
rect 3706 3097 3764 3123
rect 3806 3157 3864 3183
rect 3806 3123 3818 3157
rect 3852 3123 3864 3157
rect 3806 3097 3864 3123
rect 3906 3157 3964 3183
rect 3906 3123 3918 3157
rect 3952 3123 3964 3157
rect 3906 3097 3964 3123
rect 4006 3157 4064 3183
rect 4006 3123 4018 3157
rect 4052 3123 4064 3157
rect 4006 3097 4064 3123
rect 4106 3157 4164 3183
rect 4106 3123 4118 3157
rect 4152 3123 4164 3157
rect 4106 3097 4164 3123
rect 4206 3157 4264 3183
rect 4206 3123 4218 3157
rect 4252 3123 4264 3157
rect 4206 3097 4264 3123
rect 4306 3157 4364 3183
rect 4306 3123 4318 3157
rect 4352 3123 4364 3157
rect 4306 3097 4364 3123
rect 4406 3157 4464 3183
rect 4406 3123 4418 3157
rect 4452 3123 4464 3157
rect 4406 3097 4464 3123
rect 4506 3157 4564 3183
rect 4506 3123 4518 3157
rect 4552 3123 4564 3157
rect 4506 3097 4564 3123
rect 4606 3157 4664 3183
rect 4606 3123 4618 3157
rect 4652 3123 4664 3157
rect 4606 3097 4664 3123
rect 4706 3157 4764 3183
rect 4706 3123 4718 3157
rect 4752 3123 4764 3157
rect 4706 3097 4764 3123
rect 4806 3157 4864 3183
rect 4806 3123 4818 3157
rect 4852 3123 4864 3157
rect 4806 3097 4864 3123
rect 4906 3157 4964 3183
rect 4906 3123 4918 3157
rect 4952 3123 4964 3157
rect 4906 3097 4964 3123
rect 5006 3157 5064 3183
rect 5006 3123 5018 3157
rect 5052 3123 5064 3157
rect 5006 3097 5064 3123
rect 5106 3157 5164 3183
rect 5106 3123 5118 3157
rect 5152 3123 5164 3157
rect 5106 3097 5164 3123
rect 5206 3157 5264 3183
rect 5206 3123 5218 3157
rect 5252 3123 5264 3157
rect 5206 3097 5264 3123
rect 5306 3157 5364 3183
rect 5306 3123 5318 3157
rect 5352 3123 5364 3157
rect 5306 3097 5364 3123
rect 5406 3157 5464 3183
rect 5406 3123 5412 3157
rect 5452 3123 5464 3157
rect 5406 3097 5464 3123
rect 5506 3157 5564 3183
rect 5506 3123 5518 3157
rect 5558 3123 5564 3157
rect 5506 3097 5564 3123
rect 5606 3157 5664 3183
rect 5606 3123 5612 3157
rect 5652 3123 5664 3157
rect 5606 3097 5664 3123
rect 5706 3157 5764 3183
rect 5706 3123 5718 3157
rect 5758 3123 5764 3157
rect 5706 3097 5764 3123
rect 5806 3157 5864 3183
rect 5806 3123 5812 3157
rect 5852 3123 5864 3157
rect 5806 3097 5864 3123
rect 5906 3157 5964 3183
rect 5906 3123 5918 3157
rect 5958 3123 5964 3157
rect 5906 3097 5964 3123
rect 6006 3157 6064 3183
rect 6006 3123 6018 3157
rect 6052 3123 6064 3157
rect 6006 3097 6064 3123
rect 6106 3157 6164 3183
rect 6106 3123 6118 3157
rect 6152 3123 6164 3157
rect 6106 3097 6164 3123
rect 6206 3157 6264 3183
rect 6206 3123 6218 3157
rect 6252 3123 6264 3157
rect 6206 3097 6264 3123
rect 6306 3157 6364 3183
rect 6306 3123 6312 3157
rect 6352 3123 6364 3157
rect 6306 3097 6364 3123
rect 6406 3157 6464 3183
rect 6406 3123 6418 3157
rect 6458 3123 6464 3157
rect 6406 3097 6464 3123
rect 6506 3157 6564 3183
rect 6506 3123 6512 3157
rect 6552 3123 6564 3157
rect 6506 3097 6564 3123
rect 6606 3157 6664 3183
rect 6606 3123 6618 3157
rect 6658 3123 6664 3157
rect 6606 3097 6664 3123
rect 6706 3157 6764 3183
rect 6706 3123 6718 3157
rect 6752 3123 6764 3157
rect 6706 3097 6764 3123
rect 6806 3157 6864 3183
rect 6806 3123 6818 3157
rect 6852 3123 6864 3157
rect 6806 3097 6864 3123
rect 6906 3157 6964 3183
rect 6906 3123 6918 3157
rect 6952 3123 6964 3157
rect 6906 3097 6964 3123
rect 7006 3157 7064 3183
rect 7006 3123 7012 3157
rect 7052 3123 7064 3157
rect 7006 3097 7064 3123
rect 7106 3157 7164 3183
rect 7106 3123 7118 3157
rect 7158 3123 7164 3157
rect 7106 3097 7164 3123
rect 7206 3157 7264 3183
rect 7206 3123 7218 3157
rect 7252 3123 7264 3157
rect 7206 3097 7264 3123
rect 7306 3157 7364 3183
rect 7306 3123 7318 3157
rect 7352 3123 7364 3157
rect 7306 3097 7364 3123
rect 7406 3157 7464 3183
rect 7406 3123 7418 3157
rect 7452 3123 7464 3157
rect 7406 3097 7464 3123
rect 7506 3157 7564 3183
rect 7506 3123 7518 3157
rect 7552 3123 7564 3157
rect 7506 3097 7564 3123
rect 7606 3157 7664 3183
rect 7606 3123 7618 3157
rect 7652 3123 7664 3157
rect 7606 3097 7664 3123
rect 7706 3157 7764 3183
rect 7706 3123 7718 3157
rect 7752 3123 7764 3157
rect 7706 3097 7764 3123
rect 7806 3157 7864 3183
rect 7806 3123 7818 3157
rect 7852 3123 7864 3157
rect 7806 3097 7864 3123
rect 7906 3157 7964 3183
rect 7906 3123 7918 3157
rect 7952 3123 7964 3157
rect 7906 3097 7964 3123
rect 8006 3157 8064 3183
rect 8006 3123 8018 3157
rect 8052 3123 8064 3157
rect 8006 3097 8064 3123
rect 8106 3157 8164 3183
rect 8106 3123 8112 3157
rect 8152 3123 8164 3157
rect 8106 3097 8164 3123
rect 8206 3157 8264 3183
rect 8206 3123 8218 3157
rect 8258 3123 8264 3157
rect 8206 3097 8264 3123
rect 8306 3157 8364 3183
rect 8306 3123 8318 3157
rect 8352 3123 8364 3157
rect 8306 3097 8364 3123
rect 8406 3157 8464 3183
rect 8406 3123 8418 3157
rect 8452 3123 8464 3157
rect 8406 3097 8464 3123
rect 8506 3157 8564 3183
rect 8506 3123 8518 3157
rect 8552 3123 8564 3157
rect 8506 3097 8564 3123
rect 8606 3157 8664 3183
rect 8606 3123 8618 3157
rect 8652 3123 8664 3157
rect 8606 3097 8664 3123
rect 8706 3157 8764 3183
rect 8706 3123 8718 3157
rect 8752 3123 8764 3157
rect 8706 3097 8764 3123
rect 8806 3157 8864 3183
rect 8806 3123 8812 3157
rect 8852 3123 8864 3157
rect 8806 3097 8864 3123
rect 8906 3157 8964 3183
rect 8906 3123 8918 3157
rect 8958 3123 8964 3157
rect 8906 3097 8964 3123
rect 9006 3157 9064 3183
rect 9006 3123 9018 3157
rect 9052 3123 9064 3157
rect 9006 3097 9064 3123
rect 9106 3157 9164 3183
rect 9106 3123 9118 3157
rect 9152 3123 9164 3157
rect 9106 3097 9164 3123
rect 9206 3157 9264 3183
rect 9206 3123 9218 3157
rect 9252 3123 9264 3157
rect 9206 3097 9264 3123
rect 9306 3157 9364 3183
rect 9306 3123 9318 3157
rect 9352 3123 9364 3157
rect 9306 3097 9364 3123
rect 9406 3157 9464 3183
rect 9406 3123 9418 3157
rect 9452 3123 9464 3157
rect 9406 3097 9464 3123
rect 9506 3157 9564 3183
rect 9506 3123 9518 3157
rect 9552 3123 9564 3157
rect 9506 3097 9564 3123
rect 9606 3157 9664 3183
rect 9606 3123 9618 3157
rect 9652 3123 9664 3157
rect 9606 3097 9664 3123
rect 9706 3157 9764 3183
rect 9706 3123 9718 3157
rect 9752 3123 9764 3157
rect 9706 3097 9764 3123
rect 9806 3157 9864 3183
rect 9806 3123 9818 3157
rect 9852 3123 9864 3157
rect 9806 3097 9864 3123
rect 9906 3157 9964 3183
rect 9906 3123 9912 3157
rect 9952 3123 9964 3157
rect 9906 3097 9964 3123
rect 10006 3157 10064 3183
rect 10006 3123 10018 3157
rect 10058 3123 10064 3157
rect 10006 3097 10064 3123
rect 10106 3157 10164 3183
rect 10106 3123 10112 3157
rect 10152 3123 10164 3157
rect 10106 3097 10164 3123
rect 10206 3157 10264 3183
rect 10206 3123 10218 3157
rect 10258 3123 10264 3157
rect 10206 3097 10264 3123
rect 10306 3157 10364 3183
rect 10306 3123 10312 3157
rect 10352 3123 10364 3157
rect 10306 3097 10364 3123
rect 10406 3157 10464 3183
rect 10406 3123 10418 3157
rect 10458 3123 10464 3157
rect 10406 3097 10464 3123
rect 10506 3157 10564 3183
rect 10506 3123 10518 3157
rect 10552 3123 10564 3157
rect 10506 3097 10564 3123
rect 10606 3157 10664 3183
rect 10606 3123 10618 3157
rect 10652 3123 10664 3157
rect 10606 3097 10664 3123
rect 10706 3157 10764 3183
rect 10706 3123 10718 3157
rect 10752 3123 10764 3157
rect 10706 3097 10764 3123
rect 10806 3157 10864 3183
rect 10806 3123 10812 3157
rect 10852 3123 10864 3157
rect 10806 3097 10864 3123
rect 10906 3157 10964 3183
rect 10906 3123 10918 3157
rect 10958 3123 10964 3157
rect 10906 3097 10964 3123
rect 11006 3157 11064 3183
rect 11006 3123 11018 3157
rect 11052 3123 11064 3157
rect 11006 3097 11064 3123
rect 11106 3157 11164 3183
rect 11106 3123 11118 3157
rect 11152 3123 11164 3157
rect 11106 3097 11164 3123
rect 11206 3157 11264 3183
rect 11206 3123 11218 3157
rect 11252 3123 11264 3157
rect 11206 3097 11264 3123
rect 11306 3157 11364 3183
rect 11306 3123 11318 3157
rect 11352 3123 11364 3157
rect 11306 3097 11364 3123
rect 11406 3157 11464 3183
rect 11406 3123 11418 3157
rect 11452 3123 11464 3157
rect 11406 3097 11464 3123
rect 11506 3157 11564 3183
rect 11506 3123 11512 3157
rect 11552 3123 11564 3157
rect 11506 3097 11564 3123
rect 11606 3157 11664 3183
rect 11606 3123 11618 3157
rect 11658 3123 11664 3157
rect 11606 3097 11664 3123
rect 11706 3157 11764 3183
rect 11706 3123 11718 3157
rect 11752 3123 11764 3157
rect 11706 3097 11764 3123
rect 11806 3157 11864 3183
rect 11806 3123 11818 3157
rect 11852 3123 11864 3157
rect 11806 3097 11864 3123
rect 11906 3157 11964 3183
rect 11906 3123 11918 3157
rect 11952 3123 11964 3157
rect 11906 3097 11964 3123
rect 12006 3157 12064 3183
rect 12006 3123 12018 3157
rect 12052 3123 12064 3157
rect 12006 3097 12064 3123
rect 12106 3157 12164 3183
rect 12106 3123 12118 3157
rect 12152 3123 12164 3157
rect 12106 3097 12164 3123
rect 12206 3157 12264 3183
rect 12206 3123 12218 3157
rect 12252 3123 12264 3157
rect 12206 3097 12264 3123
rect 12306 3157 12364 3183
rect 12306 3123 12318 3157
rect 12352 3123 12364 3157
rect 12306 3097 12364 3123
rect 12406 3157 12464 3183
rect 12406 3123 12418 3157
rect 12452 3123 12464 3157
rect 12406 3097 12464 3123
rect 12506 3157 12564 3183
rect 12506 3123 12518 3157
rect 12552 3123 12564 3157
rect 12506 3097 12564 3123
rect 12606 3157 12664 3183
rect 12606 3123 12618 3157
rect 12652 3123 12664 3157
rect 12606 3097 12664 3123
rect 12706 3157 12764 3183
rect 12706 3123 12718 3157
rect 12752 3123 12764 3157
rect 12706 3097 12764 3123
rect 12806 3157 12864 3183
rect 13018 3176 13262 3210
rect 12806 3123 12818 3157
rect 12852 3123 12864 3157
rect 12908 3138 12916 3172
rect 12958 3138 12974 3172
rect 13018 3157 13052 3176
rect 12806 3097 12864 3123
rect 13228 3157 13262 3176
rect 13018 3107 13052 3123
rect 13096 3108 13112 3142
rect 13154 3108 13162 3142
rect 13228 3107 13262 3123
rect 13328 3157 13462 3173
rect 13362 3123 13428 3157
rect 13328 3107 13462 3123
rect 13528 3157 13662 3173
rect 13562 3123 13628 3157
rect 13528 3107 13662 3123
rect 6 3017 64 3043
rect 6 2983 18 3017
rect 52 2983 64 3017
rect 6 2957 64 2983
rect 106 3017 164 3043
rect 106 2983 118 3017
rect 152 2983 164 3017
rect 106 2957 164 2983
rect 206 3017 264 3043
rect 206 2983 218 3017
rect 252 2983 264 3017
rect 206 2957 264 2983
rect 306 3017 364 3043
rect 306 2983 318 3017
rect 352 2983 364 3017
rect 306 2957 364 2983
rect 406 3017 464 3043
rect 406 2983 418 3017
rect 452 2983 464 3017
rect 406 2957 464 2983
rect 506 3017 564 3043
rect 506 2983 518 3017
rect 552 2983 564 3017
rect 506 2957 564 2983
rect 606 3017 664 3043
rect 606 2983 612 3017
rect 652 2983 664 3017
rect 606 2957 664 2983
rect 706 3017 764 3043
rect 706 2983 718 3017
rect 758 2983 764 3017
rect 706 2957 764 2983
rect 806 3017 864 3043
rect 806 2983 818 3017
rect 852 2983 864 3017
rect 806 2957 864 2983
rect 906 3017 964 3043
rect 906 2983 918 3017
rect 952 2983 964 3017
rect 906 2957 964 2983
rect 1006 3017 1064 3043
rect 1006 2983 1018 3017
rect 1052 2983 1064 3017
rect 1006 2957 1064 2983
rect 1106 3017 1164 3043
rect 1106 2983 1118 3017
rect 1152 2983 1164 3017
rect 1106 2957 1164 2983
rect 1206 3017 1264 3043
rect 1206 2983 1218 3017
rect 1252 2983 1264 3017
rect 1206 2957 1264 2983
rect 1306 3017 1364 3043
rect 1306 2983 1318 3017
rect 1352 2983 1364 3017
rect 1306 2957 1364 2983
rect 1406 3017 1464 3043
rect 1406 2983 1418 3017
rect 1452 2983 1464 3017
rect 1406 2957 1464 2983
rect 1506 3017 1564 3043
rect 1506 2983 1518 3017
rect 1552 2983 1564 3017
rect 1506 2957 1564 2983
rect 1606 3017 1664 3043
rect 1606 2983 1618 3017
rect 1652 2983 1664 3017
rect 1606 2957 1664 2983
rect 1706 3017 1764 3043
rect 1706 2983 1718 3017
rect 1752 2983 1764 3017
rect 1706 2957 1764 2983
rect 1806 3017 1864 3043
rect 1806 2983 1818 3017
rect 1852 2983 1864 3017
rect 1806 2957 1864 2983
rect 1906 3017 1964 3043
rect 1906 2983 1918 3017
rect 1952 2983 1964 3017
rect 1906 2957 1964 2983
rect 2006 3017 2064 3043
rect 2006 2983 2012 3017
rect 2052 2983 2064 3017
rect 2006 2957 2064 2983
rect 2106 3017 2164 3043
rect 2106 2983 2118 3017
rect 2158 2983 2164 3017
rect 2106 2957 2164 2983
rect 2206 3017 2264 3043
rect 2206 2983 2218 3017
rect 2252 2983 2264 3017
rect 2206 2957 2264 2983
rect 2306 3017 2364 3043
rect 2306 2983 2318 3017
rect 2352 2983 2364 3017
rect 2306 2957 2364 2983
rect 2406 3017 2464 3043
rect 2406 2983 2418 3017
rect 2452 2983 2464 3017
rect 2406 2957 2464 2983
rect 2506 3017 2564 3043
rect 2506 2983 2518 3017
rect 2552 2983 2564 3017
rect 2506 2957 2564 2983
rect 2606 3017 2664 3043
rect 2606 2983 2618 3017
rect 2652 2983 2664 3017
rect 2606 2957 2664 2983
rect 2706 3017 2764 3043
rect 2706 2983 2718 3017
rect 2752 2983 2764 3017
rect 2706 2957 2764 2983
rect 2806 3017 2864 3043
rect 2806 2983 2818 3017
rect 2852 2983 2864 3017
rect 2806 2957 2864 2983
rect 2906 3017 2964 3043
rect 2906 2983 2918 3017
rect 2952 2983 2964 3017
rect 2906 2957 2964 2983
rect 3006 3017 3064 3043
rect 3006 2983 3012 3017
rect 3052 2983 3064 3017
rect 3006 2957 3064 2983
rect 3106 3017 3164 3043
rect 3106 2983 3118 3017
rect 3158 2983 3164 3017
rect 3106 2957 3164 2983
rect 3206 3017 3264 3043
rect 3206 2983 3218 3017
rect 3252 2983 3264 3017
rect 3206 2957 3264 2983
rect 3306 3017 3364 3043
rect 3306 2983 3318 3017
rect 3352 2983 3364 3017
rect 3306 2957 3364 2983
rect 3406 3017 3464 3043
rect 3406 2983 3418 3017
rect 3452 2983 3464 3017
rect 3406 2957 3464 2983
rect 3506 3017 3564 3043
rect 3506 2983 3518 3017
rect 3552 2983 3564 3017
rect 3506 2957 3564 2983
rect 3606 3017 3664 3043
rect 3606 2983 3618 3017
rect 3652 2983 3664 3017
rect 3606 2957 3664 2983
rect 3706 3017 3764 3043
rect 3706 2983 3718 3017
rect 3752 2983 3764 3017
rect 3706 2957 3764 2983
rect 3806 3017 3864 3043
rect 3806 2983 3812 3017
rect 3852 2983 3864 3017
rect 3806 2957 3864 2983
rect 3906 3017 3964 3043
rect 3906 2983 3918 3017
rect 3958 2983 3964 3017
rect 3906 2957 3964 2983
rect 4006 3017 4064 3043
rect 4006 2983 4018 3017
rect 4052 2983 4064 3017
rect 4006 2957 4064 2983
rect 4106 3017 4164 3043
rect 4106 2983 4118 3017
rect 4152 2983 4164 3017
rect 4106 2957 4164 2983
rect 4206 3017 4264 3043
rect 4206 2983 4218 3017
rect 4252 2983 4264 3017
rect 4206 2957 4264 2983
rect 4306 3017 4364 3043
rect 4306 2983 4318 3017
rect 4352 2983 4364 3017
rect 4306 2957 4364 2983
rect 4406 3017 4464 3043
rect 4406 2983 4418 3017
rect 4452 2983 4464 3017
rect 4406 2957 4464 2983
rect 4506 3017 4564 3043
rect 4506 2983 4512 3017
rect 4552 2983 4564 3017
rect 4506 2957 4564 2983
rect 4606 3017 4664 3043
rect 4606 2983 4618 3017
rect 4658 2983 4664 3017
rect 4606 2957 4664 2983
rect 4706 3017 4764 3043
rect 4706 2983 4718 3017
rect 4752 2983 4764 3017
rect 4706 2957 4764 2983
rect 4806 3017 4864 3043
rect 4806 2983 4818 3017
rect 4852 2983 4864 3017
rect 4806 2957 4864 2983
rect 4906 3017 4964 3043
rect 4906 2983 4912 3017
rect 4952 2983 4964 3017
rect 4906 2957 4964 2983
rect 5006 3017 5064 3043
rect 5006 2983 5018 3017
rect 5058 2983 5064 3017
rect 5006 2957 5064 2983
rect 5106 3017 5164 3043
rect 5106 2983 5118 3017
rect 5152 2983 5164 3017
rect 5106 2957 5164 2983
rect 5206 3017 5264 3043
rect 5206 2983 5218 3017
rect 5252 2983 5264 3017
rect 5206 2957 5264 2983
rect 5306 3017 5364 3043
rect 5306 2983 5318 3017
rect 5352 2983 5364 3017
rect 5306 2957 5364 2983
rect 5406 3017 5464 3043
rect 5406 2983 5418 3017
rect 5452 2983 5464 3017
rect 5406 2957 5464 2983
rect 5506 3017 5564 3043
rect 5506 2983 5518 3017
rect 5552 2983 5564 3017
rect 5506 2957 5564 2983
rect 5606 3017 5664 3043
rect 5606 2983 5618 3017
rect 5652 2983 5664 3017
rect 5606 2957 5664 2983
rect 5706 3017 5764 3043
rect 5706 2983 5718 3017
rect 5752 2983 5764 3017
rect 5706 2957 5764 2983
rect 5806 3017 5864 3043
rect 5806 2983 5818 3017
rect 5852 2983 5864 3017
rect 5806 2957 5864 2983
rect 5906 3017 5964 3043
rect 5906 2983 5912 3017
rect 5952 2983 5964 3017
rect 5906 2957 5964 2983
rect 6006 3017 6064 3043
rect 6006 2983 6018 3017
rect 6058 2983 6064 3017
rect 6006 2957 6064 2983
rect 6106 3017 6164 3043
rect 6106 2983 6118 3017
rect 6152 2983 6164 3017
rect 6106 2957 6164 2983
rect 6206 3017 6264 3043
rect 6206 2983 6218 3017
rect 6252 2983 6264 3017
rect 6206 2957 6264 2983
rect 6306 3017 6364 3043
rect 6306 2983 6318 3017
rect 6352 2983 6364 3017
rect 6306 2957 6364 2983
rect 6406 3017 6464 3043
rect 6406 2983 6418 3017
rect 6452 2983 6464 3017
rect 6406 2957 6464 2983
rect 6506 3017 6564 3043
rect 6506 2983 6518 3017
rect 6552 2983 6564 3017
rect 6506 2957 6564 2983
rect 6606 3017 6664 3043
rect 6606 2983 6618 3017
rect 6652 2983 6664 3017
rect 6606 2957 6664 2983
rect 6706 3017 6764 3043
rect 6706 2983 6718 3017
rect 6752 2983 6764 3017
rect 6706 2957 6764 2983
rect 6806 3017 6864 3043
rect 6806 2983 6818 3017
rect 6852 2983 6864 3017
rect 6806 2957 6864 2983
rect 6906 3017 6964 3043
rect 6906 2983 6918 3017
rect 6952 2983 6964 3017
rect 6906 2957 6964 2983
rect 7006 3017 7064 3043
rect 7006 2983 7018 3017
rect 7052 2983 7064 3017
rect 7006 2957 7064 2983
rect 7106 3017 7164 3043
rect 7106 2983 7118 3017
rect 7152 2983 7164 3017
rect 7106 2957 7164 2983
rect 7206 3017 7264 3043
rect 7206 2983 7218 3017
rect 7252 2983 7264 3017
rect 7206 2957 7264 2983
rect 7306 3017 7364 3043
rect 7306 2983 7318 3017
rect 7352 2983 7364 3017
rect 7306 2957 7364 2983
rect 7406 3017 7464 3043
rect 7406 2983 7418 3017
rect 7452 2983 7464 3017
rect 7406 2957 7464 2983
rect 7506 3017 7564 3043
rect 7506 2983 7518 3017
rect 7552 2983 7564 3017
rect 7506 2957 7564 2983
rect 7606 3017 7664 3043
rect 7606 2983 7618 3017
rect 7652 2983 7664 3017
rect 7606 2957 7664 2983
rect 7706 3017 7764 3043
rect 7706 2983 7718 3017
rect 7752 2983 7764 3017
rect 7706 2957 7764 2983
rect 7806 3017 7864 3043
rect 7806 2983 7818 3017
rect 7852 2983 7864 3017
rect 7806 2957 7864 2983
rect 7906 3017 7964 3043
rect 7906 2983 7918 3017
rect 7952 2983 7964 3017
rect 7906 2957 7964 2983
rect 8006 3017 8064 3043
rect 8006 2983 8012 3017
rect 8052 2983 8064 3017
rect 8006 2957 8064 2983
rect 8106 3017 8164 3043
rect 8106 2983 8118 3017
rect 8158 2983 8164 3017
rect 8106 2957 8164 2983
rect 8206 3017 8264 3043
rect 8206 2983 8218 3017
rect 8252 2983 8264 3017
rect 8206 2957 8264 2983
rect 8306 3017 8364 3043
rect 8306 2983 8318 3017
rect 8352 2983 8364 3017
rect 8306 2957 8364 2983
rect 8406 3017 8464 3043
rect 8406 2983 8418 3017
rect 8452 2983 8464 3017
rect 8406 2957 8464 2983
rect 8506 3017 8564 3043
rect 8506 2983 8518 3017
rect 8552 2983 8564 3017
rect 8506 2957 8564 2983
rect 8606 3017 8664 3043
rect 8606 2983 8618 3017
rect 8652 2983 8664 3017
rect 8606 2957 8664 2983
rect 8706 3017 8764 3043
rect 8706 2983 8718 3017
rect 8752 2983 8764 3017
rect 8706 2957 8764 2983
rect 8806 3017 8864 3043
rect 8806 2983 8812 3017
rect 8852 2983 8864 3017
rect 8806 2957 8864 2983
rect 8906 3017 8964 3043
rect 8906 2983 8918 3017
rect 8958 2983 8964 3017
rect 8906 2957 8964 2983
rect 9006 3017 9064 3043
rect 9006 2983 9018 3017
rect 9052 2983 9064 3017
rect 9006 2957 9064 2983
rect 9106 3017 9164 3043
rect 9106 2983 9112 3017
rect 9152 2983 9164 3017
rect 9106 2957 9164 2983
rect 9206 3017 9264 3043
rect 9206 2983 9218 3017
rect 9258 2983 9264 3017
rect 9206 2957 9264 2983
rect 9306 3017 9364 3043
rect 9306 2983 9318 3017
rect 9352 2983 9364 3017
rect 9306 2957 9364 2983
rect 9406 3017 9464 3043
rect 9406 2983 9412 3017
rect 9452 2983 9464 3017
rect 9406 2957 9464 2983
rect 9506 3017 9564 3043
rect 9506 2983 9518 3017
rect 9558 2983 9564 3017
rect 9506 2957 9564 2983
rect 9606 3017 9664 3043
rect 9606 2983 9618 3017
rect 9652 2983 9664 3017
rect 9606 2957 9664 2983
rect 9706 3017 9764 3043
rect 9706 2983 9718 3017
rect 9752 2983 9764 3017
rect 9706 2957 9764 2983
rect 9806 3017 9864 3043
rect 9806 2983 9818 3017
rect 9852 2983 9864 3017
rect 9806 2957 9864 2983
rect 9906 3017 9964 3043
rect 9906 2983 9918 3017
rect 9952 2983 9964 3017
rect 9906 2957 9964 2983
rect 10006 3017 10064 3043
rect 10006 2983 10018 3017
rect 10052 2983 10064 3017
rect 10006 2957 10064 2983
rect 10106 3017 10164 3043
rect 10106 2983 10118 3017
rect 10152 2983 10164 3017
rect 10106 2957 10164 2983
rect 10206 3017 10264 3043
rect 10206 2983 10218 3017
rect 10252 2983 10264 3017
rect 10206 2957 10264 2983
rect 10306 3017 10364 3043
rect 10306 2983 10318 3017
rect 10352 2983 10364 3017
rect 10306 2957 10364 2983
rect 10406 3017 10464 3043
rect 10406 2983 10418 3017
rect 10452 2983 10464 3017
rect 10406 2957 10464 2983
rect 10506 3017 10564 3043
rect 10506 2983 10518 3017
rect 10552 2983 10564 3017
rect 10506 2957 10564 2983
rect 10606 3017 10664 3043
rect 10606 2983 10618 3017
rect 10652 2983 10664 3017
rect 10606 2957 10664 2983
rect 10706 3017 10764 3043
rect 10706 2983 10718 3017
rect 10752 2983 10764 3017
rect 10706 2957 10764 2983
rect 10806 3017 10864 3043
rect 10806 2983 10818 3017
rect 10852 2983 10864 3017
rect 10806 2957 10864 2983
rect 10906 3017 10964 3043
rect 10906 2983 10918 3017
rect 10952 2983 10964 3017
rect 10906 2957 10964 2983
rect 11006 3017 11064 3043
rect 11006 2983 11018 3017
rect 11052 2983 11064 3017
rect 11006 2957 11064 2983
rect 11106 3017 11164 3043
rect 11106 2983 11118 3017
rect 11152 2983 11164 3017
rect 11106 2957 11164 2983
rect 11206 3017 11264 3043
rect 11206 2983 11218 3017
rect 11252 2983 11264 3017
rect 11206 2957 11264 2983
rect 11306 3017 11364 3043
rect 11306 2983 11318 3017
rect 11352 2983 11364 3017
rect 11306 2957 11364 2983
rect 11406 3017 11464 3043
rect 11406 2983 11418 3017
rect 11452 2983 11464 3017
rect 11406 2957 11464 2983
rect 11506 3017 11564 3043
rect 11506 2983 11512 3017
rect 11552 2983 11564 3017
rect 11506 2957 11564 2983
rect 11606 3017 11664 3043
rect 11606 2983 11618 3017
rect 11658 2983 11664 3017
rect 11606 2957 11664 2983
rect 11706 3017 11764 3043
rect 11706 2983 11718 3017
rect 11752 2983 11764 3017
rect 11706 2957 11764 2983
rect 11806 3017 11864 3043
rect 11806 2983 11818 3017
rect 11852 2983 11864 3017
rect 11806 2957 11864 2983
rect 11906 3017 11964 3043
rect 11906 2983 11918 3017
rect 11952 2983 11964 3017
rect 11906 2957 11964 2983
rect 12006 3017 12064 3043
rect 12006 2983 12018 3017
rect 12052 2983 12064 3017
rect 12006 2957 12064 2983
rect 12106 3017 12164 3043
rect 12106 2983 12118 3017
rect 12152 2983 12164 3017
rect 12106 2957 12164 2983
rect 12206 3017 12264 3043
rect 12206 2983 12218 3017
rect 12252 2983 12264 3017
rect 12206 2957 12264 2983
rect 12306 3017 12364 3043
rect 12306 2983 12318 3017
rect 12352 2983 12364 3017
rect 12306 2957 12364 2983
rect 12406 3017 12464 3043
rect 12406 2983 12418 3017
rect 12452 2983 12464 3017
rect 12406 2957 12464 2983
rect 12506 3017 12564 3043
rect 12506 2983 12518 3017
rect 12552 2983 12564 3017
rect 12506 2957 12564 2983
rect 12606 3017 12664 3043
rect 12606 2983 12618 3017
rect 12652 2983 12664 3017
rect 12606 2957 12664 2983
rect 12706 3017 12764 3043
rect 12706 2983 12718 3017
rect 12752 2983 12764 3017
rect 12706 2957 12764 2983
rect 12806 3017 12864 3043
rect 13018 3036 13262 3070
rect 12806 2983 12812 3017
rect 12852 2983 12864 3017
rect 12908 2998 12916 3032
rect 12958 2998 12974 3032
rect 13018 3017 13052 3036
rect 12806 2957 12864 2983
rect 13228 3033 13262 3036
rect 13228 3017 13362 3033
rect 13018 2967 13052 2983
rect 13096 2968 13112 3002
rect 13154 2968 13162 3002
rect 13262 2983 13328 3017
rect 13228 2967 13362 2983
rect 13428 3017 13562 3033
rect 13462 2983 13528 3017
rect 13428 2967 13562 2983
rect 13628 3017 13662 3033
rect 13628 2967 13662 2983
rect 6 2877 64 2903
rect 6 2843 18 2877
rect 58 2843 64 2877
rect 6 2817 64 2843
rect 106 2877 164 2903
rect 106 2843 118 2877
rect 152 2843 164 2877
rect 106 2817 164 2843
rect 206 2877 264 2903
rect 206 2843 218 2877
rect 252 2843 264 2877
rect 206 2817 264 2843
rect 306 2877 364 2903
rect 306 2843 318 2877
rect 352 2843 364 2877
rect 306 2817 364 2843
rect 406 2877 464 2903
rect 406 2843 418 2877
rect 452 2843 464 2877
rect 406 2817 464 2843
rect 506 2877 564 2903
rect 506 2843 518 2877
rect 552 2843 564 2877
rect 506 2817 564 2843
rect 606 2877 664 2903
rect 606 2843 618 2877
rect 652 2843 664 2877
rect 606 2817 664 2843
rect 706 2877 764 2903
rect 706 2843 718 2877
rect 752 2843 764 2877
rect 706 2817 764 2843
rect 806 2877 864 2903
rect 806 2843 812 2877
rect 852 2843 864 2877
rect 806 2817 864 2843
rect 906 2877 964 2903
rect 906 2843 918 2877
rect 958 2843 964 2877
rect 906 2817 964 2843
rect 1006 2877 1064 2903
rect 1006 2843 1018 2877
rect 1052 2843 1064 2877
rect 1006 2817 1064 2843
rect 1106 2877 1164 2903
rect 1106 2843 1118 2877
rect 1152 2843 1164 2877
rect 1106 2817 1164 2843
rect 1206 2877 1264 2903
rect 1206 2843 1218 2877
rect 1252 2843 1264 2877
rect 1206 2817 1264 2843
rect 1306 2877 1364 2903
rect 1306 2843 1318 2877
rect 1352 2843 1364 2877
rect 1306 2817 1364 2843
rect 1406 2877 1464 2903
rect 1406 2843 1418 2877
rect 1452 2843 1464 2877
rect 1406 2817 1464 2843
rect 1506 2877 1564 2903
rect 1506 2843 1518 2877
rect 1552 2843 1564 2877
rect 1506 2817 1564 2843
rect 1606 2877 1664 2903
rect 1606 2843 1618 2877
rect 1652 2843 1664 2877
rect 1606 2817 1664 2843
rect 1706 2877 1764 2903
rect 1706 2843 1718 2877
rect 1752 2843 1764 2877
rect 1706 2817 1764 2843
rect 1806 2877 1864 2903
rect 1806 2843 1818 2877
rect 1852 2843 1864 2877
rect 1806 2817 1864 2843
rect 1906 2877 1964 2903
rect 1906 2843 1918 2877
rect 1952 2843 1964 2877
rect 1906 2817 1964 2843
rect 2006 2877 2064 2903
rect 2006 2843 2018 2877
rect 2052 2843 2064 2877
rect 2006 2817 2064 2843
rect 2106 2877 2164 2903
rect 2106 2843 2118 2877
rect 2152 2843 2164 2877
rect 2106 2817 2164 2843
rect 2206 2877 2264 2903
rect 2206 2843 2218 2877
rect 2252 2843 2264 2877
rect 2206 2817 2264 2843
rect 2306 2877 2364 2903
rect 2306 2843 2318 2877
rect 2352 2843 2364 2877
rect 2306 2817 2364 2843
rect 2406 2877 2464 2903
rect 2406 2843 2418 2877
rect 2452 2843 2464 2877
rect 2406 2817 2464 2843
rect 2506 2877 2564 2903
rect 2506 2843 2518 2877
rect 2552 2843 2564 2877
rect 2506 2817 2564 2843
rect 2606 2877 2664 2903
rect 2606 2843 2612 2877
rect 2652 2843 2664 2877
rect 2606 2817 2664 2843
rect 2706 2877 2764 2903
rect 2706 2843 2718 2877
rect 2758 2843 2764 2877
rect 2706 2817 2764 2843
rect 2806 2877 2864 2903
rect 2806 2843 2818 2877
rect 2852 2843 2864 2877
rect 2806 2817 2864 2843
rect 2906 2877 2964 2903
rect 2906 2843 2912 2877
rect 2952 2843 2964 2877
rect 2906 2817 2964 2843
rect 3006 2877 3064 2903
rect 3006 2843 3018 2877
rect 3058 2843 3064 2877
rect 3006 2817 3064 2843
rect 3106 2877 3164 2903
rect 3106 2843 3118 2877
rect 3152 2843 3164 2877
rect 3106 2817 3164 2843
rect 3206 2877 3264 2903
rect 3206 2843 3218 2877
rect 3252 2843 3264 2877
rect 3206 2817 3264 2843
rect 3306 2877 3364 2903
rect 3306 2843 3312 2877
rect 3352 2843 3364 2877
rect 3306 2817 3364 2843
rect 3406 2877 3464 2903
rect 3406 2843 3418 2877
rect 3458 2843 3464 2877
rect 3406 2817 3464 2843
rect 3506 2877 3564 2903
rect 3506 2843 3518 2877
rect 3552 2843 3564 2877
rect 3506 2817 3564 2843
rect 3606 2877 3664 2903
rect 3606 2843 3618 2877
rect 3652 2843 3664 2877
rect 3606 2817 3664 2843
rect 3706 2877 3764 2903
rect 3706 2843 3718 2877
rect 3752 2843 3764 2877
rect 3706 2817 3764 2843
rect 3806 2877 3864 2903
rect 3806 2843 3818 2877
rect 3852 2843 3864 2877
rect 3806 2817 3864 2843
rect 3906 2877 3964 2903
rect 3906 2843 3912 2877
rect 3952 2843 3964 2877
rect 3906 2817 3964 2843
rect 4006 2877 4064 2903
rect 4006 2843 4018 2877
rect 4058 2843 4064 2877
rect 4006 2817 4064 2843
rect 4106 2877 4164 2903
rect 4106 2843 4118 2877
rect 4152 2843 4164 2877
rect 4106 2817 4164 2843
rect 4206 2877 4264 2903
rect 4206 2843 4218 2877
rect 4252 2843 4264 2877
rect 4206 2817 4264 2843
rect 4306 2877 4364 2903
rect 4306 2843 4318 2877
rect 4352 2843 4364 2877
rect 4306 2817 4364 2843
rect 4406 2877 4464 2903
rect 4406 2843 4418 2877
rect 4452 2843 4464 2877
rect 4406 2817 4464 2843
rect 4506 2877 4564 2903
rect 4506 2843 4518 2877
rect 4552 2843 4564 2877
rect 4506 2817 4564 2843
rect 4606 2877 4664 2903
rect 4606 2843 4618 2877
rect 4652 2843 4664 2877
rect 4606 2817 4664 2843
rect 4706 2877 4764 2903
rect 4706 2843 4718 2877
rect 4752 2843 4764 2877
rect 4706 2817 4764 2843
rect 4806 2877 4864 2903
rect 4806 2843 4818 2877
rect 4852 2843 4864 2877
rect 4806 2817 4864 2843
rect 4906 2877 4964 2903
rect 4906 2843 4918 2877
rect 4952 2843 4964 2877
rect 4906 2817 4964 2843
rect 5006 2877 5064 2903
rect 5006 2843 5018 2877
rect 5052 2843 5064 2877
rect 5006 2817 5064 2843
rect 5106 2877 5164 2903
rect 5106 2843 5118 2877
rect 5152 2843 5164 2877
rect 5106 2817 5164 2843
rect 5206 2877 5264 2903
rect 5206 2843 5218 2877
rect 5252 2843 5264 2877
rect 5206 2817 5264 2843
rect 5306 2877 5364 2903
rect 5306 2843 5312 2877
rect 5352 2843 5364 2877
rect 5306 2817 5364 2843
rect 5406 2877 5464 2903
rect 5406 2843 5418 2877
rect 5458 2843 5464 2877
rect 5406 2817 5464 2843
rect 5506 2877 5564 2903
rect 5506 2843 5518 2877
rect 5552 2843 5564 2877
rect 5506 2817 5564 2843
rect 5606 2877 5664 2903
rect 5606 2843 5618 2877
rect 5652 2843 5664 2877
rect 5606 2817 5664 2843
rect 5706 2877 5764 2903
rect 5706 2843 5718 2877
rect 5752 2843 5764 2877
rect 5706 2817 5764 2843
rect 5806 2877 5864 2903
rect 5806 2843 5818 2877
rect 5852 2843 5864 2877
rect 5806 2817 5864 2843
rect 5906 2877 5964 2903
rect 5906 2843 5918 2877
rect 5952 2843 5964 2877
rect 5906 2817 5964 2843
rect 6006 2877 6064 2903
rect 6006 2843 6012 2877
rect 6052 2843 6064 2877
rect 6006 2817 6064 2843
rect 6106 2877 6164 2903
rect 6106 2843 6118 2877
rect 6158 2843 6164 2877
rect 6106 2817 6164 2843
rect 6206 2877 6264 2903
rect 6206 2843 6218 2877
rect 6252 2843 6264 2877
rect 6206 2817 6264 2843
rect 6306 2877 6364 2903
rect 6306 2843 6318 2877
rect 6352 2843 6364 2877
rect 6306 2817 6364 2843
rect 6406 2877 6464 2903
rect 6406 2843 6418 2877
rect 6452 2843 6464 2877
rect 6406 2817 6464 2843
rect 6506 2877 6564 2903
rect 6506 2843 6518 2877
rect 6552 2843 6564 2877
rect 6506 2817 6564 2843
rect 6606 2877 6664 2903
rect 6606 2843 6618 2877
rect 6652 2843 6664 2877
rect 6606 2817 6664 2843
rect 6706 2877 6764 2903
rect 6706 2843 6718 2877
rect 6752 2843 6764 2877
rect 6706 2817 6764 2843
rect 6806 2877 6864 2903
rect 6806 2843 6818 2877
rect 6852 2843 6864 2877
rect 6806 2817 6864 2843
rect 6906 2877 6964 2903
rect 6906 2843 6912 2877
rect 6952 2843 6964 2877
rect 6906 2817 6964 2843
rect 7006 2877 7064 2903
rect 7006 2843 7018 2877
rect 7058 2843 7064 2877
rect 7006 2817 7064 2843
rect 7106 2877 7164 2903
rect 7106 2843 7118 2877
rect 7152 2843 7164 2877
rect 7106 2817 7164 2843
rect 7206 2877 7264 2903
rect 7206 2843 7218 2877
rect 7252 2843 7264 2877
rect 7206 2817 7264 2843
rect 7306 2877 7364 2903
rect 7306 2843 7312 2877
rect 7352 2843 7364 2877
rect 7306 2817 7364 2843
rect 7406 2877 7464 2903
rect 7406 2843 7418 2877
rect 7458 2843 7464 2877
rect 7406 2817 7464 2843
rect 7506 2877 7564 2903
rect 7506 2843 7518 2877
rect 7552 2843 7564 2877
rect 7506 2817 7564 2843
rect 7606 2877 7664 2903
rect 7606 2843 7618 2877
rect 7652 2843 7664 2877
rect 7606 2817 7664 2843
rect 7706 2877 7764 2903
rect 7706 2843 7718 2877
rect 7752 2843 7764 2877
rect 7706 2817 7764 2843
rect 7806 2877 7864 2903
rect 7806 2843 7818 2877
rect 7852 2843 7864 2877
rect 7806 2817 7864 2843
rect 7906 2877 7964 2903
rect 7906 2843 7912 2877
rect 7952 2843 7964 2877
rect 7906 2817 7964 2843
rect 8006 2877 8064 2903
rect 8006 2843 8018 2877
rect 8058 2843 8064 2877
rect 8006 2817 8064 2843
rect 8106 2877 8164 2903
rect 8106 2843 8118 2877
rect 8152 2843 8164 2877
rect 8106 2817 8164 2843
rect 8206 2877 8264 2903
rect 8206 2843 8218 2877
rect 8252 2843 8264 2877
rect 8206 2817 8264 2843
rect 8306 2877 8364 2903
rect 8306 2843 8318 2877
rect 8352 2843 8364 2877
rect 8306 2817 8364 2843
rect 8406 2877 8464 2903
rect 8406 2843 8418 2877
rect 8452 2843 8464 2877
rect 8406 2817 8464 2843
rect 8506 2877 8564 2903
rect 8506 2843 8518 2877
rect 8552 2843 8564 2877
rect 8506 2817 8564 2843
rect 8606 2877 8664 2903
rect 8606 2843 8618 2877
rect 8652 2843 8664 2877
rect 8606 2817 8664 2843
rect 8706 2877 8764 2903
rect 8706 2843 8712 2877
rect 8752 2843 8764 2877
rect 8706 2817 8764 2843
rect 8806 2877 8864 2903
rect 8806 2843 8818 2877
rect 8858 2843 8864 2877
rect 8806 2817 8864 2843
rect 8906 2877 8964 2903
rect 8906 2843 8918 2877
rect 8952 2843 8964 2877
rect 8906 2817 8964 2843
rect 9006 2877 9064 2903
rect 9006 2843 9018 2877
rect 9052 2843 9064 2877
rect 9006 2817 9064 2843
rect 9106 2877 9164 2903
rect 9106 2843 9118 2877
rect 9152 2843 9164 2877
rect 9106 2817 9164 2843
rect 9206 2877 9264 2903
rect 9206 2843 9218 2877
rect 9252 2843 9264 2877
rect 9206 2817 9264 2843
rect 9306 2877 9364 2903
rect 9306 2843 9318 2877
rect 9352 2843 9364 2877
rect 9306 2817 9364 2843
rect 9406 2877 9464 2903
rect 9406 2843 9418 2877
rect 9452 2843 9464 2877
rect 9406 2817 9464 2843
rect 9506 2877 9564 2903
rect 9506 2843 9518 2877
rect 9552 2843 9564 2877
rect 9506 2817 9564 2843
rect 9606 2877 9664 2903
rect 9606 2843 9618 2877
rect 9652 2843 9664 2877
rect 9606 2817 9664 2843
rect 9706 2877 9764 2903
rect 9706 2843 9718 2877
rect 9752 2843 9764 2877
rect 9706 2817 9764 2843
rect 9806 2877 9864 2903
rect 9806 2843 9818 2877
rect 9852 2843 9864 2877
rect 9806 2817 9864 2843
rect 9906 2877 9964 2903
rect 9906 2843 9918 2877
rect 9952 2843 9964 2877
rect 9906 2817 9964 2843
rect 10006 2877 10064 2903
rect 10006 2843 10018 2877
rect 10052 2843 10064 2877
rect 10006 2817 10064 2843
rect 10106 2877 10164 2903
rect 10106 2843 10118 2877
rect 10152 2843 10164 2877
rect 10106 2817 10164 2843
rect 10206 2877 10264 2903
rect 10206 2843 10218 2877
rect 10252 2843 10264 2877
rect 10206 2817 10264 2843
rect 10306 2877 10364 2903
rect 10306 2843 10318 2877
rect 10352 2843 10364 2877
rect 10306 2817 10364 2843
rect 10406 2877 10464 2903
rect 10406 2843 10418 2877
rect 10452 2843 10464 2877
rect 10406 2817 10464 2843
rect 10506 2877 10564 2903
rect 10506 2843 10512 2877
rect 10552 2843 10564 2877
rect 10506 2817 10564 2843
rect 10606 2877 10664 2903
rect 10606 2843 10618 2877
rect 10658 2843 10664 2877
rect 10606 2817 10664 2843
rect 10706 2877 10764 2903
rect 10706 2843 10718 2877
rect 10752 2843 10764 2877
rect 10706 2817 10764 2843
rect 10806 2877 10864 2903
rect 10806 2843 10818 2877
rect 10852 2843 10864 2877
rect 10806 2817 10864 2843
rect 10906 2877 10964 2903
rect 10906 2843 10918 2877
rect 10952 2843 10964 2877
rect 10906 2817 10964 2843
rect 11006 2877 11064 2903
rect 11006 2843 11018 2877
rect 11052 2843 11064 2877
rect 11006 2817 11064 2843
rect 11106 2877 11164 2903
rect 11106 2843 11118 2877
rect 11152 2843 11164 2877
rect 11106 2817 11164 2843
rect 11206 2877 11264 2903
rect 11206 2843 11218 2877
rect 11252 2843 11264 2877
rect 11206 2817 11264 2843
rect 11306 2877 11364 2903
rect 11306 2843 11312 2877
rect 11352 2843 11364 2877
rect 11306 2817 11364 2843
rect 11406 2877 11464 2903
rect 11406 2843 11418 2877
rect 11458 2843 11464 2877
rect 11406 2817 11464 2843
rect 11506 2877 11564 2903
rect 11506 2843 11518 2877
rect 11552 2843 11564 2877
rect 11506 2817 11564 2843
rect 11606 2877 11664 2903
rect 11606 2843 11618 2877
rect 11652 2843 11664 2877
rect 11606 2817 11664 2843
rect 11706 2877 11764 2903
rect 11706 2843 11718 2877
rect 11752 2843 11764 2877
rect 11706 2817 11764 2843
rect 11806 2877 11864 2903
rect 11806 2843 11812 2877
rect 11852 2843 11864 2877
rect 11806 2817 11864 2843
rect 11906 2877 11964 2903
rect 11906 2843 11918 2877
rect 11958 2843 11964 2877
rect 11906 2817 11964 2843
rect 12006 2877 12064 2903
rect 12006 2843 12018 2877
rect 12052 2843 12064 2877
rect 12006 2817 12064 2843
rect 12106 2877 12164 2903
rect 12106 2843 12118 2877
rect 12152 2843 12164 2877
rect 12106 2817 12164 2843
rect 12206 2877 12264 2903
rect 12206 2843 12218 2877
rect 12252 2843 12264 2877
rect 12206 2817 12264 2843
rect 12306 2877 12364 2903
rect 12306 2843 12318 2877
rect 12352 2843 12364 2877
rect 12306 2817 12364 2843
rect 12406 2877 12464 2903
rect 12406 2843 12418 2877
rect 12452 2843 12464 2877
rect 12406 2817 12464 2843
rect 12506 2877 12564 2903
rect 12506 2843 12518 2877
rect 12552 2843 12564 2877
rect 12506 2817 12564 2843
rect 12606 2877 12664 2903
rect 12606 2843 12618 2877
rect 12652 2843 12664 2877
rect 12606 2817 12664 2843
rect 12706 2877 12764 2903
rect 12706 2843 12718 2877
rect 12752 2843 12764 2877
rect 12706 2817 12764 2843
rect 12806 2877 12864 2903
rect 13018 2896 13262 2930
rect 12806 2843 12812 2877
rect 12852 2843 12864 2877
rect 12908 2858 12916 2892
rect 12958 2858 12974 2892
rect 13018 2877 13052 2896
rect 12806 2817 12864 2843
rect 13228 2877 13262 2896
rect 13018 2827 13052 2843
rect 13096 2828 13112 2862
rect 13154 2828 13162 2862
rect 13228 2827 13262 2843
rect 13328 2877 13562 2893
rect 13362 2843 13428 2877
rect 13462 2843 13528 2877
rect 13328 2827 13562 2843
rect 13628 2877 13662 2893
rect 13628 2827 13662 2843
rect 6 2737 64 2763
rect 6 2703 18 2737
rect 52 2703 64 2737
rect 6 2677 64 2703
rect 106 2737 164 2763
rect 106 2703 118 2737
rect 152 2703 164 2737
rect 106 2677 164 2703
rect 206 2737 264 2763
rect 206 2703 218 2737
rect 252 2703 264 2737
rect 206 2677 264 2703
rect 306 2737 364 2763
rect 306 2703 318 2737
rect 352 2703 364 2737
rect 306 2677 364 2703
rect 406 2737 464 2763
rect 406 2703 418 2737
rect 452 2703 464 2737
rect 406 2677 464 2703
rect 506 2737 564 2763
rect 506 2703 518 2737
rect 552 2703 564 2737
rect 506 2677 564 2703
rect 606 2737 664 2763
rect 606 2703 618 2737
rect 652 2703 664 2737
rect 606 2677 664 2703
rect 706 2737 764 2763
rect 706 2703 718 2737
rect 752 2703 764 2737
rect 706 2677 764 2703
rect 806 2737 864 2763
rect 806 2703 818 2737
rect 852 2703 864 2737
rect 806 2677 864 2703
rect 906 2737 964 2763
rect 906 2703 918 2737
rect 952 2703 964 2737
rect 906 2677 964 2703
rect 1006 2737 1064 2763
rect 1006 2703 1018 2737
rect 1052 2703 1064 2737
rect 1006 2677 1064 2703
rect 1106 2737 1164 2763
rect 1106 2703 1112 2737
rect 1152 2703 1164 2737
rect 1106 2677 1164 2703
rect 1206 2737 1264 2763
rect 1206 2703 1218 2737
rect 1258 2703 1264 2737
rect 1206 2677 1264 2703
rect 1306 2737 1364 2763
rect 1306 2703 1318 2737
rect 1352 2703 1364 2737
rect 1306 2677 1364 2703
rect 1406 2737 1464 2763
rect 1406 2703 1418 2737
rect 1452 2703 1464 2737
rect 1406 2677 1464 2703
rect 1506 2737 1564 2763
rect 1506 2703 1518 2737
rect 1552 2703 1564 2737
rect 1506 2677 1564 2703
rect 1606 2737 1664 2763
rect 1606 2703 1618 2737
rect 1652 2703 1664 2737
rect 1606 2677 1664 2703
rect 1706 2737 1764 2763
rect 1706 2703 1718 2737
rect 1752 2703 1764 2737
rect 1706 2677 1764 2703
rect 1806 2737 1864 2763
rect 1806 2703 1818 2737
rect 1852 2703 1864 2737
rect 1806 2677 1864 2703
rect 1906 2737 1964 2763
rect 1906 2703 1918 2737
rect 1952 2703 1964 2737
rect 1906 2677 1964 2703
rect 2006 2737 2064 2763
rect 2006 2703 2018 2737
rect 2052 2703 2064 2737
rect 2006 2677 2064 2703
rect 2106 2737 2164 2763
rect 2106 2703 2118 2737
rect 2152 2703 2164 2737
rect 2106 2677 2164 2703
rect 2206 2737 2264 2763
rect 2206 2703 2218 2737
rect 2252 2703 2264 2737
rect 2206 2677 2264 2703
rect 2306 2737 2364 2763
rect 2306 2703 2312 2737
rect 2352 2703 2364 2737
rect 2306 2677 2364 2703
rect 2406 2737 2464 2763
rect 2406 2703 2418 2737
rect 2458 2703 2464 2737
rect 2406 2677 2464 2703
rect 2506 2737 2564 2763
rect 2506 2703 2518 2737
rect 2552 2703 2564 2737
rect 2506 2677 2564 2703
rect 2606 2737 2664 2763
rect 2606 2703 2618 2737
rect 2652 2703 2664 2737
rect 2606 2677 2664 2703
rect 2706 2737 2764 2763
rect 2706 2703 2718 2737
rect 2752 2703 2764 2737
rect 2706 2677 2764 2703
rect 2806 2737 2864 2763
rect 2806 2703 2818 2737
rect 2852 2703 2864 2737
rect 2806 2677 2864 2703
rect 2906 2737 2964 2763
rect 2906 2703 2918 2737
rect 2952 2703 2964 2737
rect 2906 2677 2964 2703
rect 3006 2737 3064 2763
rect 3006 2703 3018 2737
rect 3052 2703 3064 2737
rect 3006 2677 3064 2703
rect 3106 2737 3164 2763
rect 3106 2703 3118 2737
rect 3152 2703 3164 2737
rect 3106 2677 3164 2703
rect 3206 2737 3264 2763
rect 3206 2703 3218 2737
rect 3252 2703 3264 2737
rect 3206 2677 3264 2703
rect 3306 2737 3364 2763
rect 3306 2703 3318 2737
rect 3352 2703 3364 2737
rect 3306 2677 3364 2703
rect 3406 2737 3464 2763
rect 3406 2703 3418 2737
rect 3452 2703 3464 2737
rect 3406 2677 3464 2703
rect 3506 2737 3564 2763
rect 3506 2703 3518 2737
rect 3552 2703 3564 2737
rect 3506 2677 3564 2703
rect 3606 2737 3664 2763
rect 3606 2703 3618 2737
rect 3652 2703 3664 2737
rect 3606 2677 3664 2703
rect 3706 2737 3764 2763
rect 3706 2703 3718 2737
rect 3752 2703 3764 2737
rect 3706 2677 3764 2703
rect 3806 2737 3864 2763
rect 3806 2703 3818 2737
rect 3852 2703 3864 2737
rect 3806 2677 3864 2703
rect 3906 2737 3964 2763
rect 3906 2703 3918 2737
rect 3952 2703 3964 2737
rect 3906 2677 3964 2703
rect 4006 2737 4064 2763
rect 4006 2703 4018 2737
rect 4052 2703 4064 2737
rect 4006 2677 4064 2703
rect 4106 2737 4164 2763
rect 4106 2703 4112 2737
rect 4152 2703 4164 2737
rect 4106 2677 4164 2703
rect 4206 2737 4264 2763
rect 4206 2703 4218 2737
rect 4258 2703 4264 2737
rect 4206 2677 4264 2703
rect 4306 2737 4364 2763
rect 4306 2703 4318 2737
rect 4352 2703 4364 2737
rect 4306 2677 4364 2703
rect 4406 2737 4464 2763
rect 4406 2703 4418 2737
rect 4452 2703 4464 2737
rect 4406 2677 4464 2703
rect 4506 2737 4564 2763
rect 4506 2703 4518 2737
rect 4552 2703 4564 2737
rect 4506 2677 4564 2703
rect 4606 2737 4664 2763
rect 4606 2703 4618 2737
rect 4652 2703 4664 2737
rect 4606 2677 4664 2703
rect 4706 2737 4764 2763
rect 4706 2703 4712 2737
rect 4752 2703 4764 2737
rect 4706 2677 4764 2703
rect 4806 2737 4864 2763
rect 4806 2703 4818 2737
rect 4858 2703 4864 2737
rect 4806 2677 4864 2703
rect 4906 2737 4964 2763
rect 4906 2703 4918 2737
rect 4952 2703 4964 2737
rect 4906 2677 4964 2703
rect 5006 2737 5064 2763
rect 5006 2703 5018 2737
rect 5052 2703 5064 2737
rect 5006 2677 5064 2703
rect 5106 2737 5164 2763
rect 5106 2703 5112 2737
rect 5152 2703 5164 2737
rect 5106 2677 5164 2703
rect 5206 2737 5264 2763
rect 5206 2703 5218 2737
rect 5258 2703 5264 2737
rect 5206 2677 5264 2703
rect 5306 2737 5364 2763
rect 5306 2703 5312 2737
rect 5352 2703 5364 2737
rect 5306 2677 5364 2703
rect 5406 2737 5464 2763
rect 5406 2703 5418 2737
rect 5458 2703 5464 2737
rect 5406 2677 5464 2703
rect 5506 2737 5564 2763
rect 5506 2703 5518 2737
rect 5552 2703 5564 2737
rect 5506 2677 5564 2703
rect 5606 2737 5664 2763
rect 5606 2703 5618 2737
rect 5652 2703 5664 2737
rect 5606 2677 5664 2703
rect 5706 2737 5764 2763
rect 5706 2703 5718 2737
rect 5752 2703 5764 2737
rect 5706 2677 5764 2703
rect 5806 2737 5864 2763
rect 5806 2703 5818 2737
rect 5852 2703 5864 2737
rect 5806 2677 5864 2703
rect 5906 2737 5964 2763
rect 5906 2703 5918 2737
rect 5952 2703 5964 2737
rect 5906 2677 5964 2703
rect 6006 2737 6064 2763
rect 6006 2703 6012 2737
rect 6052 2703 6064 2737
rect 6006 2677 6064 2703
rect 6106 2737 6164 2763
rect 6106 2703 6118 2737
rect 6158 2703 6164 2737
rect 6106 2677 6164 2703
rect 6206 2737 6264 2763
rect 6206 2703 6212 2737
rect 6252 2703 6264 2737
rect 6206 2677 6264 2703
rect 6306 2737 6364 2763
rect 6306 2703 6318 2737
rect 6358 2703 6364 2737
rect 6306 2677 6364 2703
rect 6406 2737 6464 2763
rect 6406 2703 6418 2737
rect 6452 2703 6464 2737
rect 6406 2677 6464 2703
rect 6506 2737 6564 2763
rect 6506 2703 6512 2737
rect 6552 2703 6564 2737
rect 6506 2677 6564 2703
rect 6606 2737 6664 2763
rect 6606 2703 6618 2737
rect 6658 2703 6664 2737
rect 6606 2677 6664 2703
rect 6706 2737 6764 2763
rect 6706 2703 6718 2737
rect 6752 2703 6764 2737
rect 6706 2677 6764 2703
rect 6806 2737 6864 2763
rect 6806 2703 6818 2737
rect 6852 2703 6864 2737
rect 6806 2677 6864 2703
rect 6906 2737 6964 2763
rect 6906 2703 6918 2737
rect 6952 2703 6964 2737
rect 6906 2677 6964 2703
rect 7006 2737 7064 2763
rect 7006 2703 7018 2737
rect 7052 2703 7064 2737
rect 7006 2677 7064 2703
rect 7106 2737 7164 2763
rect 7106 2703 7118 2737
rect 7152 2703 7164 2737
rect 7106 2677 7164 2703
rect 7206 2737 7264 2763
rect 7206 2703 7218 2737
rect 7252 2703 7264 2737
rect 7206 2677 7264 2703
rect 7306 2737 7364 2763
rect 7306 2703 7318 2737
rect 7352 2703 7364 2737
rect 7306 2677 7364 2703
rect 7406 2737 7464 2763
rect 7406 2703 7418 2737
rect 7452 2703 7464 2737
rect 7406 2677 7464 2703
rect 7506 2737 7564 2763
rect 7506 2703 7518 2737
rect 7552 2703 7564 2737
rect 7506 2677 7564 2703
rect 7606 2737 7664 2763
rect 7606 2703 7618 2737
rect 7652 2703 7664 2737
rect 7606 2677 7664 2703
rect 7706 2737 7764 2763
rect 7706 2703 7718 2737
rect 7752 2703 7764 2737
rect 7706 2677 7764 2703
rect 7806 2737 7864 2763
rect 7806 2703 7818 2737
rect 7852 2703 7864 2737
rect 7806 2677 7864 2703
rect 7906 2737 7964 2763
rect 7906 2703 7918 2737
rect 7952 2703 7964 2737
rect 7906 2677 7964 2703
rect 8006 2737 8064 2763
rect 8006 2703 8018 2737
rect 8052 2703 8064 2737
rect 8006 2677 8064 2703
rect 8106 2737 8164 2763
rect 8106 2703 8118 2737
rect 8152 2703 8164 2737
rect 8106 2677 8164 2703
rect 8206 2737 8264 2763
rect 8206 2703 8212 2737
rect 8252 2703 8264 2737
rect 8206 2677 8264 2703
rect 8306 2737 8364 2763
rect 8306 2703 8318 2737
rect 8358 2703 8364 2737
rect 8306 2677 8364 2703
rect 8406 2737 8464 2763
rect 8406 2703 8418 2737
rect 8452 2703 8464 2737
rect 8406 2677 8464 2703
rect 8506 2737 8564 2763
rect 8506 2703 8518 2737
rect 8552 2703 8564 2737
rect 8506 2677 8564 2703
rect 8606 2737 8664 2763
rect 8606 2703 8618 2737
rect 8652 2703 8664 2737
rect 8606 2677 8664 2703
rect 8706 2737 8764 2763
rect 8706 2703 8712 2737
rect 8752 2703 8764 2737
rect 8706 2677 8764 2703
rect 8806 2737 8864 2763
rect 8806 2703 8818 2737
rect 8858 2703 8864 2737
rect 8806 2677 8864 2703
rect 8906 2737 8964 2763
rect 8906 2703 8912 2737
rect 8952 2703 8964 2737
rect 8906 2677 8964 2703
rect 9006 2737 9064 2763
rect 9006 2703 9018 2737
rect 9058 2703 9064 2737
rect 9006 2677 9064 2703
rect 9106 2737 9164 2763
rect 9106 2703 9112 2737
rect 9152 2703 9164 2737
rect 9106 2677 9164 2703
rect 9206 2737 9264 2763
rect 9206 2703 9218 2737
rect 9258 2703 9264 2737
rect 9206 2677 9264 2703
rect 9306 2737 9364 2763
rect 9306 2703 9312 2737
rect 9352 2703 9364 2737
rect 9306 2677 9364 2703
rect 9406 2737 9464 2763
rect 9406 2703 9418 2737
rect 9458 2703 9464 2737
rect 9406 2677 9464 2703
rect 9506 2737 9564 2763
rect 9506 2703 9512 2737
rect 9552 2703 9564 2737
rect 9506 2677 9564 2703
rect 9606 2737 9664 2763
rect 9606 2703 9618 2737
rect 9658 2703 9664 2737
rect 9606 2677 9664 2703
rect 9706 2737 9764 2763
rect 9706 2703 9718 2737
rect 9752 2703 9764 2737
rect 9706 2677 9764 2703
rect 9806 2737 9864 2763
rect 9806 2703 9818 2737
rect 9852 2703 9864 2737
rect 9806 2677 9864 2703
rect 9906 2737 9964 2763
rect 9906 2703 9912 2737
rect 9952 2703 9964 2737
rect 9906 2677 9964 2703
rect 10006 2737 10064 2763
rect 10006 2703 10018 2737
rect 10058 2703 10064 2737
rect 10006 2677 10064 2703
rect 10106 2737 10164 2763
rect 10106 2703 10118 2737
rect 10152 2703 10164 2737
rect 10106 2677 10164 2703
rect 10206 2737 10264 2763
rect 10206 2703 10218 2737
rect 10252 2703 10264 2737
rect 10206 2677 10264 2703
rect 10306 2737 10364 2763
rect 10306 2703 10318 2737
rect 10352 2703 10364 2737
rect 10306 2677 10364 2703
rect 10406 2737 10464 2763
rect 10406 2703 10412 2737
rect 10452 2703 10464 2737
rect 10406 2677 10464 2703
rect 10506 2737 10564 2763
rect 10506 2703 10518 2737
rect 10558 2703 10564 2737
rect 10506 2677 10564 2703
rect 10606 2737 10664 2763
rect 10606 2703 10612 2737
rect 10652 2703 10664 2737
rect 10606 2677 10664 2703
rect 10706 2737 10764 2763
rect 10706 2703 10718 2737
rect 10758 2703 10764 2737
rect 10706 2677 10764 2703
rect 10806 2737 10864 2763
rect 10806 2703 10818 2737
rect 10852 2703 10864 2737
rect 10806 2677 10864 2703
rect 10906 2737 10964 2763
rect 10906 2703 10918 2737
rect 10952 2703 10964 2737
rect 10906 2677 10964 2703
rect 11006 2737 11064 2763
rect 11006 2703 11018 2737
rect 11052 2703 11064 2737
rect 11006 2677 11064 2703
rect 11106 2737 11164 2763
rect 11106 2703 11118 2737
rect 11152 2703 11164 2737
rect 11106 2677 11164 2703
rect 11206 2737 11264 2763
rect 11206 2703 11218 2737
rect 11252 2703 11264 2737
rect 11206 2677 11264 2703
rect 11306 2737 11364 2763
rect 11306 2703 11318 2737
rect 11352 2703 11364 2737
rect 11306 2677 11364 2703
rect 11406 2737 11464 2763
rect 11406 2703 11418 2737
rect 11452 2703 11464 2737
rect 11406 2677 11464 2703
rect 11506 2737 11564 2763
rect 11506 2703 11518 2737
rect 11552 2703 11564 2737
rect 11506 2677 11564 2703
rect 11606 2737 11664 2763
rect 11606 2703 11612 2737
rect 11652 2703 11664 2737
rect 11606 2677 11664 2703
rect 11706 2737 11764 2763
rect 11706 2703 11718 2737
rect 11758 2703 11764 2737
rect 11706 2677 11764 2703
rect 11806 2737 11864 2763
rect 11806 2703 11818 2737
rect 11852 2703 11864 2737
rect 11806 2677 11864 2703
rect 11906 2737 11964 2763
rect 11906 2703 11918 2737
rect 11952 2703 11964 2737
rect 11906 2677 11964 2703
rect 12006 2737 12064 2763
rect 12006 2703 12018 2737
rect 12052 2703 12064 2737
rect 12006 2677 12064 2703
rect 12106 2737 12164 2763
rect 12106 2703 12118 2737
rect 12152 2703 12164 2737
rect 12106 2677 12164 2703
rect 12206 2737 12264 2763
rect 12206 2703 12218 2737
rect 12252 2703 12264 2737
rect 12206 2677 12264 2703
rect 12306 2737 12364 2763
rect 12306 2703 12318 2737
rect 12352 2703 12364 2737
rect 12306 2677 12364 2703
rect 12406 2737 12464 2763
rect 12406 2703 12418 2737
rect 12452 2703 12464 2737
rect 12406 2677 12464 2703
rect 12506 2737 12564 2763
rect 12506 2703 12518 2737
rect 12552 2703 12564 2737
rect 12506 2677 12564 2703
rect 12606 2737 12664 2763
rect 12606 2703 12618 2737
rect 12652 2703 12664 2737
rect 12606 2677 12664 2703
rect 12706 2737 12764 2763
rect 12706 2703 12718 2737
rect 12752 2703 12764 2737
rect 12706 2677 12764 2703
rect 12806 2737 12864 2763
rect 13018 2756 13262 2790
rect 12806 2703 12818 2737
rect 12852 2703 12864 2737
rect 12908 2718 12916 2752
rect 12958 2718 12974 2752
rect 13018 2737 13052 2756
rect 12806 2677 12864 2703
rect 13228 2753 13262 2756
rect 13228 2737 13362 2753
rect 13018 2687 13052 2703
rect 13096 2688 13112 2722
rect 13154 2688 13162 2722
rect 13262 2703 13328 2737
rect 13228 2687 13362 2703
rect 13428 2737 13462 2753
rect 13428 2687 13462 2703
rect 13528 2737 13662 2753
rect 13562 2703 13628 2737
rect 13528 2687 13662 2703
rect 6 2597 64 2623
rect 6 2563 18 2597
rect 52 2563 64 2597
rect 6 2537 64 2563
rect 106 2597 164 2623
rect 106 2563 118 2597
rect 152 2563 164 2597
rect 106 2537 164 2563
rect 206 2597 264 2623
rect 206 2563 218 2597
rect 252 2563 264 2597
rect 206 2537 264 2563
rect 306 2597 364 2623
rect 306 2563 318 2597
rect 352 2563 364 2597
rect 306 2537 364 2563
rect 406 2597 464 2623
rect 406 2563 418 2597
rect 452 2563 464 2597
rect 406 2537 464 2563
rect 506 2597 564 2623
rect 506 2563 518 2597
rect 552 2563 564 2597
rect 506 2537 564 2563
rect 606 2597 664 2623
rect 606 2563 618 2597
rect 652 2563 664 2597
rect 606 2537 664 2563
rect 706 2597 764 2623
rect 706 2563 718 2597
rect 752 2563 764 2597
rect 706 2537 764 2563
rect 806 2597 864 2623
rect 806 2563 818 2597
rect 852 2563 864 2597
rect 806 2537 864 2563
rect 906 2597 964 2623
rect 906 2563 918 2597
rect 952 2563 964 2597
rect 906 2537 964 2563
rect 1006 2597 1064 2623
rect 1006 2563 1018 2597
rect 1052 2563 1064 2597
rect 1006 2537 1064 2563
rect 1106 2597 1164 2623
rect 1106 2563 1118 2597
rect 1152 2563 1164 2597
rect 1106 2537 1164 2563
rect 1206 2597 1264 2623
rect 1206 2563 1218 2597
rect 1252 2563 1264 2597
rect 1206 2537 1264 2563
rect 1306 2597 1364 2623
rect 1306 2563 1318 2597
rect 1352 2563 1364 2597
rect 1306 2537 1364 2563
rect 1406 2597 1464 2623
rect 1406 2563 1418 2597
rect 1452 2563 1464 2597
rect 1406 2537 1464 2563
rect 1506 2597 1564 2623
rect 1506 2563 1518 2597
rect 1552 2563 1564 2597
rect 1506 2537 1564 2563
rect 1606 2597 1664 2623
rect 1606 2563 1618 2597
rect 1652 2563 1664 2597
rect 1606 2537 1664 2563
rect 1706 2597 1764 2623
rect 1706 2563 1718 2597
rect 1752 2563 1764 2597
rect 1706 2537 1764 2563
rect 1806 2597 1864 2623
rect 1806 2563 1818 2597
rect 1852 2563 1864 2597
rect 1806 2537 1864 2563
rect 1906 2597 1964 2623
rect 1906 2563 1918 2597
rect 1952 2563 1964 2597
rect 1906 2537 1964 2563
rect 2006 2597 2064 2623
rect 2006 2563 2018 2597
rect 2052 2563 2064 2597
rect 2006 2537 2064 2563
rect 2106 2597 2164 2623
rect 2106 2563 2118 2597
rect 2152 2563 2164 2597
rect 2106 2537 2164 2563
rect 2206 2597 2264 2623
rect 2206 2563 2218 2597
rect 2252 2563 2264 2597
rect 2206 2537 2264 2563
rect 2306 2597 2364 2623
rect 2306 2563 2318 2597
rect 2352 2563 2364 2597
rect 2306 2537 2364 2563
rect 2406 2597 2464 2623
rect 2406 2563 2418 2597
rect 2452 2563 2464 2597
rect 2406 2537 2464 2563
rect 2506 2597 2564 2623
rect 2506 2563 2512 2597
rect 2552 2563 2564 2597
rect 2506 2537 2564 2563
rect 2606 2597 2664 2623
rect 2606 2563 2618 2597
rect 2658 2563 2664 2597
rect 2606 2537 2664 2563
rect 2706 2597 2764 2623
rect 2706 2563 2718 2597
rect 2752 2563 2764 2597
rect 2706 2537 2764 2563
rect 2806 2597 2864 2623
rect 2806 2563 2818 2597
rect 2852 2563 2864 2597
rect 2806 2537 2864 2563
rect 2906 2597 2964 2623
rect 2906 2563 2918 2597
rect 2952 2563 2964 2597
rect 2906 2537 2964 2563
rect 3006 2597 3064 2623
rect 3006 2563 3018 2597
rect 3052 2563 3064 2597
rect 3006 2537 3064 2563
rect 3106 2597 3164 2623
rect 3106 2563 3118 2597
rect 3152 2563 3164 2597
rect 3106 2537 3164 2563
rect 3206 2597 3264 2623
rect 3206 2563 3218 2597
rect 3252 2563 3264 2597
rect 3206 2537 3264 2563
rect 3306 2597 3364 2623
rect 3306 2563 3312 2597
rect 3352 2563 3364 2597
rect 3306 2537 3364 2563
rect 3406 2597 3464 2623
rect 3406 2563 3418 2597
rect 3458 2563 3464 2597
rect 3406 2537 3464 2563
rect 3506 2597 3564 2623
rect 3506 2563 3518 2597
rect 3552 2563 3564 2597
rect 3506 2537 3564 2563
rect 3606 2597 3664 2623
rect 3606 2563 3618 2597
rect 3652 2563 3664 2597
rect 3606 2537 3664 2563
rect 3706 2597 3764 2623
rect 3706 2563 3718 2597
rect 3752 2563 3764 2597
rect 3706 2537 3764 2563
rect 3806 2597 3864 2623
rect 3806 2563 3818 2597
rect 3852 2563 3864 2597
rect 3806 2537 3864 2563
rect 3906 2597 3964 2623
rect 3906 2563 3912 2597
rect 3952 2563 3964 2597
rect 3906 2537 3964 2563
rect 4006 2597 4064 2623
rect 4006 2563 4018 2597
rect 4058 2563 4064 2597
rect 4006 2537 4064 2563
rect 4106 2597 4164 2623
rect 4106 2563 4112 2597
rect 4152 2563 4164 2597
rect 4106 2537 4164 2563
rect 4206 2597 4264 2623
rect 4206 2563 4218 2597
rect 4258 2563 4264 2597
rect 4206 2537 4264 2563
rect 4306 2597 4364 2623
rect 4306 2563 4312 2597
rect 4352 2563 4364 2597
rect 4306 2537 4364 2563
rect 4406 2597 4464 2623
rect 4406 2563 4418 2597
rect 4458 2563 4464 2597
rect 4406 2537 4464 2563
rect 4506 2597 4564 2623
rect 4506 2563 4518 2597
rect 4552 2563 4564 2597
rect 4506 2537 4564 2563
rect 4606 2597 4664 2623
rect 4606 2563 4618 2597
rect 4652 2563 4664 2597
rect 4606 2537 4664 2563
rect 4706 2597 4764 2623
rect 4706 2563 4712 2597
rect 4752 2563 4764 2597
rect 4706 2537 4764 2563
rect 4806 2597 4864 2623
rect 4806 2563 4818 2597
rect 4858 2563 4864 2597
rect 4806 2537 4864 2563
rect 4906 2597 4964 2623
rect 4906 2563 4918 2597
rect 4952 2563 4964 2597
rect 4906 2537 4964 2563
rect 5006 2597 5064 2623
rect 5006 2563 5018 2597
rect 5052 2563 5064 2597
rect 5006 2537 5064 2563
rect 5106 2597 5164 2623
rect 5106 2563 5118 2597
rect 5152 2563 5164 2597
rect 5106 2537 5164 2563
rect 5206 2597 5264 2623
rect 5206 2563 5218 2597
rect 5252 2563 5264 2597
rect 5206 2537 5264 2563
rect 5306 2597 5364 2623
rect 5306 2563 5318 2597
rect 5352 2563 5364 2597
rect 5306 2537 5364 2563
rect 5406 2597 5464 2623
rect 5406 2563 5418 2597
rect 5452 2563 5464 2597
rect 5406 2537 5464 2563
rect 5506 2597 5564 2623
rect 5506 2563 5518 2597
rect 5552 2563 5564 2597
rect 5506 2537 5564 2563
rect 5606 2597 5664 2623
rect 5606 2563 5618 2597
rect 5652 2563 5664 2597
rect 5606 2537 5664 2563
rect 5706 2597 5764 2623
rect 5706 2563 5718 2597
rect 5752 2563 5764 2597
rect 5706 2537 5764 2563
rect 5806 2597 5864 2623
rect 5806 2563 5818 2597
rect 5852 2563 5864 2597
rect 5806 2537 5864 2563
rect 5906 2597 5964 2623
rect 5906 2563 5918 2597
rect 5952 2563 5964 2597
rect 5906 2537 5964 2563
rect 6006 2597 6064 2623
rect 6006 2563 6018 2597
rect 6052 2563 6064 2597
rect 6006 2537 6064 2563
rect 6106 2597 6164 2623
rect 6106 2563 6118 2597
rect 6152 2563 6164 2597
rect 6106 2537 6164 2563
rect 6206 2597 6264 2623
rect 6206 2563 6212 2597
rect 6252 2563 6264 2597
rect 6206 2537 6264 2563
rect 6306 2597 6364 2623
rect 6306 2563 6318 2597
rect 6358 2563 6364 2597
rect 6306 2537 6364 2563
rect 6406 2597 6464 2623
rect 6406 2563 6418 2597
rect 6452 2563 6464 2597
rect 6406 2537 6464 2563
rect 6506 2597 6564 2623
rect 6506 2563 6518 2597
rect 6552 2563 6564 2597
rect 6506 2537 6564 2563
rect 6606 2597 6664 2623
rect 6606 2563 6618 2597
rect 6652 2563 6664 2597
rect 6606 2537 6664 2563
rect 6706 2597 6764 2623
rect 6706 2563 6712 2597
rect 6752 2563 6764 2597
rect 6706 2537 6764 2563
rect 6806 2597 6864 2623
rect 6806 2563 6818 2597
rect 6858 2563 6864 2597
rect 6806 2537 6864 2563
rect 6906 2597 6964 2623
rect 6906 2563 6918 2597
rect 6952 2563 6964 2597
rect 6906 2537 6964 2563
rect 7006 2597 7064 2623
rect 7006 2563 7018 2597
rect 7052 2563 7064 2597
rect 7006 2537 7064 2563
rect 7106 2597 7164 2623
rect 7106 2563 7118 2597
rect 7152 2563 7164 2597
rect 7106 2537 7164 2563
rect 7206 2597 7264 2623
rect 7206 2563 7218 2597
rect 7252 2563 7264 2597
rect 7206 2537 7264 2563
rect 7306 2597 7364 2623
rect 7306 2563 7318 2597
rect 7352 2563 7364 2597
rect 7306 2537 7364 2563
rect 7406 2597 7464 2623
rect 7406 2563 7418 2597
rect 7452 2563 7464 2597
rect 7406 2537 7464 2563
rect 7506 2597 7564 2623
rect 7506 2563 7518 2597
rect 7552 2563 7564 2597
rect 7506 2537 7564 2563
rect 7606 2597 7664 2623
rect 7606 2563 7618 2597
rect 7652 2563 7664 2597
rect 7606 2537 7664 2563
rect 7706 2597 7764 2623
rect 7706 2563 7718 2597
rect 7752 2563 7764 2597
rect 7706 2537 7764 2563
rect 7806 2597 7864 2623
rect 7806 2563 7818 2597
rect 7852 2563 7864 2597
rect 7806 2537 7864 2563
rect 7906 2597 7964 2623
rect 7906 2563 7918 2597
rect 7952 2563 7964 2597
rect 7906 2537 7964 2563
rect 8006 2597 8064 2623
rect 8006 2563 8018 2597
rect 8052 2563 8064 2597
rect 8006 2537 8064 2563
rect 8106 2597 8164 2623
rect 8106 2563 8118 2597
rect 8152 2563 8164 2597
rect 8106 2537 8164 2563
rect 8206 2597 8264 2623
rect 8206 2563 8212 2597
rect 8252 2563 8264 2597
rect 8206 2537 8264 2563
rect 8306 2597 8364 2623
rect 8306 2563 8318 2597
rect 8358 2563 8364 2597
rect 8306 2537 8364 2563
rect 8406 2597 8464 2623
rect 8406 2563 8412 2597
rect 8452 2563 8464 2597
rect 8406 2537 8464 2563
rect 8506 2597 8564 2623
rect 8506 2563 8518 2597
rect 8558 2563 8564 2597
rect 8506 2537 8564 2563
rect 8606 2597 8664 2623
rect 8606 2563 8618 2597
rect 8652 2563 8664 2597
rect 8606 2537 8664 2563
rect 8706 2597 8764 2623
rect 8706 2563 8712 2597
rect 8752 2563 8764 2597
rect 8706 2537 8764 2563
rect 8806 2597 8864 2623
rect 8806 2563 8818 2597
rect 8858 2563 8864 2597
rect 8806 2537 8864 2563
rect 8906 2597 8964 2623
rect 8906 2563 8918 2597
rect 8952 2563 8964 2597
rect 8906 2537 8964 2563
rect 9006 2597 9064 2623
rect 9006 2563 9012 2597
rect 9052 2563 9064 2597
rect 9006 2537 9064 2563
rect 9106 2597 9164 2623
rect 9106 2563 9118 2597
rect 9158 2563 9164 2597
rect 9106 2537 9164 2563
rect 9206 2597 9264 2623
rect 9206 2563 9212 2597
rect 9252 2563 9264 2597
rect 9206 2537 9264 2563
rect 9306 2597 9364 2623
rect 9306 2563 9318 2597
rect 9358 2563 9364 2597
rect 9306 2537 9364 2563
rect 9406 2597 9464 2623
rect 9406 2563 9418 2597
rect 9452 2563 9464 2597
rect 9406 2537 9464 2563
rect 9506 2597 9564 2623
rect 9506 2563 9512 2597
rect 9552 2563 9564 2597
rect 9506 2537 9564 2563
rect 9606 2597 9664 2623
rect 9606 2563 9618 2597
rect 9658 2563 9664 2597
rect 9606 2537 9664 2563
rect 9706 2597 9764 2623
rect 9706 2563 9718 2597
rect 9752 2563 9764 2597
rect 9706 2537 9764 2563
rect 9806 2597 9864 2623
rect 9806 2563 9818 2597
rect 9852 2563 9864 2597
rect 9806 2537 9864 2563
rect 9906 2597 9964 2623
rect 9906 2563 9912 2597
rect 9952 2563 9964 2597
rect 9906 2537 9964 2563
rect 10006 2597 10064 2623
rect 10006 2563 10018 2597
rect 10058 2563 10064 2597
rect 10006 2537 10064 2563
rect 10106 2597 10164 2623
rect 10106 2563 10118 2597
rect 10152 2563 10164 2597
rect 10106 2537 10164 2563
rect 10206 2597 10264 2623
rect 10206 2563 10218 2597
rect 10252 2563 10264 2597
rect 10206 2537 10264 2563
rect 10306 2597 10364 2623
rect 10306 2563 10318 2597
rect 10352 2563 10364 2597
rect 10306 2537 10364 2563
rect 10406 2597 10464 2623
rect 10406 2563 10418 2597
rect 10452 2563 10464 2597
rect 10406 2537 10464 2563
rect 10506 2597 10564 2623
rect 10506 2563 10518 2597
rect 10552 2563 10564 2597
rect 10506 2537 10564 2563
rect 10606 2597 10664 2623
rect 10606 2563 10618 2597
rect 10652 2563 10664 2597
rect 10606 2537 10664 2563
rect 10706 2597 10764 2623
rect 10706 2563 10718 2597
rect 10752 2563 10764 2597
rect 10706 2537 10764 2563
rect 10806 2597 10864 2623
rect 10806 2563 10818 2597
rect 10852 2563 10864 2597
rect 10806 2537 10864 2563
rect 10906 2597 10964 2623
rect 10906 2563 10912 2597
rect 10952 2563 10964 2597
rect 10906 2537 10964 2563
rect 11006 2597 11064 2623
rect 11006 2563 11018 2597
rect 11058 2563 11064 2597
rect 11006 2537 11064 2563
rect 11106 2597 11164 2623
rect 11106 2563 11112 2597
rect 11152 2563 11164 2597
rect 11106 2537 11164 2563
rect 11206 2597 11264 2623
rect 11206 2563 11218 2597
rect 11258 2563 11264 2597
rect 11206 2537 11264 2563
rect 11306 2597 11364 2623
rect 11306 2563 11312 2597
rect 11352 2563 11364 2597
rect 11306 2537 11364 2563
rect 11406 2597 11464 2623
rect 11406 2563 11418 2597
rect 11458 2563 11464 2597
rect 11406 2537 11464 2563
rect 11506 2597 11564 2623
rect 11506 2563 11518 2597
rect 11552 2563 11564 2597
rect 11506 2537 11564 2563
rect 11606 2597 11664 2623
rect 11606 2563 11612 2597
rect 11652 2563 11664 2597
rect 11606 2537 11664 2563
rect 11706 2597 11764 2623
rect 11706 2563 11718 2597
rect 11758 2563 11764 2597
rect 11706 2537 11764 2563
rect 11806 2597 11864 2623
rect 11806 2563 11818 2597
rect 11852 2563 11864 2597
rect 11806 2537 11864 2563
rect 11906 2597 11964 2623
rect 11906 2563 11918 2597
rect 11952 2563 11964 2597
rect 11906 2537 11964 2563
rect 12006 2597 12064 2623
rect 12006 2563 12018 2597
rect 12052 2563 12064 2597
rect 12006 2537 12064 2563
rect 12106 2597 12164 2623
rect 12106 2563 12118 2597
rect 12152 2563 12164 2597
rect 12106 2537 12164 2563
rect 12206 2597 12264 2623
rect 12206 2563 12218 2597
rect 12252 2563 12264 2597
rect 12206 2537 12264 2563
rect 12306 2597 12364 2623
rect 12306 2563 12318 2597
rect 12352 2563 12364 2597
rect 12306 2537 12364 2563
rect 12406 2597 12464 2623
rect 12406 2563 12418 2597
rect 12452 2563 12464 2597
rect 12406 2537 12464 2563
rect 12506 2597 12564 2623
rect 12506 2563 12518 2597
rect 12552 2563 12564 2597
rect 12506 2537 12564 2563
rect 12606 2597 12664 2623
rect 12606 2563 12618 2597
rect 12652 2563 12664 2597
rect 12606 2537 12664 2563
rect 12706 2597 12764 2623
rect 12706 2563 12718 2597
rect 12752 2563 12764 2597
rect 12706 2537 12764 2563
rect 12806 2597 12864 2623
rect 13018 2616 13262 2650
rect 12806 2563 12818 2597
rect 12852 2563 12864 2597
rect 12908 2578 12916 2612
rect 12958 2578 12974 2612
rect 13018 2597 13052 2616
rect 12806 2537 12864 2563
rect 13228 2597 13262 2616
rect 13018 2547 13052 2563
rect 13096 2548 13112 2582
rect 13154 2548 13162 2582
rect 13228 2547 13262 2563
rect 13328 2597 13462 2613
rect 13362 2563 13428 2597
rect 13328 2547 13462 2563
rect 13528 2597 13662 2613
rect 13562 2563 13628 2597
rect 13528 2547 13662 2563
rect 8 2440 18 2474
rect 52 2440 118 2474
rect 152 2440 168 2474
rect 208 2456 218 2490
rect 252 2456 318 2490
rect 352 2456 368 2490
rect 408 2440 418 2474
rect 452 2440 518 2474
rect 552 2440 568 2474
rect 608 2456 618 2490
rect 652 2456 718 2490
rect 752 2456 768 2490
rect 808 2440 818 2474
rect 852 2440 918 2474
rect 952 2440 968 2474
rect 1008 2456 1018 2490
rect 1052 2456 1118 2490
rect 1152 2456 1168 2490
rect 1208 2440 1218 2474
rect 1252 2440 1318 2474
rect 1352 2440 1368 2474
rect 1408 2456 1418 2490
rect 1452 2456 1518 2490
rect 1552 2456 1568 2490
rect 1608 2440 1618 2474
rect 1652 2440 1718 2474
rect 1752 2440 1768 2474
rect 1808 2456 1818 2490
rect 1852 2456 1918 2490
rect 1952 2456 1968 2490
rect 2008 2440 2018 2474
rect 2052 2440 2118 2474
rect 2152 2440 2168 2474
rect 2208 2456 2218 2490
rect 2252 2456 2318 2490
rect 2352 2456 2368 2490
rect 2408 2440 2418 2474
rect 2452 2440 2518 2474
rect 2552 2440 2568 2474
rect 2608 2456 2618 2490
rect 2652 2456 2718 2490
rect 2752 2456 2768 2490
rect 2808 2440 2818 2474
rect 2852 2440 2918 2474
rect 2952 2440 2968 2474
rect 3008 2456 3018 2490
rect 3052 2456 3118 2490
rect 3152 2456 3168 2490
rect 3208 2440 3218 2474
rect 3252 2440 3318 2474
rect 3352 2440 3368 2474
rect 3408 2456 3418 2490
rect 3452 2456 3518 2490
rect 3552 2456 3568 2490
rect 3608 2440 3618 2474
rect 3652 2440 3718 2474
rect 3752 2440 3768 2474
rect 3808 2456 3818 2490
rect 3852 2456 3918 2490
rect 3952 2456 3968 2490
rect 4008 2440 4018 2474
rect 4052 2440 4118 2474
rect 4152 2440 4168 2474
rect 4208 2456 4218 2490
rect 4252 2456 4318 2490
rect 4352 2456 4368 2490
rect 4408 2440 4418 2474
rect 4452 2440 4518 2474
rect 4552 2440 4568 2474
rect 4608 2456 4618 2490
rect 4652 2456 4718 2490
rect 4752 2456 4768 2490
rect 4808 2440 4818 2474
rect 4852 2440 4918 2474
rect 4952 2440 4968 2474
rect 5008 2456 5018 2490
rect 5052 2456 5118 2490
rect 5152 2456 5168 2490
rect 5208 2440 5218 2474
rect 5252 2440 5318 2474
rect 5352 2440 5368 2474
rect 5408 2456 5418 2490
rect 5452 2456 5518 2490
rect 5552 2456 5568 2490
rect 5608 2440 5618 2474
rect 5652 2440 5718 2474
rect 5752 2440 5768 2474
rect 5808 2456 5818 2490
rect 5852 2456 5918 2490
rect 5952 2456 5968 2490
rect 6008 2440 6018 2474
rect 6052 2440 6118 2474
rect 6152 2440 6168 2474
rect 6208 2456 6218 2490
rect 6252 2456 6318 2490
rect 6352 2456 6368 2490
rect 6408 2440 6418 2474
rect 6452 2440 6518 2474
rect 6552 2440 6568 2474
rect 6608 2456 6618 2490
rect 6652 2456 6718 2490
rect 6752 2456 6768 2490
rect 6808 2440 6818 2474
rect 6852 2440 6918 2474
rect 6952 2440 6968 2474
rect 7008 2456 7018 2490
rect 7052 2456 7118 2490
rect 7152 2456 7168 2490
rect 7208 2440 7218 2474
rect 7252 2440 7318 2474
rect 7352 2440 7368 2474
rect 7408 2456 7418 2490
rect 7452 2456 7518 2490
rect 7552 2456 7568 2490
rect 7608 2440 7618 2474
rect 7652 2440 7718 2474
rect 7752 2440 7768 2474
rect 7808 2456 7818 2490
rect 7852 2456 7918 2490
rect 7952 2456 7968 2490
rect 8008 2440 8018 2474
rect 8052 2440 8118 2474
rect 8152 2440 8168 2474
rect 8208 2456 8218 2490
rect 8252 2456 8318 2490
rect 8352 2456 8368 2490
rect 8408 2440 8418 2474
rect 8452 2440 8518 2474
rect 8552 2440 8568 2474
rect 8608 2456 8618 2490
rect 8652 2456 8718 2490
rect 8752 2456 8768 2490
rect 8808 2440 8818 2474
rect 8852 2440 8918 2474
rect 8952 2440 8968 2474
rect 9008 2456 9018 2490
rect 9052 2456 9118 2490
rect 9152 2456 9168 2490
rect 9208 2440 9218 2474
rect 9252 2440 9318 2474
rect 9352 2440 9368 2474
rect 9408 2456 9418 2490
rect 9452 2456 9518 2490
rect 9552 2456 9568 2490
rect 9608 2440 9618 2474
rect 9652 2440 9718 2474
rect 9752 2440 9768 2474
rect 9808 2456 9818 2490
rect 9852 2456 9918 2490
rect 9952 2456 9968 2490
rect 10008 2440 10018 2474
rect 10052 2440 10118 2474
rect 10152 2440 10168 2474
rect 10208 2456 10218 2490
rect 10252 2456 10318 2490
rect 10352 2456 10368 2490
rect 10408 2440 10418 2474
rect 10452 2440 10518 2474
rect 10552 2440 10568 2474
rect 10608 2456 10618 2490
rect 10652 2456 10718 2490
rect 10752 2456 10768 2490
rect 10808 2440 10818 2474
rect 10852 2440 10918 2474
rect 10952 2440 10968 2474
rect 11008 2456 11018 2490
rect 11052 2456 11118 2490
rect 11152 2456 11168 2490
rect 11208 2440 11218 2474
rect 11252 2440 11318 2474
rect 11352 2440 11368 2474
rect 11408 2456 11418 2490
rect 11452 2456 11518 2490
rect 11552 2456 11568 2490
rect 11608 2440 11618 2474
rect 11652 2440 11718 2474
rect 11752 2440 11768 2474
rect 11808 2456 11818 2490
rect 11852 2456 11918 2490
rect 11952 2456 11968 2490
rect 12008 2440 12018 2474
rect 12052 2440 12118 2474
rect 12152 2440 12168 2474
rect 12208 2456 12218 2490
rect 12252 2456 12318 2490
rect 12352 2456 12368 2490
rect 12408 2440 12418 2474
rect 12452 2440 12518 2474
rect 12552 2440 12568 2474
rect 12608 2456 12618 2490
rect 12652 2456 12718 2490
rect 12752 2456 12768 2490
rect 12916 2471 12968 2488
rect 12950 2454 12968 2471
rect 13002 2454 13018 2488
rect 13052 2454 13068 2488
rect 13102 2459 13120 2488
rect 13102 2454 13154 2459
rect 13262 2454 13278 2488
rect 13312 2454 13328 2488
rect 13362 2454 13378 2488
rect 13412 2454 13428 2488
rect 13462 2454 13478 2488
rect 13512 2454 13528 2488
rect 13562 2454 13578 2488
rect 13612 2454 13628 2488
rect 6 2367 64 2393
rect 6 2333 18 2367
rect 58 2333 64 2367
rect 6 2307 64 2333
rect 106 2367 164 2393
rect 106 2333 112 2367
rect 152 2333 164 2367
rect 106 2307 164 2333
rect 206 2367 264 2393
rect 206 2333 218 2367
rect 258 2333 264 2367
rect 206 2307 264 2333
rect 306 2367 364 2393
rect 306 2333 318 2367
rect 352 2333 364 2367
rect 306 2307 364 2333
rect 406 2367 464 2393
rect 406 2333 412 2367
rect 452 2333 464 2367
rect 406 2307 464 2333
rect 506 2367 564 2393
rect 506 2333 518 2367
rect 558 2333 564 2367
rect 506 2307 564 2333
rect 606 2367 664 2393
rect 606 2333 612 2367
rect 652 2333 664 2367
rect 606 2307 664 2333
rect 706 2367 764 2393
rect 706 2333 718 2367
rect 758 2333 764 2367
rect 706 2307 764 2333
rect 806 2367 864 2393
rect 806 2333 818 2367
rect 852 2333 864 2367
rect 806 2307 864 2333
rect 906 2367 964 2393
rect 906 2333 918 2367
rect 952 2333 964 2367
rect 906 2307 964 2333
rect 1006 2367 1064 2393
rect 1006 2333 1018 2367
rect 1052 2333 1064 2367
rect 1006 2307 1064 2333
rect 1106 2367 1164 2393
rect 1106 2333 1118 2367
rect 1152 2333 1164 2367
rect 1106 2307 1164 2333
rect 1206 2367 1264 2393
rect 1206 2333 1218 2367
rect 1252 2333 1264 2367
rect 1206 2307 1264 2333
rect 1306 2367 1364 2393
rect 1306 2333 1318 2367
rect 1352 2333 1364 2367
rect 1306 2307 1364 2333
rect 1406 2367 1464 2393
rect 1406 2333 1418 2367
rect 1452 2333 1464 2367
rect 1406 2307 1464 2333
rect 1506 2367 1564 2393
rect 1506 2333 1518 2367
rect 1552 2333 1564 2367
rect 1506 2307 1564 2333
rect 1606 2367 1664 2393
rect 1606 2333 1618 2367
rect 1652 2333 1664 2367
rect 1606 2307 1664 2333
rect 1706 2367 1764 2393
rect 1706 2333 1718 2367
rect 1752 2333 1764 2367
rect 1706 2307 1764 2333
rect 1806 2367 1864 2393
rect 1806 2333 1818 2367
rect 1852 2333 1864 2367
rect 1806 2307 1864 2333
rect 1906 2367 1964 2393
rect 1906 2333 1918 2367
rect 1952 2333 1964 2367
rect 1906 2307 1964 2333
rect 2006 2367 2064 2393
rect 2006 2333 2018 2367
rect 2052 2333 2064 2367
rect 2006 2307 2064 2333
rect 2106 2367 2164 2393
rect 2106 2333 2118 2367
rect 2152 2333 2164 2367
rect 2106 2307 2164 2333
rect 2206 2367 2264 2393
rect 2206 2333 2218 2367
rect 2252 2333 2264 2367
rect 2206 2307 2264 2333
rect 2306 2367 2364 2393
rect 2306 2333 2312 2367
rect 2352 2333 2364 2367
rect 2306 2307 2364 2333
rect 2406 2367 2464 2393
rect 2406 2333 2418 2367
rect 2458 2333 2464 2367
rect 2406 2307 2464 2333
rect 2506 2367 2564 2393
rect 2506 2333 2518 2367
rect 2552 2333 2564 2367
rect 2506 2307 2564 2333
rect 2606 2367 2664 2393
rect 2606 2333 2612 2367
rect 2652 2333 2664 2367
rect 2606 2307 2664 2333
rect 2706 2367 2764 2393
rect 2706 2333 2718 2367
rect 2758 2333 2764 2367
rect 2706 2307 2764 2333
rect 2806 2367 2864 2393
rect 2806 2333 2818 2367
rect 2852 2333 2864 2367
rect 2806 2307 2864 2333
rect 2906 2367 2964 2393
rect 2906 2333 2918 2367
rect 2952 2333 2964 2367
rect 2906 2307 2964 2333
rect 3006 2367 3064 2393
rect 3006 2333 3018 2367
rect 3052 2333 3064 2367
rect 3006 2307 3064 2333
rect 3106 2367 3164 2393
rect 3106 2333 3118 2367
rect 3152 2333 3164 2367
rect 3106 2307 3164 2333
rect 3206 2367 3264 2393
rect 3206 2333 3218 2367
rect 3252 2333 3264 2367
rect 3206 2307 3264 2333
rect 3306 2367 3364 2393
rect 3306 2333 3318 2367
rect 3352 2333 3364 2367
rect 3306 2307 3364 2333
rect 3406 2367 3464 2393
rect 3406 2333 3418 2367
rect 3452 2333 3464 2367
rect 3406 2307 3464 2333
rect 3506 2367 3564 2393
rect 3506 2333 3518 2367
rect 3552 2333 3564 2367
rect 3506 2307 3564 2333
rect 3606 2367 3664 2393
rect 3606 2333 3618 2367
rect 3652 2333 3664 2367
rect 3606 2307 3664 2333
rect 3706 2367 3764 2393
rect 3706 2333 3718 2367
rect 3752 2333 3764 2367
rect 3706 2307 3764 2333
rect 3806 2367 3864 2393
rect 3806 2333 3818 2367
rect 3852 2333 3864 2367
rect 3806 2307 3864 2333
rect 3906 2367 3964 2393
rect 3906 2333 3918 2367
rect 3952 2333 3964 2367
rect 3906 2307 3964 2333
rect 4006 2367 4064 2393
rect 4006 2333 4018 2367
rect 4052 2333 4064 2367
rect 4006 2307 4064 2333
rect 4106 2367 4164 2393
rect 4106 2333 4118 2367
rect 4152 2333 4164 2367
rect 4106 2307 4164 2333
rect 4206 2367 4264 2393
rect 4206 2333 4218 2367
rect 4252 2333 4264 2367
rect 4206 2307 4264 2333
rect 4306 2367 4364 2393
rect 4306 2333 4318 2367
rect 4352 2333 4364 2367
rect 4306 2307 4364 2333
rect 4406 2367 4464 2393
rect 4406 2333 4418 2367
rect 4452 2333 4464 2367
rect 4406 2307 4464 2333
rect 4506 2367 4564 2393
rect 4506 2333 4518 2367
rect 4552 2333 4564 2367
rect 4506 2307 4564 2333
rect 4606 2367 4664 2393
rect 4606 2333 4618 2367
rect 4652 2333 4664 2367
rect 4606 2307 4664 2333
rect 4706 2367 4764 2393
rect 4706 2333 4718 2367
rect 4752 2333 4764 2367
rect 4706 2307 4764 2333
rect 4806 2367 4864 2393
rect 4806 2333 4818 2367
rect 4852 2333 4864 2367
rect 4806 2307 4864 2333
rect 4906 2367 4964 2393
rect 4906 2333 4918 2367
rect 4952 2333 4964 2367
rect 4906 2307 4964 2333
rect 5006 2367 5064 2393
rect 5006 2333 5018 2367
rect 5052 2333 5064 2367
rect 5006 2307 5064 2333
rect 5106 2367 5164 2393
rect 5106 2333 5118 2367
rect 5152 2333 5164 2367
rect 5106 2307 5164 2333
rect 5206 2367 5264 2393
rect 5206 2333 5218 2367
rect 5252 2333 5264 2367
rect 5206 2307 5264 2333
rect 5306 2367 5364 2393
rect 5306 2333 5318 2367
rect 5352 2333 5364 2367
rect 5306 2307 5364 2333
rect 5406 2367 5464 2393
rect 5406 2333 5418 2367
rect 5452 2333 5464 2367
rect 5406 2307 5464 2333
rect 5506 2367 5564 2393
rect 5506 2333 5518 2367
rect 5552 2333 5564 2367
rect 5506 2307 5564 2333
rect 5606 2367 5664 2393
rect 5606 2333 5618 2367
rect 5652 2333 5664 2367
rect 5606 2307 5664 2333
rect 5706 2367 5764 2393
rect 5706 2333 5718 2367
rect 5752 2333 5764 2367
rect 5706 2307 5764 2333
rect 5806 2367 5864 2393
rect 5806 2333 5818 2367
rect 5852 2333 5864 2367
rect 5806 2307 5864 2333
rect 5906 2367 5964 2393
rect 5906 2333 5918 2367
rect 5952 2333 5964 2367
rect 5906 2307 5964 2333
rect 6006 2367 6064 2393
rect 6006 2333 6018 2367
rect 6052 2333 6064 2367
rect 6006 2307 6064 2333
rect 6106 2367 6164 2393
rect 6106 2333 6118 2367
rect 6152 2333 6164 2367
rect 6106 2307 6164 2333
rect 6206 2367 6264 2393
rect 6206 2333 6218 2367
rect 6252 2333 6264 2367
rect 6206 2307 6264 2333
rect 6306 2367 6364 2393
rect 6306 2333 6318 2367
rect 6352 2333 6364 2367
rect 6306 2307 6364 2333
rect 6406 2367 6464 2393
rect 6406 2333 6418 2367
rect 6452 2333 6464 2367
rect 6406 2307 6464 2333
rect 6506 2367 6564 2393
rect 6506 2333 6518 2367
rect 6552 2333 6564 2367
rect 6506 2307 6564 2333
rect 6606 2367 6664 2393
rect 6606 2333 6618 2367
rect 6652 2333 6664 2367
rect 6606 2307 6664 2333
rect 6706 2367 6764 2393
rect 6706 2333 6718 2367
rect 6752 2333 6764 2367
rect 6706 2307 6764 2333
rect 6806 2367 6864 2393
rect 6806 2333 6818 2367
rect 6852 2333 6864 2367
rect 6806 2307 6864 2333
rect 6906 2367 6964 2393
rect 6906 2333 6912 2367
rect 6952 2333 6964 2367
rect 6906 2307 6964 2333
rect 7006 2367 7064 2393
rect 7006 2333 7018 2367
rect 7058 2333 7064 2367
rect 7006 2307 7064 2333
rect 7106 2367 7164 2393
rect 7106 2333 7118 2367
rect 7152 2333 7164 2367
rect 7106 2307 7164 2333
rect 7206 2367 7264 2393
rect 7206 2333 7212 2367
rect 7252 2333 7264 2367
rect 7206 2307 7264 2333
rect 7306 2367 7364 2393
rect 7306 2333 7318 2367
rect 7358 2333 7364 2367
rect 7306 2307 7364 2333
rect 7406 2367 7464 2393
rect 7406 2333 7418 2367
rect 7452 2333 7464 2367
rect 7406 2307 7464 2333
rect 7506 2367 7564 2393
rect 7506 2333 7518 2367
rect 7552 2333 7564 2367
rect 7506 2307 7564 2333
rect 7606 2367 7664 2393
rect 7606 2333 7618 2367
rect 7652 2333 7664 2367
rect 7606 2307 7664 2333
rect 7706 2367 7764 2393
rect 7706 2333 7718 2367
rect 7752 2333 7764 2367
rect 7706 2307 7764 2333
rect 7806 2367 7864 2393
rect 7806 2333 7818 2367
rect 7852 2333 7864 2367
rect 7806 2307 7864 2333
rect 7906 2367 7964 2393
rect 7906 2333 7918 2367
rect 7952 2333 7964 2367
rect 7906 2307 7964 2333
rect 8006 2367 8064 2393
rect 8006 2333 8018 2367
rect 8052 2333 8064 2367
rect 8006 2307 8064 2333
rect 8106 2367 8164 2393
rect 8106 2333 8118 2367
rect 8152 2333 8164 2367
rect 8106 2307 8164 2333
rect 8206 2367 8264 2393
rect 8206 2333 8218 2367
rect 8252 2333 8264 2367
rect 8206 2307 8264 2333
rect 8306 2367 8364 2393
rect 8306 2333 8318 2367
rect 8352 2333 8364 2367
rect 8306 2307 8364 2333
rect 8406 2367 8464 2393
rect 8406 2333 8418 2367
rect 8452 2333 8464 2367
rect 8406 2307 8464 2333
rect 8506 2367 8564 2393
rect 8506 2333 8512 2367
rect 8552 2333 8564 2367
rect 8506 2307 8564 2333
rect 8606 2367 8664 2393
rect 8606 2333 8618 2367
rect 8658 2333 8664 2367
rect 8606 2307 8664 2333
rect 8706 2367 8764 2393
rect 8706 2333 8718 2367
rect 8752 2333 8764 2367
rect 8706 2307 8764 2333
rect 8806 2367 8864 2393
rect 8806 2333 8818 2367
rect 8852 2333 8864 2367
rect 8806 2307 8864 2333
rect 8906 2367 8964 2393
rect 8906 2333 8918 2367
rect 8952 2333 8964 2367
rect 8906 2307 8964 2333
rect 9006 2367 9064 2393
rect 9006 2333 9018 2367
rect 9052 2333 9064 2367
rect 9006 2307 9064 2333
rect 9106 2367 9164 2393
rect 9106 2333 9118 2367
rect 9152 2333 9164 2367
rect 9106 2307 9164 2333
rect 9206 2367 9264 2393
rect 9206 2333 9218 2367
rect 9252 2333 9264 2367
rect 9206 2307 9264 2333
rect 9306 2367 9364 2393
rect 9306 2333 9318 2367
rect 9352 2333 9364 2367
rect 9306 2307 9364 2333
rect 9406 2367 9464 2393
rect 9406 2333 9418 2367
rect 9452 2333 9464 2367
rect 9406 2307 9464 2333
rect 9506 2367 9564 2393
rect 9506 2333 9518 2367
rect 9552 2333 9564 2367
rect 9506 2307 9564 2333
rect 9606 2367 9664 2393
rect 9606 2333 9612 2367
rect 9652 2333 9664 2367
rect 9606 2307 9664 2333
rect 9706 2367 9764 2393
rect 9706 2333 9718 2367
rect 9758 2333 9764 2367
rect 9706 2307 9764 2333
rect 9806 2367 9864 2393
rect 9806 2333 9818 2367
rect 9852 2333 9864 2367
rect 9806 2307 9864 2333
rect 9906 2367 9964 2393
rect 9906 2333 9918 2367
rect 9952 2333 9964 2367
rect 9906 2307 9964 2333
rect 10006 2367 10064 2393
rect 10006 2333 10018 2367
rect 10052 2333 10064 2367
rect 10006 2307 10064 2333
rect 10106 2367 10164 2393
rect 10106 2333 10118 2367
rect 10152 2333 10164 2367
rect 10106 2307 10164 2333
rect 10206 2367 10264 2393
rect 10206 2333 10218 2367
rect 10252 2333 10264 2367
rect 10206 2307 10264 2333
rect 10306 2367 10364 2393
rect 10306 2333 10318 2367
rect 10352 2333 10364 2367
rect 10306 2307 10364 2333
rect 10406 2367 10464 2393
rect 10406 2333 10418 2367
rect 10452 2333 10464 2367
rect 10406 2307 10464 2333
rect 10506 2367 10564 2393
rect 10506 2333 10518 2367
rect 10552 2333 10564 2367
rect 10506 2307 10564 2333
rect 10606 2367 10664 2393
rect 10606 2333 10618 2367
rect 10652 2333 10664 2367
rect 10606 2307 10664 2333
rect 10706 2367 10764 2393
rect 10706 2333 10718 2367
rect 10752 2333 10764 2367
rect 10706 2307 10764 2333
rect 10806 2367 10864 2393
rect 10806 2333 10818 2367
rect 10852 2333 10864 2367
rect 10806 2307 10864 2333
rect 10906 2367 10964 2393
rect 10906 2333 10918 2367
rect 10952 2333 10964 2367
rect 10906 2307 10964 2333
rect 11006 2367 11064 2393
rect 11006 2333 11018 2367
rect 11052 2333 11064 2367
rect 11006 2307 11064 2333
rect 11106 2367 11164 2393
rect 11106 2333 11118 2367
rect 11152 2333 11164 2367
rect 11106 2307 11164 2333
rect 11206 2367 11264 2393
rect 11206 2333 11218 2367
rect 11252 2333 11264 2367
rect 11206 2307 11264 2333
rect 11306 2367 11364 2393
rect 11306 2333 11318 2367
rect 11352 2333 11364 2367
rect 11306 2307 11364 2333
rect 11406 2367 11464 2393
rect 11406 2333 11418 2367
rect 11452 2333 11464 2367
rect 11406 2307 11464 2333
rect 11506 2367 11564 2393
rect 11506 2333 11518 2367
rect 11552 2333 11564 2367
rect 11506 2307 11564 2333
rect 11606 2367 11664 2393
rect 11606 2333 11618 2367
rect 11652 2333 11664 2367
rect 11606 2307 11664 2333
rect 11706 2367 11764 2393
rect 11706 2333 11712 2367
rect 11752 2333 11764 2367
rect 11706 2307 11764 2333
rect 11806 2367 11864 2393
rect 11806 2333 11818 2367
rect 11858 2333 11864 2367
rect 11806 2307 11864 2333
rect 11906 2367 11964 2393
rect 11906 2333 11912 2367
rect 11952 2333 11964 2367
rect 11906 2307 11964 2333
rect 12006 2367 12064 2393
rect 12006 2333 12018 2367
rect 12058 2333 12064 2367
rect 12006 2307 12064 2333
rect 12106 2367 12164 2393
rect 12106 2333 12118 2367
rect 12152 2333 12164 2367
rect 12106 2307 12164 2333
rect 12206 2367 12264 2393
rect 12206 2333 12218 2367
rect 12252 2333 12264 2367
rect 12206 2307 12264 2333
rect 12306 2367 12364 2393
rect 12306 2333 12318 2367
rect 12352 2333 12364 2367
rect 12306 2307 12364 2333
rect 12406 2367 12464 2393
rect 12406 2333 12418 2367
rect 12452 2333 12464 2367
rect 12406 2307 12464 2333
rect 12506 2367 12564 2393
rect 12506 2333 12512 2367
rect 12552 2333 12564 2367
rect 12506 2307 12564 2333
rect 12606 2367 12664 2393
rect 12606 2333 12618 2367
rect 12658 2333 12664 2367
rect 12606 2307 12664 2333
rect 12706 2367 12764 2393
rect 12706 2333 12718 2367
rect 12752 2333 12764 2367
rect 12706 2307 12764 2333
rect 12806 2367 12864 2393
rect 13018 2386 13262 2420
rect 12806 2333 12818 2367
rect 12852 2333 12864 2367
rect 12908 2348 12916 2382
rect 12958 2348 12974 2382
rect 13018 2367 13052 2386
rect 12806 2307 12864 2333
rect 13228 2383 13262 2386
rect 13228 2367 13362 2383
rect 13018 2317 13052 2333
rect 13096 2318 13112 2352
rect 13154 2318 13162 2352
rect 13262 2333 13328 2367
rect 13228 2317 13362 2333
rect 13428 2367 13562 2383
rect 13462 2333 13528 2367
rect 13428 2317 13562 2333
rect 13628 2367 13662 2383
rect 13628 2317 13662 2333
rect 6 2227 64 2253
rect 6 2193 18 2227
rect 58 2193 64 2227
rect 6 2167 64 2193
rect 106 2227 164 2253
rect 106 2193 118 2227
rect 152 2193 164 2227
rect 106 2167 164 2193
rect 206 2227 264 2253
rect 206 2193 218 2227
rect 252 2193 264 2227
rect 206 2167 264 2193
rect 306 2227 364 2253
rect 306 2193 318 2227
rect 352 2193 364 2227
rect 306 2167 364 2193
rect 406 2227 464 2253
rect 406 2193 418 2227
rect 452 2193 464 2227
rect 406 2167 464 2193
rect 506 2227 564 2253
rect 506 2193 518 2227
rect 552 2193 564 2227
rect 506 2167 564 2193
rect 606 2227 664 2253
rect 606 2193 618 2227
rect 652 2193 664 2227
rect 606 2167 664 2193
rect 706 2227 764 2253
rect 706 2193 718 2227
rect 752 2193 764 2227
rect 706 2167 764 2193
rect 806 2227 864 2253
rect 806 2193 812 2227
rect 852 2193 864 2227
rect 806 2167 864 2193
rect 906 2227 964 2253
rect 906 2193 918 2227
rect 958 2193 964 2227
rect 906 2167 964 2193
rect 1006 2227 1064 2253
rect 1006 2193 1012 2227
rect 1052 2193 1064 2227
rect 1006 2167 1064 2193
rect 1106 2227 1164 2253
rect 1106 2193 1118 2227
rect 1158 2193 1164 2227
rect 1106 2167 1164 2193
rect 1206 2227 1264 2253
rect 1206 2193 1218 2227
rect 1252 2193 1264 2227
rect 1206 2167 1264 2193
rect 1306 2227 1364 2253
rect 1306 2193 1318 2227
rect 1352 2193 1364 2227
rect 1306 2167 1364 2193
rect 1406 2227 1464 2253
rect 1406 2193 1418 2227
rect 1452 2193 1464 2227
rect 1406 2167 1464 2193
rect 1506 2227 1564 2253
rect 1506 2193 1518 2227
rect 1552 2193 1564 2227
rect 1506 2167 1564 2193
rect 1606 2227 1664 2253
rect 1606 2193 1618 2227
rect 1652 2193 1664 2227
rect 1606 2167 1664 2193
rect 1706 2227 1764 2253
rect 1706 2193 1718 2227
rect 1752 2193 1764 2227
rect 1706 2167 1764 2193
rect 1806 2227 1864 2253
rect 1806 2193 1818 2227
rect 1852 2193 1864 2227
rect 1806 2167 1864 2193
rect 1906 2227 1964 2253
rect 1906 2193 1918 2227
rect 1952 2193 1964 2227
rect 1906 2167 1964 2193
rect 2006 2227 2064 2253
rect 2006 2193 2018 2227
rect 2052 2193 2064 2227
rect 2006 2167 2064 2193
rect 2106 2227 2164 2253
rect 2106 2193 2118 2227
rect 2152 2193 2164 2227
rect 2106 2167 2164 2193
rect 2206 2227 2264 2253
rect 2206 2193 2218 2227
rect 2252 2193 2264 2227
rect 2206 2167 2264 2193
rect 2306 2227 2364 2253
rect 2306 2193 2318 2227
rect 2352 2193 2364 2227
rect 2306 2167 2364 2193
rect 2406 2227 2464 2253
rect 2406 2193 2418 2227
rect 2452 2193 2464 2227
rect 2406 2167 2464 2193
rect 2506 2227 2564 2253
rect 2506 2193 2518 2227
rect 2552 2193 2564 2227
rect 2506 2167 2564 2193
rect 2606 2227 2664 2253
rect 2606 2193 2612 2227
rect 2652 2193 2664 2227
rect 2606 2167 2664 2193
rect 2706 2227 2764 2253
rect 2706 2193 2718 2227
rect 2758 2193 2764 2227
rect 2706 2167 2764 2193
rect 2806 2227 2864 2253
rect 2806 2193 2812 2227
rect 2852 2193 2864 2227
rect 2806 2167 2864 2193
rect 2906 2227 2964 2253
rect 2906 2193 2918 2227
rect 2958 2193 2964 2227
rect 2906 2167 2964 2193
rect 3006 2227 3064 2253
rect 3006 2193 3012 2227
rect 3052 2193 3064 2227
rect 3006 2167 3064 2193
rect 3106 2227 3164 2253
rect 3106 2193 3118 2227
rect 3158 2193 3164 2227
rect 3106 2167 3164 2193
rect 3206 2227 3264 2253
rect 3206 2193 3218 2227
rect 3252 2193 3264 2227
rect 3206 2167 3264 2193
rect 3306 2227 3364 2253
rect 3306 2193 3312 2227
rect 3352 2193 3364 2227
rect 3306 2167 3364 2193
rect 3406 2227 3464 2253
rect 3406 2193 3418 2227
rect 3458 2193 3464 2227
rect 3406 2167 3464 2193
rect 3506 2227 3564 2253
rect 3506 2193 3518 2227
rect 3552 2193 3564 2227
rect 3506 2167 3564 2193
rect 3606 2227 3664 2253
rect 3606 2193 3612 2227
rect 3652 2193 3664 2227
rect 3606 2167 3664 2193
rect 3706 2227 3764 2253
rect 3706 2193 3718 2227
rect 3758 2193 3764 2227
rect 3706 2167 3764 2193
rect 3806 2227 3864 2253
rect 3806 2193 3812 2227
rect 3852 2193 3864 2227
rect 3806 2167 3864 2193
rect 3906 2227 3964 2253
rect 3906 2193 3918 2227
rect 3958 2193 3964 2227
rect 3906 2167 3964 2193
rect 4006 2227 4064 2253
rect 4006 2193 4018 2227
rect 4052 2193 4064 2227
rect 4006 2167 4064 2193
rect 4106 2227 4164 2253
rect 4106 2193 4118 2227
rect 4152 2193 4164 2227
rect 4106 2167 4164 2193
rect 4206 2227 4264 2253
rect 4206 2193 4218 2227
rect 4252 2193 4264 2227
rect 4206 2167 4264 2193
rect 4306 2227 4364 2253
rect 4306 2193 4312 2227
rect 4352 2193 4364 2227
rect 4306 2167 4364 2193
rect 4406 2227 4464 2253
rect 4406 2193 4418 2227
rect 4458 2193 4464 2227
rect 4406 2167 4464 2193
rect 4506 2227 4564 2253
rect 4506 2193 4518 2227
rect 4552 2193 4564 2227
rect 4506 2167 4564 2193
rect 4606 2227 4664 2253
rect 4606 2193 4618 2227
rect 4652 2193 4664 2227
rect 4606 2167 4664 2193
rect 4706 2227 4764 2253
rect 4706 2193 4718 2227
rect 4752 2193 4764 2227
rect 4706 2167 4764 2193
rect 4806 2227 4864 2253
rect 4806 2193 4818 2227
rect 4852 2193 4864 2227
rect 4806 2167 4864 2193
rect 4906 2227 4964 2253
rect 4906 2193 4918 2227
rect 4952 2193 4964 2227
rect 4906 2167 4964 2193
rect 5006 2227 5064 2253
rect 5006 2193 5018 2227
rect 5052 2193 5064 2227
rect 5006 2167 5064 2193
rect 5106 2227 5164 2253
rect 5106 2193 5118 2227
rect 5152 2193 5164 2227
rect 5106 2167 5164 2193
rect 5206 2227 5264 2253
rect 5206 2193 5218 2227
rect 5252 2193 5264 2227
rect 5206 2167 5264 2193
rect 5306 2227 5364 2253
rect 5306 2193 5318 2227
rect 5352 2193 5364 2227
rect 5306 2167 5364 2193
rect 5406 2227 5464 2253
rect 5406 2193 5418 2227
rect 5452 2193 5464 2227
rect 5406 2167 5464 2193
rect 5506 2227 5564 2253
rect 5506 2193 5518 2227
rect 5552 2193 5564 2227
rect 5506 2167 5564 2193
rect 5606 2227 5664 2253
rect 5606 2193 5618 2227
rect 5652 2193 5664 2227
rect 5606 2167 5664 2193
rect 5706 2227 5764 2253
rect 5706 2193 5718 2227
rect 5752 2193 5764 2227
rect 5706 2167 5764 2193
rect 5806 2227 5864 2253
rect 5806 2193 5818 2227
rect 5852 2193 5864 2227
rect 5806 2167 5864 2193
rect 5906 2227 5964 2253
rect 5906 2193 5918 2227
rect 5952 2193 5964 2227
rect 5906 2167 5964 2193
rect 6006 2227 6064 2253
rect 6006 2193 6018 2227
rect 6052 2193 6064 2227
rect 6006 2167 6064 2193
rect 6106 2227 6164 2253
rect 6106 2193 6112 2227
rect 6152 2193 6164 2227
rect 6106 2167 6164 2193
rect 6206 2227 6264 2253
rect 6206 2193 6218 2227
rect 6258 2193 6264 2227
rect 6206 2167 6264 2193
rect 6306 2227 6364 2253
rect 6306 2193 6318 2227
rect 6352 2193 6364 2227
rect 6306 2167 6364 2193
rect 6406 2227 6464 2253
rect 6406 2193 6412 2227
rect 6452 2193 6464 2227
rect 6406 2167 6464 2193
rect 6506 2227 6564 2253
rect 6506 2193 6518 2227
rect 6558 2193 6564 2227
rect 6506 2167 6564 2193
rect 6606 2227 6664 2253
rect 6606 2193 6618 2227
rect 6652 2193 6664 2227
rect 6606 2167 6664 2193
rect 6706 2227 6764 2253
rect 6706 2193 6712 2227
rect 6752 2193 6764 2227
rect 6706 2167 6764 2193
rect 6806 2227 6864 2253
rect 6806 2193 6818 2227
rect 6858 2193 6864 2227
rect 6806 2167 6864 2193
rect 6906 2227 6964 2253
rect 6906 2193 6912 2227
rect 6952 2193 6964 2227
rect 6906 2167 6964 2193
rect 7006 2227 7064 2253
rect 7006 2193 7018 2227
rect 7058 2193 7064 2227
rect 7006 2167 7064 2193
rect 7106 2227 7164 2253
rect 7106 2193 7118 2227
rect 7152 2193 7164 2227
rect 7106 2167 7164 2193
rect 7206 2227 7264 2253
rect 7206 2193 7218 2227
rect 7252 2193 7264 2227
rect 7206 2167 7264 2193
rect 7306 2227 7364 2253
rect 7306 2193 7318 2227
rect 7352 2193 7364 2227
rect 7306 2167 7364 2193
rect 7406 2227 7464 2253
rect 7406 2193 7418 2227
rect 7452 2193 7464 2227
rect 7406 2167 7464 2193
rect 7506 2227 7564 2253
rect 7506 2193 7512 2227
rect 7552 2193 7564 2227
rect 7506 2167 7564 2193
rect 7606 2227 7664 2253
rect 7606 2193 7618 2227
rect 7658 2193 7664 2227
rect 7606 2167 7664 2193
rect 7706 2227 7764 2253
rect 7706 2193 7712 2227
rect 7752 2193 7764 2227
rect 7706 2167 7764 2193
rect 7806 2227 7864 2253
rect 7806 2193 7818 2227
rect 7858 2193 7864 2227
rect 7806 2167 7864 2193
rect 7906 2227 7964 2253
rect 7906 2193 7918 2227
rect 7952 2193 7964 2227
rect 7906 2167 7964 2193
rect 8006 2227 8064 2253
rect 8006 2193 8018 2227
rect 8052 2193 8064 2227
rect 8006 2167 8064 2193
rect 8106 2227 8164 2253
rect 8106 2193 8118 2227
rect 8152 2193 8164 2227
rect 8106 2167 8164 2193
rect 8206 2227 8264 2253
rect 8206 2193 8218 2227
rect 8252 2193 8264 2227
rect 8206 2167 8264 2193
rect 8306 2227 8364 2253
rect 8306 2193 8318 2227
rect 8352 2193 8364 2227
rect 8306 2167 8364 2193
rect 8406 2227 8464 2253
rect 8406 2193 8418 2227
rect 8452 2193 8464 2227
rect 8406 2167 8464 2193
rect 8506 2227 8564 2253
rect 8506 2193 8518 2227
rect 8552 2193 8564 2227
rect 8506 2167 8564 2193
rect 8606 2227 8664 2253
rect 8606 2193 8618 2227
rect 8652 2193 8664 2227
rect 8606 2167 8664 2193
rect 8706 2227 8764 2253
rect 8706 2193 8718 2227
rect 8752 2193 8764 2227
rect 8706 2167 8764 2193
rect 8806 2227 8864 2253
rect 8806 2193 8812 2227
rect 8852 2193 8864 2227
rect 8806 2167 8864 2193
rect 8906 2227 8964 2253
rect 8906 2193 8918 2227
rect 8958 2193 8964 2227
rect 8906 2167 8964 2193
rect 9006 2227 9064 2253
rect 9006 2193 9012 2227
rect 9052 2193 9064 2227
rect 9006 2167 9064 2193
rect 9106 2227 9164 2253
rect 9106 2193 9118 2227
rect 9158 2193 9164 2227
rect 9106 2167 9164 2193
rect 9206 2227 9264 2253
rect 9206 2193 9212 2227
rect 9252 2193 9264 2227
rect 9206 2167 9264 2193
rect 9306 2227 9364 2253
rect 9306 2193 9318 2227
rect 9358 2193 9364 2227
rect 9306 2167 9364 2193
rect 9406 2227 9464 2253
rect 9406 2193 9418 2227
rect 9452 2193 9464 2227
rect 9406 2167 9464 2193
rect 9506 2227 9564 2253
rect 9506 2193 9512 2227
rect 9552 2193 9564 2227
rect 9506 2167 9564 2193
rect 9606 2227 9664 2253
rect 9606 2193 9618 2227
rect 9658 2193 9664 2227
rect 9606 2167 9664 2193
rect 9706 2227 9764 2253
rect 9706 2193 9718 2227
rect 9752 2193 9764 2227
rect 9706 2167 9764 2193
rect 9806 2227 9864 2253
rect 9806 2193 9818 2227
rect 9852 2193 9864 2227
rect 9806 2167 9864 2193
rect 9906 2227 9964 2253
rect 9906 2193 9918 2227
rect 9952 2193 9964 2227
rect 9906 2167 9964 2193
rect 10006 2227 10064 2253
rect 10006 2193 10018 2227
rect 10052 2193 10064 2227
rect 10006 2167 10064 2193
rect 10106 2227 10164 2253
rect 10106 2193 10118 2227
rect 10152 2193 10164 2227
rect 10106 2167 10164 2193
rect 10206 2227 10264 2253
rect 10206 2193 10218 2227
rect 10252 2193 10264 2227
rect 10206 2167 10264 2193
rect 10306 2227 10364 2253
rect 10306 2193 10318 2227
rect 10352 2193 10364 2227
rect 10306 2167 10364 2193
rect 10406 2227 10464 2253
rect 10406 2193 10418 2227
rect 10452 2193 10464 2227
rect 10406 2167 10464 2193
rect 10506 2227 10564 2253
rect 10506 2193 10512 2227
rect 10552 2193 10564 2227
rect 10506 2167 10564 2193
rect 10606 2227 10664 2253
rect 10606 2193 10618 2227
rect 10658 2193 10664 2227
rect 10606 2167 10664 2193
rect 10706 2227 10764 2253
rect 10706 2193 10718 2227
rect 10752 2193 10764 2227
rect 10706 2167 10764 2193
rect 10806 2227 10864 2253
rect 10806 2193 10818 2227
rect 10852 2193 10864 2227
rect 10806 2167 10864 2193
rect 10906 2227 10964 2253
rect 10906 2193 10918 2227
rect 10952 2193 10964 2227
rect 10906 2167 10964 2193
rect 11006 2227 11064 2253
rect 11006 2193 11018 2227
rect 11052 2193 11064 2227
rect 11006 2167 11064 2193
rect 11106 2227 11164 2253
rect 11106 2193 11118 2227
rect 11152 2193 11164 2227
rect 11106 2167 11164 2193
rect 11206 2227 11264 2253
rect 11206 2193 11218 2227
rect 11252 2193 11264 2227
rect 11206 2167 11264 2193
rect 11306 2227 11364 2253
rect 11306 2193 11318 2227
rect 11352 2193 11364 2227
rect 11306 2167 11364 2193
rect 11406 2227 11464 2253
rect 11406 2193 11418 2227
rect 11452 2193 11464 2227
rect 11406 2167 11464 2193
rect 11506 2227 11564 2253
rect 11506 2193 11518 2227
rect 11552 2193 11564 2227
rect 11506 2167 11564 2193
rect 11606 2227 11664 2253
rect 11606 2193 11618 2227
rect 11652 2193 11664 2227
rect 11606 2167 11664 2193
rect 11706 2227 11764 2253
rect 11706 2193 11718 2227
rect 11752 2193 11764 2227
rect 11706 2167 11764 2193
rect 11806 2227 11864 2253
rect 11806 2193 11818 2227
rect 11852 2193 11864 2227
rect 11806 2167 11864 2193
rect 11906 2227 11964 2253
rect 11906 2193 11918 2227
rect 11952 2193 11964 2227
rect 11906 2167 11964 2193
rect 12006 2227 12064 2253
rect 12006 2193 12012 2227
rect 12052 2193 12064 2227
rect 12006 2167 12064 2193
rect 12106 2227 12164 2253
rect 12106 2193 12118 2227
rect 12158 2193 12164 2227
rect 12106 2167 12164 2193
rect 12206 2227 12264 2253
rect 12206 2193 12218 2227
rect 12252 2193 12264 2227
rect 12206 2167 12264 2193
rect 12306 2227 12364 2253
rect 12306 2193 12312 2227
rect 12352 2193 12364 2227
rect 12306 2167 12364 2193
rect 12406 2227 12464 2253
rect 12406 2193 12418 2227
rect 12458 2193 12464 2227
rect 12406 2167 12464 2193
rect 12506 2227 12564 2253
rect 12506 2193 12518 2227
rect 12552 2193 12564 2227
rect 12506 2167 12564 2193
rect 12606 2227 12664 2253
rect 12606 2193 12612 2227
rect 12652 2193 12664 2227
rect 12606 2167 12664 2193
rect 12706 2227 12764 2253
rect 12706 2193 12718 2227
rect 12758 2193 12764 2227
rect 12706 2167 12764 2193
rect 12806 2227 12864 2253
rect 13018 2246 13262 2280
rect 12806 2193 12812 2227
rect 12852 2193 12864 2227
rect 12908 2208 12916 2242
rect 12958 2208 12974 2242
rect 13018 2227 13052 2246
rect 12806 2167 12864 2193
rect 13228 2227 13262 2246
rect 13018 2177 13052 2193
rect 13096 2178 13112 2212
rect 13154 2178 13162 2212
rect 13228 2177 13262 2193
rect 13328 2227 13562 2243
rect 13362 2193 13428 2227
rect 13462 2193 13528 2227
rect 13328 2177 13562 2193
rect 13628 2227 13662 2243
rect 13628 2177 13662 2193
rect 6 2087 64 2113
rect 6 2053 18 2087
rect 52 2053 64 2087
rect 6 2027 64 2053
rect 106 2087 164 2113
rect 106 2053 118 2087
rect 152 2053 164 2087
rect 106 2027 164 2053
rect 206 2087 264 2113
rect 206 2053 218 2087
rect 252 2053 264 2087
rect 206 2027 264 2053
rect 306 2087 364 2113
rect 306 2053 318 2087
rect 352 2053 364 2087
rect 306 2027 364 2053
rect 406 2087 464 2113
rect 406 2053 418 2087
rect 452 2053 464 2087
rect 406 2027 464 2053
rect 506 2087 564 2113
rect 506 2053 518 2087
rect 552 2053 564 2087
rect 506 2027 564 2053
rect 606 2087 664 2113
rect 606 2053 618 2087
rect 652 2053 664 2087
rect 606 2027 664 2053
rect 706 2087 764 2113
rect 706 2053 712 2087
rect 752 2053 764 2087
rect 706 2027 764 2053
rect 806 2087 864 2113
rect 806 2053 818 2087
rect 858 2053 864 2087
rect 806 2027 864 2053
rect 906 2087 964 2113
rect 906 2053 918 2087
rect 952 2053 964 2087
rect 906 2027 964 2053
rect 1006 2087 1064 2113
rect 1006 2053 1018 2087
rect 1052 2053 1064 2087
rect 1006 2027 1064 2053
rect 1106 2087 1164 2113
rect 1106 2053 1118 2087
rect 1152 2053 1164 2087
rect 1106 2027 1164 2053
rect 1206 2087 1264 2113
rect 1206 2053 1218 2087
rect 1252 2053 1264 2087
rect 1206 2027 1264 2053
rect 1306 2087 1364 2113
rect 1306 2053 1318 2087
rect 1352 2053 1364 2087
rect 1306 2027 1364 2053
rect 1406 2087 1464 2113
rect 1406 2053 1412 2087
rect 1452 2053 1464 2087
rect 1406 2027 1464 2053
rect 1506 2087 1564 2113
rect 1506 2053 1518 2087
rect 1558 2053 1564 2087
rect 1506 2027 1564 2053
rect 1606 2087 1664 2113
rect 1606 2053 1618 2087
rect 1652 2053 1664 2087
rect 1606 2027 1664 2053
rect 1706 2087 1764 2113
rect 1706 2053 1718 2087
rect 1752 2053 1764 2087
rect 1706 2027 1764 2053
rect 1806 2087 1864 2113
rect 1806 2053 1818 2087
rect 1852 2053 1864 2087
rect 1806 2027 1864 2053
rect 1906 2087 1964 2113
rect 1906 2053 1918 2087
rect 1952 2053 1964 2087
rect 1906 2027 1964 2053
rect 2006 2087 2064 2113
rect 2006 2053 2018 2087
rect 2052 2053 2064 2087
rect 2006 2027 2064 2053
rect 2106 2087 2164 2113
rect 2106 2053 2118 2087
rect 2152 2053 2164 2087
rect 2106 2027 2164 2053
rect 2206 2087 2264 2113
rect 2206 2053 2218 2087
rect 2252 2053 2264 2087
rect 2206 2027 2264 2053
rect 2306 2087 2364 2113
rect 2306 2053 2318 2087
rect 2352 2053 2364 2087
rect 2306 2027 2364 2053
rect 2406 2087 2464 2113
rect 2406 2053 2418 2087
rect 2452 2053 2464 2087
rect 2406 2027 2464 2053
rect 2506 2087 2564 2113
rect 2506 2053 2518 2087
rect 2552 2053 2564 2087
rect 2506 2027 2564 2053
rect 2606 2087 2664 2113
rect 2606 2053 2618 2087
rect 2652 2053 2664 2087
rect 2606 2027 2664 2053
rect 2706 2087 2764 2113
rect 2706 2053 2712 2087
rect 2752 2053 2764 2087
rect 2706 2027 2764 2053
rect 2806 2087 2864 2113
rect 2806 2053 2818 2087
rect 2858 2053 2864 2087
rect 2806 2027 2864 2053
rect 2906 2087 2964 2113
rect 2906 2053 2912 2087
rect 2952 2053 2964 2087
rect 2906 2027 2964 2053
rect 3006 2087 3064 2113
rect 3006 2053 3018 2087
rect 3058 2053 3064 2087
rect 3006 2027 3064 2053
rect 3106 2087 3164 2113
rect 3106 2053 3118 2087
rect 3152 2053 3164 2087
rect 3106 2027 3164 2053
rect 3206 2087 3264 2113
rect 3206 2053 3218 2087
rect 3252 2053 3264 2087
rect 3206 2027 3264 2053
rect 3306 2087 3364 2113
rect 3306 2053 3318 2087
rect 3352 2053 3364 2087
rect 3306 2027 3364 2053
rect 3406 2087 3464 2113
rect 3406 2053 3418 2087
rect 3452 2053 3464 2087
rect 3406 2027 3464 2053
rect 3506 2087 3564 2113
rect 3506 2053 3512 2087
rect 3552 2053 3564 2087
rect 3506 2027 3564 2053
rect 3606 2087 3664 2113
rect 3606 2053 3618 2087
rect 3658 2053 3664 2087
rect 3606 2027 3664 2053
rect 3706 2087 3764 2113
rect 3706 2053 3718 2087
rect 3752 2053 3764 2087
rect 3706 2027 3764 2053
rect 3806 2087 3864 2113
rect 3806 2053 3818 2087
rect 3852 2053 3864 2087
rect 3806 2027 3864 2053
rect 3906 2087 3964 2113
rect 3906 2053 3918 2087
rect 3952 2053 3964 2087
rect 3906 2027 3964 2053
rect 4006 2087 4064 2113
rect 4006 2053 4018 2087
rect 4052 2053 4064 2087
rect 4006 2027 4064 2053
rect 4106 2087 4164 2113
rect 4106 2053 4118 2087
rect 4152 2053 4164 2087
rect 4106 2027 4164 2053
rect 4206 2087 4264 2113
rect 4206 2053 4218 2087
rect 4252 2053 4264 2087
rect 4206 2027 4264 2053
rect 4306 2087 4364 2113
rect 4306 2053 4318 2087
rect 4352 2053 4364 2087
rect 4306 2027 4364 2053
rect 4406 2087 4464 2113
rect 4406 2053 4418 2087
rect 4452 2053 4464 2087
rect 4406 2027 4464 2053
rect 4506 2087 4564 2113
rect 4506 2053 4518 2087
rect 4552 2053 4564 2087
rect 4506 2027 4564 2053
rect 4606 2087 4664 2113
rect 4606 2053 4612 2087
rect 4652 2053 4664 2087
rect 4606 2027 4664 2053
rect 4706 2087 4764 2113
rect 4706 2053 4718 2087
rect 4758 2053 4764 2087
rect 4706 2027 4764 2053
rect 4806 2087 4864 2113
rect 4806 2053 4818 2087
rect 4852 2053 4864 2087
rect 4806 2027 4864 2053
rect 4906 2087 4964 2113
rect 4906 2053 4912 2087
rect 4952 2053 4964 2087
rect 4906 2027 4964 2053
rect 5006 2087 5064 2113
rect 5006 2053 5018 2087
rect 5058 2053 5064 2087
rect 5006 2027 5064 2053
rect 5106 2087 5164 2113
rect 5106 2053 5118 2087
rect 5152 2053 5164 2087
rect 5106 2027 5164 2053
rect 5206 2087 5264 2113
rect 5206 2053 5218 2087
rect 5252 2053 5264 2087
rect 5206 2027 5264 2053
rect 5306 2087 5364 2113
rect 5306 2053 5318 2087
rect 5352 2053 5364 2087
rect 5306 2027 5364 2053
rect 5406 2087 5464 2113
rect 5406 2053 5418 2087
rect 5452 2053 5464 2087
rect 5406 2027 5464 2053
rect 5506 2087 5564 2113
rect 5506 2053 5518 2087
rect 5552 2053 5564 2087
rect 5506 2027 5564 2053
rect 5606 2087 5664 2113
rect 5606 2053 5618 2087
rect 5652 2053 5664 2087
rect 5606 2027 5664 2053
rect 5706 2087 5764 2113
rect 5706 2053 5712 2087
rect 5752 2053 5764 2087
rect 5706 2027 5764 2053
rect 5806 2087 5864 2113
rect 5806 2053 5818 2087
rect 5858 2053 5864 2087
rect 5806 2027 5864 2053
rect 5906 2087 5964 2113
rect 5906 2053 5918 2087
rect 5952 2053 5964 2087
rect 5906 2027 5964 2053
rect 6006 2087 6064 2113
rect 6006 2053 6018 2087
rect 6052 2053 6064 2087
rect 6006 2027 6064 2053
rect 6106 2087 6164 2113
rect 6106 2053 6118 2087
rect 6152 2053 6164 2087
rect 6106 2027 6164 2053
rect 6206 2087 6264 2113
rect 6206 2053 6218 2087
rect 6252 2053 6264 2087
rect 6206 2027 6264 2053
rect 6306 2087 6364 2113
rect 6306 2053 6318 2087
rect 6352 2053 6364 2087
rect 6306 2027 6364 2053
rect 6406 2087 6464 2113
rect 6406 2053 6418 2087
rect 6452 2053 6464 2087
rect 6406 2027 6464 2053
rect 6506 2087 6564 2113
rect 6506 2053 6518 2087
rect 6552 2053 6564 2087
rect 6506 2027 6564 2053
rect 6606 2087 6664 2113
rect 6606 2053 6612 2087
rect 6652 2053 6664 2087
rect 6606 2027 6664 2053
rect 6706 2087 6764 2113
rect 6706 2053 6718 2087
rect 6758 2053 6764 2087
rect 6706 2027 6764 2053
rect 6806 2087 6864 2113
rect 6806 2053 6812 2087
rect 6852 2053 6864 2087
rect 6806 2027 6864 2053
rect 6906 2087 6964 2113
rect 6906 2053 6918 2087
rect 6958 2053 6964 2087
rect 6906 2027 6964 2053
rect 7006 2087 7064 2113
rect 7006 2053 7018 2087
rect 7052 2053 7064 2087
rect 7006 2027 7064 2053
rect 7106 2087 7164 2113
rect 7106 2053 7118 2087
rect 7152 2053 7164 2087
rect 7106 2027 7164 2053
rect 7206 2087 7264 2113
rect 7206 2053 7218 2087
rect 7252 2053 7264 2087
rect 7206 2027 7264 2053
rect 7306 2087 7364 2113
rect 7306 2053 7318 2087
rect 7352 2053 7364 2087
rect 7306 2027 7364 2053
rect 7406 2087 7464 2113
rect 7406 2053 7418 2087
rect 7452 2053 7464 2087
rect 7406 2027 7464 2053
rect 7506 2087 7564 2113
rect 7506 2053 7518 2087
rect 7552 2053 7564 2087
rect 7506 2027 7564 2053
rect 7606 2087 7664 2113
rect 7606 2053 7618 2087
rect 7652 2053 7664 2087
rect 7606 2027 7664 2053
rect 7706 2087 7764 2113
rect 7706 2053 7718 2087
rect 7752 2053 7764 2087
rect 7706 2027 7764 2053
rect 7806 2087 7864 2113
rect 7806 2053 7818 2087
rect 7852 2053 7864 2087
rect 7806 2027 7864 2053
rect 7906 2087 7964 2113
rect 7906 2053 7918 2087
rect 7952 2053 7964 2087
rect 7906 2027 7964 2053
rect 8006 2087 8064 2113
rect 8006 2053 8018 2087
rect 8052 2053 8064 2087
rect 8006 2027 8064 2053
rect 8106 2087 8164 2113
rect 8106 2053 8112 2087
rect 8152 2053 8164 2087
rect 8106 2027 8164 2053
rect 8206 2087 8264 2113
rect 8206 2053 8218 2087
rect 8258 2053 8264 2087
rect 8206 2027 8264 2053
rect 8306 2087 8364 2113
rect 8306 2053 8312 2087
rect 8352 2053 8364 2087
rect 8306 2027 8364 2053
rect 8406 2087 8464 2113
rect 8406 2053 8418 2087
rect 8458 2053 8464 2087
rect 8406 2027 8464 2053
rect 8506 2087 8564 2113
rect 8506 2053 8518 2087
rect 8552 2053 8564 2087
rect 8506 2027 8564 2053
rect 8606 2087 8664 2113
rect 8606 2053 8618 2087
rect 8652 2053 8664 2087
rect 8606 2027 8664 2053
rect 8706 2087 8764 2113
rect 8706 2053 8712 2087
rect 8752 2053 8764 2087
rect 8706 2027 8764 2053
rect 8806 2087 8864 2113
rect 8806 2053 8818 2087
rect 8858 2053 8864 2087
rect 8806 2027 8864 2053
rect 8906 2087 8964 2113
rect 8906 2053 8912 2087
rect 8952 2053 8964 2087
rect 8906 2027 8964 2053
rect 9006 2087 9064 2113
rect 9006 2053 9018 2087
rect 9058 2053 9064 2087
rect 9006 2027 9064 2053
rect 9106 2087 9164 2113
rect 9106 2053 9118 2087
rect 9152 2053 9164 2087
rect 9106 2027 9164 2053
rect 9206 2087 9264 2113
rect 9206 2053 9212 2087
rect 9252 2053 9264 2087
rect 9206 2027 9264 2053
rect 9306 2087 9364 2113
rect 9306 2053 9318 2087
rect 9358 2053 9364 2087
rect 9306 2027 9364 2053
rect 9406 2087 9464 2113
rect 9406 2053 9418 2087
rect 9452 2053 9464 2087
rect 9406 2027 9464 2053
rect 9506 2087 9564 2113
rect 9506 2053 9518 2087
rect 9552 2053 9564 2087
rect 9506 2027 9564 2053
rect 9606 2087 9664 2113
rect 9606 2053 9618 2087
rect 9652 2053 9664 2087
rect 9606 2027 9664 2053
rect 9706 2087 9764 2113
rect 9706 2053 9718 2087
rect 9752 2053 9764 2087
rect 9706 2027 9764 2053
rect 9806 2087 9864 2113
rect 9806 2053 9818 2087
rect 9852 2053 9864 2087
rect 9806 2027 9864 2053
rect 9906 2087 9964 2113
rect 9906 2053 9918 2087
rect 9952 2053 9964 2087
rect 9906 2027 9964 2053
rect 10006 2087 10064 2113
rect 10006 2053 10018 2087
rect 10052 2053 10064 2087
rect 10006 2027 10064 2053
rect 10106 2087 10164 2113
rect 10106 2053 10118 2087
rect 10152 2053 10164 2087
rect 10106 2027 10164 2053
rect 10206 2087 10264 2113
rect 10206 2053 10218 2087
rect 10252 2053 10264 2087
rect 10206 2027 10264 2053
rect 10306 2087 10364 2113
rect 10306 2053 10318 2087
rect 10352 2053 10364 2087
rect 10306 2027 10364 2053
rect 10406 2087 10464 2113
rect 10406 2053 10418 2087
rect 10452 2053 10464 2087
rect 10406 2027 10464 2053
rect 10506 2087 10564 2113
rect 10506 2053 10518 2087
rect 10552 2053 10564 2087
rect 10506 2027 10564 2053
rect 10606 2087 10664 2113
rect 10606 2053 10618 2087
rect 10652 2053 10664 2087
rect 10606 2027 10664 2053
rect 10706 2087 10764 2113
rect 10706 2053 10718 2087
rect 10752 2053 10764 2087
rect 10706 2027 10764 2053
rect 10806 2087 10864 2113
rect 10806 2053 10818 2087
rect 10852 2053 10864 2087
rect 10806 2027 10864 2053
rect 10906 2087 10964 2113
rect 10906 2053 10918 2087
rect 10952 2053 10964 2087
rect 10906 2027 10964 2053
rect 11006 2087 11064 2113
rect 11006 2053 11018 2087
rect 11052 2053 11064 2087
rect 11006 2027 11064 2053
rect 11106 2087 11164 2113
rect 11106 2053 11118 2087
rect 11152 2053 11164 2087
rect 11106 2027 11164 2053
rect 11206 2087 11264 2113
rect 11206 2053 11212 2087
rect 11252 2053 11264 2087
rect 11206 2027 11264 2053
rect 11306 2087 11364 2113
rect 11306 2053 11318 2087
rect 11358 2053 11364 2087
rect 11306 2027 11364 2053
rect 11406 2087 11464 2113
rect 11406 2053 11412 2087
rect 11452 2053 11464 2087
rect 11406 2027 11464 2053
rect 11506 2087 11564 2113
rect 11506 2053 11518 2087
rect 11558 2053 11564 2087
rect 11506 2027 11564 2053
rect 11606 2087 11664 2113
rect 11606 2053 11618 2087
rect 11652 2053 11664 2087
rect 11606 2027 11664 2053
rect 11706 2087 11764 2113
rect 11706 2053 11718 2087
rect 11752 2053 11764 2087
rect 11706 2027 11764 2053
rect 11806 2087 11864 2113
rect 11806 2053 11818 2087
rect 11852 2053 11864 2087
rect 11806 2027 11864 2053
rect 11906 2087 11964 2113
rect 11906 2053 11918 2087
rect 11952 2053 11964 2087
rect 11906 2027 11964 2053
rect 12006 2087 12064 2113
rect 12006 2053 12018 2087
rect 12052 2053 12064 2087
rect 12006 2027 12064 2053
rect 12106 2087 12164 2113
rect 12106 2053 12118 2087
rect 12152 2053 12164 2087
rect 12106 2027 12164 2053
rect 12206 2087 12264 2113
rect 12206 2053 12218 2087
rect 12252 2053 12264 2087
rect 12206 2027 12264 2053
rect 12306 2087 12364 2113
rect 12306 2053 12318 2087
rect 12352 2053 12364 2087
rect 12306 2027 12364 2053
rect 12406 2087 12464 2113
rect 12406 2053 12418 2087
rect 12452 2053 12464 2087
rect 12406 2027 12464 2053
rect 12506 2087 12564 2113
rect 12506 2053 12518 2087
rect 12552 2053 12564 2087
rect 12506 2027 12564 2053
rect 12606 2087 12664 2113
rect 12606 2053 12612 2087
rect 12652 2053 12664 2087
rect 12606 2027 12664 2053
rect 12706 2087 12764 2113
rect 12706 2053 12718 2087
rect 12758 2053 12764 2087
rect 12706 2027 12764 2053
rect 12806 2087 12864 2113
rect 13018 2106 13262 2140
rect 12806 2053 12812 2087
rect 12852 2053 12864 2087
rect 12908 2068 12916 2102
rect 12958 2068 12974 2102
rect 13018 2087 13052 2106
rect 12806 2027 12864 2053
rect 13228 2103 13262 2106
rect 13228 2087 13362 2103
rect 13018 2037 13052 2053
rect 13096 2038 13112 2072
rect 13154 2038 13162 2072
rect 13262 2053 13328 2087
rect 13228 2037 13362 2053
rect 13428 2087 13462 2103
rect 13428 2037 13462 2053
rect 13528 2087 13662 2103
rect 13562 2053 13628 2087
rect 13528 2037 13662 2053
rect 6 1947 64 1973
rect 6 1913 18 1947
rect 52 1913 64 1947
rect 6 1887 64 1913
rect 106 1947 164 1973
rect 106 1913 118 1947
rect 152 1913 164 1947
rect 106 1887 164 1913
rect 206 1947 264 1973
rect 206 1913 218 1947
rect 252 1913 264 1947
rect 206 1887 264 1913
rect 306 1947 364 1973
rect 306 1913 318 1947
rect 352 1913 364 1947
rect 306 1887 364 1913
rect 406 1947 464 1973
rect 406 1913 418 1947
rect 452 1913 464 1947
rect 406 1887 464 1913
rect 506 1947 564 1973
rect 506 1913 518 1947
rect 552 1913 564 1947
rect 506 1887 564 1913
rect 606 1947 664 1973
rect 606 1913 618 1947
rect 652 1913 664 1947
rect 606 1887 664 1913
rect 706 1947 764 1973
rect 706 1913 718 1947
rect 752 1913 764 1947
rect 706 1887 764 1913
rect 806 1947 864 1973
rect 806 1913 818 1947
rect 852 1913 864 1947
rect 806 1887 864 1913
rect 906 1947 964 1973
rect 906 1913 912 1947
rect 952 1913 964 1947
rect 906 1887 964 1913
rect 1006 1947 1064 1973
rect 1006 1913 1018 1947
rect 1058 1913 1064 1947
rect 1006 1887 1064 1913
rect 1106 1947 1164 1973
rect 1106 1913 1118 1947
rect 1152 1913 1164 1947
rect 1106 1887 1164 1913
rect 1206 1947 1264 1973
rect 1206 1913 1218 1947
rect 1252 1913 1264 1947
rect 1206 1887 1264 1913
rect 1306 1947 1364 1973
rect 1306 1913 1318 1947
rect 1352 1913 1364 1947
rect 1306 1887 1364 1913
rect 1406 1947 1464 1973
rect 1406 1913 1418 1947
rect 1452 1913 1464 1947
rect 1406 1887 1464 1913
rect 1506 1947 1564 1973
rect 1506 1913 1512 1947
rect 1552 1913 1564 1947
rect 1506 1887 1564 1913
rect 1606 1947 1664 1973
rect 1606 1913 1618 1947
rect 1658 1913 1664 1947
rect 1606 1887 1664 1913
rect 1706 1947 1764 1973
rect 1706 1913 1718 1947
rect 1752 1913 1764 1947
rect 1706 1887 1764 1913
rect 1806 1947 1864 1973
rect 1806 1913 1818 1947
rect 1852 1913 1864 1947
rect 1806 1887 1864 1913
rect 1906 1947 1964 1973
rect 1906 1913 1918 1947
rect 1952 1913 1964 1947
rect 1906 1887 1964 1913
rect 2006 1947 2064 1973
rect 2006 1913 2018 1947
rect 2052 1913 2064 1947
rect 2006 1887 2064 1913
rect 2106 1947 2164 1973
rect 2106 1913 2118 1947
rect 2152 1913 2164 1947
rect 2106 1887 2164 1913
rect 2206 1947 2264 1973
rect 2206 1913 2218 1947
rect 2252 1913 2264 1947
rect 2206 1887 2264 1913
rect 2306 1947 2364 1973
rect 2306 1913 2318 1947
rect 2352 1913 2364 1947
rect 2306 1887 2364 1913
rect 2406 1947 2464 1973
rect 2406 1913 2418 1947
rect 2452 1913 2464 1947
rect 2406 1887 2464 1913
rect 2506 1947 2564 1973
rect 2506 1913 2518 1947
rect 2552 1913 2564 1947
rect 2506 1887 2564 1913
rect 2606 1947 2664 1973
rect 2606 1913 2618 1947
rect 2652 1913 2664 1947
rect 2606 1887 2664 1913
rect 2706 1947 2764 1973
rect 2706 1913 2718 1947
rect 2752 1913 2764 1947
rect 2706 1887 2764 1913
rect 2806 1947 2864 1973
rect 2806 1913 2818 1947
rect 2852 1913 2864 1947
rect 2806 1887 2864 1913
rect 2906 1947 2964 1973
rect 2906 1913 2918 1947
rect 2952 1913 2964 1947
rect 2906 1887 2964 1913
rect 3006 1947 3064 1973
rect 3006 1913 3018 1947
rect 3052 1913 3064 1947
rect 3006 1887 3064 1913
rect 3106 1947 3164 1973
rect 3106 1913 3118 1947
rect 3152 1913 3164 1947
rect 3106 1887 3164 1913
rect 3206 1947 3264 1973
rect 3206 1913 3218 1947
rect 3252 1913 3264 1947
rect 3206 1887 3264 1913
rect 3306 1947 3364 1973
rect 3306 1913 3318 1947
rect 3352 1913 3364 1947
rect 3306 1887 3364 1913
rect 3406 1947 3464 1973
rect 3406 1913 3418 1947
rect 3452 1913 3464 1947
rect 3406 1887 3464 1913
rect 3506 1947 3564 1973
rect 3506 1913 3518 1947
rect 3552 1913 3564 1947
rect 3506 1887 3564 1913
rect 3606 1947 3664 1973
rect 3606 1913 3612 1947
rect 3652 1913 3664 1947
rect 3606 1887 3664 1913
rect 3706 1947 3764 1973
rect 3706 1913 3718 1947
rect 3758 1913 3764 1947
rect 3706 1887 3764 1913
rect 3806 1947 3864 1973
rect 3806 1913 3818 1947
rect 3852 1913 3864 1947
rect 3806 1887 3864 1913
rect 3906 1947 3964 1973
rect 3906 1913 3918 1947
rect 3952 1913 3964 1947
rect 3906 1887 3964 1913
rect 4006 1947 4064 1973
rect 4006 1913 4018 1947
rect 4052 1913 4064 1947
rect 4006 1887 4064 1913
rect 4106 1947 4164 1973
rect 4106 1913 4118 1947
rect 4152 1913 4164 1947
rect 4106 1887 4164 1913
rect 4206 1947 4264 1973
rect 4206 1913 4212 1947
rect 4252 1913 4264 1947
rect 4206 1887 4264 1913
rect 4306 1947 4364 1973
rect 4306 1913 4318 1947
rect 4358 1913 4364 1947
rect 4306 1887 4364 1913
rect 4406 1947 4464 1973
rect 4406 1913 4412 1947
rect 4452 1913 4464 1947
rect 4406 1887 4464 1913
rect 4506 1947 4564 1973
rect 4506 1913 4518 1947
rect 4558 1913 4564 1947
rect 4506 1887 4564 1913
rect 4606 1947 4664 1973
rect 4606 1913 4612 1947
rect 4652 1913 4664 1947
rect 4606 1887 4664 1913
rect 4706 1947 4764 1973
rect 4706 1913 4718 1947
rect 4758 1913 4764 1947
rect 4706 1887 4764 1913
rect 4806 1947 4864 1973
rect 4806 1913 4818 1947
rect 4852 1913 4864 1947
rect 4806 1887 4864 1913
rect 4906 1947 4964 1973
rect 4906 1913 4918 1947
rect 4952 1913 4964 1947
rect 4906 1887 4964 1913
rect 5006 1947 5064 1973
rect 5006 1913 5018 1947
rect 5052 1913 5064 1947
rect 5006 1887 5064 1913
rect 5106 1947 5164 1973
rect 5106 1913 5112 1947
rect 5152 1913 5164 1947
rect 5106 1887 5164 1913
rect 5206 1947 5264 1973
rect 5206 1913 5218 1947
rect 5258 1913 5264 1947
rect 5206 1887 5264 1913
rect 5306 1947 5364 1973
rect 5306 1913 5318 1947
rect 5352 1913 5364 1947
rect 5306 1887 5364 1913
rect 5406 1947 5464 1973
rect 5406 1913 5418 1947
rect 5452 1913 5464 1947
rect 5406 1887 5464 1913
rect 5506 1947 5564 1973
rect 5506 1913 5518 1947
rect 5552 1913 5564 1947
rect 5506 1887 5564 1913
rect 5606 1947 5664 1973
rect 5606 1913 5618 1947
rect 5652 1913 5664 1947
rect 5606 1887 5664 1913
rect 5706 1947 5764 1973
rect 5706 1913 5712 1947
rect 5752 1913 5764 1947
rect 5706 1887 5764 1913
rect 5806 1947 5864 1973
rect 5806 1913 5818 1947
rect 5858 1913 5864 1947
rect 5806 1887 5864 1913
rect 5906 1947 5964 1973
rect 5906 1913 5918 1947
rect 5952 1913 5964 1947
rect 5906 1887 5964 1913
rect 6006 1947 6064 1973
rect 6006 1913 6018 1947
rect 6052 1913 6064 1947
rect 6006 1887 6064 1913
rect 6106 1947 6164 1973
rect 6106 1913 6118 1947
rect 6152 1913 6164 1947
rect 6106 1887 6164 1913
rect 6206 1947 6264 1973
rect 6206 1913 6218 1947
rect 6252 1913 6264 1947
rect 6206 1887 6264 1913
rect 6306 1947 6364 1973
rect 6306 1913 6318 1947
rect 6352 1913 6364 1947
rect 6306 1887 6364 1913
rect 6406 1947 6464 1973
rect 6406 1913 6418 1947
rect 6452 1913 6464 1947
rect 6406 1887 6464 1913
rect 6506 1947 6564 1973
rect 6506 1913 6518 1947
rect 6552 1913 6564 1947
rect 6506 1887 6564 1913
rect 6606 1947 6664 1973
rect 6606 1913 6618 1947
rect 6652 1913 6664 1947
rect 6606 1887 6664 1913
rect 6706 1947 6764 1973
rect 6706 1913 6712 1947
rect 6752 1913 6764 1947
rect 6706 1887 6764 1913
rect 6806 1947 6864 1973
rect 6806 1913 6818 1947
rect 6858 1913 6864 1947
rect 6806 1887 6864 1913
rect 6906 1947 6964 1973
rect 6906 1913 6912 1947
rect 6952 1913 6964 1947
rect 6906 1887 6964 1913
rect 7006 1947 7064 1973
rect 7006 1913 7018 1947
rect 7058 1913 7064 1947
rect 7006 1887 7064 1913
rect 7106 1947 7164 1973
rect 7106 1913 7118 1947
rect 7152 1913 7164 1947
rect 7106 1887 7164 1913
rect 7206 1947 7264 1973
rect 7206 1913 7218 1947
rect 7252 1913 7264 1947
rect 7206 1887 7264 1913
rect 7306 1947 7364 1973
rect 7306 1913 7318 1947
rect 7352 1913 7364 1947
rect 7306 1887 7364 1913
rect 7406 1947 7464 1973
rect 7406 1913 7418 1947
rect 7452 1913 7464 1947
rect 7406 1887 7464 1913
rect 7506 1947 7564 1973
rect 7506 1913 7518 1947
rect 7552 1913 7564 1947
rect 7506 1887 7564 1913
rect 7606 1947 7664 1973
rect 7606 1913 7618 1947
rect 7652 1913 7664 1947
rect 7606 1887 7664 1913
rect 7706 1947 7764 1973
rect 7706 1913 7718 1947
rect 7752 1913 7764 1947
rect 7706 1887 7764 1913
rect 7806 1947 7864 1973
rect 7806 1913 7818 1947
rect 7852 1913 7864 1947
rect 7806 1887 7864 1913
rect 7906 1947 7964 1973
rect 7906 1913 7918 1947
rect 7952 1913 7964 1947
rect 7906 1887 7964 1913
rect 8006 1947 8064 1973
rect 8006 1913 8018 1947
rect 8052 1913 8064 1947
rect 8006 1887 8064 1913
rect 8106 1947 8164 1973
rect 8106 1913 8118 1947
rect 8152 1913 8164 1947
rect 8106 1887 8164 1913
rect 8206 1947 8264 1973
rect 8206 1913 8218 1947
rect 8252 1913 8264 1947
rect 8206 1887 8264 1913
rect 8306 1947 8364 1973
rect 8306 1913 8318 1947
rect 8352 1913 8364 1947
rect 8306 1887 8364 1913
rect 8406 1947 8464 1973
rect 8406 1913 8418 1947
rect 8452 1913 8464 1947
rect 8406 1887 8464 1913
rect 8506 1947 8564 1973
rect 8506 1913 8518 1947
rect 8552 1913 8564 1947
rect 8506 1887 8564 1913
rect 8606 1947 8664 1973
rect 8606 1913 8618 1947
rect 8652 1913 8664 1947
rect 8606 1887 8664 1913
rect 8706 1947 8764 1973
rect 8706 1913 8718 1947
rect 8752 1913 8764 1947
rect 8706 1887 8764 1913
rect 8806 1947 8864 1973
rect 8806 1913 8818 1947
rect 8852 1913 8864 1947
rect 8806 1887 8864 1913
rect 8906 1947 8964 1973
rect 8906 1913 8918 1947
rect 8952 1913 8964 1947
rect 8906 1887 8964 1913
rect 9006 1947 9064 1973
rect 9006 1913 9018 1947
rect 9052 1913 9064 1947
rect 9006 1887 9064 1913
rect 9106 1947 9164 1973
rect 9106 1913 9118 1947
rect 9152 1913 9164 1947
rect 9106 1887 9164 1913
rect 9206 1947 9264 1973
rect 9206 1913 9218 1947
rect 9252 1913 9264 1947
rect 9206 1887 9264 1913
rect 9306 1947 9364 1973
rect 9306 1913 9318 1947
rect 9352 1913 9364 1947
rect 9306 1887 9364 1913
rect 9406 1947 9464 1973
rect 9406 1913 9418 1947
rect 9452 1913 9464 1947
rect 9406 1887 9464 1913
rect 9506 1947 9564 1973
rect 9506 1913 9518 1947
rect 9552 1913 9564 1947
rect 9506 1887 9564 1913
rect 9606 1947 9664 1973
rect 9606 1913 9618 1947
rect 9652 1913 9664 1947
rect 9606 1887 9664 1913
rect 9706 1947 9764 1973
rect 9706 1913 9718 1947
rect 9752 1913 9764 1947
rect 9706 1887 9764 1913
rect 9806 1947 9864 1973
rect 9806 1913 9818 1947
rect 9852 1913 9864 1947
rect 9806 1887 9864 1913
rect 9906 1947 9964 1973
rect 9906 1913 9918 1947
rect 9952 1913 9964 1947
rect 9906 1887 9964 1913
rect 10006 1947 10064 1973
rect 10006 1913 10018 1947
rect 10052 1913 10064 1947
rect 10006 1887 10064 1913
rect 10106 1947 10164 1973
rect 10106 1913 10118 1947
rect 10152 1913 10164 1947
rect 10106 1887 10164 1913
rect 10206 1947 10264 1973
rect 10206 1913 10218 1947
rect 10252 1913 10264 1947
rect 10206 1887 10264 1913
rect 10306 1947 10364 1973
rect 10306 1913 10318 1947
rect 10352 1913 10364 1947
rect 10306 1887 10364 1913
rect 10406 1947 10464 1973
rect 10406 1913 10418 1947
rect 10452 1913 10464 1947
rect 10406 1887 10464 1913
rect 10506 1947 10564 1973
rect 10506 1913 10518 1947
rect 10552 1913 10564 1947
rect 10506 1887 10564 1913
rect 10606 1947 10664 1973
rect 10606 1913 10618 1947
rect 10652 1913 10664 1947
rect 10606 1887 10664 1913
rect 10706 1947 10764 1973
rect 10706 1913 10718 1947
rect 10752 1913 10764 1947
rect 10706 1887 10764 1913
rect 10806 1947 10864 1973
rect 10806 1913 10818 1947
rect 10852 1913 10864 1947
rect 10806 1887 10864 1913
rect 10906 1947 10964 1973
rect 10906 1913 10918 1947
rect 10952 1913 10964 1947
rect 10906 1887 10964 1913
rect 11006 1947 11064 1973
rect 11006 1913 11012 1947
rect 11052 1913 11064 1947
rect 11006 1887 11064 1913
rect 11106 1947 11164 1973
rect 11106 1913 11118 1947
rect 11158 1913 11164 1947
rect 11106 1887 11164 1913
rect 11206 1947 11264 1973
rect 11206 1913 11212 1947
rect 11252 1913 11264 1947
rect 11206 1887 11264 1913
rect 11306 1947 11364 1973
rect 11306 1913 11318 1947
rect 11358 1913 11364 1947
rect 11306 1887 11364 1913
rect 11406 1947 11464 1973
rect 11406 1913 11418 1947
rect 11452 1913 11464 1947
rect 11406 1887 11464 1913
rect 11506 1947 11564 1973
rect 11506 1913 11518 1947
rect 11552 1913 11564 1947
rect 11506 1887 11564 1913
rect 11606 1947 11664 1973
rect 11606 1913 11618 1947
rect 11652 1913 11664 1947
rect 11606 1887 11664 1913
rect 11706 1947 11764 1973
rect 11706 1913 11718 1947
rect 11752 1913 11764 1947
rect 11706 1887 11764 1913
rect 11806 1947 11864 1973
rect 11806 1913 11818 1947
rect 11852 1913 11864 1947
rect 11806 1887 11864 1913
rect 11906 1947 11964 1973
rect 11906 1913 11918 1947
rect 11952 1913 11964 1947
rect 11906 1887 11964 1913
rect 12006 1947 12064 1973
rect 12006 1913 12018 1947
rect 12052 1913 12064 1947
rect 12006 1887 12064 1913
rect 12106 1947 12164 1973
rect 12106 1913 12118 1947
rect 12152 1913 12164 1947
rect 12106 1887 12164 1913
rect 12206 1947 12264 1973
rect 12206 1913 12218 1947
rect 12252 1913 12264 1947
rect 12206 1887 12264 1913
rect 12306 1947 12364 1973
rect 12306 1913 12318 1947
rect 12352 1913 12364 1947
rect 12306 1887 12364 1913
rect 12406 1947 12464 1973
rect 12406 1913 12418 1947
rect 12452 1913 12464 1947
rect 12406 1887 12464 1913
rect 12506 1947 12564 1973
rect 12506 1913 12518 1947
rect 12552 1913 12564 1947
rect 12506 1887 12564 1913
rect 12606 1947 12664 1973
rect 12606 1913 12612 1947
rect 12652 1913 12664 1947
rect 12606 1887 12664 1913
rect 12706 1947 12764 1973
rect 12706 1913 12718 1947
rect 12758 1913 12764 1947
rect 12706 1887 12764 1913
rect 12806 1947 12864 1973
rect 13018 1966 13262 2000
rect 12806 1913 12812 1947
rect 12852 1913 12864 1947
rect 12908 1928 12916 1962
rect 12958 1928 12974 1962
rect 13018 1947 13052 1966
rect 12806 1887 12864 1913
rect 13228 1947 13262 1966
rect 13018 1897 13052 1913
rect 13096 1898 13112 1932
rect 13154 1898 13162 1932
rect 13228 1897 13262 1913
rect 13328 1947 13462 1963
rect 13362 1913 13428 1947
rect 13328 1897 13462 1913
rect 13528 1947 13662 1963
rect 13562 1913 13628 1947
rect 13528 1897 13662 1913
rect 6 1807 64 1833
rect 6 1773 18 1807
rect 52 1773 64 1807
rect 6 1747 64 1773
rect 106 1807 164 1833
rect 106 1773 118 1807
rect 152 1773 164 1807
rect 106 1747 164 1773
rect 206 1807 264 1833
rect 206 1773 218 1807
rect 252 1773 264 1807
rect 206 1747 264 1773
rect 306 1807 364 1833
rect 306 1773 318 1807
rect 352 1773 364 1807
rect 306 1747 364 1773
rect 406 1807 464 1833
rect 406 1773 418 1807
rect 452 1773 464 1807
rect 406 1747 464 1773
rect 506 1807 564 1833
rect 506 1773 518 1807
rect 552 1773 564 1807
rect 506 1747 564 1773
rect 606 1807 664 1833
rect 606 1773 618 1807
rect 652 1773 664 1807
rect 606 1747 664 1773
rect 706 1807 764 1833
rect 706 1773 718 1807
rect 752 1773 764 1807
rect 706 1747 764 1773
rect 806 1807 864 1833
rect 806 1773 818 1807
rect 852 1773 864 1807
rect 806 1747 864 1773
rect 906 1807 964 1833
rect 906 1773 918 1807
rect 952 1773 964 1807
rect 906 1747 964 1773
rect 1006 1807 1064 1833
rect 1006 1773 1018 1807
rect 1052 1773 1064 1807
rect 1006 1747 1064 1773
rect 1106 1807 1164 1833
rect 1106 1773 1118 1807
rect 1152 1773 1164 1807
rect 1106 1747 1164 1773
rect 1206 1807 1264 1833
rect 1206 1773 1218 1807
rect 1252 1773 1264 1807
rect 1206 1747 1264 1773
rect 1306 1807 1364 1833
rect 1306 1773 1318 1807
rect 1352 1773 1364 1807
rect 1306 1747 1364 1773
rect 1406 1807 1464 1833
rect 1406 1773 1418 1807
rect 1452 1773 1464 1807
rect 1406 1747 1464 1773
rect 1506 1807 1564 1833
rect 1506 1773 1518 1807
rect 1552 1773 1564 1807
rect 1506 1747 1564 1773
rect 1606 1807 1664 1833
rect 1606 1773 1618 1807
rect 1652 1773 1664 1807
rect 1606 1747 1664 1773
rect 1706 1807 1764 1833
rect 1706 1773 1718 1807
rect 1752 1773 1764 1807
rect 1706 1747 1764 1773
rect 1806 1807 1864 1833
rect 1806 1773 1818 1807
rect 1852 1773 1864 1807
rect 1806 1747 1864 1773
rect 1906 1807 1964 1833
rect 1906 1773 1918 1807
rect 1952 1773 1964 1807
rect 1906 1747 1964 1773
rect 2006 1807 2064 1833
rect 2006 1773 2018 1807
rect 2052 1773 2064 1807
rect 2006 1747 2064 1773
rect 2106 1807 2164 1833
rect 2106 1773 2118 1807
rect 2152 1773 2164 1807
rect 2106 1747 2164 1773
rect 2206 1807 2264 1833
rect 2206 1773 2218 1807
rect 2252 1773 2264 1807
rect 2206 1747 2264 1773
rect 2306 1807 2364 1833
rect 2306 1773 2318 1807
rect 2352 1773 2364 1807
rect 2306 1747 2364 1773
rect 2406 1807 2464 1833
rect 2406 1773 2418 1807
rect 2452 1773 2464 1807
rect 2406 1747 2464 1773
rect 2506 1807 2564 1833
rect 2506 1773 2518 1807
rect 2552 1773 2564 1807
rect 2506 1747 2564 1773
rect 2606 1807 2664 1833
rect 2606 1773 2618 1807
rect 2652 1773 2664 1807
rect 2606 1747 2664 1773
rect 2706 1807 2764 1833
rect 2706 1773 2718 1807
rect 2752 1773 2764 1807
rect 2706 1747 2764 1773
rect 2806 1807 2864 1833
rect 2806 1773 2818 1807
rect 2852 1773 2864 1807
rect 2806 1747 2864 1773
rect 2906 1807 2964 1833
rect 2906 1773 2918 1807
rect 2952 1773 2964 1807
rect 2906 1747 2964 1773
rect 3006 1807 3064 1833
rect 3006 1773 3018 1807
rect 3052 1773 3064 1807
rect 3006 1747 3064 1773
rect 3106 1807 3164 1833
rect 3106 1773 3112 1807
rect 3152 1773 3164 1807
rect 3106 1747 3164 1773
rect 3206 1807 3264 1833
rect 3206 1773 3218 1807
rect 3258 1773 3264 1807
rect 3206 1747 3264 1773
rect 3306 1807 3364 1833
rect 3306 1773 3312 1807
rect 3352 1773 3364 1807
rect 3306 1747 3364 1773
rect 3406 1807 3464 1833
rect 3406 1773 3418 1807
rect 3458 1773 3464 1807
rect 3406 1747 3464 1773
rect 3506 1807 3564 1833
rect 3506 1773 3518 1807
rect 3552 1773 3564 1807
rect 3506 1747 3564 1773
rect 3606 1807 3664 1833
rect 3606 1773 3618 1807
rect 3652 1773 3664 1807
rect 3606 1747 3664 1773
rect 3706 1807 3764 1833
rect 3706 1773 3718 1807
rect 3752 1773 3764 1807
rect 3706 1747 3764 1773
rect 3806 1807 3864 1833
rect 3806 1773 3818 1807
rect 3852 1773 3864 1807
rect 3806 1747 3864 1773
rect 3906 1807 3964 1833
rect 3906 1773 3912 1807
rect 3952 1773 3964 1807
rect 3906 1747 3964 1773
rect 4006 1807 4064 1833
rect 4006 1773 4018 1807
rect 4058 1773 4064 1807
rect 4006 1747 4064 1773
rect 4106 1807 4164 1833
rect 4106 1773 4112 1807
rect 4152 1773 4164 1807
rect 4106 1747 4164 1773
rect 4206 1807 4264 1833
rect 4206 1773 4218 1807
rect 4258 1773 4264 1807
rect 4206 1747 4264 1773
rect 4306 1807 4364 1833
rect 4306 1773 4318 1807
rect 4352 1773 4364 1807
rect 4306 1747 4364 1773
rect 4406 1807 4464 1833
rect 4406 1773 4418 1807
rect 4452 1773 4464 1807
rect 4406 1747 4464 1773
rect 4506 1807 4564 1833
rect 4506 1773 4518 1807
rect 4552 1773 4564 1807
rect 4506 1747 4564 1773
rect 4606 1807 4664 1833
rect 4606 1773 4618 1807
rect 4652 1773 4664 1807
rect 4606 1747 4664 1773
rect 4706 1807 4764 1833
rect 4706 1773 4718 1807
rect 4752 1773 4764 1807
rect 4706 1747 4764 1773
rect 4806 1807 4864 1833
rect 4806 1773 4812 1807
rect 4852 1773 4864 1807
rect 4806 1747 4864 1773
rect 4906 1807 4964 1833
rect 4906 1773 4918 1807
rect 4958 1773 4964 1807
rect 4906 1747 4964 1773
rect 5006 1807 5064 1833
rect 5006 1773 5018 1807
rect 5052 1773 5064 1807
rect 5006 1747 5064 1773
rect 5106 1807 5164 1833
rect 5106 1773 5118 1807
rect 5152 1773 5164 1807
rect 5106 1747 5164 1773
rect 5206 1807 5264 1833
rect 5206 1773 5218 1807
rect 5252 1773 5264 1807
rect 5206 1747 5264 1773
rect 5306 1807 5364 1833
rect 5306 1773 5318 1807
rect 5352 1773 5364 1807
rect 5306 1747 5364 1773
rect 5406 1807 5464 1833
rect 5406 1773 5418 1807
rect 5452 1773 5464 1807
rect 5406 1747 5464 1773
rect 5506 1807 5564 1833
rect 5506 1773 5518 1807
rect 5552 1773 5564 1807
rect 5506 1747 5564 1773
rect 5606 1807 5664 1833
rect 5606 1773 5618 1807
rect 5652 1773 5664 1807
rect 5606 1747 5664 1773
rect 5706 1807 5764 1833
rect 5706 1773 5718 1807
rect 5752 1773 5764 1807
rect 5706 1747 5764 1773
rect 5806 1807 5864 1833
rect 5806 1773 5818 1807
rect 5852 1773 5864 1807
rect 5806 1747 5864 1773
rect 5906 1807 5964 1833
rect 5906 1773 5918 1807
rect 5952 1773 5964 1807
rect 5906 1747 5964 1773
rect 6006 1807 6064 1833
rect 6006 1773 6018 1807
rect 6052 1773 6064 1807
rect 6006 1747 6064 1773
rect 6106 1807 6164 1833
rect 6106 1773 6118 1807
rect 6152 1773 6164 1807
rect 6106 1747 6164 1773
rect 6206 1807 6264 1833
rect 6206 1773 6218 1807
rect 6252 1773 6264 1807
rect 6206 1747 6264 1773
rect 6306 1807 6364 1833
rect 6306 1773 6312 1807
rect 6352 1773 6364 1807
rect 6306 1747 6364 1773
rect 6406 1807 6464 1833
rect 6406 1773 6418 1807
rect 6458 1773 6464 1807
rect 6406 1747 6464 1773
rect 6506 1807 6564 1833
rect 6506 1773 6518 1807
rect 6552 1773 6564 1807
rect 6506 1747 6564 1773
rect 6606 1807 6664 1833
rect 6606 1773 6618 1807
rect 6652 1773 6664 1807
rect 6606 1747 6664 1773
rect 6706 1807 6764 1833
rect 6706 1773 6718 1807
rect 6752 1773 6764 1807
rect 6706 1747 6764 1773
rect 6806 1807 6864 1833
rect 6806 1773 6818 1807
rect 6852 1773 6864 1807
rect 6806 1747 6864 1773
rect 6906 1807 6964 1833
rect 6906 1773 6918 1807
rect 6952 1773 6964 1807
rect 6906 1747 6964 1773
rect 7006 1807 7064 1833
rect 7006 1773 7018 1807
rect 7052 1773 7064 1807
rect 7006 1747 7064 1773
rect 7106 1807 7164 1833
rect 7106 1773 7112 1807
rect 7152 1773 7164 1807
rect 7106 1747 7164 1773
rect 7206 1807 7264 1833
rect 7206 1773 7218 1807
rect 7258 1773 7264 1807
rect 7206 1747 7264 1773
rect 7306 1807 7364 1833
rect 7306 1773 7318 1807
rect 7352 1773 7364 1807
rect 7306 1747 7364 1773
rect 7406 1807 7464 1833
rect 7406 1773 7412 1807
rect 7452 1773 7464 1807
rect 7406 1747 7464 1773
rect 7506 1807 7564 1833
rect 7506 1773 7518 1807
rect 7558 1773 7564 1807
rect 7506 1747 7564 1773
rect 7606 1807 7664 1833
rect 7606 1773 7618 1807
rect 7652 1773 7664 1807
rect 7606 1747 7664 1773
rect 7706 1807 7764 1833
rect 7706 1773 7712 1807
rect 7752 1773 7764 1807
rect 7706 1747 7764 1773
rect 7806 1807 7864 1833
rect 7806 1773 7818 1807
rect 7858 1773 7864 1807
rect 7806 1747 7864 1773
rect 7906 1807 7964 1833
rect 7906 1773 7918 1807
rect 7952 1773 7964 1807
rect 7906 1747 7964 1773
rect 8006 1807 8064 1833
rect 8006 1773 8012 1807
rect 8052 1773 8064 1807
rect 8006 1747 8064 1773
rect 8106 1807 8164 1833
rect 8106 1773 8118 1807
rect 8158 1773 8164 1807
rect 8106 1747 8164 1773
rect 8206 1807 8264 1833
rect 8206 1773 8218 1807
rect 8252 1773 8264 1807
rect 8206 1747 8264 1773
rect 8306 1807 8364 1833
rect 8306 1773 8318 1807
rect 8352 1773 8364 1807
rect 8306 1747 8364 1773
rect 8406 1807 8464 1833
rect 8406 1773 8418 1807
rect 8452 1773 8464 1807
rect 8406 1747 8464 1773
rect 8506 1807 8564 1833
rect 8506 1773 8518 1807
rect 8552 1773 8564 1807
rect 8506 1747 8564 1773
rect 8606 1807 8664 1833
rect 8606 1773 8612 1807
rect 8652 1773 8664 1807
rect 8606 1747 8664 1773
rect 8706 1807 8764 1833
rect 8706 1773 8718 1807
rect 8758 1773 8764 1807
rect 8706 1747 8764 1773
rect 8806 1807 8864 1833
rect 8806 1773 8818 1807
rect 8852 1773 8864 1807
rect 8806 1747 8864 1773
rect 8906 1807 8964 1833
rect 8906 1773 8918 1807
rect 8952 1773 8964 1807
rect 8906 1747 8964 1773
rect 9006 1807 9064 1833
rect 9006 1773 9018 1807
rect 9052 1773 9064 1807
rect 9006 1747 9064 1773
rect 9106 1807 9164 1833
rect 9106 1773 9118 1807
rect 9152 1773 9164 1807
rect 9106 1747 9164 1773
rect 9206 1807 9264 1833
rect 9206 1773 9218 1807
rect 9252 1773 9264 1807
rect 9206 1747 9264 1773
rect 9306 1807 9364 1833
rect 9306 1773 9318 1807
rect 9352 1773 9364 1807
rect 9306 1747 9364 1773
rect 9406 1807 9464 1833
rect 9406 1773 9418 1807
rect 9452 1773 9464 1807
rect 9406 1747 9464 1773
rect 9506 1807 9564 1833
rect 9506 1773 9518 1807
rect 9552 1773 9564 1807
rect 9506 1747 9564 1773
rect 9606 1807 9664 1833
rect 9606 1773 9618 1807
rect 9652 1773 9664 1807
rect 9606 1747 9664 1773
rect 9706 1807 9764 1833
rect 9706 1773 9718 1807
rect 9752 1773 9764 1807
rect 9706 1747 9764 1773
rect 9806 1807 9864 1833
rect 9806 1773 9812 1807
rect 9852 1773 9864 1807
rect 9806 1747 9864 1773
rect 9906 1807 9964 1833
rect 9906 1773 9918 1807
rect 9958 1773 9964 1807
rect 9906 1747 9964 1773
rect 10006 1807 10064 1833
rect 10006 1773 10012 1807
rect 10052 1773 10064 1807
rect 10006 1747 10064 1773
rect 10106 1807 10164 1833
rect 10106 1773 10118 1807
rect 10158 1773 10164 1807
rect 10106 1747 10164 1773
rect 10206 1807 10264 1833
rect 10206 1773 10212 1807
rect 10252 1773 10264 1807
rect 10206 1747 10264 1773
rect 10306 1807 10364 1833
rect 10306 1773 10318 1807
rect 10358 1773 10364 1807
rect 10306 1747 10364 1773
rect 10406 1807 10464 1833
rect 10406 1773 10412 1807
rect 10452 1773 10464 1807
rect 10406 1747 10464 1773
rect 10506 1807 10564 1833
rect 10506 1773 10518 1807
rect 10558 1773 10564 1807
rect 10506 1747 10564 1773
rect 10606 1807 10664 1833
rect 10606 1773 10618 1807
rect 10652 1773 10664 1807
rect 10606 1747 10664 1773
rect 10706 1807 10764 1833
rect 10706 1773 10712 1807
rect 10752 1773 10764 1807
rect 10706 1747 10764 1773
rect 10806 1807 10864 1833
rect 10806 1773 10818 1807
rect 10858 1773 10864 1807
rect 10806 1747 10864 1773
rect 10906 1807 10964 1833
rect 10906 1773 10918 1807
rect 10952 1773 10964 1807
rect 10906 1747 10964 1773
rect 11006 1807 11064 1833
rect 11006 1773 11018 1807
rect 11052 1773 11064 1807
rect 11006 1747 11064 1773
rect 11106 1807 11164 1833
rect 11106 1773 11118 1807
rect 11152 1773 11164 1807
rect 11106 1747 11164 1773
rect 11206 1807 11264 1833
rect 11206 1773 11218 1807
rect 11252 1773 11264 1807
rect 11206 1747 11264 1773
rect 11306 1807 11364 1833
rect 11306 1773 11318 1807
rect 11352 1773 11364 1807
rect 11306 1747 11364 1773
rect 11406 1807 11464 1833
rect 11406 1773 11418 1807
rect 11452 1773 11464 1807
rect 11406 1747 11464 1773
rect 11506 1807 11564 1833
rect 11506 1773 11518 1807
rect 11552 1773 11564 1807
rect 11506 1747 11564 1773
rect 11606 1807 11664 1833
rect 11606 1773 11612 1807
rect 11652 1773 11664 1807
rect 11606 1747 11664 1773
rect 11706 1807 11764 1833
rect 11706 1773 11718 1807
rect 11758 1773 11764 1807
rect 11706 1747 11764 1773
rect 11806 1807 11864 1833
rect 11806 1773 11818 1807
rect 11852 1773 11864 1807
rect 11806 1747 11864 1773
rect 11906 1807 11964 1833
rect 11906 1773 11912 1807
rect 11952 1773 11964 1807
rect 11906 1747 11964 1773
rect 12006 1807 12064 1833
rect 12006 1773 12018 1807
rect 12058 1773 12064 1807
rect 12006 1747 12064 1773
rect 12106 1807 12164 1833
rect 12106 1773 12118 1807
rect 12152 1773 12164 1807
rect 12106 1747 12164 1773
rect 12206 1807 12264 1833
rect 12206 1773 12218 1807
rect 12252 1773 12264 1807
rect 12206 1747 12264 1773
rect 12306 1807 12364 1833
rect 12306 1773 12318 1807
rect 12352 1773 12364 1807
rect 12306 1747 12364 1773
rect 12406 1807 12464 1833
rect 12406 1773 12418 1807
rect 12452 1773 12464 1807
rect 12406 1747 12464 1773
rect 12506 1807 12564 1833
rect 12506 1773 12518 1807
rect 12552 1773 12564 1807
rect 12506 1747 12564 1773
rect 12606 1807 12664 1833
rect 12606 1773 12618 1807
rect 12652 1773 12664 1807
rect 12606 1747 12664 1773
rect 12706 1807 12764 1833
rect 12706 1773 12718 1807
rect 12752 1773 12764 1807
rect 12706 1747 12764 1773
rect 12806 1807 12864 1833
rect 13018 1826 13262 1860
rect 12806 1773 12812 1807
rect 12852 1773 12864 1807
rect 12908 1788 12916 1822
rect 12958 1788 12974 1822
rect 13018 1807 13052 1826
rect 12806 1747 12864 1773
rect 13228 1823 13262 1826
rect 13228 1807 13362 1823
rect 13018 1757 13052 1773
rect 13096 1758 13112 1792
rect 13154 1758 13162 1792
rect 13262 1773 13328 1807
rect 13228 1757 13362 1773
rect 13428 1807 13562 1823
rect 13462 1773 13528 1807
rect 13428 1757 13562 1773
rect 13628 1807 13662 1823
rect 13628 1757 13662 1773
rect 6 1667 64 1693
rect 6 1633 18 1667
rect 52 1633 64 1667
rect 6 1607 64 1633
rect 106 1667 164 1693
rect 106 1633 118 1667
rect 152 1633 164 1667
rect 106 1607 164 1633
rect 206 1667 264 1693
rect 206 1633 218 1667
rect 252 1633 264 1667
rect 206 1607 264 1633
rect 306 1667 364 1693
rect 306 1633 318 1667
rect 352 1633 364 1667
rect 306 1607 364 1633
rect 406 1667 464 1693
rect 406 1633 418 1667
rect 452 1633 464 1667
rect 406 1607 464 1633
rect 506 1667 564 1693
rect 506 1633 518 1667
rect 552 1633 564 1667
rect 506 1607 564 1633
rect 606 1667 664 1693
rect 606 1633 612 1667
rect 652 1633 664 1667
rect 606 1607 664 1633
rect 706 1667 764 1693
rect 706 1633 718 1667
rect 758 1633 764 1667
rect 706 1607 764 1633
rect 806 1667 864 1693
rect 806 1633 818 1667
rect 852 1633 864 1667
rect 806 1607 864 1633
rect 906 1667 964 1693
rect 906 1633 918 1667
rect 952 1633 964 1667
rect 906 1607 964 1633
rect 1006 1667 1064 1693
rect 1006 1633 1012 1667
rect 1052 1633 1064 1667
rect 1006 1607 1064 1633
rect 1106 1667 1164 1693
rect 1106 1633 1118 1667
rect 1158 1633 1164 1667
rect 1106 1607 1164 1633
rect 1206 1667 1264 1693
rect 1206 1633 1212 1667
rect 1252 1633 1264 1667
rect 1206 1607 1264 1633
rect 1306 1667 1364 1693
rect 1306 1633 1318 1667
rect 1358 1633 1364 1667
rect 1306 1607 1364 1633
rect 1406 1667 1464 1693
rect 1406 1633 1418 1667
rect 1452 1633 1464 1667
rect 1406 1607 1464 1633
rect 1506 1667 1564 1693
rect 1506 1633 1512 1667
rect 1552 1633 1564 1667
rect 1506 1607 1564 1633
rect 1606 1667 1664 1693
rect 1606 1633 1618 1667
rect 1658 1633 1664 1667
rect 1606 1607 1664 1633
rect 1706 1667 1764 1693
rect 1706 1633 1718 1667
rect 1752 1633 1764 1667
rect 1706 1607 1764 1633
rect 1806 1667 1864 1693
rect 1806 1633 1818 1667
rect 1852 1633 1864 1667
rect 1806 1607 1864 1633
rect 1906 1667 1964 1693
rect 1906 1633 1918 1667
rect 1952 1633 1964 1667
rect 1906 1607 1964 1633
rect 2006 1667 2064 1693
rect 2006 1633 2018 1667
rect 2052 1633 2064 1667
rect 2006 1607 2064 1633
rect 2106 1667 2164 1693
rect 2106 1633 2118 1667
rect 2152 1633 2164 1667
rect 2106 1607 2164 1633
rect 2206 1667 2264 1693
rect 2206 1633 2218 1667
rect 2252 1633 2264 1667
rect 2206 1607 2264 1633
rect 2306 1667 2364 1693
rect 2306 1633 2318 1667
rect 2352 1633 2364 1667
rect 2306 1607 2364 1633
rect 2406 1667 2464 1693
rect 2406 1633 2418 1667
rect 2452 1633 2464 1667
rect 2406 1607 2464 1633
rect 2506 1667 2564 1693
rect 2506 1633 2518 1667
rect 2552 1633 2564 1667
rect 2506 1607 2564 1633
rect 2606 1667 2664 1693
rect 2606 1633 2612 1667
rect 2652 1633 2664 1667
rect 2606 1607 2664 1633
rect 2706 1667 2764 1693
rect 2706 1633 2718 1667
rect 2758 1633 2764 1667
rect 2706 1607 2764 1633
rect 2806 1667 2864 1693
rect 2806 1633 2818 1667
rect 2852 1633 2864 1667
rect 2806 1607 2864 1633
rect 2906 1667 2964 1693
rect 2906 1633 2918 1667
rect 2952 1633 2964 1667
rect 2906 1607 2964 1633
rect 3006 1667 3064 1693
rect 3006 1633 3018 1667
rect 3052 1633 3064 1667
rect 3006 1607 3064 1633
rect 3106 1667 3164 1693
rect 3106 1633 3118 1667
rect 3152 1633 3164 1667
rect 3106 1607 3164 1633
rect 3206 1667 3264 1693
rect 3206 1633 3218 1667
rect 3252 1633 3264 1667
rect 3206 1607 3264 1633
rect 3306 1667 3364 1693
rect 3306 1633 3318 1667
rect 3352 1633 3364 1667
rect 3306 1607 3364 1633
rect 3406 1667 3464 1693
rect 3406 1633 3418 1667
rect 3452 1633 3464 1667
rect 3406 1607 3464 1633
rect 3506 1667 3564 1693
rect 3506 1633 3518 1667
rect 3552 1633 3564 1667
rect 3506 1607 3564 1633
rect 3606 1667 3664 1693
rect 3606 1633 3618 1667
rect 3652 1633 3664 1667
rect 3606 1607 3664 1633
rect 3706 1667 3764 1693
rect 3706 1633 3712 1667
rect 3752 1633 3764 1667
rect 3706 1607 3764 1633
rect 3806 1667 3864 1693
rect 3806 1633 3818 1667
rect 3858 1633 3864 1667
rect 3806 1607 3864 1633
rect 3906 1667 3964 1693
rect 3906 1633 3912 1667
rect 3952 1633 3964 1667
rect 3906 1607 3964 1633
rect 4006 1667 4064 1693
rect 4006 1633 4018 1667
rect 4058 1633 4064 1667
rect 4006 1607 4064 1633
rect 4106 1667 4164 1693
rect 4106 1633 4112 1667
rect 4152 1633 4164 1667
rect 4106 1607 4164 1633
rect 4206 1667 4264 1693
rect 4206 1633 4218 1667
rect 4258 1633 4264 1667
rect 4206 1607 4264 1633
rect 4306 1667 4364 1693
rect 4306 1633 4318 1667
rect 4352 1633 4364 1667
rect 4306 1607 4364 1633
rect 4406 1667 4464 1693
rect 4406 1633 4412 1667
rect 4452 1633 4464 1667
rect 4406 1607 4464 1633
rect 4506 1667 4564 1693
rect 4506 1633 4518 1667
rect 4558 1633 4564 1667
rect 4506 1607 4564 1633
rect 4606 1667 4664 1693
rect 4606 1633 4618 1667
rect 4652 1633 4664 1667
rect 4606 1607 4664 1633
rect 4706 1667 4764 1693
rect 4706 1633 4718 1667
rect 4752 1633 4764 1667
rect 4706 1607 4764 1633
rect 4806 1667 4864 1693
rect 4806 1633 4818 1667
rect 4852 1633 4864 1667
rect 4806 1607 4864 1633
rect 4906 1667 4964 1693
rect 4906 1633 4912 1667
rect 4952 1633 4964 1667
rect 4906 1607 4964 1633
rect 5006 1667 5064 1693
rect 5006 1633 5018 1667
rect 5058 1633 5064 1667
rect 5006 1607 5064 1633
rect 5106 1667 5164 1693
rect 5106 1633 5118 1667
rect 5152 1633 5164 1667
rect 5106 1607 5164 1633
rect 5206 1667 5264 1693
rect 5206 1633 5212 1667
rect 5252 1633 5264 1667
rect 5206 1607 5264 1633
rect 5306 1667 5364 1693
rect 5306 1633 5318 1667
rect 5358 1633 5364 1667
rect 5306 1607 5364 1633
rect 5406 1667 5464 1693
rect 5406 1633 5418 1667
rect 5452 1633 5464 1667
rect 5406 1607 5464 1633
rect 5506 1667 5564 1693
rect 5506 1633 5518 1667
rect 5552 1633 5564 1667
rect 5506 1607 5564 1633
rect 5606 1667 5664 1693
rect 5606 1633 5612 1667
rect 5652 1633 5664 1667
rect 5606 1607 5664 1633
rect 5706 1667 5764 1693
rect 5706 1633 5718 1667
rect 5758 1633 5764 1667
rect 5706 1607 5764 1633
rect 5806 1667 5864 1693
rect 5806 1633 5818 1667
rect 5852 1633 5864 1667
rect 5806 1607 5864 1633
rect 5906 1667 5964 1693
rect 5906 1633 5912 1667
rect 5952 1633 5964 1667
rect 5906 1607 5964 1633
rect 6006 1667 6064 1693
rect 6006 1633 6018 1667
rect 6058 1633 6064 1667
rect 6006 1607 6064 1633
rect 6106 1667 6164 1693
rect 6106 1633 6112 1667
rect 6152 1633 6164 1667
rect 6106 1607 6164 1633
rect 6206 1667 6264 1693
rect 6206 1633 6218 1667
rect 6258 1633 6264 1667
rect 6206 1607 6264 1633
rect 6306 1667 6364 1693
rect 6306 1633 6318 1667
rect 6352 1633 6364 1667
rect 6306 1607 6364 1633
rect 6406 1667 6464 1693
rect 6406 1633 6418 1667
rect 6452 1633 6464 1667
rect 6406 1607 6464 1633
rect 6506 1667 6564 1693
rect 6506 1633 6512 1667
rect 6552 1633 6564 1667
rect 6506 1607 6564 1633
rect 6606 1667 6664 1693
rect 6606 1633 6618 1667
rect 6658 1633 6664 1667
rect 6606 1607 6664 1633
rect 6706 1667 6764 1693
rect 6706 1633 6718 1667
rect 6752 1633 6764 1667
rect 6706 1607 6764 1633
rect 6806 1667 6864 1693
rect 6806 1633 6818 1667
rect 6852 1633 6864 1667
rect 6806 1607 6864 1633
rect 6906 1667 6964 1693
rect 6906 1633 6918 1667
rect 6952 1633 6964 1667
rect 6906 1607 6964 1633
rect 7006 1667 7064 1693
rect 7006 1633 7018 1667
rect 7052 1633 7064 1667
rect 7006 1607 7064 1633
rect 7106 1667 7164 1693
rect 7106 1633 7118 1667
rect 7152 1633 7164 1667
rect 7106 1607 7164 1633
rect 7206 1667 7264 1693
rect 7206 1633 7218 1667
rect 7252 1633 7264 1667
rect 7206 1607 7264 1633
rect 7306 1667 7364 1693
rect 7306 1633 7318 1667
rect 7352 1633 7364 1667
rect 7306 1607 7364 1633
rect 7406 1667 7464 1693
rect 7406 1633 7418 1667
rect 7452 1633 7464 1667
rect 7406 1607 7464 1633
rect 7506 1667 7564 1693
rect 7506 1633 7518 1667
rect 7552 1633 7564 1667
rect 7506 1607 7564 1633
rect 7606 1667 7664 1693
rect 7606 1633 7618 1667
rect 7652 1633 7664 1667
rect 7606 1607 7664 1633
rect 7706 1667 7764 1693
rect 7706 1633 7718 1667
rect 7752 1633 7764 1667
rect 7706 1607 7764 1633
rect 7806 1667 7864 1693
rect 7806 1633 7818 1667
rect 7852 1633 7864 1667
rect 7806 1607 7864 1633
rect 7906 1667 7964 1693
rect 7906 1633 7918 1667
rect 7952 1633 7964 1667
rect 7906 1607 7964 1633
rect 8006 1667 8064 1693
rect 8006 1633 8018 1667
rect 8052 1633 8064 1667
rect 8006 1607 8064 1633
rect 8106 1667 8164 1693
rect 8106 1633 8118 1667
rect 8152 1633 8164 1667
rect 8106 1607 8164 1633
rect 8206 1667 8264 1693
rect 8206 1633 8218 1667
rect 8252 1633 8264 1667
rect 8206 1607 8264 1633
rect 8306 1667 8364 1693
rect 8306 1633 8318 1667
rect 8352 1633 8364 1667
rect 8306 1607 8364 1633
rect 8406 1667 8464 1693
rect 8406 1633 8418 1667
rect 8452 1633 8464 1667
rect 8406 1607 8464 1633
rect 8506 1667 8564 1693
rect 8506 1633 8518 1667
rect 8552 1633 8564 1667
rect 8506 1607 8564 1633
rect 8606 1667 8664 1693
rect 8606 1633 8618 1667
rect 8652 1633 8664 1667
rect 8606 1607 8664 1633
rect 8706 1667 8764 1693
rect 8706 1633 8718 1667
rect 8752 1633 8764 1667
rect 8706 1607 8764 1633
rect 8806 1667 8864 1693
rect 8806 1633 8818 1667
rect 8852 1633 8864 1667
rect 8806 1607 8864 1633
rect 8906 1667 8964 1693
rect 8906 1633 8918 1667
rect 8952 1633 8964 1667
rect 8906 1607 8964 1633
rect 9006 1667 9064 1693
rect 9006 1633 9018 1667
rect 9052 1633 9064 1667
rect 9006 1607 9064 1633
rect 9106 1667 9164 1693
rect 9106 1633 9118 1667
rect 9152 1633 9164 1667
rect 9106 1607 9164 1633
rect 9206 1667 9264 1693
rect 9206 1633 9218 1667
rect 9252 1633 9264 1667
rect 9206 1607 9264 1633
rect 9306 1667 9364 1693
rect 9306 1633 9318 1667
rect 9352 1633 9364 1667
rect 9306 1607 9364 1633
rect 9406 1667 9464 1693
rect 9406 1633 9418 1667
rect 9452 1633 9464 1667
rect 9406 1607 9464 1633
rect 9506 1667 9564 1693
rect 9506 1633 9512 1667
rect 9552 1633 9564 1667
rect 9506 1607 9564 1633
rect 9606 1667 9664 1693
rect 9606 1633 9618 1667
rect 9658 1633 9664 1667
rect 9606 1607 9664 1633
rect 9706 1667 9764 1693
rect 9706 1633 9718 1667
rect 9752 1633 9764 1667
rect 9706 1607 9764 1633
rect 9806 1667 9864 1693
rect 9806 1633 9818 1667
rect 9852 1633 9864 1667
rect 9806 1607 9864 1633
rect 9906 1667 9964 1693
rect 9906 1633 9918 1667
rect 9952 1633 9964 1667
rect 9906 1607 9964 1633
rect 10006 1667 10064 1693
rect 10006 1633 10018 1667
rect 10052 1633 10064 1667
rect 10006 1607 10064 1633
rect 10106 1667 10164 1693
rect 10106 1633 10118 1667
rect 10152 1633 10164 1667
rect 10106 1607 10164 1633
rect 10206 1667 10264 1693
rect 10206 1633 10218 1667
rect 10252 1633 10264 1667
rect 10206 1607 10264 1633
rect 10306 1667 10364 1693
rect 10306 1633 10318 1667
rect 10352 1633 10364 1667
rect 10306 1607 10364 1633
rect 10406 1667 10464 1693
rect 10406 1633 10418 1667
rect 10452 1633 10464 1667
rect 10406 1607 10464 1633
rect 10506 1667 10564 1693
rect 10506 1633 10518 1667
rect 10552 1633 10564 1667
rect 10506 1607 10564 1633
rect 10606 1667 10664 1693
rect 10606 1633 10618 1667
rect 10652 1633 10664 1667
rect 10606 1607 10664 1633
rect 10706 1667 10764 1693
rect 10706 1633 10718 1667
rect 10752 1633 10764 1667
rect 10706 1607 10764 1633
rect 10806 1667 10864 1693
rect 10806 1633 10818 1667
rect 10852 1633 10864 1667
rect 10806 1607 10864 1633
rect 10906 1667 10964 1693
rect 10906 1633 10912 1667
rect 10952 1633 10964 1667
rect 10906 1607 10964 1633
rect 11006 1667 11064 1693
rect 11006 1633 11018 1667
rect 11058 1633 11064 1667
rect 11006 1607 11064 1633
rect 11106 1667 11164 1693
rect 11106 1633 11118 1667
rect 11152 1633 11164 1667
rect 11106 1607 11164 1633
rect 11206 1667 11264 1693
rect 11206 1633 11218 1667
rect 11252 1633 11264 1667
rect 11206 1607 11264 1633
rect 11306 1667 11364 1693
rect 11306 1633 11318 1667
rect 11352 1633 11364 1667
rect 11306 1607 11364 1633
rect 11406 1667 11464 1693
rect 11406 1633 11418 1667
rect 11452 1633 11464 1667
rect 11406 1607 11464 1633
rect 11506 1667 11564 1693
rect 11506 1633 11518 1667
rect 11552 1633 11564 1667
rect 11506 1607 11564 1633
rect 11606 1667 11664 1693
rect 11606 1633 11618 1667
rect 11652 1633 11664 1667
rect 11606 1607 11664 1633
rect 11706 1667 11764 1693
rect 11706 1633 11712 1667
rect 11752 1633 11764 1667
rect 11706 1607 11764 1633
rect 11806 1667 11864 1693
rect 11806 1633 11818 1667
rect 11858 1633 11864 1667
rect 11806 1607 11864 1633
rect 11906 1667 11964 1693
rect 11906 1633 11918 1667
rect 11952 1633 11964 1667
rect 11906 1607 11964 1633
rect 12006 1667 12064 1693
rect 12006 1633 12018 1667
rect 12052 1633 12064 1667
rect 12006 1607 12064 1633
rect 12106 1667 12164 1693
rect 12106 1633 12118 1667
rect 12152 1633 12164 1667
rect 12106 1607 12164 1633
rect 12206 1667 12264 1693
rect 12206 1633 12218 1667
rect 12252 1633 12264 1667
rect 12206 1607 12264 1633
rect 12306 1667 12364 1693
rect 12306 1633 12318 1667
rect 12352 1633 12364 1667
rect 12306 1607 12364 1633
rect 12406 1667 12464 1693
rect 12406 1633 12418 1667
rect 12452 1633 12464 1667
rect 12406 1607 12464 1633
rect 12506 1667 12564 1693
rect 12506 1633 12518 1667
rect 12552 1633 12564 1667
rect 12506 1607 12564 1633
rect 12606 1667 12664 1693
rect 12606 1633 12618 1667
rect 12652 1633 12664 1667
rect 12606 1607 12664 1633
rect 12706 1667 12764 1693
rect 12706 1633 12718 1667
rect 12752 1633 12764 1667
rect 12706 1607 12764 1633
rect 12806 1667 12864 1693
rect 13018 1686 13262 1720
rect 12806 1633 12818 1667
rect 12852 1633 12864 1667
rect 12908 1648 12916 1682
rect 12958 1648 12974 1682
rect 13018 1667 13052 1686
rect 12806 1607 12864 1633
rect 13228 1667 13262 1686
rect 13018 1617 13052 1633
rect 13096 1618 13112 1652
rect 13154 1618 13162 1652
rect 13228 1617 13262 1633
rect 13328 1667 13562 1683
rect 13362 1633 13428 1667
rect 13462 1633 13528 1667
rect 13328 1617 13562 1633
rect 13628 1667 13662 1683
rect 13628 1617 13662 1633
rect 6 1527 64 1553
rect 6 1493 18 1527
rect 52 1493 64 1527
rect 6 1467 64 1493
rect 106 1527 164 1553
rect 106 1493 118 1527
rect 152 1493 164 1527
rect 106 1467 164 1493
rect 206 1527 264 1553
rect 206 1493 218 1527
rect 252 1493 264 1527
rect 206 1467 264 1493
rect 306 1527 364 1553
rect 306 1493 318 1527
rect 352 1493 364 1527
rect 306 1467 364 1493
rect 406 1527 464 1553
rect 406 1493 412 1527
rect 452 1493 464 1527
rect 406 1467 464 1493
rect 506 1527 564 1553
rect 506 1493 518 1527
rect 558 1493 564 1527
rect 506 1467 564 1493
rect 606 1527 664 1553
rect 606 1493 618 1527
rect 652 1493 664 1527
rect 606 1467 664 1493
rect 706 1527 764 1553
rect 706 1493 718 1527
rect 752 1493 764 1527
rect 706 1467 764 1493
rect 806 1527 864 1553
rect 806 1493 818 1527
rect 852 1493 864 1527
rect 806 1467 864 1493
rect 906 1527 964 1553
rect 906 1493 918 1527
rect 952 1493 964 1527
rect 906 1467 964 1493
rect 1006 1527 1064 1553
rect 1006 1493 1018 1527
rect 1052 1493 1064 1527
rect 1006 1467 1064 1493
rect 1106 1527 1164 1553
rect 1106 1493 1118 1527
rect 1152 1493 1164 1527
rect 1106 1467 1164 1493
rect 1206 1527 1264 1553
rect 1206 1493 1218 1527
rect 1252 1493 1264 1527
rect 1206 1467 1264 1493
rect 1306 1527 1364 1553
rect 1306 1493 1318 1527
rect 1352 1493 1364 1527
rect 1306 1467 1364 1493
rect 1406 1527 1464 1553
rect 1406 1493 1418 1527
rect 1452 1493 1464 1527
rect 1406 1467 1464 1493
rect 1506 1527 1564 1553
rect 1506 1493 1518 1527
rect 1552 1493 1564 1527
rect 1506 1467 1564 1493
rect 1606 1527 1664 1553
rect 1606 1493 1618 1527
rect 1652 1493 1664 1527
rect 1606 1467 1664 1493
rect 1706 1527 1764 1553
rect 1706 1493 1718 1527
rect 1752 1493 1764 1527
rect 1706 1467 1764 1493
rect 1806 1527 1864 1553
rect 1806 1493 1818 1527
rect 1852 1493 1864 1527
rect 1806 1467 1864 1493
rect 1906 1527 1964 1553
rect 1906 1493 1918 1527
rect 1952 1493 1964 1527
rect 1906 1467 1964 1493
rect 2006 1527 2064 1553
rect 2006 1493 2018 1527
rect 2052 1493 2064 1527
rect 2006 1467 2064 1493
rect 2106 1527 2164 1553
rect 2106 1493 2118 1527
rect 2152 1493 2164 1527
rect 2106 1467 2164 1493
rect 2206 1527 2264 1553
rect 2206 1493 2218 1527
rect 2252 1493 2264 1527
rect 2206 1467 2264 1493
rect 2306 1527 2364 1553
rect 2306 1493 2318 1527
rect 2352 1493 2364 1527
rect 2306 1467 2364 1493
rect 2406 1527 2464 1553
rect 2406 1493 2418 1527
rect 2452 1493 2464 1527
rect 2406 1467 2464 1493
rect 2506 1527 2564 1553
rect 2506 1493 2512 1527
rect 2552 1493 2564 1527
rect 2506 1467 2564 1493
rect 2606 1527 2664 1553
rect 2606 1493 2618 1527
rect 2658 1493 2664 1527
rect 2606 1467 2664 1493
rect 2706 1527 2764 1553
rect 2706 1493 2718 1527
rect 2752 1493 2764 1527
rect 2706 1467 2764 1493
rect 2806 1527 2864 1553
rect 2806 1493 2818 1527
rect 2852 1493 2864 1527
rect 2806 1467 2864 1493
rect 2906 1527 2964 1553
rect 2906 1493 2918 1527
rect 2952 1493 2964 1527
rect 2906 1467 2964 1493
rect 3006 1527 3064 1553
rect 3006 1493 3018 1527
rect 3052 1493 3064 1527
rect 3006 1467 3064 1493
rect 3106 1527 3164 1553
rect 3106 1493 3112 1527
rect 3152 1493 3164 1527
rect 3106 1467 3164 1493
rect 3206 1527 3264 1553
rect 3206 1493 3218 1527
rect 3258 1493 3264 1527
rect 3206 1467 3264 1493
rect 3306 1527 3364 1553
rect 3306 1493 3318 1527
rect 3352 1493 3364 1527
rect 3306 1467 3364 1493
rect 3406 1527 3464 1553
rect 3406 1493 3418 1527
rect 3452 1493 3464 1527
rect 3406 1467 3464 1493
rect 3506 1527 3564 1553
rect 3506 1493 3512 1527
rect 3552 1493 3564 1527
rect 3506 1467 3564 1493
rect 3606 1527 3664 1553
rect 3606 1493 3618 1527
rect 3658 1493 3664 1527
rect 3606 1467 3664 1493
rect 3706 1527 3764 1553
rect 3706 1493 3718 1527
rect 3752 1493 3764 1527
rect 3706 1467 3764 1493
rect 3806 1527 3864 1553
rect 3806 1493 3818 1527
rect 3852 1493 3864 1527
rect 3806 1467 3864 1493
rect 3906 1527 3964 1553
rect 3906 1493 3918 1527
rect 3952 1493 3964 1527
rect 3906 1467 3964 1493
rect 4006 1527 4064 1553
rect 4006 1493 4012 1527
rect 4052 1493 4064 1527
rect 4006 1467 4064 1493
rect 4106 1527 4164 1553
rect 4106 1493 4118 1527
rect 4158 1493 4164 1527
rect 4106 1467 4164 1493
rect 4206 1527 4264 1553
rect 4206 1493 4218 1527
rect 4252 1493 4264 1527
rect 4206 1467 4264 1493
rect 4306 1527 4364 1553
rect 4306 1493 4318 1527
rect 4352 1493 4364 1527
rect 4306 1467 4364 1493
rect 4406 1527 4464 1553
rect 4406 1493 4418 1527
rect 4452 1493 4464 1527
rect 4406 1467 4464 1493
rect 4506 1527 4564 1553
rect 4506 1493 4518 1527
rect 4552 1493 4564 1527
rect 4506 1467 4564 1493
rect 4606 1527 4664 1553
rect 4606 1493 4618 1527
rect 4652 1493 4664 1527
rect 4606 1467 4664 1493
rect 4706 1527 4764 1553
rect 4706 1493 4718 1527
rect 4752 1493 4764 1527
rect 4706 1467 4764 1493
rect 4806 1527 4864 1553
rect 4806 1493 4812 1527
rect 4852 1493 4864 1527
rect 4806 1467 4864 1493
rect 4906 1527 4964 1553
rect 4906 1493 4918 1527
rect 4958 1493 4964 1527
rect 4906 1467 4964 1493
rect 5006 1527 5064 1553
rect 5006 1493 5018 1527
rect 5052 1493 5064 1527
rect 5006 1467 5064 1493
rect 5106 1527 5164 1553
rect 5106 1493 5118 1527
rect 5152 1493 5164 1527
rect 5106 1467 5164 1493
rect 5206 1527 5264 1553
rect 5206 1493 5218 1527
rect 5252 1493 5264 1527
rect 5206 1467 5264 1493
rect 5306 1527 5364 1553
rect 5306 1493 5318 1527
rect 5352 1493 5364 1527
rect 5306 1467 5364 1493
rect 5406 1527 5464 1553
rect 5406 1493 5418 1527
rect 5452 1493 5464 1527
rect 5406 1467 5464 1493
rect 5506 1527 5564 1553
rect 5506 1493 5518 1527
rect 5552 1493 5564 1527
rect 5506 1467 5564 1493
rect 5606 1527 5664 1553
rect 5606 1493 5618 1527
rect 5652 1493 5664 1527
rect 5606 1467 5664 1493
rect 5706 1527 5764 1553
rect 5706 1493 5718 1527
rect 5752 1493 5764 1527
rect 5706 1467 5764 1493
rect 5806 1527 5864 1553
rect 5806 1493 5812 1527
rect 5852 1493 5864 1527
rect 5806 1467 5864 1493
rect 5906 1527 5964 1553
rect 5906 1493 5918 1527
rect 5958 1493 5964 1527
rect 5906 1467 5964 1493
rect 6006 1527 6064 1553
rect 6006 1493 6012 1527
rect 6052 1493 6064 1527
rect 6006 1467 6064 1493
rect 6106 1527 6164 1553
rect 6106 1493 6118 1527
rect 6158 1493 6164 1527
rect 6106 1467 6164 1493
rect 6206 1527 6264 1553
rect 6206 1493 6218 1527
rect 6252 1493 6264 1527
rect 6206 1467 6264 1493
rect 6306 1527 6364 1553
rect 6306 1493 6312 1527
rect 6352 1493 6364 1527
rect 6306 1467 6364 1493
rect 6406 1527 6464 1553
rect 6406 1493 6418 1527
rect 6458 1493 6464 1527
rect 6406 1467 6464 1493
rect 6506 1527 6564 1553
rect 6506 1493 6518 1527
rect 6552 1493 6564 1527
rect 6506 1467 6564 1493
rect 6606 1527 6664 1553
rect 6606 1493 6618 1527
rect 6652 1493 6664 1527
rect 6606 1467 6664 1493
rect 6706 1527 6764 1553
rect 6706 1493 6718 1527
rect 6752 1493 6764 1527
rect 6706 1467 6764 1493
rect 6806 1527 6864 1553
rect 6806 1493 6818 1527
rect 6852 1493 6864 1527
rect 6806 1467 6864 1493
rect 6906 1527 6964 1553
rect 6906 1493 6918 1527
rect 6952 1493 6964 1527
rect 6906 1467 6964 1493
rect 7006 1527 7064 1553
rect 7006 1493 7018 1527
rect 7052 1493 7064 1527
rect 7006 1467 7064 1493
rect 7106 1527 7164 1553
rect 7106 1493 7118 1527
rect 7152 1493 7164 1527
rect 7106 1467 7164 1493
rect 7206 1527 7264 1553
rect 7206 1493 7218 1527
rect 7252 1493 7264 1527
rect 7206 1467 7264 1493
rect 7306 1527 7364 1553
rect 7306 1493 7318 1527
rect 7352 1493 7364 1527
rect 7306 1467 7364 1493
rect 7406 1527 7464 1553
rect 7406 1493 7418 1527
rect 7452 1493 7464 1527
rect 7406 1467 7464 1493
rect 7506 1527 7564 1553
rect 7506 1493 7518 1527
rect 7552 1493 7564 1527
rect 7506 1467 7564 1493
rect 7606 1527 7664 1553
rect 7606 1493 7618 1527
rect 7652 1493 7664 1527
rect 7606 1467 7664 1493
rect 7706 1527 7764 1553
rect 7706 1493 7712 1527
rect 7752 1493 7764 1527
rect 7706 1467 7764 1493
rect 7806 1527 7864 1553
rect 7806 1493 7818 1527
rect 7858 1493 7864 1527
rect 7806 1467 7864 1493
rect 7906 1527 7964 1553
rect 7906 1493 7912 1527
rect 7952 1493 7964 1527
rect 7906 1467 7964 1493
rect 8006 1527 8064 1553
rect 8006 1493 8018 1527
rect 8058 1493 8064 1527
rect 8006 1467 8064 1493
rect 8106 1527 8164 1553
rect 8106 1493 8118 1527
rect 8152 1493 8164 1527
rect 8106 1467 8164 1493
rect 8206 1527 8264 1553
rect 8206 1493 8218 1527
rect 8252 1493 8264 1527
rect 8206 1467 8264 1493
rect 8306 1527 8364 1553
rect 8306 1493 8318 1527
rect 8352 1493 8364 1527
rect 8306 1467 8364 1493
rect 8406 1527 8464 1553
rect 8406 1493 8418 1527
rect 8452 1493 8464 1527
rect 8406 1467 8464 1493
rect 8506 1527 8564 1553
rect 8506 1493 8512 1527
rect 8552 1493 8564 1527
rect 8506 1467 8564 1493
rect 8606 1527 8664 1553
rect 8606 1493 8618 1527
rect 8658 1493 8664 1527
rect 8606 1467 8664 1493
rect 8706 1527 8764 1553
rect 8706 1493 8718 1527
rect 8752 1493 8764 1527
rect 8706 1467 8764 1493
rect 8806 1527 8864 1553
rect 8806 1493 8818 1527
rect 8852 1493 8864 1527
rect 8806 1467 8864 1493
rect 8906 1527 8964 1553
rect 8906 1493 8918 1527
rect 8952 1493 8964 1527
rect 8906 1467 8964 1493
rect 9006 1527 9064 1553
rect 9006 1493 9018 1527
rect 9052 1493 9064 1527
rect 9006 1467 9064 1493
rect 9106 1527 9164 1553
rect 9106 1493 9118 1527
rect 9152 1493 9164 1527
rect 9106 1467 9164 1493
rect 9206 1527 9264 1553
rect 9206 1493 9218 1527
rect 9252 1493 9264 1527
rect 9206 1467 9264 1493
rect 9306 1527 9364 1553
rect 9306 1493 9312 1527
rect 9352 1493 9364 1527
rect 9306 1467 9364 1493
rect 9406 1527 9464 1553
rect 9406 1493 9418 1527
rect 9458 1493 9464 1527
rect 9406 1467 9464 1493
rect 9506 1527 9564 1553
rect 9506 1493 9518 1527
rect 9552 1493 9564 1527
rect 9506 1467 9564 1493
rect 9606 1527 9664 1553
rect 9606 1493 9618 1527
rect 9652 1493 9664 1527
rect 9606 1467 9664 1493
rect 9706 1527 9764 1553
rect 9706 1493 9718 1527
rect 9752 1493 9764 1527
rect 9706 1467 9764 1493
rect 9806 1527 9864 1553
rect 9806 1493 9818 1527
rect 9852 1493 9864 1527
rect 9806 1467 9864 1493
rect 9906 1527 9964 1553
rect 9906 1493 9918 1527
rect 9952 1493 9964 1527
rect 9906 1467 9964 1493
rect 10006 1527 10064 1553
rect 10006 1493 10018 1527
rect 10052 1493 10064 1527
rect 10006 1467 10064 1493
rect 10106 1527 10164 1553
rect 10106 1493 10118 1527
rect 10152 1493 10164 1527
rect 10106 1467 10164 1493
rect 10206 1527 10264 1553
rect 10206 1493 10218 1527
rect 10252 1493 10264 1527
rect 10206 1467 10264 1493
rect 10306 1527 10364 1553
rect 10306 1493 10318 1527
rect 10352 1493 10364 1527
rect 10306 1467 10364 1493
rect 10406 1527 10464 1553
rect 10406 1493 10418 1527
rect 10452 1493 10464 1527
rect 10406 1467 10464 1493
rect 10506 1527 10564 1553
rect 10506 1493 10518 1527
rect 10552 1493 10564 1527
rect 10506 1467 10564 1493
rect 10606 1527 10664 1553
rect 10606 1493 10618 1527
rect 10652 1493 10664 1527
rect 10606 1467 10664 1493
rect 10706 1527 10764 1553
rect 10706 1493 10718 1527
rect 10752 1493 10764 1527
rect 10706 1467 10764 1493
rect 10806 1527 10864 1553
rect 10806 1493 10818 1527
rect 10852 1493 10864 1527
rect 10806 1467 10864 1493
rect 10906 1527 10964 1553
rect 10906 1493 10912 1527
rect 10952 1493 10964 1527
rect 10906 1467 10964 1493
rect 11006 1527 11064 1553
rect 11006 1493 11018 1527
rect 11058 1493 11064 1527
rect 11006 1467 11064 1493
rect 11106 1527 11164 1553
rect 11106 1493 11112 1527
rect 11152 1493 11164 1527
rect 11106 1467 11164 1493
rect 11206 1527 11264 1553
rect 11206 1493 11218 1527
rect 11258 1493 11264 1527
rect 11206 1467 11264 1493
rect 11306 1527 11364 1553
rect 11306 1493 11318 1527
rect 11352 1493 11364 1527
rect 11306 1467 11364 1493
rect 11406 1527 11464 1553
rect 11406 1493 11418 1527
rect 11452 1493 11464 1527
rect 11406 1467 11464 1493
rect 11506 1527 11564 1553
rect 11506 1493 11518 1527
rect 11552 1493 11564 1527
rect 11506 1467 11564 1493
rect 11606 1527 11664 1553
rect 11606 1493 11618 1527
rect 11652 1493 11664 1527
rect 11606 1467 11664 1493
rect 11706 1527 11764 1553
rect 11706 1493 11718 1527
rect 11752 1493 11764 1527
rect 11706 1467 11764 1493
rect 11806 1527 11864 1553
rect 11806 1493 11818 1527
rect 11852 1493 11864 1527
rect 11806 1467 11864 1493
rect 11906 1527 11964 1553
rect 11906 1493 11918 1527
rect 11952 1493 11964 1527
rect 11906 1467 11964 1493
rect 12006 1527 12064 1553
rect 12006 1493 12012 1527
rect 12052 1493 12064 1527
rect 12006 1467 12064 1493
rect 12106 1527 12164 1553
rect 12106 1493 12118 1527
rect 12158 1493 12164 1527
rect 12106 1467 12164 1493
rect 12206 1527 12264 1553
rect 12206 1493 12218 1527
rect 12252 1493 12264 1527
rect 12206 1467 12264 1493
rect 12306 1527 12364 1553
rect 12306 1493 12318 1527
rect 12352 1493 12364 1527
rect 12306 1467 12364 1493
rect 12406 1527 12464 1553
rect 12406 1493 12412 1527
rect 12452 1493 12464 1527
rect 12406 1467 12464 1493
rect 12506 1527 12564 1553
rect 12506 1493 12518 1527
rect 12558 1493 12564 1527
rect 12506 1467 12564 1493
rect 12606 1527 12664 1553
rect 12606 1493 12618 1527
rect 12652 1493 12664 1527
rect 12606 1467 12664 1493
rect 12706 1527 12764 1553
rect 12706 1493 12718 1527
rect 12752 1493 12764 1527
rect 12706 1467 12764 1493
rect 12806 1527 12864 1553
rect 13018 1546 13262 1580
rect 12806 1493 12818 1527
rect 12852 1493 12864 1527
rect 12908 1508 12916 1542
rect 12958 1508 12974 1542
rect 13018 1527 13052 1546
rect 12806 1467 12864 1493
rect 13228 1543 13262 1546
rect 13228 1527 13362 1543
rect 13018 1477 13052 1493
rect 13096 1478 13112 1512
rect 13154 1478 13162 1512
rect 13262 1493 13328 1527
rect 13228 1477 13362 1493
rect 13428 1527 13462 1543
rect 13428 1477 13462 1493
rect 13528 1527 13662 1543
rect 13562 1493 13628 1527
rect 13528 1477 13662 1493
rect 6 1387 64 1413
rect 6 1353 18 1387
rect 52 1353 64 1387
rect 6 1327 64 1353
rect 106 1387 164 1413
rect 106 1353 118 1387
rect 152 1353 164 1387
rect 106 1327 164 1353
rect 206 1387 264 1413
rect 206 1353 218 1387
rect 252 1353 264 1387
rect 206 1327 264 1353
rect 306 1387 364 1413
rect 306 1353 318 1387
rect 352 1353 364 1387
rect 306 1327 364 1353
rect 406 1387 464 1413
rect 406 1353 418 1387
rect 452 1353 464 1387
rect 406 1327 464 1353
rect 506 1387 564 1413
rect 506 1353 518 1387
rect 552 1353 564 1387
rect 506 1327 564 1353
rect 606 1387 664 1413
rect 606 1353 618 1387
rect 652 1353 664 1387
rect 606 1327 664 1353
rect 706 1387 764 1413
rect 706 1353 718 1387
rect 752 1353 764 1387
rect 706 1327 764 1353
rect 806 1387 864 1413
rect 806 1353 812 1387
rect 852 1353 864 1387
rect 806 1327 864 1353
rect 906 1387 964 1413
rect 906 1353 918 1387
rect 958 1353 964 1387
rect 906 1327 964 1353
rect 1006 1387 1064 1413
rect 1006 1353 1018 1387
rect 1052 1353 1064 1387
rect 1006 1327 1064 1353
rect 1106 1387 1164 1413
rect 1106 1353 1118 1387
rect 1152 1353 1164 1387
rect 1106 1327 1164 1353
rect 1206 1387 1264 1413
rect 1206 1353 1218 1387
rect 1252 1353 1264 1387
rect 1206 1327 1264 1353
rect 1306 1387 1364 1413
rect 1306 1353 1318 1387
rect 1352 1353 1364 1387
rect 1306 1327 1364 1353
rect 1406 1387 1464 1413
rect 1406 1353 1418 1387
rect 1452 1353 1464 1387
rect 1406 1327 1464 1353
rect 1506 1387 1564 1413
rect 1506 1353 1518 1387
rect 1552 1353 1564 1387
rect 1506 1327 1564 1353
rect 1606 1387 1664 1413
rect 1606 1353 1618 1387
rect 1652 1353 1664 1387
rect 1606 1327 1664 1353
rect 1706 1387 1764 1413
rect 1706 1353 1718 1387
rect 1752 1353 1764 1387
rect 1706 1327 1764 1353
rect 1806 1387 1864 1413
rect 1806 1353 1818 1387
rect 1852 1353 1864 1387
rect 1806 1327 1864 1353
rect 1906 1387 1964 1413
rect 1906 1353 1918 1387
rect 1952 1353 1964 1387
rect 1906 1327 1964 1353
rect 2006 1387 2064 1413
rect 2006 1353 2018 1387
rect 2052 1353 2064 1387
rect 2006 1327 2064 1353
rect 2106 1387 2164 1413
rect 2106 1353 2118 1387
rect 2152 1353 2164 1387
rect 2106 1327 2164 1353
rect 2206 1387 2264 1413
rect 2206 1353 2218 1387
rect 2252 1353 2264 1387
rect 2206 1327 2264 1353
rect 2306 1387 2364 1413
rect 2306 1353 2318 1387
rect 2352 1353 2364 1387
rect 2306 1327 2364 1353
rect 2406 1387 2464 1413
rect 2406 1353 2418 1387
rect 2452 1353 2464 1387
rect 2406 1327 2464 1353
rect 2506 1387 2564 1413
rect 2506 1353 2518 1387
rect 2552 1353 2564 1387
rect 2506 1327 2564 1353
rect 2606 1387 2664 1413
rect 2606 1353 2618 1387
rect 2652 1353 2664 1387
rect 2606 1327 2664 1353
rect 2706 1387 2764 1413
rect 2706 1353 2718 1387
rect 2752 1353 2764 1387
rect 2706 1327 2764 1353
rect 2806 1387 2864 1413
rect 2806 1353 2812 1387
rect 2852 1353 2864 1387
rect 2806 1327 2864 1353
rect 2906 1387 2964 1413
rect 2906 1353 2918 1387
rect 2958 1353 2964 1387
rect 2906 1327 2964 1353
rect 3006 1387 3064 1413
rect 3006 1353 3018 1387
rect 3052 1353 3064 1387
rect 3006 1327 3064 1353
rect 3106 1387 3164 1413
rect 3106 1353 3118 1387
rect 3152 1353 3164 1387
rect 3106 1327 3164 1353
rect 3206 1387 3264 1413
rect 3206 1353 3218 1387
rect 3252 1353 3264 1387
rect 3206 1327 3264 1353
rect 3306 1387 3364 1413
rect 3306 1353 3318 1387
rect 3352 1353 3364 1387
rect 3306 1327 3364 1353
rect 3406 1387 3464 1413
rect 3406 1353 3418 1387
rect 3452 1353 3464 1387
rect 3406 1327 3464 1353
rect 3506 1387 3564 1413
rect 3506 1353 3518 1387
rect 3552 1353 3564 1387
rect 3506 1327 3564 1353
rect 3606 1387 3664 1413
rect 3606 1353 3618 1387
rect 3652 1353 3664 1387
rect 3606 1327 3664 1353
rect 3706 1387 3764 1413
rect 3706 1353 3718 1387
rect 3752 1353 3764 1387
rect 3706 1327 3764 1353
rect 3806 1387 3864 1413
rect 3806 1353 3818 1387
rect 3852 1353 3864 1387
rect 3806 1327 3864 1353
rect 3906 1387 3964 1413
rect 3906 1353 3918 1387
rect 3952 1353 3964 1387
rect 3906 1327 3964 1353
rect 4006 1387 4064 1413
rect 4006 1353 4018 1387
rect 4052 1353 4064 1387
rect 4006 1327 4064 1353
rect 4106 1387 4164 1413
rect 4106 1353 4118 1387
rect 4152 1353 4164 1387
rect 4106 1327 4164 1353
rect 4206 1387 4264 1413
rect 4206 1353 4218 1387
rect 4252 1353 4264 1387
rect 4206 1327 4264 1353
rect 4306 1387 4364 1413
rect 4306 1353 4318 1387
rect 4352 1353 4364 1387
rect 4306 1327 4364 1353
rect 4406 1387 4464 1413
rect 4406 1353 4418 1387
rect 4452 1353 4464 1387
rect 4406 1327 4464 1353
rect 4506 1387 4564 1413
rect 4506 1353 4518 1387
rect 4552 1353 4564 1387
rect 4506 1327 4564 1353
rect 4606 1387 4664 1413
rect 4606 1353 4612 1387
rect 4652 1353 4664 1387
rect 4606 1327 4664 1353
rect 4706 1387 4764 1413
rect 4706 1353 4718 1387
rect 4758 1353 4764 1387
rect 4706 1327 4764 1353
rect 4806 1387 4864 1413
rect 4806 1353 4812 1387
rect 4852 1353 4864 1387
rect 4806 1327 4864 1353
rect 4906 1387 4964 1413
rect 4906 1353 4918 1387
rect 4958 1353 4964 1387
rect 4906 1327 4964 1353
rect 5006 1387 5064 1413
rect 5006 1353 5018 1387
rect 5052 1353 5064 1387
rect 5006 1327 5064 1353
rect 5106 1387 5164 1413
rect 5106 1353 5112 1387
rect 5152 1353 5164 1387
rect 5106 1327 5164 1353
rect 5206 1387 5264 1413
rect 5206 1353 5218 1387
rect 5258 1353 5264 1387
rect 5206 1327 5264 1353
rect 5306 1387 5364 1413
rect 5306 1353 5318 1387
rect 5352 1353 5364 1387
rect 5306 1327 5364 1353
rect 5406 1387 5464 1413
rect 5406 1353 5418 1387
rect 5452 1353 5464 1387
rect 5406 1327 5464 1353
rect 5506 1387 5564 1413
rect 5506 1353 5518 1387
rect 5552 1353 5564 1387
rect 5506 1327 5564 1353
rect 5606 1387 5664 1413
rect 5606 1353 5618 1387
rect 5652 1353 5664 1387
rect 5606 1327 5664 1353
rect 5706 1387 5764 1413
rect 5706 1353 5718 1387
rect 5752 1353 5764 1387
rect 5706 1327 5764 1353
rect 5806 1387 5864 1413
rect 5806 1353 5818 1387
rect 5852 1353 5864 1387
rect 5806 1327 5864 1353
rect 5906 1387 5964 1413
rect 5906 1353 5918 1387
rect 5952 1353 5964 1387
rect 5906 1327 5964 1353
rect 6006 1387 6064 1413
rect 6006 1353 6018 1387
rect 6052 1353 6064 1387
rect 6006 1327 6064 1353
rect 6106 1387 6164 1413
rect 6106 1353 6118 1387
rect 6152 1353 6164 1387
rect 6106 1327 6164 1353
rect 6206 1387 6264 1413
rect 6206 1353 6212 1387
rect 6252 1353 6264 1387
rect 6206 1327 6264 1353
rect 6306 1387 6364 1413
rect 6306 1353 6318 1387
rect 6358 1353 6364 1387
rect 6306 1327 6364 1353
rect 6406 1387 6464 1413
rect 6406 1353 6412 1387
rect 6452 1353 6464 1387
rect 6406 1327 6464 1353
rect 6506 1387 6564 1413
rect 6506 1353 6518 1387
rect 6558 1353 6564 1387
rect 6506 1327 6564 1353
rect 6606 1387 6664 1413
rect 6606 1353 6618 1387
rect 6652 1353 6664 1387
rect 6606 1327 6664 1353
rect 6706 1387 6764 1413
rect 6706 1353 6712 1387
rect 6752 1353 6764 1387
rect 6706 1327 6764 1353
rect 6806 1387 6864 1413
rect 6806 1353 6818 1387
rect 6858 1353 6864 1387
rect 6806 1327 6864 1353
rect 6906 1387 6964 1413
rect 6906 1353 6912 1387
rect 6952 1353 6964 1387
rect 6906 1327 6964 1353
rect 7006 1387 7064 1413
rect 7006 1353 7018 1387
rect 7058 1353 7064 1387
rect 7006 1327 7064 1353
rect 7106 1387 7164 1413
rect 7106 1353 7118 1387
rect 7152 1353 7164 1387
rect 7106 1327 7164 1353
rect 7206 1387 7264 1413
rect 7206 1353 7218 1387
rect 7252 1353 7264 1387
rect 7206 1327 7264 1353
rect 7306 1387 7364 1413
rect 7306 1353 7318 1387
rect 7352 1353 7364 1387
rect 7306 1327 7364 1353
rect 7406 1387 7464 1413
rect 7406 1353 7418 1387
rect 7452 1353 7464 1387
rect 7406 1327 7464 1353
rect 7506 1387 7564 1413
rect 7506 1353 7518 1387
rect 7552 1353 7564 1387
rect 7506 1327 7564 1353
rect 7606 1387 7664 1413
rect 7606 1353 7618 1387
rect 7652 1353 7664 1387
rect 7606 1327 7664 1353
rect 7706 1387 7764 1413
rect 7706 1353 7718 1387
rect 7752 1353 7764 1387
rect 7706 1327 7764 1353
rect 7806 1387 7864 1413
rect 7806 1353 7818 1387
rect 7852 1353 7864 1387
rect 7806 1327 7864 1353
rect 7906 1387 7964 1413
rect 7906 1353 7912 1387
rect 7952 1353 7964 1387
rect 7906 1327 7964 1353
rect 8006 1387 8064 1413
rect 8006 1353 8018 1387
rect 8058 1353 8064 1387
rect 8006 1327 8064 1353
rect 8106 1387 8164 1413
rect 8106 1353 8118 1387
rect 8152 1353 8164 1387
rect 8106 1327 8164 1353
rect 8206 1387 8264 1413
rect 8206 1353 8218 1387
rect 8252 1353 8264 1387
rect 8206 1327 8264 1353
rect 8306 1387 8364 1413
rect 8306 1353 8318 1387
rect 8352 1353 8364 1387
rect 8306 1327 8364 1353
rect 8406 1387 8464 1413
rect 8406 1353 8418 1387
rect 8452 1353 8464 1387
rect 8406 1327 8464 1353
rect 8506 1387 8564 1413
rect 8506 1353 8518 1387
rect 8552 1353 8564 1387
rect 8506 1327 8564 1353
rect 8606 1387 8664 1413
rect 8606 1353 8618 1387
rect 8652 1353 8664 1387
rect 8606 1327 8664 1353
rect 8706 1387 8764 1413
rect 8706 1353 8718 1387
rect 8752 1353 8764 1387
rect 8706 1327 8764 1353
rect 8806 1387 8864 1413
rect 8806 1353 8818 1387
rect 8852 1353 8864 1387
rect 8806 1327 8864 1353
rect 8906 1387 8964 1413
rect 8906 1353 8918 1387
rect 8952 1353 8964 1387
rect 8906 1327 8964 1353
rect 9006 1387 9064 1413
rect 9006 1353 9018 1387
rect 9052 1353 9064 1387
rect 9006 1327 9064 1353
rect 9106 1387 9164 1413
rect 9106 1353 9118 1387
rect 9152 1353 9164 1387
rect 9106 1327 9164 1353
rect 9206 1387 9264 1413
rect 9206 1353 9218 1387
rect 9252 1353 9264 1387
rect 9206 1327 9264 1353
rect 9306 1387 9364 1413
rect 9306 1353 9312 1387
rect 9352 1353 9364 1387
rect 9306 1327 9364 1353
rect 9406 1387 9464 1413
rect 9406 1353 9418 1387
rect 9458 1353 9464 1387
rect 9406 1327 9464 1353
rect 9506 1387 9564 1413
rect 9506 1353 9518 1387
rect 9552 1353 9564 1387
rect 9506 1327 9564 1353
rect 9606 1387 9664 1413
rect 9606 1353 9618 1387
rect 9652 1353 9664 1387
rect 9606 1327 9664 1353
rect 9706 1387 9764 1413
rect 9706 1353 9718 1387
rect 9752 1353 9764 1387
rect 9706 1327 9764 1353
rect 9806 1387 9864 1413
rect 9806 1353 9818 1387
rect 9852 1353 9864 1387
rect 9806 1327 9864 1353
rect 9906 1387 9964 1413
rect 9906 1353 9918 1387
rect 9952 1353 9964 1387
rect 9906 1327 9964 1353
rect 10006 1387 10064 1413
rect 10006 1353 10018 1387
rect 10052 1353 10064 1387
rect 10006 1327 10064 1353
rect 10106 1387 10164 1413
rect 10106 1353 10118 1387
rect 10152 1353 10164 1387
rect 10106 1327 10164 1353
rect 10206 1387 10264 1413
rect 10206 1353 10212 1387
rect 10252 1353 10264 1387
rect 10206 1327 10264 1353
rect 10306 1387 10364 1413
rect 10306 1353 10318 1387
rect 10358 1353 10364 1387
rect 10306 1327 10364 1353
rect 10406 1387 10464 1413
rect 10406 1353 10418 1387
rect 10452 1353 10464 1387
rect 10406 1327 10464 1353
rect 10506 1387 10564 1413
rect 10506 1353 10518 1387
rect 10552 1353 10564 1387
rect 10506 1327 10564 1353
rect 10606 1387 10664 1413
rect 10606 1353 10618 1387
rect 10652 1353 10664 1387
rect 10606 1327 10664 1353
rect 10706 1387 10764 1413
rect 10706 1353 10718 1387
rect 10752 1353 10764 1387
rect 10706 1327 10764 1353
rect 10806 1387 10864 1413
rect 10806 1353 10818 1387
rect 10852 1353 10864 1387
rect 10806 1327 10864 1353
rect 10906 1387 10964 1413
rect 10906 1353 10918 1387
rect 10952 1353 10964 1387
rect 10906 1327 10964 1353
rect 11006 1387 11064 1413
rect 11006 1353 11018 1387
rect 11052 1353 11064 1387
rect 11006 1327 11064 1353
rect 11106 1387 11164 1413
rect 11106 1353 11112 1387
rect 11152 1353 11164 1387
rect 11106 1327 11164 1353
rect 11206 1387 11264 1413
rect 11206 1353 11218 1387
rect 11258 1353 11264 1387
rect 11206 1327 11264 1353
rect 11306 1387 11364 1413
rect 11306 1353 11318 1387
rect 11352 1353 11364 1387
rect 11306 1327 11364 1353
rect 11406 1387 11464 1413
rect 11406 1353 11418 1387
rect 11452 1353 11464 1387
rect 11406 1327 11464 1353
rect 11506 1387 11564 1413
rect 11506 1353 11518 1387
rect 11552 1353 11564 1387
rect 11506 1327 11564 1353
rect 11606 1387 11664 1413
rect 11606 1353 11618 1387
rect 11652 1353 11664 1387
rect 11606 1327 11664 1353
rect 11706 1387 11764 1413
rect 11706 1353 11712 1387
rect 11752 1353 11764 1387
rect 11706 1327 11764 1353
rect 11806 1387 11864 1413
rect 11806 1353 11818 1387
rect 11858 1353 11864 1387
rect 11806 1327 11864 1353
rect 11906 1387 11964 1413
rect 11906 1353 11918 1387
rect 11952 1353 11964 1387
rect 11906 1327 11964 1353
rect 12006 1387 12064 1413
rect 12006 1353 12018 1387
rect 12052 1353 12064 1387
rect 12006 1327 12064 1353
rect 12106 1387 12164 1413
rect 12106 1353 12118 1387
rect 12152 1353 12164 1387
rect 12106 1327 12164 1353
rect 12206 1387 12264 1413
rect 12206 1353 12218 1387
rect 12252 1353 12264 1387
rect 12206 1327 12264 1353
rect 12306 1387 12364 1413
rect 12306 1353 12318 1387
rect 12352 1353 12364 1387
rect 12306 1327 12364 1353
rect 12406 1387 12464 1413
rect 12406 1353 12412 1387
rect 12452 1353 12464 1387
rect 12406 1327 12464 1353
rect 12506 1387 12564 1413
rect 12506 1353 12518 1387
rect 12558 1353 12564 1387
rect 12506 1327 12564 1353
rect 12606 1387 12664 1413
rect 12606 1353 12618 1387
rect 12652 1353 12664 1387
rect 12606 1327 12664 1353
rect 12706 1387 12764 1413
rect 12706 1353 12718 1387
rect 12752 1353 12764 1387
rect 12706 1327 12764 1353
rect 12806 1387 12864 1413
rect 13018 1406 13262 1440
rect 12806 1353 12818 1387
rect 12852 1353 12864 1387
rect 12908 1368 12916 1402
rect 12958 1368 12974 1402
rect 13018 1387 13052 1406
rect 12806 1327 12864 1353
rect 13228 1387 13262 1406
rect 13018 1337 13052 1353
rect 13096 1338 13112 1372
rect 13154 1338 13162 1372
rect 13228 1337 13262 1353
rect 13328 1387 13462 1403
rect 13362 1353 13428 1387
rect 13328 1337 13462 1353
rect 13528 1387 13662 1403
rect 13562 1353 13628 1387
rect 13528 1337 13662 1353
rect 8 1230 18 1264
rect 52 1230 118 1264
rect 152 1230 168 1264
rect 208 1246 218 1280
rect 252 1246 318 1280
rect 352 1246 368 1280
rect 408 1230 418 1264
rect 452 1230 518 1264
rect 552 1230 568 1264
rect 608 1246 618 1280
rect 652 1246 718 1280
rect 752 1246 768 1280
rect 808 1230 818 1264
rect 852 1230 918 1264
rect 952 1230 968 1264
rect 1008 1246 1018 1280
rect 1052 1246 1118 1280
rect 1152 1246 1168 1280
rect 1208 1230 1218 1264
rect 1252 1230 1318 1264
rect 1352 1230 1368 1264
rect 1408 1246 1418 1280
rect 1452 1246 1518 1280
rect 1552 1246 1568 1280
rect 1608 1230 1618 1264
rect 1652 1230 1718 1264
rect 1752 1230 1768 1264
rect 1808 1246 1818 1280
rect 1852 1246 1918 1280
rect 1952 1246 1968 1280
rect 2008 1230 2018 1264
rect 2052 1230 2118 1264
rect 2152 1230 2168 1264
rect 2208 1246 2218 1280
rect 2252 1246 2318 1280
rect 2352 1246 2368 1280
rect 2408 1230 2418 1264
rect 2452 1230 2518 1264
rect 2552 1230 2568 1264
rect 2608 1246 2618 1280
rect 2652 1246 2718 1280
rect 2752 1246 2768 1280
rect 2808 1230 2818 1264
rect 2852 1230 2918 1264
rect 2952 1230 2968 1264
rect 3008 1246 3018 1280
rect 3052 1246 3118 1280
rect 3152 1246 3168 1280
rect 3208 1230 3218 1264
rect 3252 1230 3318 1264
rect 3352 1230 3368 1264
rect 3408 1246 3418 1280
rect 3452 1246 3518 1280
rect 3552 1246 3568 1280
rect 3608 1230 3618 1264
rect 3652 1230 3718 1264
rect 3752 1230 3768 1264
rect 3808 1246 3818 1280
rect 3852 1246 3918 1280
rect 3952 1246 3968 1280
rect 4008 1230 4018 1264
rect 4052 1230 4118 1264
rect 4152 1230 4168 1264
rect 4208 1246 4218 1280
rect 4252 1246 4318 1280
rect 4352 1246 4368 1280
rect 4408 1230 4418 1264
rect 4452 1230 4518 1264
rect 4552 1230 4568 1264
rect 4608 1246 4618 1280
rect 4652 1246 4718 1280
rect 4752 1246 4768 1280
rect 4808 1230 4818 1264
rect 4852 1230 4918 1264
rect 4952 1230 4968 1264
rect 5008 1246 5018 1280
rect 5052 1246 5118 1280
rect 5152 1246 5168 1280
rect 5208 1230 5218 1264
rect 5252 1230 5318 1264
rect 5352 1230 5368 1264
rect 5408 1246 5418 1280
rect 5452 1246 5518 1280
rect 5552 1246 5568 1280
rect 5608 1230 5618 1264
rect 5652 1230 5718 1264
rect 5752 1230 5768 1264
rect 5808 1246 5818 1280
rect 5852 1246 5918 1280
rect 5952 1246 5968 1280
rect 6008 1230 6018 1264
rect 6052 1230 6118 1264
rect 6152 1230 6168 1264
rect 6208 1246 6218 1280
rect 6252 1246 6318 1280
rect 6352 1246 6368 1280
rect 6408 1230 6418 1264
rect 6452 1230 6518 1264
rect 6552 1230 6568 1264
rect 6608 1246 6618 1280
rect 6652 1246 6718 1280
rect 6752 1246 6768 1280
rect 6808 1230 6818 1264
rect 6852 1230 6918 1264
rect 6952 1230 6968 1264
rect 7008 1246 7018 1280
rect 7052 1246 7118 1280
rect 7152 1246 7168 1280
rect 7208 1230 7218 1264
rect 7252 1230 7318 1264
rect 7352 1230 7368 1264
rect 7408 1246 7418 1280
rect 7452 1246 7518 1280
rect 7552 1246 7568 1280
rect 7608 1230 7618 1264
rect 7652 1230 7718 1264
rect 7752 1230 7768 1264
rect 7808 1246 7818 1280
rect 7852 1246 7918 1280
rect 7952 1246 7968 1280
rect 8008 1230 8018 1264
rect 8052 1230 8118 1264
rect 8152 1230 8168 1264
rect 8208 1246 8218 1280
rect 8252 1246 8318 1280
rect 8352 1246 8368 1280
rect 8408 1230 8418 1264
rect 8452 1230 8518 1264
rect 8552 1230 8568 1264
rect 8608 1246 8618 1280
rect 8652 1246 8718 1280
rect 8752 1246 8768 1280
rect 8808 1230 8818 1264
rect 8852 1230 8918 1264
rect 8952 1230 8968 1264
rect 9008 1246 9018 1280
rect 9052 1246 9118 1280
rect 9152 1246 9168 1280
rect 9208 1230 9218 1264
rect 9252 1230 9318 1264
rect 9352 1230 9368 1264
rect 9408 1246 9418 1280
rect 9452 1246 9518 1280
rect 9552 1246 9568 1280
rect 9608 1230 9618 1264
rect 9652 1230 9718 1264
rect 9752 1230 9768 1264
rect 9808 1246 9818 1280
rect 9852 1246 9918 1280
rect 9952 1246 9968 1280
rect 10008 1230 10018 1264
rect 10052 1230 10118 1264
rect 10152 1230 10168 1264
rect 10208 1246 10218 1280
rect 10252 1246 10318 1280
rect 10352 1246 10368 1280
rect 10408 1230 10418 1264
rect 10452 1230 10518 1264
rect 10552 1230 10568 1264
rect 10608 1246 10618 1280
rect 10652 1246 10718 1280
rect 10752 1246 10768 1280
rect 10808 1230 10818 1264
rect 10852 1230 10918 1264
rect 10952 1230 10968 1264
rect 11008 1246 11018 1280
rect 11052 1246 11118 1280
rect 11152 1246 11168 1280
rect 11208 1230 11218 1264
rect 11252 1230 11318 1264
rect 11352 1230 11368 1264
rect 11408 1246 11418 1280
rect 11452 1246 11518 1280
rect 11552 1246 11568 1280
rect 11608 1230 11618 1264
rect 11652 1230 11718 1264
rect 11752 1230 11768 1264
rect 11808 1246 11818 1280
rect 11852 1246 11918 1280
rect 11952 1246 11968 1280
rect 12008 1230 12018 1264
rect 12052 1230 12118 1264
rect 12152 1230 12168 1264
rect 12208 1246 12218 1280
rect 12252 1246 12318 1280
rect 12352 1246 12368 1280
rect 12408 1230 12418 1264
rect 12452 1230 12518 1264
rect 12552 1230 12568 1264
rect 12608 1246 12618 1280
rect 12652 1246 12718 1280
rect 12752 1246 12768 1280
rect 12916 1261 12968 1278
rect 12950 1244 12968 1261
rect 13002 1244 13018 1278
rect 13052 1244 13068 1278
rect 13102 1249 13120 1278
rect 13102 1244 13154 1249
rect 13262 1244 13278 1278
rect 13312 1244 13328 1278
rect 13362 1244 13378 1278
rect 13412 1244 13428 1278
rect 13462 1244 13478 1278
rect 13512 1244 13528 1278
rect 13562 1244 13578 1278
rect 13612 1244 13628 1278
rect 6 1157 64 1183
rect 6 1123 18 1157
rect 52 1123 64 1157
rect 6 1097 64 1123
rect 106 1157 164 1183
rect 106 1123 118 1157
rect 152 1123 164 1157
rect 106 1097 164 1123
rect 206 1157 264 1183
rect 206 1123 218 1157
rect 252 1123 264 1157
rect 206 1097 264 1123
rect 306 1157 364 1183
rect 306 1123 318 1157
rect 352 1123 364 1157
rect 306 1097 364 1123
rect 406 1157 464 1183
rect 406 1123 418 1157
rect 452 1123 464 1157
rect 406 1097 464 1123
rect 506 1157 564 1183
rect 506 1123 518 1157
rect 552 1123 564 1157
rect 506 1097 564 1123
rect 606 1157 664 1183
rect 606 1123 618 1157
rect 652 1123 664 1157
rect 606 1097 664 1123
rect 706 1157 764 1183
rect 706 1123 718 1157
rect 752 1123 764 1157
rect 706 1097 764 1123
rect 806 1157 864 1183
rect 806 1123 818 1157
rect 852 1123 864 1157
rect 806 1097 864 1123
rect 906 1157 964 1183
rect 906 1123 918 1157
rect 952 1123 964 1157
rect 906 1097 964 1123
rect 1006 1157 1064 1183
rect 1006 1123 1018 1157
rect 1052 1123 1064 1157
rect 1006 1097 1064 1123
rect 1106 1157 1164 1183
rect 1106 1123 1118 1157
rect 1152 1123 1164 1157
rect 1106 1097 1164 1123
rect 1206 1157 1264 1183
rect 1206 1123 1218 1157
rect 1252 1123 1264 1157
rect 1206 1097 1264 1123
rect 1306 1157 1364 1183
rect 1306 1123 1318 1157
rect 1352 1123 1364 1157
rect 1306 1097 1364 1123
rect 1406 1157 1464 1183
rect 1406 1123 1418 1157
rect 1452 1123 1464 1157
rect 1406 1097 1464 1123
rect 1506 1157 1564 1183
rect 1506 1123 1518 1157
rect 1552 1123 1564 1157
rect 1506 1097 1564 1123
rect 1606 1157 1664 1183
rect 1606 1123 1618 1157
rect 1652 1123 1664 1157
rect 1606 1097 1664 1123
rect 1706 1157 1764 1183
rect 1706 1123 1712 1157
rect 1752 1123 1764 1157
rect 1706 1097 1764 1123
rect 1806 1157 1864 1183
rect 1806 1123 1818 1157
rect 1858 1123 1864 1157
rect 1806 1097 1864 1123
rect 1906 1157 1964 1183
rect 1906 1123 1918 1157
rect 1952 1123 1964 1157
rect 1906 1097 1964 1123
rect 2006 1157 2064 1183
rect 2006 1123 2012 1157
rect 2052 1123 2064 1157
rect 2006 1097 2064 1123
rect 2106 1157 2164 1183
rect 2106 1123 2118 1157
rect 2158 1123 2164 1157
rect 2106 1097 2164 1123
rect 2206 1157 2264 1183
rect 2206 1123 2218 1157
rect 2252 1123 2264 1157
rect 2206 1097 2264 1123
rect 2306 1157 2364 1183
rect 2306 1123 2318 1157
rect 2352 1123 2364 1157
rect 2306 1097 2364 1123
rect 2406 1157 2464 1183
rect 2406 1123 2418 1157
rect 2452 1123 2464 1157
rect 2406 1097 2464 1123
rect 2506 1157 2564 1183
rect 2506 1123 2518 1157
rect 2552 1123 2564 1157
rect 2506 1097 2564 1123
rect 2606 1157 2664 1183
rect 2606 1123 2618 1157
rect 2652 1123 2664 1157
rect 2606 1097 2664 1123
rect 2706 1157 2764 1183
rect 2706 1123 2718 1157
rect 2752 1123 2764 1157
rect 2706 1097 2764 1123
rect 2806 1157 2864 1183
rect 2806 1123 2818 1157
rect 2852 1123 2864 1157
rect 2806 1097 2864 1123
rect 2906 1157 2964 1183
rect 2906 1123 2918 1157
rect 2952 1123 2964 1157
rect 2906 1097 2964 1123
rect 3006 1157 3064 1183
rect 3006 1123 3012 1157
rect 3052 1123 3064 1157
rect 3006 1097 3064 1123
rect 3106 1157 3164 1183
rect 3106 1123 3118 1157
rect 3158 1123 3164 1157
rect 3106 1097 3164 1123
rect 3206 1157 3264 1183
rect 3206 1123 3212 1157
rect 3252 1123 3264 1157
rect 3206 1097 3264 1123
rect 3306 1157 3364 1183
rect 3306 1123 3318 1157
rect 3358 1123 3364 1157
rect 3306 1097 3364 1123
rect 3406 1157 3464 1183
rect 3406 1123 3418 1157
rect 3452 1123 3464 1157
rect 3406 1097 3464 1123
rect 3506 1157 3564 1183
rect 3506 1123 3518 1157
rect 3552 1123 3564 1157
rect 3506 1097 3564 1123
rect 3606 1157 3664 1183
rect 3606 1123 3618 1157
rect 3652 1123 3664 1157
rect 3606 1097 3664 1123
rect 3706 1157 3764 1183
rect 3706 1123 3712 1157
rect 3752 1123 3764 1157
rect 3706 1097 3764 1123
rect 3806 1157 3864 1183
rect 3806 1123 3818 1157
rect 3858 1123 3864 1157
rect 3806 1097 3864 1123
rect 3906 1157 3964 1183
rect 3906 1123 3918 1157
rect 3952 1123 3964 1157
rect 3906 1097 3964 1123
rect 4006 1157 4064 1183
rect 4006 1123 4018 1157
rect 4052 1123 4064 1157
rect 4006 1097 4064 1123
rect 4106 1157 4164 1183
rect 4106 1123 4118 1157
rect 4152 1123 4164 1157
rect 4106 1097 4164 1123
rect 4206 1157 4264 1183
rect 4206 1123 4218 1157
rect 4252 1123 4264 1157
rect 4206 1097 4264 1123
rect 4306 1157 4364 1183
rect 4306 1123 4318 1157
rect 4352 1123 4364 1157
rect 4306 1097 4364 1123
rect 4406 1157 4464 1183
rect 4406 1123 4412 1157
rect 4452 1123 4464 1157
rect 4406 1097 4464 1123
rect 4506 1157 4564 1183
rect 4506 1123 4518 1157
rect 4558 1123 4564 1157
rect 4506 1097 4564 1123
rect 4606 1157 4664 1183
rect 4606 1123 4612 1157
rect 4652 1123 4664 1157
rect 4606 1097 4664 1123
rect 4706 1157 4764 1183
rect 4706 1123 4718 1157
rect 4758 1123 4764 1157
rect 4706 1097 4764 1123
rect 4806 1157 4864 1183
rect 4806 1123 4818 1157
rect 4852 1123 4864 1157
rect 4806 1097 4864 1123
rect 4906 1157 4964 1183
rect 4906 1123 4918 1157
rect 4952 1123 4964 1157
rect 4906 1097 4964 1123
rect 5006 1157 5064 1183
rect 5006 1123 5018 1157
rect 5052 1123 5064 1157
rect 5006 1097 5064 1123
rect 5106 1157 5164 1183
rect 5106 1123 5118 1157
rect 5152 1123 5164 1157
rect 5106 1097 5164 1123
rect 5206 1157 5264 1183
rect 5206 1123 5218 1157
rect 5252 1123 5264 1157
rect 5206 1097 5264 1123
rect 5306 1157 5364 1183
rect 5306 1123 5318 1157
rect 5352 1123 5364 1157
rect 5306 1097 5364 1123
rect 5406 1157 5464 1183
rect 5406 1123 5412 1157
rect 5452 1123 5464 1157
rect 5406 1097 5464 1123
rect 5506 1157 5564 1183
rect 5506 1123 5518 1157
rect 5558 1123 5564 1157
rect 5506 1097 5564 1123
rect 5606 1157 5664 1183
rect 5606 1123 5618 1157
rect 5652 1123 5664 1157
rect 5606 1097 5664 1123
rect 5706 1157 5764 1183
rect 5706 1123 5718 1157
rect 5752 1123 5764 1157
rect 5706 1097 5764 1123
rect 5806 1157 5864 1183
rect 5806 1123 5818 1157
rect 5852 1123 5864 1157
rect 5806 1097 5864 1123
rect 5906 1157 5964 1183
rect 5906 1123 5918 1157
rect 5952 1123 5964 1157
rect 5906 1097 5964 1123
rect 6006 1157 6064 1183
rect 6006 1123 6018 1157
rect 6052 1123 6064 1157
rect 6006 1097 6064 1123
rect 6106 1157 6164 1183
rect 6106 1123 6118 1157
rect 6152 1123 6164 1157
rect 6106 1097 6164 1123
rect 6206 1157 6264 1183
rect 6206 1123 6218 1157
rect 6252 1123 6264 1157
rect 6206 1097 6264 1123
rect 6306 1157 6364 1183
rect 6306 1123 6318 1157
rect 6352 1123 6364 1157
rect 6306 1097 6364 1123
rect 6406 1157 6464 1183
rect 6406 1123 6418 1157
rect 6452 1123 6464 1157
rect 6406 1097 6464 1123
rect 6506 1157 6564 1183
rect 6506 1123 6518 1157
rect 6552 1123 6564 1157
rect 6506 1097 6564 1123
rect 6606 1157 6664 1183
rect 6606 1123 6618 1157
rect 6652 1123 6664 1157
rect 6606 1097 6664 1123
rect 6706 1157 6764 1183
rect 6706 1123 6712 1157
rect 6752 1123 6764 1157
rect 6706 1097 6764 1123
rect 6806 1157 6864 1183
rect 6806 1123 6818 1157
rect 6858 1123 6864 1157
rect 6806 1097 6864 1123
rect 6906 1157 6964 1183
rect 6906 1123 6918 1157
rect 6952 1123 6964 1157
rect 6906 1097 6964 1123
rect 7006 1157 7064 1183
rect 7006 1123 7018 1157
rect 7052 1123 7064 1157
rect 7006 1097 7064 1123
rect 7106 1157 7164 1183
rect 7106 1123 7118 1157
rect 7152 1123 7164 1157
rect 7106 1097 7164 1123
rect 7206 1157 7264 1183
rect 7206 1123 7218 1157
rect 7252 1123 7264 1157
rect 7206 1097 7264 1123
rect 7306 1157 7364 1183
rect 7306 1123 7318 1157
rect 7352 1123 7364 1157
rect 7306 1097 7364 1123
rect 7406 1157 7464 1183
rect 7406 1123 7418 1157
rect 7452 1123 7464 1157
rect 7406 1097 7464 1123
rect 7506 1157 7564 1183
rect 7506 1123 7518 1157
rect 7552 1123 7564 1157
rect 7506 1097 7564 1123
rect 7606 1157 7664 1183
rect 7606 1123 7618 1157
rect 7652 1123 7664 1157
rect 7606 1097 7664 1123
rect 7706 1157 7764 1183
rect 7706 1123 7718 1157
rect 7752 1123 7764 1157
rect 7706 1097 7764 1123
rect 7806 1157 7864 1183
rect 7806 1123 7818 1157
rect 7852 1123 7864 1157
rect 7806 1097 7864 1123
rect 7906 1157 7964 1183
rect 7906 1123 7918 1157
rect 7952 1123 7964 1157
rect 7906 1097 7964 1123
rect 8006 1157 8064 1183
rect 8006 1123 8018 1157
rect 8052 1123 8064 1157
rect 8006 1097 8064 1123
rect 8106 1157 8164 1183
rect 8106 1123 8118 1157
rect 8152 1123 8164 1157
rect 8106 1097 8164 1123
rect 8206 1157 8264 1183
rect 8206 1123 8218 1157
rect 8252 1123 8264 1157
rect 8206 1097 8264 1123
rect 8306 1157 8364 1183
rect 8306 1123 8318 1157
rect 8352 1123 8364 1157
rect 8306 1097 8364 1123
rect 8406 1157 8464 1183
rect 8406 1123 8418 1157
rect 8452 1123 8464 1157
rect 8406 1097 8464 1123
rect 8506 1157 8564 1183
rect 8506 1123 8518 1157
rect 8552 1123 8564 1157
rect 8506 1097 8564 1123
rect 8606 1157 8664 1183
rect 8606 1123 8618 1157
rect 8652 1123 8664 1157
rect 8606 1097 8664 1123
rect 8706 1157 8764 1183
rect 8706 1123 8718 1157
rect 8752 1123 8764 1157
rect 8706 1097 8764 1123
rect 8806 1157 8864 1183
rect 8806 1123 8818 1157
rect 8852 1123 8864 1157
rect 8806 1097 8864 1123
rect 8906 1157 8964 1183
rect 8906 1123 8918 1157
rect 8952 1123 8964 1157
rect 8906 1097 8964 1123
rect 9006 1157 9064 1183
rect 9006 1123 9018 1157
rect 9052 1123 9064 1157
rect 9006 1097 9064 1123
rect 9106 1157 9164 1183
rect 9106 1123 9118 1157
rect 9152 1123 9164 1157
rect 9106 1097 9164 1123
rect 9206 1157 9264 1183
rect 9206 1123 9218 1157
rect 9252 1123 9264 1157
rect 9206 1097 9264 1123
rect 9306 1157 9364 1183
rect 9306 1123 9318 1157
rect 9352 1123 9364 1157
rect 9306 1097 9364 1123
rect 9406 1157 9464 1183
rect 9406 1123 9418 1157
rect 9452 1123 9464 1157
rect 9406 1097 9464 1123
rect 9506 1157 9564 1183
rect 9506 1123 9518 1157
rect 9552 1123 9564 1157
rect 9506 1097 9564 1123
rect 9606 1157 9664 1183
rect 9606 1123 9612 1157
rect 9652 1123 9664 1157
rect 9606 1097 9664 1123
rect 9706 1157 9764 1183
rect 9706 1123 9718 1157
rect 9758 1123 9764 1157
rect 9706 1097 9764 1123
rect 9806 1157 9864 1183
rect 9806 1123 9818 1157
rect 9852 1123 9864 1157
rect 9806 1097 9864 1123
rect 9906 1157 9964 1183
rect 9906 1123 9918 1157
rect 9952 1123 9964 1157
rect 9906 1097 9964 1123
rect 10006 1157 10064 1183
rect 10006 1123 10018 1157
rect 10052 1123 10064 1157
rect 10006 1097 10064 1123
rect 10106 1157 10164 1183
rect 10106 1123 10118 1157
rect 10152 1123 10164 1157
rect 10106 1097 10164 1123
rect 10206 1157 10264 1183
rect 10206 1123 10218 1157
rect 10252 1123 10264 1157
rect 10206 1097 10264 1123
rect 10306 1157 10364 1183
rect 10306 1123 10318 1157
rect 10352 1123 10364 1157
rect 10306 1097 10364 1123
rect 10406 1157 10464 1183
rect 10406 1123 10418 1157
rect 10452 1123 10464 1157
rect 10406 1097 10464 1123
rect 10506 1157 10564 1183
rect 10506 1123 10518 1157
rect 10552 1123 10564 1157
rect 10506 1097 10564 1123
rect 10606 1157 10664 1183
rect 10606 1123 10618 1157
rect 10652 1123 10664 1157
rect 10606 1097 10664 1123
rect 10706 1157 10764 1183
rect 10706 1123 10718 1157
rect 10752 1123 10764 1157
rect 10706 1097 10764 1123
rect 10806 1157 10864 1183
rect 10806 1123 10818 1157
rect 10852 1123 10864 1157
rect 10806 1097 10864 1123
rect 10906 1157 10964 1183
rect 10906 1123 10918 1157
rect 10952 1123 10964 1157
rect 10906 1097 10964 1123
rect 11006 1157 11064 1183
rect 11006 1123 11012 1157
rect 11052 1123 11064 1157
rect 11006 1097 11064 1123
rect 11106 1157 11164 1183
rect 11106 1123 11118 1157
rect 11158 1123 11164 1157
rect 11106 1097 11164 1123
rect 11206 1157 11264 1183
rect 11206 1123 11212 1157
rect 11252 1123 11264 1157
rect 11206 1097 11264 1123
rect 11306 1157 11364 1183
rect 11306 1123 11318 1157
rect 11358 1123 11364 1157
rect 11306 1097 11364 1123
rect 11406 1157 11464 1183
rect 11406 1123 11412 1157
rect 11452 1123 11464 1157
rect 11406 1097 11464 1123
rect 11506 1157 11564 1183
rect 11506 1123 11518 1157
rect 11558 1123 11564 1157
rect 11506 1097 11564 1123
rect 11606 1157 11664 1183
rect 11606 1123 11618 1157
rect 11652 1123 11664 1157
rect 11606 1097 11664 1123
rect 11706 1157 11764 1183
rect 11706 1123 11718 1157
rect 11752 1123 11764 1157
rect 11706 1097 11764 1123
rect 11806 1157 11864 1183
rect 11806 1123 11818 1157
rect 11852 1123 11864 1157
rect 11806 1097 11864 1123
rect 11906 1157 11964 1183
rect 11906 1123 11918 1157
rect 11952 1123 11964 1157
rect 11906 1097 11964 1123
rect 12006 1157 12064 1183
rect 12006 1123 12012 1157
rect 12052 1123 12064 1157
rect 12006 1097 12064 1123
rect 12106 1157 12164 1183
rect 12106 1123 12118 1157
rect 12158 1123 12164 1157
rect 12106 1097 12164 1123
rect 12206 1157 12264 1183
rect 12206 1123 12218 1157
rect 12252 1123 12264 1157
rect 12206 1097 12264 1123
rect 12306 1157 12364 1183
rect 12306 1123 12318 1157
rect 12352 1123 12364 1157
rect 12306 1097 12364 1123
rect 12406 1157 12464 1183
rect 12406 1123 12418 1157
rect 12452 1123 12464 1157
rect 12406 1097 12464 1123
rect 12506 1157 12564 1183
rect 12506 1123 12518 1157
rect 12552 1123 12564 1157
rect 12506 1097 12564 1123
rect 12606 1157 12664 1183
rect 12606 1123 12612 1157
rect 12652 1123 12664 1157
rect 12606 1097 12664 1123
rect 12706 1157 12764 1183
rect 12706 1123 12718 1157
rect 12758 1123 12764 1157
rect 12706 1097 12764 1123
rect 12806 1157 12864 1183
rect 13018 1176 13262 1210
rect 12806 1123 12812 1157
rect 12852 1123 12864 1157
rect 12908 1138 12916 1172
rect 12958 1138 12974 1172
rect 13018 1157 13052 1176
rect 12806 1097 12864 1123
rect 13228 1173 13262 1176
rect 13228 1157 13362 1173
rect 13018 1107 13052 1123
rect 13096 1108 13112 1142
rect 13154 1108 13162 1142
rect 13262 1123 13328 1157
rect 13228 1107 13362 1123
rect 13428 1157 13562 1173
rect 13462 1123 13528 1157
rect 13428 1107 13562 1123
rect 13628 1157 13662 1173
rect 13628 1107 13662 1123
rect 6 1017 64 1043
rect 6 983 18 1017
rect 58 983 64 1017
rect 6 957 64 983
rect 106 1017 164 1043
rect 106 983 112 1017
rect 152 983 164 1017
rect 106 957 164 983
rect 206 1017 264 1043
rect 206 983 218 1017
rect 258 983 264 1017
rect 206 957 264 983
rect 306 1017 364 1043
rect 306 983 318 1017
rect 352 983 364 1017
rect 306 957 364 983
rect 406 1017 464 1043
rect 406 983 418 1017
rect 452 983 464 1017
rect 406 957 464 983
rect 506 1017 564 1043
rect 506 983 518 1017
rect 552 983 564 1017
rect 506 957 564 983
rect 606 1017 664 1043
rect 606 983 612 1017
rect 652 983 664 1017
rect 606 957 664 983
rect 706 1017 764 1043
rect 706 983 718 1017
rect 758 983 764 1017
rect 706 957 764 983
rect 806 1017 864 1043
rect 806 983 818 1017
rect 852 983 864 1017
rect 806 957 864 983
rect 906 1017 964 1043
rect 906 983 918 1017
rect 952 983 964 1017
rect 906 957 964 983
rect 1006 1017 1064 1043
rect 1006 983 1018 1017
rect 1052 983 1064 1017
rect 1006 957 1064 983
rect 1106 1017 1164 1043
rect 1106 983 1118 1017
rect 1152 983 1164 1017
rect 1106 957 1164 983
rect 1206 1017 1264 1043
rect 1206 983 1212 1017
rect 1252 983 1264 1017
rect 1206 957 1264 983
rect 1306 1017 1364 1043
rect 1306 983 1318 1017
rect 1358 983 1364 1017
rect 1306 957 1364 983
rect 1406 1017 1464 1043
rect 1406 983 1418 1017
rect 1452 983 1464 1017
rect 1406 957 1464 983
rect 1506 1017 1564 1043
rect 1506 983 1518 1017
rect 1552 983 1564 1017
rect 1506 957 1564 983
rect 1606 1017 1664 1043
rect 1606 983 1618 1017
rect 1652 983 1664 1017
rect 1606 957 1664 983
rect 1706 1017 1764 1043
rect 1706 983 1718 1017
rect 1752 983 1764 1017
rect 1706 957 1764 983
rect 1806 1017 1864 1043
rect 1806 983 1818 1017
rect 1852 983 1864 1017
rect 1806 957 1864 983
rect 1906 1017 1964 1043
rect 1906 983 1918 1017
rect 1952 983 1964 1017
rect 1906 957 1964 983
rect 2006 1017 2064 1043
rect 2006 983 2018 1017
rect 2052 983 2064 1017
rect 2006 957 2064 983
rect 2106 1017 2164 1043
rect 2106 983 2118 1017
rect 2152 983 2164 1017
rect 2106 957 2164 983
rect 2206 1017 2264 1043
rect 2206 983 2218 1017
rect 2252 983 2264 1017
rect 2206 957 2264 983
rect 2306 1017 2364 1043
rect 2306 983 2318 1017
rect 2352 983 2364 1017
rect 2306 957 2364 983
rect 2406 1017 2464 1043
rect 2406 983 2418 1017
rect 2452 983 2464 1017
rect 2406 957 2464 983
rect 2506 1017 2564 1043
rect 2506 983 2518 1017
rect 2552 983 2564 1017
rect 2506 957 2564 983
rect 2606 1017 2664 1043
rect 2606 983 2612 1017
rect 2652 983 2664 1017
rect 2606 957 2664 983
rect 2706 1017 2764 1043
rect 2706 983 2718 1017
rect 2758 983 2764 1017
rect 2706 957 2764 983
rect 2806 1017 2864 1043
rect 2806 983 2812 1017
rect 2852 983 2864 1017
rect 2806 957 2864 983
rect 2906 1017 2964 1043
rect 2906 983 2918 1017
rect 2958 983 2964 1017
rect 2906 957 2964 983
rect 3006 1017 3064 1043
rect 3006 983 3018 1017
rect 3052 983 3064 1017
rect 3006 957 3064 983
rect 3106 1017 3164 1043
rect 3106 983 3112 1017
rect 3152 983 3164 1017
rect 3106 957 3164 983
rect 3206 1017 3264 1043
rect 3206 983 3218 1017
rect 3258 983 3264 1017
rect 3206 957 3264 983
rect 3306 1017 3364 1043
rect 3306 983 3312 1017
rect 3352 983 3364 1017
rect 3306 957 3364 983
rect 3406 1017 3464 1043
rect 3406 983 3418 1017
rect 3458 983 3464 1017
rect 3406 957 3464 983
rect 3506 1017 3564 1043
rect 3506 983 3518 1017
rect 3552 983 3564 1017
rect 3506 957 3564 983
rect 3606 1017 3664 1043
rect 3606 983 3612 1017
rect 3652 983 3664 1017
rect 3606 957 3664 983
rect 3706 1017 3764 1043
rect 3706 983 3718 1017
rect 3758 983 3764 1017
rect 3706 957 3764 983
rect 3806 1017 3864 1043
rect 3806 983 3812 1017
rect 3852 983 3864 1017
rect 3806 957 3864 983
rect 3906 1017 3964 1043
rect 3906 983 3918 1017
rect 3958 983 3964 1017
rect 3906 957 3964 983
rect 4006 1017 4064 1043
rect 4006 983 4018 1017
rect 4052 983 4064 1017
rect 4006 957 4064 983
rect 4106 1017 4164 1043
rect 4106 983 4118 1017
rect 4152 983 4164 1017
rect 4106 957 4164 983
rect 4206 1017 4264 1043
rect 4206 983 4218 1017
rect 4252 983 4264 1017
rect 4206 957 4264 983
rect 4306 1017 4364 1043
rect 4306 983 4318 1017
rect 4352 983 4364 1017
rect 4306 957 4364 983
rect 4406 1017 4464 1043
rect 4406 983 4418 1017
rect 4452 983 4464 1017
rect 4406 957 4464 983
rect 4506 1017 4564 1043
rect 4506 983 4518 1017
rect 4552 983 4564 1017
rect 4506 957 4564 983
rect 4606 1017 4664 1043
rect 4606 983 4618 1017
rect 4652 983 4664 1017
rect 4606 957 4664 983
rect 4706 1017 4764 1043
rect 4706 983 4718 1017
rect 4752 983 4764 1017
rect 4706 957 4764 983
rect 4806 1017 4864 1043
rect 4806 983 4812 1017
rect 4852 983 4864 1017
rect 4806 957 4864 983
rect 4906 1017 4964 1043
rect 4906 983 4918 1017
rect 4958 983 4964 1017
rect 4906 957 4964 983
rect 5006 1017 5064 1043
rect 5006 983 5018 1017
rect 5052 983 5064 1017
rect 5006 957 5064 983
rect 5106 1017 5164 1043
rect 5106 983 5118 1017
rect 5152 983 5164 1017
rect 5106 957 5164 983
rect 5206 1017 5264 1043
rect 5206 983 5218 1017
rect 5252 983 5264 1017
rect 5206 957 5264 983
rect 5306 1017 5364 1043
rect 5306 983 5312 1017
rect 5352 983 5364 1017
rect 5306 957 5364 983
rect 5406 1017 5464 1043
rect 5406 983 5418 1017
rect 5458 983 5464 1017
rect 5406 957 5464 983
rect 5506 1017 5564 1043
rect 5506 983 5518 1017
rect 5552 983 5564 1017
rect 5506 957 5564 983
rect 5606 1017 5664 1043
rect 5606 983 5618 1017
rect 5652 983 5664 1017
rect 5606 957 5664 983
rect 5706 1017 5764 1043
rect 5706 983 5718 1017
rect 5752 983 5764 1017
rect 5706 957 5764 983
rect 5806 1017 5864 1043
rect 5806 983 5818 1017
rect 5852 983 5864 1017
rect 5806 957 5864 983
rect 5906 1017 5964 1043
rect 5906 983 5918 1017
rect 5952 983 5964 1017
rect 5906 957 5964 983
rect 6006 1017 6064 1043
rect 6006 983 6018 1017
rect 6052 983 6064 1017
rect 6006 957 6064 983
rect 6106 1017 6164 1043
rect 6106 983 6118 1017
rect 6152 983 6164 1017
rect 6106 957 6164 983
rect 6206 1017 6264 1043
rect 6206 983 6218 1017
rect 6252 983 6264 1017
rect 6206 957 6264 983
rect 6306 1017 6364 1043
rect 6306 983 6318 1017
rect 6352 983 6364 1017
rect 6306 957 6364 983
rect 6406 1017 6464 1043
rect 6406 983 6412 1017
rect 6452 983 6464 1017
rect 6406 957 6464 983
rect 6506 1017 6564 1043
rect 6506 983 6518 1017
rect 6558 983 6564 1017
rect 6506 957 6564 983
rect 6606 1017 6664 1043
rect 6606 983 6618 1017
rect 6652 983 6664 1017
rect 6606 957 6664 983
rect 6706 1017 6764 1043
rect 6706 983 6718 1017
rect 6752 983 6764 1017
rect 6706 957 6764 983
rect 6806 1017 6864 1043
rect 6806 983 6818 1017
rect 6852 983 6864 1017
rect 6806 957 6864 983
rect 6906 1017 6964 1043
rect 6906 983 6912 1017
rect 6952 983 6964 1017
rect 6906 957 6964 983
rect 7006 1017 7064 1043
rect 7006 983 7018 1017
rect 7058 983 7064 1017
rect 7006 957 7064 983
rect 7106 1017 7164 1043
rect 7106 983 7112 1017
rect 7152 983 7164 1017
rect 7106 957 7164 983
rect 7206 1017 7264 1043
rect 7206 983 7218 1017
rect 7258 983 7264 1017
rect 7206 957 7264 983
rect 7306 1017 7364 1043
rect 7306 983 7312 1017
rect 7352 983 7364 1017
rect 7306 957 7364 983
rect 7406 1017 7464 1043
rect 7406 983 7418 1017
rect 7458 983 7464 1017
rect 7406 957 7464 983
rect 7506 1017 7564 1043
rect 7506 983 7518 1017
rect 7552 983 7564 1017
rect 7506 957 7564 983
rect 7606 1017 7664 1043
rect 7606 983 7618 1017
rect 7652 983 7664 1017
rect 7606 957 7664 983
rect 7706 1017 7764 1043
rect 7706 983 7718 1017
rect 7752 983 7764 1017
rect 7706 957 7764 983
rect 7806 1017 7864 1043
rect 7806 983 7818 1017
rect 7852 983 7864 1017
rect 7806 957 7864 983
rect 7906 1017 7964 1043
rect 7906 983 7918 1017
rect 7952 983 7964 1017
rect 7906 957 7964 983
rect 8006 1017 8064 1043
rect 8006 983 8018 1017
rect 8052 983 8064 1017
rect 8006 957 8064 983
rect 8106 1017 8164 1043
rect 8106 983 8118 1017
rect 8152 983 8164 1017
rect 8106 957 8164 983
rect 8206 1017 8264 1043
rect 8206 983 8218 1017
rect 8252 983 8264 1017
rect 8206 957 8264 983
rect 8306 1017 8364 1043
rect 8306 983 8318 1017
rect 8352 983 8364 1017
rect 8306 957 8364 983
rect 8406 1017 8464 1043
rect 8406 983 8418 1017
rect 8452 983 8464 1017
rect 8406 957 8464 983
rect 8506 1017 8564 1043
rect 8506 983 8518 1017
rect 8552 983 8564 1017
rect 8506 957 8564 983
rect 8606 1017 8664 1043
rect 8606 983 8612 1017
rect 8652 983 8664 1017
rect 8606 957 8664 983
rect 8706 1017 8764 1043
rect 8706 983 8718 1017
rect 8758 983 8764 1017
rect 8706 957 8764 983
rect 8806 1017 8864 1043
rect 8806 983 8812 1017
rect 8852 983 8864 1017
rect 8806 957 8864 983
rect 8906 1017 8964 1043
rect 8906 983 8918 1017
rect 8958 983 8964 1017
rect 8906 957 8964 983
rect 9006 1017 9064 1043
rect 9006 983 9018 1017
rect 9052 983 9064 1017
rect 9006 957 9064 983
rect 9106 1017 9164 1043
rect 9106 983 9118 1017
rect 9152 983 9164 1017
rect 9106 957 9164 983
rect 9206 1017 9264 1043
rect 9206 983 9218 1017
rect 9252 983 9264 1017
rect 9206 957 9264 983
rect 9306 1017 9364 1043
rect 9306 983 9318 1017
rect 9352 983 9364 1017
rect 9306 957 9364 983
rect 9406 1017 9464 1043
rect 9406 983 9418 1017
rect 9452 983 9464 1017
rect 9406 957 9464 983
rect 9506 1017 9564 1043
rect 9506 983 9512 1017
rect 9552 983 9564 1017
rect 9506 957 9564 983
rect 9606 1017 9664 1043
rect 9606 983 9618 1017
rect 9658 983 9664 1017
rect 9606 957 9664 983
rect 9706 1017 9764 1043
rect 9706 983 9718 1017
rect 9752 983 9764 1017
rect 9706 957 9764 983
rect 9806 1017 9864 1043
rect 9806 983 9818 1017
rect 9852 983 9864 1017
rect 9806 957 9864 983
rect 9906 1017 9964 1043
rect 9906 983 9912 1017
rect 9952 983 9964 1017
rect 9906 957 9964 983
rect 10006 1017 10064 1043
rect 10006 983 10018 1017
rect 10058 983 10064 1017
rect 10006 957 10064 983
rect 10106 1017 10164 1043
rect 10106 983 10118 1017
rect 10152 983 10164 1017
rect 10106 957 10164 983
rect 10206 1017 10264 1043
rect 10206 983 10218 1017
rect 10252 983 10264 1017
rect 10206 957 10264 983
rect 10306 1017 10364 1043
rect 10306 983 10312 1017
rect 10352 983 10364 1017
rect 10306 957 10364 983
rect 10406 1017 10464 1043
rect 10406 983 10418 1017
rect 10458 983 10464 1017
rect 10406 957 10464 983
rect 10506 1017 10564 1043
rect 10506 983 10518 1017
rect 10552 983 10564 1017
rect 10506 957 10564 983
rect 10606 1017 10664 1043
rect 10606 983 10618 1017
rect 10652 983 10664 1017
rect 10606 957 10664 983
rect 10706 1017 10764 1043
rect 10706 983 10718 1017
rect 10752 983 10764 1017
rect 10706 957 10764 983
rect 10806 1017 10864 1043
rect 10806 983 10818 1017
rect 10852 983 10864 1017
rect 10806 957 10864 983
rect 10906 1017 10964 1043
rect 10906 983 10918 1017
rect 10952 983 10964 1017
rect 10906 957 10964 983
rect 11006 1017 11064 1043
rect 11006 983 11018 1017
rect 11052 983 11064 1017
rect 11006 957 11064 983
rect 11106 1017 11164 1043
rect 11106 983 11118 1017
rect 11152 983 11164 1017
rect 11106 957 11164 983
rect 11206 1017 11264 1043
rect 11206 983 11218 1017
rect 11252 983 11264 1017
rect 11206 957 11264 983
rect 11306 1017 11364 1043
rect 11306 983 11312 1017
rect 11352 983 11364 1017
rect 11306 957 11364 983
rect 11406 1017 11464 1043
rect 11406 983 11418 1017
rect 11458 983 11464 1017
rect 11406 957 11464 983
rect 11506 1017 11564 1043
rect 11506 983 11518 1017
rect 11552 983 11564 1017
rect 11506 957 11564 983
rect 11606 1017 11664 1043
rect 11606 983 11612 1017
rect 11652 983 11664 1017
rect 11606 957 11664 983
rect 11706 1017 11764 1043
rect 11706 983 11718 1017
rect 11758 983 11764 1017
rect 11706 957 11764 983
rect 11806 1017 11864 1043
rect 11806 983 11818 1017
rect 11852 983 11864 1017
rect 11806 957 11864 983
rect 11906 1017 11964 1043
rect 11906 983 11912 1017
rect 11952 983 11964 1017
rect 11906 957 11964 983
rect 12006 1017 12064 1043
rect 12006 983 12018 1017
rect 12058 983 12064 1017
rect 12006 957 12064 983
rect 12106 1017 12164 1043
rect 12106 983 12118 1017
rect 12152 983 12164 1017
rect 12106 957 12164 983
rect 12206 1017 12264 1043
rect 12206 983 12218 1017
rect 12252 983 12264 1017
rect 12206 957 12264 983
rect 12306 1017 12364 1043
rect 12306 983 12318 1017
rect 12352 983 12364 1017
rect 12306 957 12364 983
rect 12406 1017 12464 1043
rect 12406 983 12418 1017
rect 12452 983 12464 1017
rect 12406 957 12464 983
rect 12506 1017 12564 1043
rect 12506 983 12518 1017
rect 12552 983 12564 1017
rect 12506 957 12564 983
rect 12606 1017 12664 1043
rect 12606 983 12618 1017
rect 12652 983 12664 1017
rect 12606 957 12664 983
rect 12706 1017 12764 1043
rect 12706 983 12718 1017
rect 12752 983 12764 1017
rect 12706 957 12764 983
rect 12806 1017 12864 1043
rect 13018 1036 13262 1070
rect 12806 983 12812 1017
rect 12852 983 12864 1017
rect 12908 998 12916 1032
rect 12958 998 12974 1032
rect 13018 1017 13052 1036
rect 12806 957 12864 983
rect 13228 1017 13262 1036
rect 13018 967 13052 983
rect 13096 968 13112 1002
rect 13154 968 13162 1002
rect 13228 967 13262 983
rect 13328 1017 13562 1033
rect 13362 983 13428 1017
rect 13462 983 13528 1017
rect 13328 967 13562 983
rect 13628 1017 13662 1033
rect 13628 967 13662 983
rect 6 877 64 903
rect 6 843 18 877
rect 58 843 64 877
rect 6 817 64 843
rect 106 877 164 903
rect 106 843 112 877
rect 152 843 164 877
rect 106 817 164 843
rect 206 877 264 903
rect 206 843 218 877
rect 258 843 264 877
rect 206 817 264 843
rect 306 877 364 903
rect 306 843 318 877
rect 352 843 364 877
rect 306 817 364 843
rect 406 877 464 903
rect 406 843 418 877
rect 452 843 464 877
rect 406 817 464 843
rect 506 877 564 903
rect 506 843 518 877
rect 552 843 564 877
rect 506 817 564 843
rect 606 877 664 903
rect 606 843 618 877
rect 652 843 664 877
rect 606 817 664 843
rect 706 877 764 903
rect 706 843 718 877
rect 752 843 764 877
rect 706 817 764 843
rect 806 877 864 903
rect 806 843 818 877
rect 852 843 864 877
rect 806 817 864 843
rect 906 877 964 903
rect 906 843 918 877
rect 952 843 964 877
rect 906 817 964 843
rect 1006 877 1064 903
rect 1006 843 1018 877
rect 1052 843 1064 877
rect 1006 817 1064 843
rect 1106 877 1164 903
rect 1106 843 1118 877
rect 1152 843 1164 877
rect 1106 817 1164 843
rect 1206 877 1264 903
rect 1206 843 1218 877
rect 1252 843 1264 877
rect 1206 817 1264 843
rect 1306 877 1364 903
rect 1306 843 1318 877
rect 1352 843 1364 877
rect 1306 817 1364 843
rect 1406 877 1464 903
rect 1406 843 1418 877
rect 1452 843 1464 877
rect 1406 817 1464 843
rect 1506 877 1564 903
rect 1506 843 1518 877
rect 1552 843 1564 877
rect 1506 817 1564 843
rect 1606 877 1664 903
rect 1606 843 1618 877
rect 1652 843 1664 877
rect 1606 817 1664 843
rect 1706 877 1764 903
rect 1706 843 1718 877
rect 1752 843 1764 877
rect 1706 817 1764 843
rect 1806 877 1864 903
rect 1806 843 1818 877
rect 1852 843 1864 877
rect 1806 817 1864 843
rect 1906 877 1964 903
rect 1906 843 1918 877
rect 1952 843 1964 877
rect 1906 817 1964 843
rect 2006 877 2064 903
rect 2006 843 2018 877
rect 2052 843 2064 877
rect 2006 817 2064 843
rect 2106 877 2164 903
rect 2106 843 2118 877
rect 2152 843 2164 877
rect 2106 817 2164 843
rect 2206 877 2264 903
rect 2206 843 2218 877
rect 2252 843 2264 877
rect 2206 817 2264 843
rect 2306 877 2364 903
rect 2306 843 2318 877
rect 2352 843 2364 877
rect 2306 817 2364 843
rect 2406 877 2464 903
rect 2406 843 2418 877
rect 2452 843 2464 877
rect 2406 817 2464 843
rect 2506 877 2564 903
rect 2506 843 2518 877
rect 2552 843 2564 877
rect 2506 817 2564 843
rect 2606 877 2664 903
rect 2606 843 2618 877
rect 2652 843 2664 877
rect 2606 817 2664 843
rect 2706 877 2764 903
rect 2706 843 2718 877
rect 2752 843 2764 877
rect 2706 817 2764 843
rect 2806 877 2864 903
rect 2806 843 2818 877
rect 2852 843 2864 877
rect 2806 817 2864 843
rect 2906 877 2964 903
rect 2906 843 2912 877
rect 2952 843 2964 877
rect 2906 817 2964 843
rect 3006 877 3064 903
rect 3006 843 3018 877
rect 3058 843 3064 877
rect 3006 817 3064 843
rect 3106 877 3164 903
rect 3106 843 3118 877
rect 3152 843 3164 877
rect 3106 817 3164 843
rect 3206 877 3264 903
rect 3206 843 3218 877
rect 3252 843 3264 877
rect 3206 817 3264 843
rect 3306 877 3364 903
rect 3306 843 3318 877
rect 3352 843 3364 877
rect 3306 817 3364 843
rect 3406 877 3464 903
rect 3406 843 3418 877
rect 3452 843 3464 877
rect 3406 817 3464 843
rect 3506 877 3564 903
rect 3506 843 3518 877
rect 3552 843 3564 877
rect 3506 817 3564 843
rect 3606 877 3664 903
rect 3606 843 3618 877
rect 3652 843 3664 877
rect 3606 817 3664 843
rect 3706 877 3764 903
rect 3706 843 3718 877
rect 3752 843 3764 877
rect 3706 817 3764 843
rect 3806 877 3864 903
rect 3806 843 3812 877
rect 3852 843 3864 877
rect 3806 817 3864 843
rect 3906 877 3964 903
rect 3906 843 3918 877
rect 3958 843 3964 877
rect 3906 817 3964 843
rect 4006 877 4064 903
rect 4006 843 4018 877
rect 4052 843 4064 877
rect 4006 817 4064 843
rect 4106 877 4164 903
rect 4106 843 4118 877
rect 4152 843 4164 877
rect 4106 817 4164 843
rect 4206 877 4264 903
rect 4206 843 4218 877
rect 4252 843 4264 877
rect 4206 817 4264 843
rect 4306 877 4364 903
rect 4306 843 4318 877
rect 4352 843 4364 877
rect 4306 817 4364 843
rect 4406 877 4464 903
rect 4406 843 4418 877
rect 4452 843 4464 877
rect 4406 817 4464 843
rect 4506 877 4564 903
rect 4506 843 4518 877
rect 4552 843 4564 877
rect 4506 817 4564 843
rect 4606 877 4664 903
rect 4606 843 4618 877
rect 4652 843 4664 877
rect 4606 817 4664 843
rect 4706 877 4764 903
rect 4706 843 4718 877
rect 4752 843 4764 877
rect 4706 817 4764 843
rect 4806 877 4864 903
rect 4806 843 4818 877
rect 4852 843 4864 877
rect 4806 817 4864 843
rect 4906 877 4964 903
rect 4906 843 4918 877
rect 4952 843 4964 877
rect 4906 817 4964 843
rect 5006 877 5064 903
rect 5006 843 5018 877
rect 5052 843 5064 877
rect 5006 817 5064 843
rect 5106 877 5164 903
rect 5106 843 5118 877
rect 5152 843 5164 877
rect 5106 817 5164 843
rect 5206 877 5264 903
rect 5206 843 5218 877
rect 5252 843 5264 877
rect 5206 817 5264 843
rect 5306 877 5364 903
rect 5306 843 5318 877
rect 5352 843 5364 877
rect 5306 817 5364 843
rect 5406 877 5464 903
rect 5406 843 5418 877
rect 5452 843 5464 877
rect 5406 817 5464 843
rect 5506 877 5564 903
rect 5506 843 5518 877
rect 5552 843 5564 877
rect 5506 817 5564 843
rect 5606 877 5664 903
rect 5606 843 5618 877
rect 5652 843 5664 877
rect 5606 817 5664 843
rect 5706 877 5764 903
rect 5706 843 5718 877
rect 5752 843 5764 877
rect 5706 817 5764 843
rect 5806 877 5864 903
rect 5806 843 5818 877
rect 5852 843 5864 877
rect 5806 817 5864 843
rect 5906 877 5964 903
rect 5906 843 5918 877
rect 5952 843 5964 877
rect 5906 817 5964 843
rect 6006 877 6064 903
rect 6006 843 6018 877
rect 6052 843 6064 877
rect 6006 817 6064 843
rect 6106 877 6164 903
rect 6106 843 6118 877
rect 6152 843 6164 877
rect 6106 817 6164 843
rect 6206 877 6264 903
rect 6206 843 6218 877
rect 6252 843 6264 877
rect 6206 817 6264 843
rect 6306 877 6364 903
rect 6306 843 6318 877
rect 6352 843 6364 877
rect 6306 817 6364 843
rect 6406 877 6464 903
rect 6406 843 6418 877
rect 6452 843 6464 877
rect 6406 817 6464 843
rect 6506 877 6564 903
rect 6506 843 6518 877
rect 6552 843 6564 877
rect 6506 817 6564 843
rect 6606 877 6664 903
rect 6606 843 6612 877
rect 6652 843 6664 877
rect 6606 817 6664 843
rect 6706 877 6764 903
rect 6706 843 6718 877
rect 6758 843 6764 877
rect 6706 817 6764 843
rect 6806 877 6864 903
rect 6806 843 6818 877
rect 6852 843 6864 877
rect 6806 817 6864 843
rect 6906 877 6964 903
rect 6906 843 6918 877
rect 6952 843 6964 877
rect 6906 817 6964 843
rect 7006 877 7064 903
rect 7006 843 7018 877
rect 7052 843 7064 877
rect 7006 817 7064 843
rect 7106 877 7164 903
rect 7106 843 7118 877
rect 7152 843 7164 877
rect 7106 817 7164 843
rect 7206 877 7264 903
rect 7206 843 7218 877
rect 7252 843 7264 877
rect 7206 817 7264 843
rect 7306 877 7364 903
rect 7306 843 7312 877
rect 7352 843 7364 877
rect 7306 817 7364 843
rect 7406 877 7464 903
rect 7406 843 7418 877
rect 7458 843 7464 877
rect 7406 817 7464 843
rect 7506 877 7564 903
rect 7506 843 7512 877
rect 7552 843 7564 877
rect 7506 817 7564 843
rect 7606 877 7664 903
rect 7606 843 7618 877
rect 7658 843 7664 877
rect 7606 817 7664 843
rect 7706 877 7764 903
rect 7706 843 7712 877
rect 7752 843 7764 877
rect 7706 817 7764 843
rect 7806 877 7864 903
rect 7806 843 7818 877
rect 7858 843 7864 877
rect 7806 817 7864 843
rect 7906 877 7964 903
rect 7906 843 7912 877
rect 7952 843 7964 877
rect 7906 817 7964 843
rect 8006 877 8064 903
rect 8006 843 8018 877
rect 8058 843 8064 877
rect 8006 817 8064 843
rect 8106 877 8164 903
rect 8106 843 8118 877
rect 8152 843 8164 877
rect 8106 817 8164 843
rect 8206 877 8264 903
rect 8206 843 8218 877
rect 8252 843 8264 877
rect 8206 817 8264 843
rect 8306 877 8364 903
rect 8306 843 8318 877
rect 8352 843 8364 877
rect 8306 817 8364 843
rect 8406 877 8464 903
rect 8406 843 8418 877
rect 8452 843 8464 877
rect 8406 817 8464 843
rect 8506 877 8564 903
rect 8506 843 8518 877
rect 8552 843 8564 877
rect 8506 817 8564 843
rect 8606 877 8664 903
rect 8606 843 8612 877
rect 8652 843 8664 877
rect 8606 817 8664 843
rect 8706 877 8764 903
rect 8706 843 8718 877
rect 8758 843 8764 877
rect 8706 817 8764 843
rect 8806 877 8864 903
rect 8806 843 8812 877
rect 8852 843 8864 877
rect 8806 817 8864 843
rect 8906 877 8964 903
rect 8906 843 8918 877
rect 8958 843 8964 877
rect 8906 817 8964 843
rect 9006 877 9064 903
rect 9006 843 9018 877
rect 9052 843 9064 877
rect 9006 817 9064 843
rect 9106 877 9164 903
rect 9106 843 9118 877
rect 9152 843 9164 877
rect 9106 817 9164 843
rect 9206 877 9264 903
rect 9206 843 9218 877
rect 9252 843 9264 877
rect 9206 817 9264 843
rect 9306 877 9364 903
rect 9306 843 9318 877
rect 9352 843 9364 877
rect 9306 817 9364 843
rect 9406 877 9464 903
rect 9406 843 9418 877
rect 9452 843 9464 877
rect 9406 817 9464 843
rect 9506 877 9564 903
rect 9506 843 9518 877
rect 9552 843 9564 877
rect 9506 817 9564 843
rect 9606 877 9664 903
rect 9606 843 9618 877
rect 9652 843 9664 877
rect 9606 817 9664 843
rect 9706 877 9764 903
rect 9706 843 9718 877
rect 9752 843 9764 877
rect 9706 817 9764 843
rect 9806 877 9864 903
rect 9806 843 9818 877
rect 9852 843 9864 877
rect 9806 817 9864 843
rect 9906 877 9964 903
rect 9906 843 9912 877
rect 9952 843 9964 877
rect 9906 817 9964 843
rect 10006 877 10064 903
rect 10006 843 10018 877
rect 10058 843 10064 877
rect 10006 817 10064 843
rect 10106 877 10164 903
rect 10106 843 10118 877
rect 10152 843 10164 877
rect 10106 817 10164 843
rect 10206 877 10264 903
rect 10206 843 10218 877
rect 10252 843 10264 877
rect 10206 817 10264 843
rect 10306 877 10364 903
rect 10306 843 10318 877
rect 10352 843 10364 877
rect 10306 817 10364 843
rect 10406 877 10464 903
rect 10406 843 10418 877
rect 10452 843 10464 877
rect 10406 817 10464 843
rect 10506 877 10564 903
rect 10506 843 10518 877
rect 10552 843 10564 877
rect 10506 817 10564 843
rect 10606 877 10664 903
rect 10606 843 10618 877
rect 10652 843 10664 877
rect 10606 817 10664 843
rect 10706 877 10764 903
rect 10706 843 10712 877
rect 10752 843 10764 877
rect 10706 817 10764 843
rect 10806 877 10864 903
rect 10806 843 10818 877
rect 10858 843 10864 877
rect 10806 817 10864 843
rect 10906 877 10964 903
rect 10906 843 10912 877
rect 10952 843 10964 877
rect 10906 817 10964 843
rect 11006 877 11064 903
rect 11006 843 11018 877
rect 11058 843 11064 877
rect 11006 817 11064 843
rect 11106 877 11164 903
rect 11106 843 11118 877
rect 11152 843 11164 877
rect 11106 817 11164 843
rect 11206 877 11264 903
rect 11206 843 11218 877
rect 11252 843 11264 877
rect 11206 817 11264 843
rect 11306 877 11364 903
rect 11306 843 11318 877
rect 11352 843 11364 877
rect 11306 817 11364 843
rect 11406 877 11464 903
rect 11406 843 11418 877
rect 11452 843 11464 877
rect 11406 817 11464 843
rect 11506 877 11564 903
rect 11506 843 11518 877
rect 11552 843 11564 877
rect 11506 817 11564 843
rect 11606 877 11664 903
rect 11606 843 11618 877
rect 11652 843 11664 877
rect 11606 817 11664 843
rect 11706 877 11764 903
rect 11706 843 11718 877
rect 11752 843 11764 877
rect 11706 817 11764 843
rect 11806 877 11864 903
rect 11806 843 11818 877
rect 11852 843 11864 877
rect 11806 817 11864 843
rect 11906 877 11964 903
rect 11906 843 11912 877
rect 11952 843 11964 877
rect 11906 817 11964 843
rect 12006 877 12064 903
rect 12006 843 12018 877
rect 12058 843 12064 877
rect 12006 817 12064 843
rect 12106 877 12164 903
rect 12106 843 12118 877
rect 12152 843 12164 877
rect 12106 817 12164 843
rect 12206 877 12264 903
rect 12206 843 12218 877
rect 12252 843 12264 877
rect 12206 817 12264 843
rect 12306 877 12364 903
rect 12306 843 12312 877
rect 12352 843 12364 877
rect 12306 817 12364 843
rect 12406 877 12464 903
rect 12406 843 12418 877
rect 12458 843 12464 877
rect 12406 817 12464 843
rect 12506 877 12564 903
rect 12506 843 12512 877
rect 12552 843 12564 877
rect 12506 817 12564 843
rect 12606 877 12664 903
rect 12606 843 12618 877
rect 12658 843 12664 877
rect 12606 817 12664 843
rect 12706 877 12764 903
rect 12706 843 12718 877
rect 12752 843 12764 877
rect 12706 817 12764 843
rect 12806 877 12864 903
rect 13018 896 13262 930
rect 12806 843 12818 877
rect 12852 843 12864 877
rect 12908 858 12916 892
rect 12958 858 12974 892
rect 13018 877 13052 896
rect 12806 817 12864 843
rect 13228 893 13262 896
rect 13228 877 13362 893
rect 13018 827 13052 843
rect 13096 828 13112 862
rect 13154 828 13162 862
rect 13262 843 13328 877
rect 13228 827 13362 843
rect 13428 877 13462 893
rect 13428 827 13462 843
rect 13528 877 13662 893
rect 13562 843 13628 877
rect 13528 827 13662 843
rect 6 737 64 763
rect 6 703 18 737
rect 52 703 64 737
rect 6 677 64 703
rect 106 737 164 763
rect 106 703 118 737
rect 152 703 164 737
rect 106 677 164 703
rect 206 737 264 763
rect 206 703 218 737
rect 252 703 264 737
rect 206 677 264 703
rect 306 737 364 763
rect 306 703 318 737
rect 352 703 364 737
rect 306 677 364 703
rect 406 737 464 763
rect 406 703 418 737
rect 452 703 464 737
rect 406 677 464 703
rect 506 737 564 763
rect 506 703 512 737
rect 552 703 564 737
rect 506 677 564 703
rect 606 737 664 763
rect 606 703 618 737
rect 658 703 664 737
rect 606 677 664 703
rect 706 737 764 763
rect 706 703 712 737
rect 752 703 764 737
rect 706 677 764 703
rect 806 737 864 763
rect 806 703 818 737
rect 858 703 864 737
rect 806 677 864 703
rect 906 737 964 763
rect 906 703 918 737
rect 952 703 964 737
rect 906 677 964 703
rect 1006 737 1064 763
rect 1006 703 1018 737
rect 1052 703 1064 737
rect 1006 677 1064 703
rect 1106 737 1164 763
rect 1106 703 1118 737
rect 1152 703 1164 737
rect 1106 677 1164 703
rect 1206 737 1264 763
rect 1206 703 1212 737
rect 1252 703 1264 737
rect 1206 677 1264 703
rect 1306 737 1364 763
rect 1306 703 1318 737
rect 1358 703 1364 737
rect 1306 677 1364 703
rect 1406 737 1464 763
rect 1406 703 1412 737
rect 1452 703 1464 737
rect 1406 677 1464 703
rect 1506 737 1564 763
rect 1506 703 1518 737
rect 1558 703 1564 737
rect 1506 677 1564 703
rect 1606 737 1664 763
rect 1606 703 1618 737
rect 1652 703 1664 737
rect 1606 677 1664 703
rect 1706 737 1764 763
rect 1706 703 1718 737
rect 1752 703 1764 737
rect 1706 677 1764 703
rect 1806 737 1864 763
rect 1806 703 1818 737
rect 1852 703 1864 737
rect 1806 677 1864 703
rect 1906 737 1964 763
rect 1906 703 1918 737
rect 1952 703 1964 737
rect 1906 677 1964 703
rect 2006 737 2064 763
rect 2006 703 2012 737
rect 2052 703 2064 737
rect 2006 677 2064 703
rect 2106 737 2164 763
rect 2106 703 2118 737
rect 2158 703 2164 737
rect 2106 677 2164 703
rect 2206 737 2264 763
rect 2206 703 2218 737
rect 2252 703 2264 737
rect 2206 677 2264 703
rect 2306 737 2364 763
rect 2306 703 2318 737
rect 2352 703 2364 737
rect 2306 677 2364 703
rect 2406 737 2464 763
rect 2406 703 2412 737
rect 2452 703 2464 737
rect 2406 677 2464 703
rect 2506 737 2564 763
rect 2506 703 2518 737
rect 2558 703 2564 737
rect 2506 677 2564 703
rect 2606 737 2664 763
rect 2606 703 2618 737
rect 2652 703 2664 737
rect 2606 677 2664 703
rect 2706 737 2764 763
rect 2706 703 2718 737
rect 2752 703 2764 737
rect 2706 677 2764 703
rect 2806 737 2864 763
rect 2806 703 2812 737
rect 2852 703 2864 737
rect 2806 677 2864 703
rect 2906 737 2964 763
rect 2906 703 2918 737
rect 2958 703 2964 737
rect 2906 677 2964 703
rect 3006 737 3064 763
rect 3006 703 3012 737
rect 3052 703 3064 737
rect 3006 677 3064 703
rect 3106 737 3164 763
rect 3106 703 3118 737
rect 3158 703 3164 737
rect 3106 677 3164 703
rect 3206 737 3264 763
rect 3206 703 3218 737
rect 3252 703 3264 737
rect 3206 677 3264 703
rect 3306 737 3364 763
rect 3306 703 3312 737
rect 3352 703 3364 737
rect 3306 677 3364 703
rect 3406 737 3464 763
rect 3406 703 3418 737
rect 3458 703 3464 737
rect 3406 677 3464 703
rect 3506 737 3564 763
rect 3506 703 3518 737
rect 3552 703 3564 737
rect 3506 677 3564 703
rect 3606 737 3664 763
rect 3606 703 3612 737
rect 3652 703 3664 737
rect 3606 677 3664 703
rect 3706 737 3764 763
rect 3706 703 3718 737
rect 3758 703 3764 737
rect 3706 677 3764 703
rect 3806 737 3864 763
rect 3806 703 3818 737
rect 3852 703 3864 737
rect 3806 677 3864 703
rect 3906 737 3964 763
rect 3906 703 3918 737
rect 3952 703 3964 737
rect 3906 677 3964 703
rect 4006 737 4064 763
rect 4006 703 4018 737
rect 4052 703 4064 737
rect 4006 677 4064 703
rect 4106 737 4164 763
rect 4106 703 4118 737
rect 4152 703 4164 737
rect 4106 677 4164 703
rect 4206 737 4264 763
rect 4206 703 4218 737
rect 4252 703 4264 737
rect 4206 677 4264 703
rect 4306 737 4364 763
rect 4306 703 4318 737
rect 4352 703 4364 737
rect 4306 677 4364 703
rect 4406 737 4464 763
rect 4406 703 4418 737
rect 4452 703 4464 737
rect 4406 677 4464 703
rect 4506 737 4564 763
rect 4506 703 4518 737
rect 4552 703 4564 737
rect 4506 677 4564 703
rect 4606 737 4664 763
rect 4606 703 4612 737
rect 4652 703 4664 737
rect 4606 677 4664 703
rect 4706 737 4764 763
rect 4706 703 4718 737
rect 4758 703 4764 737
rect 4706 677 4764 703
rect 4806 737 4864 763
rect 4806 703 4818 737
rect 4852 703 4864 737
rect 4806 677 4864 703
rect 4906 737 4964 763
rect 4906 703 4918 737
rect 4952 703 4964 737
rect 4906 677 4964 703
rect 5006 737 5064 763
rect 5006 703 5018 737
rect 5052 703 5064 737
rect 5006 677 5064 703
rect 5106 737 5164 763
rect 5106 703 5112 737
rect 5152 703 5164 737
rect 5106 677 5164 703
rect 5206 737 5264 763
rect 5206 703 5218 737
rect 5258 703 5264 737
rect 5206 677 5264 703
rect 5306 737 5364 763
rect 5306 703 5318 737
rect 5352 703 5364 737
rect 5306 677 5364 703
rect 5406 737 5464 763
rect 5406 703 5418 737
rect 5452 703 5464 737
rect 5406 677 5464 703
rect 5506 737 5564 763
rect 5506 703 5518 737
rect 5552 703 5564 737
rect 5506 677 5564 703
rect 5606 737 5664 763
rect 5606 703 5618 737
rect 5652 703 5664 737
rect 5606 677 5664 703
rect 5706 737 5764 763
rect 5706 703 5712 737
rect 5752 703 5764 737
rect 5706 677 5764 703
rect 5806 737 5864 763
rect 5806 703 5818 737
rect 5858 703 5864 737
rect 5806 677 5864 703
rect 5906 737 5964 763
rect 5906 703 5918 737
rect 5952 703 5964 737
rect 5906 677 5964 703
rect 6006 737 6064 763
rect 6006 703 6018 737
rect 6052 703 6064 737
rect 6006 677 6064 703
rect 6106 737 6164 763
rect 6106 703 6118 737
rect 6152 703 6164 737
rect 6106 677 6164 703
rect 6206 737 6264 763
rect 6206 703 6212 737
rect 6252 703 6264 737
rect 6206 677 6264 703
rect 6306 737 6364 763
rect 6306 703 6318 737
rect 6358 703 6364 737
rect 6306 677 6364 703
rect 6406 737 6464 763
rect 6406 703 6412 737
rect 6452 703 6464 737
rect 6406 677 6464 703
rect 6506 737 6564 763
rect 6506 703 6518 737
rect 6558 703 6564 737
rect 6506 677 6564 703
rect 6606 737 6664 763
rect 6606 703 6618 737
rect 6652 703 6664 737
rect 6606 677 6664 703
rect 6706 737 6764 763
rect 6706 703 6718 737
rect 6752 703 6764 737
rect 6706 677 6764 703
rect 6806 737 6864 763
rect 6806 703 6818 737
rect 6852 703 6864 737
rect 6806 677 6864 703
rect 6906 737 6964 763
rect 6906 703 6918 737
rect 6952 703 6964 737
rect 6906 677 6964 703
rect 7006 737 7064 763
rect 7006 703 7012 737
rect 7052 703 7064 737
rect 7006 677 7064 703
rect 7106 737 7164 763
rect 7106 703 7118 737
rect 7158 703 7164 737
rect 7106 677 7164 703
rect 7206 737 7264 763
rect 7206 703 7218 737
rect 7252 703 7264 737
rect 7206 677 7264 703
rect 7306 737 7364 763
rect 7306 703 7318 737
rect 7352 703 7364 737
rect 7306 677 7364 703
rect 7406 737 7464 763
rect 7406 703 7418 737
rect 7452 703 7464 737
rect 7406 677 7464 703
rect 7506 737 7564 763
rect 7506 703 7518 737
rect 7552 703 7564 737
rect 7506 677 7564 703
rect 7606 737 7664 763
rect 7606 703 7618 737
rect 7652 703 7664 737
rect 7606 677 7664 703
rect 7706 737 7764 763
rect 7706 703 7718 737
rect 7752 703 7764 737
rect 7706 677 7764 703
rect 7806 737 7864 763
rect 7806 703 7818 737
rect 7852 703 7864 737
rect 7806 677 7864 703
rect 7906 737 7964 763
rect 7906 703 7918 737
rect 7952 703 7964 737
rect 7906 677 7964 703
rect 8006 737 8064 763
rect 8006 703 8018 737
rect 8052 703 8064 737
rect 8006 677 8064 703
rect 8106 737 8164 763
rect 8106 703 8118 737
rect 8152 703 8164 737
rect 8106 677 8164 703
rect 8206 737 8264 763
rect 8206 703 8218 737
rect 8252 703 8264 737
rect 8206 677 8264 703
rect 8306 737 8364 763
rect 8306 703 8318 737
rect 8352 703 8364 737
rect 8306 677 8364 703
rect 8406 737 8464 763
rect 8406 703 8418 737
rect 8452 703 8464 737
rect 8406 677 8464 703
rect 8506 737 8564 763
rect 8506 703 8518 737
rect 8552 703 8564 737
rect 8506 677 8564 703
rect 8606 737 8664 763
rect 8606 703 8618 737
rect 8652 703 8664 737
rect 8606 677 8664 703
rect 8706 737 8764 763
rect 8706 703 8718 737
rect 8752 703 8764 737
rect 8706 677 8764 703
rect 8806 737 8864 763
rect 8806 703 8818 737
rect 8852 703 8864 737
rect 8806 677 8864 703
rect 8906 737 8964 763
rect 8906 703 8918 737
rect 8952 703 8964 737
rect 8906 677 8964 703
rect 9006 737 9064 763
rect 9006 703 9018 737
rect 9052 703 9064 737
rect 9006 677 9064 703
rect 9106 737 9164 763
rect 9106 703 9112 737
rect 9152 703 9164 737
rect 9106 677 9164 703
rect 9206 737 9264 763
rect 9206 703 9218 737
rect 9258 703 9264 737
rect 9206 677 9264 703
rect 9306 737 9364 763
rect 9306 703 9312 737
rect 9352 703 9364 737
rect 9306 677 9364 703
rect 9406 737 9464 763
rect 9406 703 9418 737
rect 9458 703 9464 737
rect 9406 677 9464 703
rect 9506 737 9564 763
rect 9506 703 9518 737
rect 9552 703 9564 737
rect 9506 677 9564 703
rect 9606 737 9664 763
rect 9606 703 9612 737
rect 9652 703 9664 737
rect 9606 677 9664 703
rect 9706 737 9764 763
rect 9706 703 9718 737
rect 9758 703 9764 737
rect 9706 677 9764 703
rect 9806 737 9864 763
rect 9806 703 9812 737
rect 9852 703 9864 737
rect 9806 677 9864 703
rect 9906 737 9964 763
rect 9906 703 9918 737
rect 9958 703 9964 737
rect 9906 677 9964 703
rect 10006 737 10064 763
rect 10006 703 10018 737
rect 10052 703 10064 737
rect 10006 677 10064 703
rect 10106 737 10164 763
rect 10106 703 10112 737
rect 10152 703 10164 737
rect 10106 677 10164 703
rect 10206 737 10264 763
rect 10206 703 10218 737
rect 10258 703 10264 737
rect 10206 677 10264 703
rect 10306 737 10364 763
rect 10306 703 10318 737
rect 10352 703 10364 737
rect 10306 677 10364 703
rect 10406 737 10464 763
rect 10406 703 10418 737
rect 10452 703 10464 737
rect 10406 677 10464 703
rect 10506 737 10564 763
rect 10506 703 10518 737
rect 10552 703 10564 737
rect 10506 677 10564 703
rect 10606 737 10664 763
rect 10606 703 10618 737
rect 10652 703 10664 737
rect 10606 677 10664 703
rect 10706 737 10764 763
rect 10706 703 10718 737
rect 10752 703 10764 737
rect 10706 677 10764 703
rect 10806 737 10864 763
rect 10806 703 10818 737
rect 10852 703 10864 737
rect 10806 677 10864 703
rect 10906 737 10964 763
rect 10906 703 10912 737
rect 10952 703 10964 737
rect 10906 677 10964 703
rect 11006 737 11064 763
rect 11006 703 11018 737
rect 11058 703 11064 737
rect 11006 677 11064 703
rect 11106 737 11164 763
rect 11106 703 11118 737
rect 11152 703 11164 737
rect 11106 677 11164 703
rect 11206 737 11264 763
rect 11206 703 11218 737
rect 11252 703 11264 737
rect 11206 677 11264 703
rect 11306 737 11364 763
rect 11306 703 11318 737
rect 11352 703 11364 737
rect 11306 677 11364 703
rect 11406 737 11464 763
rect 11406 703 11418 737
rect 11452 703 11464 737
rect 11406 677 11464 703
rect 11506 737 11564 763
rect 11506 703 11518 737
rect 11552 703 11564 737
rect 11506 677 11564 703
rect 11606 737 11664 763
rect 11606 703 11618 737
rect 11652 703 11664 737
rect 11606 677 11664 703
rect 11706 737 11764 763
rect 11706 703 11712 737
rect 11752 703 11764 737
rect 11706 677 11764 703
rect 11806 737 11864 763
rect 11806 703 11818 737
rect 11858 703 11864 737
rect 11806 677 11864 703
rect 11906 737 11964 763
rect 11906 703 11918 737
rect 11952 703 11964 737
rect 11906 677 11964 703
rect 12006 737 12064 763
rect 12006 703 12018 737
rect 12052 703 12064 737
rect 12006 677 12064 703
rect 12106 737 12164 763
rect 12106 703 12112 737
rect 12152 703 12164 737
rect 12106 677 12164 703
rect 12206 737 12264 763
rect 12206 703 12218 737
rect 12258 703 12264 737
rect 12206 677 12264 703
rect 12306 737 12364 763
rect 12306 703 12318 737
rect 12352 703 12364 737
rect 12306 677 12364 703
rect 12406 737 12464 763
rect 12406 703 12418 737
rect 12452 703 12464 737
rect 12406 677 12464 703
rect 12506 737 12564 763
rect 12506 703 12518 737
rect 12552 703 12564 737
rect 12506 677 12564 703
rect 12606 737 12664 763
rect 12606 703 12618 737
rect 12652 703 12664 737
rect 12606 677 12664 703
rect 12706 737 12764 763
rect 12706 703 12718 737
rect 12752 703 12764 737
rect 12706 677 12764 703
rect 12806 737 12864 763
rect 13018 756 13262 790
rect 12806 703 12818 737
rect 12852 703 12864 737
rect 12908 718 12916 752
rect 12958 718 12974 752
rect 13018 737 13052 756
rect 12806 677 12864 703
rect 13228 737 13262 756
rect 13018 687 13052 703
rect 13096 688 13112 722
rect 13154 688 13162 722
rect 13228 687 13262 703
rect 13328 737 13462 753
rect 13362 703 13428 737
rect 13328 687 13462 703
rect 13528 737 13662 753
rect 13562 703 13628 737
rect 13528 687 13662 703
rect 6 597 64 623
rect 6 563 18 597
rect 52 563 64 597
rect 6 537 64 563
rect 106 597 164 623
rect 106 563 118 597
rect 152 563 164 597
rect 106 537 164 563
rect 206 597 264 623
rect 206 563 218 597
rect 252 563 264 597
rect 206 537 264 563
rect 306 597 364 623
rect 306 563 318 597
rect 352 563 364 597
rect 306 537 364 563
rect 406 597 464 623
rect 406 563 418 597
rect 452 563 464 597
rect 406 537 464 563
rect 506 597 564 623
rect 506 563 518 597
rect 552 563 564 597
rect 506 537 564 563
rect 606 597 664 623
rect 606 563 618 597
rect 652 563 664 597
rect 606 537 664 563
rect 706 597 764 623
rect 706 563 712 597
rect 752 563 764 597
rect 706 537 764 563
rect 806 597 864 623
rect 806 563 818 597
rect 858 563 864 597
rect 806 537 864 563
rect 906 597 964 623
rect 906 563 918 597
rect 952 563 964 597
rect 906 537 964 563
rect 1006 597 1064 623
rect 1006 563 1018 597
rect 1052 563 1064 597
rect 1006 537 1064 563
rect 1106 597 1164 623
rect 1106 563 1118 597
rect 1152 563 1164 597
rect 1106 537 1164 563
rect 1206 597 1264 623
rect 1206 563 1212 597
rect 1252 563 1264 597
rect 1206 537 1264 563
rect 1306 597 1364 623
rect 1306 563 1318 597
rect 1358 563 1364 597
rect 1306 537 1364 563
rect 1406 597 1464 623
rect 1406 563 1418 597
rect 1452 563 1464 597
rect 1406 537 1464 563
rect 1506 597 1564 623
rect 1506 563 1518 597
rect 1552 563 1564 597
rect 1506 537 1564 563
rect 1606 597 1664 623
rect 1606 563 1618 597
rect 1652 563 1664 597
rect 1606 537 1664 563
rect 1706 597 1764 623
rect 1706 563 1718 597
rect 1752 563 1764 597
rect 1706 537 1764 563
rect 1806 597 1864 623
rect 1806 563 1818 597
rect 1852 563 1864 597
rect 1806 537 1864 563
rect 1906 597 1964 623
rect 1906 563 1918 597
rect 1952 563 1964 597
rect 1906 537 1964 563
rect 2006 597 2064 623
rect 2006 563 2018 597
rect 2052 563 2064 597
rect 2006 537 2064 563
rect 2106 597 2164 623
rect 2106 563 2112 597
rect 2152 563 2164 597
rect 2106 537 2164 563
rect 2206 597 2264 623
rect 2206 563 2218 597
rect 2258 563 2264 597
rect 2206 537 2264 563
rect 2306 597 2364 623
rect 2306 563 2318 597
rect 2352 563 2364 597
rect 2306 537 2364 563
rect 2406 597 2464 623
rect 2406 563 2418 597
rect 2452 563 2464 597
rect 2406 537 2464 563
rect 2506 597 2564 623
rect 2506 563 2518 597
rect 2552 563 2564 597
rect 2506 537 2564 563
rect 2606 597 2664 623
rect 2606 563 2618 597
rect 2652 563 2664 597
rect 2606 537 2664 563
rect 2706 597 2764 623
rect 2706 563 2712 597
rect 2752 563 2764 597
rect 2706 537 2764 563
rect 2806 597 2864 623
rect 2806 563 2818 597
rect 2858 563 2864 597
rect 2806 537 2864 563
rect 2906 597 2964 623
rect 2906 563 2918 597
rect 2952 563 2964 597
rect 2906 537 2964 563
rect 3006 597 3064 623
rect 3006 563 3018 597
rect 3052 563 3064 597
rect 3006 537 3064 563
rect 3106 597 3164 623
rect 3106 563 3118 597
rect 3152 563 3164 597
rect 3106 537 3164 563
rect 3206 597 3264 623
rect 3206 563 3218 597
rect 3252 563 3264 597
rect 3206 537 3264 563
rect 3306 597 3364 623
rect 3306 563 3318 597
rect 3352 563 3364 597
rect 3306 537 3364 563
rect 3406 597 3464 623
rect 3406 563 3418 597
rect 3452 563 3464 597
rect 3406 537 3464 563
rect 3506 597 3564 623
rect 3506 563 3518 597
rect 3552 563 3564 597
rect 3506 537 3564 563
rect 3606 597 3664 623
rect 3606 563 3618 597
rect 3652 563 3664 597
rect 3606 537 3664 563
rect 3706 597 3764 623
rect 3706 563 3718 597
rect 3752 563 3764 597
rect 3706 537 3764 563
rect 3806 597 3864 623
rect 3806 563 3818 597
rect 3852 563 3864 597
rect 3806 537 3864 563
rect 3906 597 3964 623
rect 3906 563 3912 597
rect 3952 563 3964 597
rect 3906 537 3964 563
rect 4006 597 4064 623
rect 4006 563 4018 597
rect 4058 563 4064 597
rect 4006 537 4064 563
rect 4106 597 4164 623
rect 4106 563 4112 597
rect 4152 563 4164 597
rect 4106 537 4164 563
rect 4206 597 4264 623
rect 4206 563 4218 597
rect 4258 563 4264 597
rect 4206 537 4264 563
rect 4306 597 4364 623
rect 4306 563 4318 597
rect 4352 563 4364 597
rect 4306 537 4364 563
rect 4406 597 4464 623
rect 4406 563 4418 597
rect 4452 563 4464 597
rect 4406 537 4464 563
rect 4506 597 4564 623
rect 4506 563 4518 597
rect 4552 563 4564 597
rect 4506 537 4564 563
rect 4606 597 4664 623
rect 4606 563 4618 597
rect 4652 563 4664 597
rect 4606 537 4664 563
rect 4706 597 4764 623
rect 4706 563 4718 597
rect 4752 563 4764 597
rect 4706 537 4764 563
rect 4806 597 4864 623
rect 4806 563 4812 597
rect 4852 563 4864 597
rect 4806 537 4864 563
rect 4906 597 4964 623
rect 4906 563 4918 597
rect 4958 563 4964 597
rect 4906 537 4964 563
rect 5006 597 5064 623
rect 5006 563 5012 597
rect 5052 563 5064 597
rect 5006 537 5064 563
rect 5106 597 5164 623
rect 5106 563 5118 597
rect 5158 563 5164 597
rect 5106 537 5164 563
rect 5206 597 5264 623
rect 5206 563 5212 597
rect 5252 563 5264 597
rect 5206 537 5264 563
rect 5306 597 5364 623
rect 5306 563 5318 597
rect 5358 563 5364 597
rect 5306 537 5364 563
rect 5406 597 5464 623
rect 5406 563 5418 597
rect 5452 563 5464 597
rect 5406 537 5464 563
rect 5506 597 5564 623
rect 5506 563 5518 597
rect 5552 563 5564 597
rect 5506 537 5564 563
rect 5606 597 5664 623
rect 5606 563 5618 597
rect 5652 563 5664 597
rect 5606 537 5664 563
rect 5706 597 5764 623
rect 5706 563 5718 597
rect 5752 563 5764 597
rect 5706 537 5764 563
rect 5806 597 5864 623
rect 5806 563 5818 597
rect 5852 563 5864 597
rect 5806 537 5864 563
rect 5906 597 5964 623
rect 5906 563 5918 597
rect 5952 563 5964 597
rect 5906 537 5964 563
rect 6006 597 6064 623
rect 6006 563 6018 597
rect 6052 563 6064 597
rect 6006 537 6064 563
rect 6106 597 6164 623
rect 6106 563 6118 597
rect 6152 563 6164 597
rect 6106 537 6164 563
rect 6206 597 6264 623
rect 6206 563 6218 597
rect 6252 563 6264 597
rect 6206 537 6264 563
rect 6306 597 6364 623
rect 6306 563 6318 597
rect 6352 563 6364 597
rect 6306 537 6364 563
rect 6406 597 6464 623
rect 6406 563 6418 597
rect 6452 563 6464 597
rect 6406 537 6464 563
rect 6506 597 6564 623
rect 6506 563 6518 597
rect 6552 563 6564 597
rect 6506 537 6564 563
rect 6606 597 6664 623
rect 6606 563 6618 597
rect 6652 563 6664 597
rect 6606 537 6664 563
rect 6706 597 6764 623
rect 6706 563 6718 597
rect 6752 563 6764 597
rect 6706 537 6764 563
rect 6806 597 6864 623
rect 6806 563 6818 597
rect 6852 563 6864 597
rect 6806 537 6864 563
rect 6906 597 6964 623
rect 6906 563 6918 597
rect 6952 563 6964 597
rect 6906 537 6964 563
rect 7006 597 7064 623
rect 7006 563 7018 597
rect 7052 563 7064 597
rect 7006 537 7064 563
rect 7106 597 7164 623
rect 7106 563 7118 597
rect 7152 563 7164 597
rect 7106 537 7164 563
rect 7206 597 7264 623
rect 7206 563 7218 597
rect 7252 563 7264 597
rect 7206 537 7264 563
rect 7306 597 7364 623
rect 7306 563 7318 597
rect 7352 563 7364 597
rect 7306 537 7364 563
rect 7406 597 7464 623
rect 7406 563 7418 597
rect 7452 563 7464 597
rect 7406 537 7464 563
rect 7506 597 7564 623
rect 7506 563 7518 597
rect 7552 563 7564 597
rect 7506 537 7564 563
rect 7606 597 7664 623
rect 7606 563 7618 597
rect 7652 563 7664 597
rect 7606 537 7664 563
rect 7706 597 7764 623
rect 7706 563 7718 597
rect 7752 563 7764 597
rect 7706 537 7764 563
rect 7806 597 7864 623
rect 7806 563 7818 597
rect 7852 563 7864 597
rect 7806 537 7864 563
rect 7906 597 7964 623
rect 7906 563 7918 597
rect 7952 563 7964 597
rect 7906 537 7964 563
rect 8006 597 8064 623
rect 8006 563 8018 597
rect 8052 563 8064 597
rect 8006 537 8064 563
rect 8106 597 8164 623
rect 8106 563 8118 597
rect 8152 563 8164 597
rect 8106 537 8164 563
rect 8206 597 8264 623
rect 8206 563 8218 597
rect 8252 563 8264 597
rect 8206 537 8264 563
rect 8306 597 8364 623
rect 8306 563 8312 597
rect 8352 563 8364 597
rect 8306 537 8364 563
rect 8406 597 8464 623
rect 8406 563 8418 597
rect 8458 563 8464 597
rect 8406 537 8464 563
rect 8506 597 8564 623
rect 8506 563 8518 597
rect 8552 563 8564 597
rect 8506 537 8564 563
rect 8606 597 8664 623
rect 8606 563 8618 597
rect 8652 563 8664 597
rect 8606 537 8664 563
rect 8706 597 8764 623
rect 8706 563 8718 597
rect 8752 563 8764 597
rect 8706 537 8764 563
rect 8806 597 8864 623
rect 8806 563 8818 597
rect 8852 563 8864 597
rect 8806 537 8864 563
rect 8906 597 8964 623
rect 8906 563 8918 597
rect 8952 563 8964 597
rect 8906 537 8964 563
rect 9006 597 9064 623
rect 9006 563 9018 597
rect 9052 563 9064 597
rect 9006 537 9064 563
rect 9106 597 9164 623
rect 9106 563 9118 597
rect 9152 563 9164 597
rect 9106 537 9164 563
rect 9206 597 9264 623
rect 9206 563 9218 597
rect 9252 563 9264 597
rect 9206 537 9264 563
rect 9306 597 9364 623
rect 9306 563 9318 597
rect 9352 563 9364 597
rect 9306 537 9364 563
rect 9406 597 9464 623
rect 9406 563 9418 597
rect 9452 563 9464 597
rect 9406 537 9464 563
rect 9506 597 9564 623
rect 9506 563 9518 597
rect 9552 563 9564 597
rect 9506 537 9564 563
rect 9606 597 9664 623
rect 9606 563 9618 597
rect 9652 563 9664 597
rect 9606 537 9664 563
rect 9706 597 9764 623
rect 9706 563 9718 597
rect 9752 563 9764 597
rect 9706 537 9764 563
rect 9806 597 9864 623
rect 9806 563 9818 597
rect 9852 563 9864 597
rect 9806 537 9864 563
rect 9906 597 9964 623
rect 9906 563 9918 597
rect 9952 563 9964 597
rect 9906 537 9964 563
rect 10006 597 10064 623
rect 10006 563 10018 597
rect 10052 563 10064 597
rect 10006 537 10064 563
rect 10106 597 10164 623
rect 10106 563 10118 597
rect 10152 563 10164 597
rect 10106 537 10164 563
rect 10206 597 10264 623
rect 10206 563 10212 597
rect 10252 563 10264 597
rect 10206 537 10264 563
rect 10306 597 10364 623
rect 10306 563 10318 597
rect 10358 563 10364 597
rect 10306 537 10364 563
rect 10406 597 10464 623
rect 10406 563 10412 597
rect 10452 563 10464 597
rect 10406 537 10464 563
rect 10506 597 10564 623
rect 10506 563 10518 597
rect 10558 563 10564 597
rect 10506 537 10564 563
rect 10606 597 10664 623
rect 10606 563 10618 597
rect 10652 563 10664 597
rect 10606 537 10664 563
rect 10706 597 10764 623
rect 10706 563 10718 597
rect 10752 563 10764 597
rect 10706 537 10764 563
rect 10806 597 10864 623
rect 10806 563 10818 597
rect 10852 563 10864 597
rect 10806 537 10864 563
rect 10906 597 10964 623
rect 10906 563 10918 597
rect 10952 563 10964 597
rect 10906 537 10964 563
rect 11006 597 11064 623
rect 11006 563 11018 597
rect 11052 563 11064 597
rect 11006 537 11064 563
rect 11106 597 11164 623
rect 11106 563 11118 597
rect 11152 563 11164 597
rect 11106 537 11164 563
rect 11206 597 11264 623
rect 11206 563 11212 597
rect 11252 563 11264 597
rect 11206 537 11264 563
rect 11306 597 11364 623
rect 11306 563 11318 597
rect 11358 563 11364 597
rect 11306 537 11364 563
rect 11406 597 11464 623
rect 11406 563 11418 597
rect 11452 563 11464 597
rect 11406 537 11464 563
rect 11506 597 11564 623
rect 11506 563 11518 597
rect 11552 563 11564 597
rect 11506 537 11564 563
rect 11606 597 11664 623
rect 11606 563 11618 597
rect 11652 563 11664 597
rect 11606 537 11664 563
rect 11706 597 11764 623
rect 11706 563 11718 597
rect 11752 563 11764 597
rect 11706 537 11764 563
rect 11806 597 11864 623
rect 11806 563 11818 597
rect 11852 563 11864 597
rect 11806 537 11864 563
rect 11906 597 11964 623
rect 11906 563 11918 597
rect 11952 563 11964 597
rect 11906 537 11964 563
rect 12006 597 12064 623
rect 12006 563 12018 597
rect 12052 563 12064 597
rect 12006 537 12064 563
rect 12106 597 12164 623
rect 12106 563 12118 597
rect 12152 563 12164 597
rect 12106 537 12164 563
rect 12206 597 12264 623
rect 12206 563 12218 597
rect 12252 563 12264 597
rect 12206 537 12264 563
rect 12306 597 12364 623
rect 12306 563 12318 597
rect 12352 563 12364 597
rect 12306 537 12364 563
rect 12406 597 12464 623
rect 12406 563 12418 597
rect 12452 563 12464 597
rect 12406 537 12464 563
rect 12506 597 12564 623
rect 12506 563 12518 597
rect 12552 563 12564 597
rect 12506 537 12564 563
rect 12606 597 12664 623
rect 12606 563 12618 597
rect 12652 563 12664 597
rect 12606 537 12664 563
rect 12706 597 12764 623
rect 12706 563 12718 597
rect 12752 563 12764 597
rect 12706 537 12764 563
rect 12806 597 12864 623
rect 13018 616 13262 650
rect 12806 563 12812 597
rect 12852 563 12864 597
rect 12908 578 12916 612
rect 12958 578 12974 612
rect 13018 597 13052 616
rect 12806 537 12864 563
rect 13228 613 13262 616
rect 13228 597 13362 613
rect 13018 547 13052 563
rect 13096 548 13112 582
rect 13154 548 13162 582
rect 13262 563 13328 597
rect 13228 547 13362 563
rect 13428 597 13562 613
rect 13462 563 13528 597
rect 13428 547 13562 563
rect 13628 597 13662 613
rect 13628 547 13662 563
rect 6 457 64 483
rect 6 423 18 457
rect 52 423 64 457
rect 6 397 64 423
rect 106 457 164 483
rect 106 423 118 457
rect 152 423 164 457
rect 106 397 164 423
rect 206 457 264 483
rect 206 423 218 457
rect 252 423 264 457
rect 206 397 264 423
rect 306 457 364 483
rect 306 423 312 457
rect 352 423 364 457
rect 306 397 364 423
rect 406 457 464 483
rect 406 423 418 457
rect 458 423 464 457
rect 406 397 464 423
rect 506 457 564 483
rect 506 423 518 457
rect 552 423 564 457
rect 506 397 564 423
rect 606 457 664 483
rect 606 423 618 457
rect 652 423 664 457
rect 606 397 664 423
rect 706 457 764 483
rect 706 423 718 457
rect 752 423 764 457
rect 706 397 764 423
rect 806 457 864 483
rect 806 423 818 457
rect 852 423 864 457
rect 806 397 864 423
rect 906 457 964 483
rect 906 423 918 457
rect 952 423 964 457
rect 906 397 964 423
rect 1006 457 1064 483
rect 1006 423 1018 457
rect 1052 423 1064 457
rect 1006 397 1064 423
rect 1106 457 1164 483
rect 1106 423 1112 457
rect 1152 423 1164 457
rect 1106 397 1164 423
rect 1206 457 1264 483
rect 1206 423 1218 457
rect 1258 423 1264 457
rect 1206 397 1264 423
rect 1306 457 1364 483
rect 1306 423 1318 457
rect 1352 423 1364 457
rect 1306 397 1364 423
rect 1406 457 1464 483
rect 1406 423 1418 457
rect 1452 423 1464 457
rect 1406 397 1464 423
rect 1506 457 1564 483
rect 1506 423 1518 457
rect 1552 423 1564 457
rect 1506 397 1564 423
rect 1606 457 1664 483
rect 1606 423 1618 457
rect 1652 423 1664 457
rect 1606 397 1664 423
rect 1706 457 1764 483
rect 1706 423 1718 457
rect 1752 423 1764 457
rect 1706 397 1764 423
rect 1806 457 1864 483
rect 1806 423 1812 457
rect 1852 423 1864 457
rect 1806 397 1864 423
rect 1906 457 1964 483
rect 1906 423 1918 457
rect 1958 423 1964 457
rect 1906 397 1964 423
rect 2006 457 2064 483
rect 2006 423 2018 457
rect 2052 423 2064 457
rect 2006 397 2064 423
rect 2106 457 2164 483
rect 2106 423 2118 457
rect 2152 423 2164 457
rect 2106 397 2164 423
rect 2206 457 2264 483
rect 2206 423 2218 457
rect 2252 423 2264 457
rect 2206 397 2264 423
rect 2306 457 2364 483
rect 2306 423 2312 457
rect 2352 423 2364 457
rect 2306 397 2364 423
rect 2406 457 2464 483
rect 2406 423 2418 457
rect 2458 423 2464 457
rect 2406 397 2464 423
rect 2506 457 2564 483
rect 2506 423 2518 457
rect 2552 423 2564 457
rect 2506 397 2564 423
rect 2606 457 2664 483
rect 2606 423 2612 457
rect 2652 423 2664 457
rect 2606 397 2664 423
rect 2706 457 2764 483
rect 2706 423 2718 457
rect 2758 423 2764 457
rect 2706 397 2764 423
rect 2806 457 2864 483
rect 2806 423 2818 457
rect 2852 423 2864 457
rect 2806 397 2864 423
rect 2906 457 2964 483
rect 2906 423 2918 457
rect 2952 423 2964 457
rect 2906 397 2964 423
rect 3006 457 3064 483
rect 3006 423 3018 457
rect 3052 423 3064 457
rect 3006 397 3064 423
rect 3106 457 3164 483
rect 3106 423 3118 457
rect 3152 423 3164 457
rect 3106 397 3164 423
rect 3206 457 3264 483
rect 3206 423 3218 457
rect 3252 423 3264 457
rect 3206 397 3264 423
rect 3306 457 3364 483
rect 3306 423 3318 457
rect 3352 423 3364 457
rect 3306 397 3364 423
rect 3406 457 3464 483
rect 3406 423 3418 457
rect 3452 423 3464 457
rect 3406 397 3464 423
rect 3506 457 3564 483
rect 3506 423 3518 457
rect 3552 423 3564 457
rect 3506 397 3564 423
rect 3606 457 3664 483
rect 3606 423 3618 457
rect 3652 423 3664 457
rect 3606 397 3664 423
rect 3706 457 3764 483
rect 3706 423 3718 457
rect 3752 423 3764 457
rect 3706 397 3764 423
rect 3806 457 3864 483
rect 3806 423 3818 457
rect 3852 423 3864 457
rect 3806 397 3864 423
rect 3906 457 3964 483
rect 3906 423 3918 457
rect 3952 423 3964 457
rect 3906 397 3964 423
rect 4006 457 4064 483
rect 4006 423 4018 457
rect 4052 423 4064 457
rect 4006 397 4064 423
rect 4106 457 4164 483
rect 4106 423 4118 457
rect 4152 423 4164 457
rect 4106 397 4164 423
rect 4206 457 4264 483
rect 4206 423 4218 457
rect 4252 423 4264 457
rect 4206 397 4264 423
rect 4306 457 4364 483
rect 4306 423 4318 457
rect 4352 423 4364 457
rect 4306 397 4364 423
rect 4406 457 4464 483
rect 4406 423 4412 457
rect 4452 423 4464 457
rect 4406 397 4464 423
rect 4506 457 4564 483
rect 4506 423 4518 457
rect 4558 423 4564 457
rect 4506 397 4564 423
rect 4606 457 4664 483
rect 4606 423 4618 457
rect 4652 423 4664 457
rect 4606 397 4664 423
rect 4706 457 4764 483
rect 4706 423 4718 457
rect 4752 423 4764 457
rect 4706 397 4764 423
rect 4806 457 4864 483
rect 4806 423 4818 457
rect 4852 423 4864 457
rect 4806 397 4864 423
rect 4906 457 4964 483
rect 4906 423 4918 457
rect 4952 423 4964 457
rect 4906 397 4964 423
rect 5006 457 5064 483
rect 5006 423 5018 457
rect 5052 423 5064 457
rect 5006 397 5064 423
rect 5106 457 5164 483
rect 5106 423 5112 457
rect 5152 423 5164 457
rect 5106 397 5164 423
rect 5206 457 5264 483
rect 5206 423 5218 457
rect 5258 423 5264 457
rect 5206 397 5264 423
rect 5306 457 5364 483
rect 5306 423 5312 457
rect 5352 423 5364 457
rect 5306 397 5364 423
rect 5406 457 5464 483
rect 5406 423 5418 457
rect 5458 423 5464 457
rect 5406 397 5464 423
rect 5506 457 5564 483
rect 5506 423 5518 457
rect 5552 423 5564 457
rect 5506 397 5564 423
rect 5606 457 5664 483
rect 5606 423 5618 457
rect 5652 423 5664 457
rect 5606 397 5664 423
rect 5706 457 5764 483
rect 5706 423 5718 457
rect 5752 423 5764 457
rect 5706 397 5764 423
rect 5806 457 5864 483
rect 5806 423 5818 457
rect 5852 423 5864 457
rect 5806 397 5864 423
rect 5906 457 5964 483
rect 5906 423 5918 457
rect 5952 423 5964 457
rect 5906 397 5964 423
rect 6006 457 6064 483
rect 6006 423 6018 457
rect 6052 423 6064 457
rect 6006 397 6064 423
rect 6106 457 6164 483
rect 6106 423 6112 457
rect 6152 423 6164 457
rect 6106 397 6164 423
rect 6206 457 6264 483
rect 6206 423 6218 457
rect 6258 423 6264 457
rect 6206 397 6264 423
rect 6306 457 6364 483
rect 6306 423 6318 457
rect 6352 423 6364 457
rect 6306 397 6364 423
rect 6406 457 6464 483
rect 6406 423 6412 457
rect 6452 423 6464 457
rect 6406 397 6464 423
rect 6506 457 6564 483
rect 6506 423 6518 457
rect 6558 423 6564 457
rect 6506 397 6564 423
rect 6606 457 6664 483
rect 6606 423 6618 457
rect 6652 423 6664 457
rect 6606 397 6664 423
rect 6706 457 6764 483
rect 6706 423 6718 457
rect 6752 423 6764 457
rect 6706 397 6764 423
rect 6806 457 6864 483
rect 6806 423 6818 457
rect 6852 423 6864 457
rect 6806 397 6864 423
rect 6906 457 6964 483
rect 6906 423 6918 457
rect 6952 423 6964 457
rect 6906 397 6964 423
rect 7006 457 7064 483
rect 7006 423 7018 457
rect 7052 423 7064 457
rect 7006 397 7064 423
rect 7106 457 7164 483
rect 7106 423 7112 457
rect 7152 423 7164 457
rect 7106 397 7164 423
rect 7206 457 7264 483
rect 7206 423 7218 457
rect 7258 423 7264 457
rect 7206 397 7264 423
rect 7306 457 7364 483
rect 7306 423 7312 457
rect 7352 423 7364 457
rect 7306 397 7364 423
rect 7406 457 7464 483
rect 7406 423 7418 457
rect 7458 423 7464 457
rect 7406 397 7464 423
rect 7506 457 7564 483
rect 7506 423 7512 457
rect 7552 423 7564 457
rect 7506 397 7564 423
rect 7606 457 7664 483
rect 7606 423 7618 457
rect 7658 423 7664 457
rect 7606 397 7664 423
rect 7706 457 7764 483
rect 7706 423 7718 457
rect 7752 423 7764 457
rect 7706 397 7764 423
rect 7806 457 7864 483
rect 7806 423 7818 457
rect 7852 423 7864 457
rect 7806 397 7864 423
rect 7906 457 7964 483
rect 7906 423 7918 457
rect 7952 423 7964 457
rect 7906 397 7964 423
rect 8006 457 8064 483
rect 8006 423 8018 457
rect 8052 423 8064 457
rect 8006 397 8064 423
rect 8106 457 8164 483
rect 8106 423 8118 457
rect 8152 423 8164 457
rect 8106 397 8164 423
rect 8206 457 8264 483
rect 8206 423 8218 457
rect 8252 423 8264 457
rect 8206 397 8264 423
rect 8306 457 8364 483
rect 8306 423 8312 457
rect 8352 423 8364 457
rect 8306 397 8364 423
rect 8406 457 8464 483
rect 8406 423 8418 457
rect 8458 423 8464 457
rect 8406 397 8464 423
rect 8506 457 8564 483
rect 8506 423 8518 457
rect 8552 423 8564 457
rect 8506 397 8564 423
rect 8606 457 8664 483
rect 8606 423 8618 457
rect 8652 423 8664 457
rect 8606 397 8664 423
rect 8706 457 8764 483
rect 8706 423 8718 457
rect 8752 423 8764 457
rect 8706 397 8764 423
rect 8806 457 8864 483
rect 8806 423 8818 457
rect 8852 423 8864 457
rect 8806 397 8864 423
rect 8906 457 8964 483
rect 8906 423 8918 457
rect 8952 423 8964 457
rect 8906 397 8964 423
rect 9006 457 9064 483
rect 9006 423 9018 457
rect 9052 423 9064 457
rect 9006 397 9064 423
rect 9106 457 9164 483
rect 9106 423 9118 457
rect 9152 423 9164 457
rect 9106 397 9164 423
rect 9206 457 9264 483
rect 9206 423 9218 457
rect 9252 423 9264 457
rect 9206 397 9264 423
rect 9306 457 9364 483
rect 9306 423 9318 457
rect 9352 423 9364 457
rect 9306 397 9364 423
rect 9406 457 9464 483
rect 9406 423 9418 457
rect 9452 423 9464 457
rect 9406 397 9464 423
rect 9506 457 9564 483
rect 9506 423 9518 457
rect 9552 423 9564 457
rect 9506 397 9564 423
rect 9606 457 9664 483
rect 9606 423 9618 457
rect 9652 423 9664 457
rect 9606 397 9664 423
rect 9706 457 9764 483
rect 9706 423 9718 457
rect 9752 423 9764 457
rect 9706 397 9764 423
rect 9806 457 9864 483
rect 9806 423 9818 457
rect 9852 423 9864 457
rect 9806 397 9864 423
rect 9906 457 9964 483
rect 9906 423 9912 457
rect 9952 423 9964 457
rect 9906 397 9964 423
rect 10006 457 10064 483
rect 10006 423 10018 457
rect 10058 423 10064 457
rect 10006 397 10064 423
rect 10106 457 10164 483
rect 10106 423 10118 457
rect 10152 423 10164 457
rect 10106 397 10164 423
rect 10206 457 10264 483
rect 10206 423 10212 457
rect 10252 423 10264 457
rect 10206 397 10264 423
rect 10306 457 10364 483
rect 10306 423 10318 457
rect 10358 423 10364 457
rect 10306 397 10364 423
rect 10406 457 10464 483
rect 10406 423 10418 457
rect 10452 423 10464 457
rect 10406 397 10464 423
rect 10506 457 10564 483
rect 10506 423 10518 457
rect 10552 423 10564 457
rect 10506 397 10564 423
rect 10606 457 10664 483
rect 10606 423 10618 457
rect 10652 423 10664 457
rect 10606 397 10664 423
rect 10706 457 10764 483
rect 10706 423 10718 457
rect 10752 423 10764 457
rect 10706 397 10764 423
rect 10806 457 10864 483
rect 10806 423 10812 457
rect 10852 423 10864 457
rect 10806 397 10864 423
rect 10906 457 10964 483
rect 10906 423 10918 457
rect 10958 423 10964 457
rect 10906 397 10964 423
rect 11006 457 11064 483
rect 11006 423 11018 457
rect 11052 423 11064 457
rect 11006 397 11064 423
rect 11106 457 11164 483
rect 11106 423 11112 457
rect 11152 423 11164 457
rect 11106 397 11164 423
rect 11206 457 11264 483
rect 11206 423 11218 457
rect 11258 423 11264 457
rect 11206 397 11264 423
rect 11306 457 11364 483
rect 11306 423 11312 457
rect 11352 423 11364 457
rect 11306 397 11364 423
rect 11406 457 11464 483
rect 11406 423 11418 457
rect 11458 423 11464 457
rect 11406 397 11464 423
rect 11506 457 11564 483
rect 11506 423 11518 457
rect 11552 423 11564 457
rect 11506 397 11564 423
rect 11606 457 11664 483
rect 11606 423 11618 457
rect 11652 423 11664 457
rect 11606 397 11664 423
rect 11706 457 11764 483
rect 11706 423 11718 457
rect 11752 423 11764 457
rect 11706 397 11764 423
rect 11806 457 11864 483
rect 11806 423 11818 457
rect 11852 423 11864 457
rect 11806 397 11864 423
rect 11906 457 11964 483
rect 11906 423 11918 457
rect 11952 423 11964 457
rect 11906 397 11964 423
rect 12006 457 12064 483
rect 12006 423 12018 457
rect 12052 423 12064 457
rect 12006 397 12064 423
rect 12106 457 12164 483
rect 12106 423 12118 457
rect 12152 423 12164 457
rect 12106 397 12164 423
rect 12206 457 12264 483
rect 12206 423 12218 457
rect 12252 423 12264 457
rect 12206 397 12264 423
rect 12306 457 12364 483
rect 12306 423 12312 457
rect 12352 423 12364 457
rect 12306 397 12364 423
rect 12406 457 12464 483
rect 12406 423 12418 457
rect 12458 423 12464 457
rect 12406 397 12464 423
rect 12506 457 12564 483
rect 12506 423 12518 457
rect 12552 423 12564 457
rect 12506 397 12564 423
rect 12606 457 12664 483
rect 12606 423 12618 457
rect 12652 423 12664 457
rect 12606 397 12664 423
rect 12706 457 12764 483
rect 12706 423 12718 457
rect 12752 423 12764 457
rect 12706 397 12764 423
rect 12806 457 12864 483
rect 13018 476 13262 510
rect 12806 423 12812 457
rect 12852 423 12864 457
rect 12908 438 12916 472
rect 12958 438 12974 472
rect 13018 457 13052 476
rect 12806 397 12864 423
rect 13228 457 13262 476
rect 13018 407 13052 423
rect 13096 408 13112 442
rect 13154 408 13162 442
rect 13228 407 13262 423
rect 13328 457 13562 473
rect 13362 423 13428 457
rect 13462 423 13528 457
rect 13328 407 13562 423
rect 13628 457 13662 473
rect 13628 407 13662 423
rect 6 317 64 343
rect 6 283 18 317
rect 52 283 64 317
rect 6 257 64 283
rect 106 317 164 343
rect 106 283 118 317
rect 152 283 164 317
rect 106 257 164 283
rect 206 317 264 343
rect 206 283 218 317
rect 252 283 264 317
rect 206 257 264 283
rect 306 317 364 343
rect 306 283 318 317
rect 352 283 364 317
rect 306 257 364 283
rect 406 317 464 343
rect 406 283 418 317
rect 452 283 464 317
rect 406 257 464 283
rect 506 317 564 343
rect 506 283 518 317
rect 552 283 564 317
rect 506 257 564 283
rect 606 317 664 343
rect 606 283 618 317
rect 652 283 664 317
rect 606 257 664 283
rect 706 317 764 343
rect 706 283 718 317
rect 752 283 764 317
rect 706 257 764 283
rect 806 317 864 343
rect 806 283 818 317
rect 852 283 864 317
rect 806 257 864 283
rect 906 317 964 343
rect 906 283 918 317
rect 952 283 964 317
rect 906 257 964 283
rect 1006 317 1064 343
rect 1006 283 1018 317
rect 1052 283 1064 317
rect 1006 257 1064 283
rect 1106 317 1164 343
rect 1106 283 1118 317
rect 1152 283 1164 317
rect 1106 257 1164 283
rect 1206 317 1264 343
rect 1206 283 1218 317
rect 1252 283 1264 317
rect 1206 257 1264 283
rect 1306 317 1364 343
rect 1306 283 1318 317
rect 1352 283 1364 317
rect 1306 257 1364 283
rect 1406 317 1464 343
rect 1406 283 1418 317
rect 1452 283 1464 317
rect 1406 257 1464 283
rect 1506 317 1564 343
rect 1506 283 1518 317
rect 1552 283 1564 317
rect 1506 257 1564 283
rect 1606 317 1664 343
rect 1606 283 1618 317
rect 1652 283 1664 317
rect 1606 257 1664 283
rect 1706 317 1764 343
rect 1706 283 1712 317
rect 1752 283 1764 317
rect 1706 257 1764 283
rect 1806 317 1864 343
rect 1806 283 1818 317
rect 1858 283 1864 317
rect 1806 257 1864 283
rect 1906 317 1964 343
rect 1906 283 1918 317
rect 1952 283 1964 317
rect 1906 257 1964 283
rect 2006 317 2064 343
rect 2006 283 2018 317
rect 2052 283 2064 317
rect 2006 257 2064 283
rect 2106 317 2164 343
rect 2106 283 2118 317
rect 2152 283 2164 317
rect 2106 257 2164 283
rect 2206 317 2264 343
rect 2206 283 2218 317
rect 2252 283 2264 317
rect 2206 257 2264 283
rect 2306 317 2364 343
rect 2306 283 2318 317
rect 2352 283 2364 317
rect 2306 257 2364 283
rect 2406 317 2464 343
rect 2406 283 2418 317
rect 2452 283 2464 317
rect 2406 257 2464 283
rect 2506 317 2564 343
rect 2506 283 2518 317
rect 2552 283 2564 317
rect 2506 257 2564 283
rect 2606 317 2664 343
rect 2606 283 2618 317
rect 2652 283 2664 317
rect 2606 257 2664 283
rect 2706 317 2764 343
rect 2706 283 2718 317
rect 2752 283 2764 317
rect 2706 257 2764 283
rect 2806 317 2864 343
rect 2806 283 2812 317
rect 2852 283 2864 317
rect 2806 257 2864 283
rect 2906 317 2964 343
rect 2906 283 2918 317
rect 2958 283 2964 317
rect 2906 257 2964 283
rect 3006 317 3064 343
rect 3006 283 3012 317
rect 3052 283 3064 317
rect 3006 257 3064 283
rect 3106 317 3164 343
rect 3106 283 3118 317
rect 3158 283 3164 317
rect 3106 257 3164 283
rect 3206 317 3264 343
rect 3206 283 3218 317
rect 3252 283 3264 317
rect 3206 257 3264 283
rect 3306 317 3364 343
rect 3306 283 3318 317
rect 3352 283 3364 317
rect 3306 257 3364 283
rect 3406 317 3464 343
rect 3406 283 3418 317
rect 3452 283 3464 317
rect 3406 257 3464 283
rect 3506 317 3564 343
rect 3506 283 3518 317
rect 3552 283 3564 317
rect 3506 257 3564 283
rect 3606 317 3664 343
rect 3606 283 3618 317
rect 3652 283 3664 317
rect 3606 257 3664 283
rect 3706 317 3764 343
rect 3706 283 3718 317
rect 3752 283 3764 317
rect 3706 257 3764 283
rect 3806 317 3864 343
rect 3806 283 3818 317
rect 3852 283 3864 317
rect 3806 257 3864 283
rect 3906 317 3964 343
rect 3906 283 3918 317
rect 3952 283 3964 317
rect 3906 257 3964 283
rect 4006 317 4064 343
rect 4006 283 4018 317
rect 4052 283 4064 317
rect 4006 257 4064 283
rect 4106 317 4164 343
rect 4106 283 4118 317
rect 4152 283 4164 317
rect 4106 257 4164 283
rect 4206 317 4264 343
rect 4206 283 4218 317
rect 4252 283 4264 317
rect 4206 257 4264 283
rect 4306 317 4364 343
rect 4306 283 4318 317
rect 4352 283 4364 317
rect 4306 257 4364 283
rect 4406 317 4464 343
rect 4406 283 4418 317
rect 4452 283 4464 317
rect 4406 257 4464 283
rect 4506 317 4564 343
rect 4506 283 4512 317
rect 4552 283 4564 317
rect 4506 257 4564 283
rect 4606 317 4664 343
rect 4606 283 4618 317
rect 4658 283 4664 317
rect 4606 257 4664 283
rect 4706 317 4764 343
rect 4706 283 4718 317
rect 4752 283 4764 317
rect 4706 257 4764 283
rect 4806 317 4864 343
rect 4806 283 4812 317
rect 4852 283 4864 317
rect 4806 257 4864 283
rect 4906 317 4964 343
rect 4906 283 4918 317
rect 4958 283 4964 317
rect 4906 257 4964 283
rect 5006 317 5064 343
rect 5006 283 5012 317
rect 5052 283 5064 317
rect 5006 257 5064 283
rect 5106 317 5164 343
rect 5106 283 5118 317
rect 5158 283 5164 317
rect 5106 257 5164 283
rect 5206 317 5264 343
rect 5206 283 5218 317
rect 5252 283 5264 317
rect 5206 257 5264 283
rect 5306 317 5364 343
rect 5306 283 5318 317
rect 5352 283 5364 317
rect 5306 257 5364 283
rect 5406 317 5464 343
rect 5406 283 5418 317
rect 5452 283 5464 317
rect 5406 257 5464 283
rect 5506 317 5564 343
rect 5506 283 5518 317
rect 5552 283 5564 317
rect 5506 257 5564 283
rect 5606 317 5664 343
rect 5606 283 5618 317
rect 5652 283 5664 317
rect 5606 257 5664 283
rect 5706 317 5764 343
rect 5706 283 5718 317
rect 5752 283 5764 317
rect 5706 257 5764 283
rect 5806 317 5864 343
rect 5806 283 5812 317
rect 5852 283 5864 317
rect 5806 257 5864 283
rect 5906 317 5964 343
rect 5906 283 5918 317
rect 5958 283 5964 317
rect 5906 257 5964 283
rect 6006 317 6064 343
rect 6006 283 6012 317
rect 6052 283 6064 317
rect 6006 257 6064 283
rect 6106 317 6164 343
rect 6106 283 6118 317
rect 6158 283 6164 317
rect 6106 257 6164 283
rect 6206 317 6264 343
rect 6206 283 6212 317
rect 6252 283 6264 317
rect 6206 257 6264 283
rect 6306 317 6364 343
rect 6306 283 6318 317
rect 6358 283 6364 317
rect 6306 257 6364 283
rect 6406 317 6464 343
rect 6406 283 6412 317
rect 6452 283 6464 317
rect 6406 257 6464 283
rect 6506 317 6564 343
rect 6506 283 6518 317
rect 6558 283 6564 317
rect 6506 257 6564 283
rect 6606 317 6664 343
rect 6606 283 6612 317
rect 6652 283 6664 317
rect 6606 257 6664 283
rect 6706 317 6764 343
rect 6706 283 6718 317
rect 6758 283 6764 317
rect 6706 257 6764 283
rect 6806 317 6864 343
rect 6806 283 6812 317
rect 6852 283 6864 317
rect 6806 257 6864 283
rect 6906 317 6964 343
rect 6906 283 6918 317
rect 6958 283 6964 317
rect 6906 257 6964 283
rect 7006 317 7064 343
rect 7006 283 7018 317
rect 7052 283 7064 317
rect 7006 257 7064 283
rect 7106 317 7164 343
rect 7106 283 7118 317
rect 7152 283 7164 317
rect 7106 257 7164 283
rect 7206 317 7264 343
rect 7206 283 7218 317
rect 7252 283 7264 317
rect 7206 257 7264 283
rect 7306 317 7364 343
rect 7306 283 7318 317
rect 7352 283 7364 317
rect 7306 257 7364 283
rect 7406 317 7464 343
rect 7406 283 7418 317
rect 7452 283 7464 317
rect 7406 257 7464 283
rect 7506 317 7564 343
rect 7506 283 7518 317
rect 7552 283 7564 317
rect 7506 257 7564 283
rect 7606 317 7664 343
rect 7606 283 7618 317
rect 7652 283 7664 317
rect 7606 257 7664 283
rect 7706 317 7764 343
rect 7706 283 7718 317
rect 7752 283 7764 317
rect 7706 257 7764 283
rect 7806 317 7864 343
rect 7806 283 7812 317
rect 7852 283 7864 317
rect 7806 257 7864 283
rect 7906 317 7964 343
rect 7906 283 7918 317
rect 7958 283 7964 317
rect 7906 257 7964 283
rect 8006 317 8064 343
rect 8006 283 8012 317
rect 8052 283 8064 317
rect 8006 257 8064 283
rect 8106 317 8164 343
rect 8106 283 8118 317
rect 8158 283 8164 317
rect 8106 257 8164 283
rect 8206 317 8264 343
rect 8206 283 8218 317
rect 8252 283 8264 317
rect 8206 257 8264 283
rect 8306 317 8364 343
rect 8306 283 8318 317
rect 8352 283 8364 317
rect 8306 257 8364 283
rect 8406 317 8464 343
rect 8406 283 8418 317
rect 8452 283 8464 317
rect 8406 257 8464 283
rect 8506 317 8564 343
rect 8506 283 8518 317
rect 8552 283 8564 317
rect 8506 257 8564 283
rect 8606 317 8664 343
rect 8606 283 8618 317
rect 8652 283 8664 317
rect 8606 257 8664 283
rect 8706 317 8764 343
rect 8706 283 8712 317
rect 8752 283 8764 317
rect 8706 257 8764 283
rect 8806 317 8864 343
rect 8806 283 8818 317
rect 8858 283 8864 317
rect 8806 257 8864 283
rect 8906 317 8964 343
rect 8906 283 8918 317
rect 8952 283 8964 317
rect 8906 257 8964 283
rect 9006 317 9064 343
rect 9006 283 9012 317
rect 9052 283 9064 317
rect 9006 257 9064 283
rect 9106 317 9164 343
rect 9106 283 9118 317
rect 9158 283 9164 317
rect 9106 257 9164 283
rect 9206 317 9264 343
rect 9206 283 9212 317
rect 9252 283 9264 317
rect 9206 257 9264 283
rect 9306 317 9364 343
rect 9306 283 9318 317
rect 9358 283 9364 317
rect 9306 257 9364 283
rect 9406 317 9464 343
rect 9406 283 9418 317
rect 9452 283 9464 317
rect 9406 257 9464 283
rect 9506 317 9564 343
rect 9506 283 9518 317
rect 9552 283 9564 317
rect 9506 257 9564 283
rect 9606 317 9664 343
rect 9606 283 9618 317
rect 9652 283 9664 317
rect 9606 257 9664 283
rect 9706 317 9764 343
rect 9706 283 9718 317
rect 9752 283 9764 317
rect 9706 257 9764 283
rect 9806 317 9864 343
rect 9806 283 9818 317
rect 9852 283 9864 317
rect 9806 257 9864 283
rect 9906 317 9964 343
rect 9906 283 9918 317
rect 9952 283 9964 317
rect 9906 257 9964 283
rect 10006 317 10064 343
rect 10006 283 10018 317
rect 10052 283 10064 317
rect 10006 257 10064 283
rect 10106 317 10164 343
rect 10106 283 10112 317
rect 10152 283 10164 317
rect 10106 257 10164 283
rect 10206 317 10264 343
rect 10206 283 10218 317
rect 10258 283 10264 317
rect 10206 257 10264 283
rect 10306 317 10364 343
rect 10306 283 10318 317
rect 10352 283 10364 317
rect 10306 257 10364 283
rect 10406 317 10464 343
rect 10406 283 10418 317
rect 10452 283 10464 317
rect 10406 257 10464 283
rect 10506 317 10564 343
rect 10506 283 10518 317
rect 10552 283 10564 317
rect 10506 257 10564 283
rect 10606 317 10664 343
rect 10606 283 10618 317
rect 10652 283 10664 317
rect 10606 257 10664 283
rect 10706 317 10764 343
rect 10706 283 10718 317
rect 10752 283 10764 317
rect 10706 257 10764 283
rect 10806 317 10864 343
rect 10806 283 10818 317
rect 10852 283 10864 317
rect 10806 257 10864 283
rect 10906 317 10964 343
rect 10906 283 10918 317
rect 10952 283 10964 317
rect 10906 257 10964 283
rect 11006 317 11064 343
rect 11006 283 11018 317
rect 11052 283 11064 317
rect 11006 257 11064 283
rect 11106 317 11164 343
rect 11106 283 11118 317
rect 11152 283 11164 317
rect 11106 257 11164 283
rect 11206 317 11264 343
rect 11206 283 11218 317
rect 11252 283 11264 317
rect 11206 257 11264 283
rect 11306 317 11364 343
rect 11306 283 11318 317
rect 11352 283 11364 317
rect 11306 257 11364 283
rect 11406 317 11464 343
rect 11406 283 11412 317
rect 11452 283 11464 317
rect 11406 257 11464 283
rect 11506 317 11564 343
rect 11506 283 11518 317
rect 11558 283 11564 317
rect 11506 257 11564 283
rect 11606 317 11664 343
rect 11606 283 11618 317
rect 11652 283 11664 317
rect 11606 257 11664 283
rect 11706 317 11764 343
rect 11706 283 11718 317
rect 11752 283 11764 317
rect 11706 257 11764 283
rect 11806 317 11864 343
rect 11806 283 11818 317
rect 11852 283 11864 317
rect 11806 257 11864 283
rect 11906 317 11964 343
rect 11906 283 11918 317
rect 11952 283 11964 317
rect 11906 257 11964 283
rect 12006 317 12064 343
rect 12006 283 12018 317
rect 12052 283 12064 317
rect 12006 257 12064 283
rect 12106 317 12164 343
rect 12106 283 12118 317
rect 12152 283 12164 317
rect 12106 257 12164 283
rect 12206 317 12264 343
rect 12206 283 12212 317
rect 12252 283 12264 317
rect 12206 257 12264 283
rect 12306 317 12364 343
rect 12306 283 12318 317
rect 12358 283 12364 317
rect 12306 257 12364 283
rect 12406 317 12464 343
rect 12406 283 12418 317
rect 12452 283 12464 317
rect 12406 257 12464 283
rect 12506 317 12564 343
rect 12506 283 12518 317
rect 12552 283 12564 317
rect 12506 257 12564 283
rect 12606 317 12664 343
rect 12606 283 12618 317
rect 12652 283 12664 317
rect 12606 257 12664 283
rect 12706 317 12764 343
rect 12706 283 12718 317
rect 12752 283 12764 317
rect 12706 257 12764 283
rect 12806 317 12864 343
rect 13018 336 13262 370
rect 12806 283 12818 317
rect 12852 283 12864 317
rect 12908 298 12916 332
rect 12958 298 12974 332
rect 13018 317 13052 336
rect 12806 257 12864 283
rect 13228 333 13262 336
rect 13228 317 13362 333
rect 13018 267 13052 283
rect 13096 268 13112 302
rect 13154 268 13162 302
rect 13262 283 13328 317
rect 13228 267 13362 283
rect 13428 317 13462 333
rect 13428 267 13462 283
rect 13528 317 13662 333
rect 13562 283 13628 317
rect 13528 267 13662 283
rect 6 177 64 203
rect 6 143 18 177
rect 58 143 64 177
rect 6 117 64 143
rect 106 177 164 203
rect 106 143 118 177
rect 152 143 164 177
rect 106 117 164 143
rect 206 177 264 203
rect 206 143 218 177
rect 252 143 264 177
rect 206 117 264 143
rect 306 177 364 203
rect 306 143 318 177
rect 352 143 364 177
rect 306 117 364 143
rect 406 177 464 203
rect 406 143 418 177
rect 452 143 464 177
rect 406 117 464 143
rect 506 177 564 203
rect 506 143 518 177
rect 552 143 564 177
rect 506 117 564 143
rect 606 177 664 203
rect 606 143 618 177
rect 652 143 664 177
rect 606 117 664 143
rect 706 177 764 203
rect 706 143 718 177
rect 752 143 764 177
rect 706 117 764 143
rect 806 177 864 203
rect 806 143 818 177
rect 852 143 864 177
rect 806 117 864 143
rect 906 177 964 203
rect 906 143 918 177
rect 952 143 964 177
rect 906 117 964 143
rect 1006 177 1064 203
rect 1006 143 1018 177
rect 1052 143 1064 177
rect 1006 117 1064 143
rect 1106 177 1164 203
rect 1106 143 1118 177
rect 1152 143 1164 177
rect 1106 117 1164 143
rect 1206 177 1264 203
rect 1206 143 1218 177
rect 1252 143 1264 177
rect 1206 117 1264 143
rect 1306 177 1364 203
rect 1306 143 1318 177
rect 1352 143 1364 177
rect 1306 117 1364 143
rect 1406 177 1464 203
rect 1406 143 1418 177
rect 1452 143 1464 177
rect 1406 117 1464 143
rect 1506 177 1564 203
rect 1506 143 1518 177
rect 1552 143 1564 177
rect 1506 117 1564 143
rect 1606 177 1664 203
rect 1606 143 1612 177
rect 1652 143 1664 177
rect 1606 117 1664 143
rect 1706 177 1764 203
rect 1706 143 1718 177
rect 1758 143 1764 177
rect 1706 117 1764 143
rect 1806 177 1864 203
rect 1806 143 1812 177
rect 1852 143 1864 177
rect 1806 117 1864 143
rect 1906 177 1964 203
rect 1906 143 1918 177
rect 1958 143 1964 177
rect 1906 117 1964 143
rect 2006 177 2064 203
rect 2006 143 2018 177
rect 2052 143 2064 177
rect 2006 117 2064 143
rect 2106 177 2164 203
rect 2106 143 2118 177
rect 2152 143 2164 177
rect 2106 117 2164 143
rect 2206 177 2264 203
rect 2206 143 2218 177
rect 2252 143 2264 177
rect 2206 117 2264 143
rect 2306 177 2364 203
rect 2306 143 2318 177
rect 2352 143 2364 177
rect 2306 117 2364 143
rect 2406 177 2464 203
rect 2406 143 2418 177
rect 2452 143 2464 177
rect 2406 117 2464 143
rect 2506 177 2564 203
rect 2506 143 2518 177
rect 2552 143 2564 177
rect 2506 117 2564 143
rect 2606 177 2664 203
rect 2606 143 2618 177
rect 2652 143 2664 177
rect 2606 117 2664 143
rect 2706 177 2764 203
rect 2706 143 2718 177
rect 2752 143 2764 177
rect 2706 117 2764 143
rect 2806 177 2864 203
rect 2806 143 2818 177
rect 2852 143 2864 177
rect 2806 117 2864 143
rect 2906 177 2964 203
rect 2906 143 2918 177
rect 2952 143 2964 177
rect 2906 117 2964 143
rect 3006 177 3064 203
rect 3006 143 3018 177
rect 3052 143 3064 177
rect 3006 117 3064 143
rect 3106 177 3164 203
rect 3106 143 3118 177
rect 3152 143 3164 177
rect 3106 117 3164 143
rect 3206 177 3264 203
rect 3206 143 3218 177
rect 3252 143 3264 177
rect 3206 117 3264 143
rect 3306 177 3364 203
rect 3306 143 3318 177
rect 3352 143 3364 177
rect 3306 117 3364 143
rect 3406 177 3464 203
rect 3406 143 3418 177
rect 3452 143 3464 177
rect 3406 117 3464 143
rect 3506 177 3564 203
rect 3506 143 3518 177
rect 3552 143 3564 177
rect 3506 117 3564 143
rect 3606 177 3664 203
rect 3606 143 3618 177
rect 3652 143 3664 177
rect 3606 117 3664 143
rect 3706 177 3764 203
rect 3706 143 3718 177
rect 3752 143 3764 177
rect 3706 117 3764 143
rect 3806 177 3864 203
rect 3806 143 3818 177
rect 3852 143 3864 177
rect 3806 117 3864 143
rect 3906 177 3964 203
rect 3906 143 3918 177
rect 3952 143 3964 177
rect 3906 117 3964 143
rect 4006 177 4064 203
rect 4006 143 4018 177
rect 4052 143 4064 177
rect 4006 117 4064 143
rect 4106 177 4164 203
rect 4106 143 4118 177
rect 4152 143 4164 177
rect 4106 117 4164 143
rect 4206 177 4264 203
rect 4206 143 4218 177
rect 4252 143 4264 177
rect 4206 117 4264 143
rect 4306 177 4364 203
rect 4306 143 4318 177
rect 4352 143 4364 177
rect 4306 117 4364 143
rect 4406 177 4464 203
rect 4406 143 4418 177
rect 4452 143 4464 177
rect 4406 117 4464 143
rect 4506 177 4564 203
rect 4506 143 4518 177
rect 4552 143 4564 177
rect 4506 117 4564 143
rect 4606 177 4664 203
rect 4606 143 4618 177
rect 4652 143 4664 177
rect 4606 117 4664 143
rect 4706 177 4764 203
rect 4706 143 4718 177
rect 4752 143 4764 177
rect 4706 117 4764 143
rect 4806 177 4864 203
rect 4806 143 4818 177
rect 4852 143 4864 177
rect 4806 117 4864 143
rect 4906 177 4964 203
rect 4906 143 4918 177
rect 4952 143 4964 177
rect 4906 117 4964 143
rect 5006 177 5064 203
rect 5006 143 5018 177
rect 5052 143 5064 177
rect 5006 117 5064 143
rect 5106 177 5164 203
rect 5106 143 5118 177
rect 5152 143 5164 177
rect 5106 117 5164 143
rect 5206 177 5264 203
rect 5206 143 5218 177
rect 5252 143 5264 177
rect 5206 117 5264 143
rect 5306 177 5364 203
rect 5306 143 5318 177
rect 5352 143 5364 177
rect 5306 117 5364 143
rect 5406 177 5464 203
rect 5406 143 5418 177
rect 5452 143 5464 177
rect 5406 117 5464 143
rect 5506 177 5564 203
rect 5506 143 5518 177
rect 5552 143 5564 177
rect 5506 117 5564 143
rect 5606 177 5664 203
rect 5606 143 5618 177
rect 5652 143 5664 177
rect 5606 117 5664 143
rect 5706 177 5764 203
rect 5706 143 5718 177
rect 5752 143 5764 177
rect 5706 117 5764 143
rect 5806 177 5864 203
rect 5806 143 5818 177
rect 5852 143 5864 177
rect 5806 117 5864 143
rect 5906 177 5964 203
rect 5906 143 5918 177
rect 5952 143 5964 177
rect 5906 117 5964 143
rect 6006 177 6064 203
rect 6006 143 6018 177
rect 6052 143 6064 177
rect 6006 117 6064 143
rect 6106 177 6164 203
rect 6106 143 6118 177
rect 6152 143 6164 177
rect 6106 117 6164 143
rect 6206 177 6264 203
rect 6206 143 6218 177
rect 6252 143 6264 177
rect 6206 117 6264 143
rect 6306 177 6364 203
rect 6306 143 6318 177
rect 6352 143 6364 177
rect 6306 117 6364 143
rect 6406 177 6464 203
rect 6406 143 6418 177
rect 6452 143 6464 177
rect 6406 117 6464 143
rect 6506 177 6564 203
rect 6506 143 6518 177
rect 6552 143 6564 177
rect 6506 117 6564 143
rect 6606 177 6664 203
rect 6606 143 6618 177
rect 6652 143 6664 177
rect 6606 117 6664 143
rect 6706 177 6764 203
rect 6706 143 6718 177
rect 6752 143 6764 177
rect 6706 117 6764 143
rect 6806 177 6864 203
rect 6806 143 6818 177
rect 6852 143 6864 177
rect 6806 117 6864 143
rect 6906 177 6964 203
rect 6906 143 6918 177
rect 6952 143 6964 177
rect 6906 117 6964 143
rect 7006 177 7064 203
rect 7006 143 7012 177
rect 7052 143 7064 177
rect 7006 117 7064 143
rect 7106 177 7164 203
rect 7106 143 7118 177
rect 7158 143 7164 177
rect 7106 117 7164 143
rect 7206 177 7264 203
rect 7206 143 7218 177
rect 7252 143 7264 177
rect 7206 117 7264 143
rect 7306 177 7364 203
rect 7306 143 7318 177
rect 7352 143 7364 177
rect 7306 117 7364 143
rect 7406 177 7464 203
rect 7406 143 7418 177
rect 7452 143 7464 177
rect 7406 117 7464 143
rect 7506 177 7564 203
rect 7506 143 7518 177
rect 7552 143 7564 177
rect 7506 117 7564 143
rect 7606 177 7664 203
rect 7606 143 7618 177
rect 7652 143 7664 177
rect 7606 117 7664 143
rect 7706 177 7764 203
rect 7706 143 7718 177
rect 7752 143 7764 177
rect 7706 117 7764 143
rect 7806 177 7864 203
rect 7806 143 7818 177
rect 7852 143 7864 177
rect 7806 117 7864 143
rect 7906 177 7964 203
rect 7906 143 7918 177
rect 7952 143 7964 177
rect 7906 117 7964 143
rect 8006 177 8064 203
rect 8006 143 8018 177
rect 8052 143 8064 177
rect 8006 117 8064 143
rect 8106 177 8164 203
rect 8106 143 8118 177
rect 8152 143 8164 177
rect 8106 117 8164 143
rect 8206 177 8264 203
rect 8206 143 8218 177
rect 8252 143 8264 177
rect 8206 117 8264 143
rect 8306 177 8364 203
rect 8306 143 8318 177
rect 8352 143 8364 177
rect 8306 117 8364 143
rect 8406 177 8464 203
rect 8406 143 8418 177
rect 8452 143 8464 177
rect 8406 117 8464 143
rect 8506 177 8564 203
rect 8506 143 8518 177
rect 8552 143 8564 177
rect 8506 117 8564 143
rect 8606 177 8664 203
rect 8606 143 8618 177
rect 8652 143 8664 177
rect 8606 117 8664 143
rect 8706 177 8764 203
rect 8706 143 8718 177
rect 8752 143 8764 177
rect 8706 117 8764 143
rect 8806 177 8864 203
rect 8806 143 8818 177
rect 8852 143 8864 177
rect 8806 117 8864 143
rect 8906 177 8964 203
rect 8906 143 8918 177
rect 8952 143 8964 177
rect 8906 117 8964 143
rect 9006 177 9064 203
rect 9006 143 9018 177
rect 9052 143 9064 177
rect 9006 117 9064 143
rect 9106 177 9164 203
rect 9106 143 9118 177
rect 9152 143 9164 177
rect 9106 117 9164 143
rect 9206 177 9264 203
rect 9206 143 9218 177
rect 9252 143 9264 177
rect 9206 117 9264 143
rect 9306 177 9364 203
rect 9306 143 9318 177
rect 9352 143 9364 177
rect 9306 117 9364 143
rect 9406 177 9464 203
rect 9406 143 9418 177
rect 9452 143 9464 177
rect 9406 117 9464 143
rect 9506 177 9564 203
rect 9506 143 9518 177
rect 9552 143 9564 177
rect 9506 117 9564 143
rect 9606 177 9664 203
rect 9606 143 9618 177
rect 9652 143 9664 177
rect 9606 117 9664 143
rect 9706 177 9764 203
rect 9706 143 9718 177
rect 9752 143 9764 177
rect 9706 117 9764 143
rect 9806 177 9864 203
rect 9806 143 9818 177
rect 9852 143 9864 177
rect 9806 117 9864 143
rect 9906 177 9964 203
rect 9906 143 9918 177
rect 9952 143 9964 177
rect 9906 117 9964 143
rect 10006 177 10064 203
rect 10006 143 10018 177
rect 10052 143 10064 177
rect 10006 117 10064 143
rect 10106 177 10164 203
rect 10106 143 10118 177
rect 10152 143 10164 177
rect 10106 117 10164 143
rect 10206 177 10264 203
rect 10206 143 10218 177
rect 10252 143 10264 177
rect 10206 117 10264 143
rect 10306 177 10364 203
rect 10306 143 10318 177
rect 10352 143 10364 177
rect 10306 117 10364 143
rect 10406 177 10464 203
rect 10406 143 10418 177
rect 10452 143 10464 177
rect 10406 117 10464 143
rect 10506 177 10564 203
rect 10506 143 10518 177
rect 10552 143 10564 177
rect 10506 117 10564 143
rect 10606 177 10664 203
rect 10606 143 10618 177
rect 10652 143 10664 177
rect 10606 117 10664 143
rect 10706 177 10764 203
rect 10706 143 10718 177
rect 10752 143 10764 177
rect 10706 117 10764 143
rect 10806 177 10864 203
rect 10806 143 10818 177
rect 10852 143 10864 177
rect 10806 117 10864 143
rect 10906 177 10964 203
rect 10906 143 10918 177
rect 10952 143 10964 177
rect 10906 117 10964 143
rect 11006 177 11064 203
rect 11006 143 11018 177
rect 11052 143 11064 177
rect 11006 117 11064 143
rect 11106 177 11164 203
rect 11106 143 11118 177
rect 11152 143 11164 177
rect 11106 117 11164 143
rect 11206 177 11264 203
rect 11206 143 11218 177
rect 11252 143 11264 177
rect 11206 117 11264 143
rect 11306 177 11364 203
rect 11306 143 11318 177
rect 11352 143 11364 177
rect 11306 117 11364 143
rect 11406 177 11464 203
rect 11406 143 11412 177
rect 11452 143 11464 177
rect 11406 117 11464 143
rect 11506 177 11564 203
rect 11506 143 11518 177
rect 11558 143 11564 177
rect 11506 117 11564 143
rect 11606 177 11664 203
rect 11606 143 11618 177
rect 11652 143 11664 177
rect 11606 117 11664 143
rect 11706 177 11764 203
rect 11706 143 11718 177
rect 11752 143 11764 177
rect 11706 117 11764 143
rect 11806 177 11864 203
rect 11806 143 11818 177
rect 11852 143 11864 177
rect 11806 117 11864 143
rect 11906 177 11964 203
rect 11906 143 11918 177
rect 11952 143 11964 177
rect 11906 117 11964 143
rect 12006 177 12064 203
rect 12006 143 12018 177
rect 12052 143 12064 177
rect 12006 117 12064 143
rect 12106 177 12164 203
rect 12106 143 12118 177
rect 12152 143 12164 177
rect 12106 117 12164 143
rect 12206 177 12264 203
rect 12206 143 12218 177
rect 12252 143 12264 177
rect 12206 117 12264 143
rect 12306 177 12364 203
rect 12306 143 12318 177
rect 12352 143 12364 177
rect 12306 117 12364 143
rect 12406 177 12464 203
rect 12406 143 12418 177
rect 12452 143 12464 177
rect 12406 117 12464 143
rect 12506 177 12564 203
rect 12506 143 12518 177
rect 12552 143 12564 177
rect 12506 117 12564 143
rect 12606 177 12664 203
rect 12606 143 12618 177
rect 12652 143 12664 177
rect 12606 117 12664 143
rect 12706 177 12764 203
rect 12706 143 12718 177
rect 12752 143 12764 177
rect 12706 117 12764 143
rect 12806 177 12864 203
rect 13018 196 13262 230
rect 12806 143 12818 177
rect 12852 143 12864 177
rect 12908 158 12916 192
rect 12958 158 12974 192
rect 13018 177 13052 196
rect 12806 117 12864 143
rect 13228 177 13262 196
rect 13018 127 13052 143
rect 13096 128 13112 162
rect 13154 128 13162 162
rect 13228 127 13262 143
rect 13328 177 13462 193
rect 13362 143 13428 177
rect 13328 127 13462 143
rect 13528 177 13662 193
rect 13562 143 13628 177
rect 13528 127 13662 143
rect 8 20 18 54
rect 52 20 118 54
rect 152 20 168 54
rect 208 36 218 70
rect 252 36 318 70
rect 352 36 368 70
rect 408 20 418 54
rect 452 20 518 54
rect 552 20 568 54
rect 608 36 618 70
rect 652 36 718 70
rect 752 36 768 70
rect 808 20 818 54
rect 852 20 918 54
rect 952 20 968 54
rect 1008 36 1018 70
rect 1052 36 1118 70
rect 1152 36 1168 70
rect 1208 20 1218 54
rect 1252 20 1318 54
rect 1352 20 1368 54
rect 1408 36 1418 70
rect 1452 36 1518 70
rect 1552 36 1568 70
rect 1608 20 1618 54
rect 1652 20 1718 54
rect 1752 20 1768 54
rect 1808 36 1818 70
rect 1852 36 1918 70
rect 1952 36 1968 70
rect 2008 20 2018 54
rect 2052 20 2118 54
rect 2152 20 2168 54
rect 2208 36 2218 70
rect 2252 36 2318 70
rect 2352 36 2368 70
rect 2408 20 2418 54
rect 2452 20 2518 54
rect 2552 20 2568 54
rect 2608 36 2618 70
rect 2652 36 2718 70
rect 2752 36 2768 70
rect 2808 20 2818 54
rect 2852 20 2918 54
rect 2952 20 2968 54
rect 3008 36 3018 70
rect 3052 36 3118 70
rect 3152 36 3168 70
rect 3208 20 3218 54
rect 3252 20 3318 54
rect 3352 20 3368 54
rect 3408 36 3418 70
rect 3452 36 3518 70
rect 3552 36 3568 70
rect 3608 20 3618 54
rect 3652 20 3718 54
rect 3752 20 3768 54
rect 3808 36 3818 70
rect 3852 36 3918 70
rect 3952 36 3968 70
rect 4008 20 4018 54
rect 4052 20 4118 54
rect 4152 20 4168 54
rect 4208 36 4218 70
rect 4252 36 4318 70
rect 4352 36 4368 70
rect 4408 20 4418 54
rect 4452 20 4518 54
rect 4552 20 4568 54
rect 4608 36 4618 70
rect 4652 36 4718 70
rect 4752 36 4768 70
rect 4808 20 4818 54
rect 4852 20 4918 54
rect 4952 20 4968 54
rect 5008 36 5018 70
rect 5052 36 5118 70
rect 5152 36 5168 70
rect 5208 20 5218 54
rect 5252 20 5318 54
rect 5352 20 5368 54
rect 5408 36 5418 70
rect 5452 36 5518 70
rect 5552 36 5568 70
rect 5608 20 5618 54
rect 5652 20 5718 54
rect 5752 20 5768 54
rect 5808 36 5818 70
rect 5852 36 5918 70
rect 5952 36 5968 70
rect 6008 20 6018 54
rect 6052 20 6118 54
rect 6152 20 6168 54
rect 6208 36 6218 70
rect 6252 36 6318 70
rect 6352 36 6368 70
rect 6408 20 6418 54
rect 6452 20 6518 54
rect 6552 20 6568 54
rect 6608 36 6618 70
rect 6652 36 6718 70
rect 6752 36 6768 70
rect 6808 20 6818 54
rect 6852 20 6918 54
rect 6952 20 6968 54
rect 7008 36 7018 70
rect 7052 36 7118 70
rect 7152 36 7168 70
rect 7208 20 7218 54
rect 7252 20 7318 54
rect 7352 20 7368 54
rect 7408 36 7418 70
rect 7452 36 7518 70
rect 7552 36 7568 70
rect 7608 20 7618 54
rect 7652 20 7718 54
rect 7752 20 7768 54
rect 7808 36 7818 70
rect 7852 36 7918 70
rect 7952 36 7968 70
rect 8008 20 8018 54
rect 8052 20 8118 54
rect 8152 20 8168 54
rect 8208 36 8218 70
rect 8252 36 8318 70
rect 8352 36 8368 70
rect 8408 20 8418 54
rect 8452 20 8518 54
rect 8552 20 8568 54
rect 8608 36 8618 70
rect 8652 36 8718 70
rect 8752 36 8768 70
rect 8808 20 8818 54
rect 8852 20 8918 54
rect 8952 20 8968 54
rect 9008 36 9018 70
rect 9052 36 9118 70
rect 9152 36 9168 70
rect 9208 20 9218 54
rect 9252 20 9318 54
rect 9352 20 9368 54
rect 9408 36 9418 70
rect 9452 36 9518 70
rect 9552 36 9568 70
rect 9608 20 9618 54
rect 9652 20 9718 54
rect 9752 20 9768 54
rect 9808 36 9818 70
rect 9852 36 9918 70
rect 9952 36 9968 70
rect 10008 20 10018 54
rect 10052 20 10118 54
rect 10152 20 10168 54
rect 10208 36 10218 70
rect 10252 36 10318 70
rect 10352 36 10368 70
rect 10408 20 10418 54
rect 10452 20 10518 54
rect 10552 20 10568 54
rect 10608 36 10618 70
rect 10652 36 10718 70
rect 10752 36 10768 70
rect 10808 20 10818 54
rect 10852 20 10918 54
rect 10952 20 10968 54
rect 11008 36 11018 70
rect 11052 36 11118 70
rect 11152 36 11168 70
rect 11208 20 11218 54
rect 11252 20 11318 54
rect 11352 20 11368 54
rect 11408 36 11418 70
rect 11452 36 11518 70
rect 11552 36 11568 70
rect 11608 20 11618 54
rect 11652 20 11718 54
rect 11752 20 11768 54
rect 11808 36 11818 70
rect 11852 36 11918 70
rect 11952 36 11968 70
rect 12008 20 12018 54
rect 12052 20 12118 54
rect 12152 20 12168 54
rect 12208 36 12218 70
rect 12252 36 12318 70
rect 12352 36 12368 70
rect 12408 20 12418 54
rect 12452 20 12518 54
rect 12552 20 12568 54
rect 12608 36 12618 70
rect 12652 36 12718 70
rect 12752 36 12768 70
rect 12916 51 12968 68
rect 12950 34 12968 51
rect 13002 34 13018 68
rect 13052 34 13068 68
rect 13102 39 13120 68
rect 13102 34 13154 39
rect 13262 34 13278 68
rect 13312 34 13328 68
rect 13362 34 13378 68
rect 13412 34 13428 68
rect 13462 34 13478 68
rect 13512 34 13528 68
rect 13562 34 13578 68
rect 13612 34 13628 68
rect -132 -61 -116 -27
rect -82 -60 -48 -27
rect -14 -61 84 -27
rect 118 -60 152 -27
rect -82 -132 -48 -94
rect 186 -61 284 -27
rect 318 -60 352 -27
rect -82 -214 -48 -183
rect 18 -133 52 -95
rect 18 -214 52 -183
rect 118 -132 152 -94
rect 386 -61 484 -27
rect 518 -60 552 -27
rect 118 -214 152 -183
rect 218 -133 252 -95
rect 218 -214 252 -183
rect 318 -132 352 -94
rect 586 -61 684 -27
rect 718 -60 752 -27
rect 318 -214 352 -183
rect 418 -133 452 -95
rect 418 -214 452 -183
rect 518 -132 552 -94
rect 786 -61 884 -27
rect 918 -60 952 -27
rect 518 -214 552 -183
rect 618 -133 652 -95
rect 618 -214 652 -183
rect 718 -132 752 -94
rect 986 -61 1084 -27
rect 1118 -60 1152 -27
rect 718 -214 752 -183
rect 818 -133 852 -95
rect 818 -214 852 -183
rect 918 -132 952 -94
rect 1186 -61 1284 -27
rect 1318 -60 1352 -27
rect 918 -214 952 -183
rect 1018 -133 1052 -95
rect 1018 -214 1052 -183
rect 1118 -132 1152 -94
rect 1386 -61 1484 -27
rect 1518 -60 1552 -27
rect 1118 -214 1152 -183
rect 1218 -133 1252 -95
rect 1218 -214 1252 -183
rect 1318 -132 1352 -94
rect 1586 -61 1684 -27
rect 1718 -60 1752 -27
rect 1318 -214 1352 -183
rect 1418 -133 1452 -95
rect 1418 -214 1452 -183
rect 1518 -132 1552 -94
rect 1786 -61 1884 -27
rect 1918 -60 1952 -27
rect 1518 -214 1552 -183
rect 1618 -133 1652 -95
rect 1618 -214 1652 -183
rect 1718 -132 1752 -94
rect 1986 -61 2084 -27
rect 2118 -60 2152 -27
rect 1718 -214 1752 -183
rect 1818 -133 1852 -95
rect 1818 -214 1852 -183
rect 1918 -132 1952 -94
rect 2186 -61 2284 -27
rect 2318 -60 2352 -27
rect 1918 -214 1952 -183
rect 2018 -133 2052 -95
rect 2018 -214 2052 -183
rect 2118 -132 2152 -94
rect 2386 -61 2484 -27
rect 2518 -60 2552 -27
rect 2118 -214 2152 -183
rect 2218 -133 2252 -95
rect 2218 -214 2252 -183
rect 2318 -132 2352 -94
rect 2586 -61 2684 -27
rect 2718 -60 2752 -27
rect 2318 -214 2352 -183
rect 2418 -133 2452 -95
rect 2418 -214 2452 -183
rect 2518 -132 2552 -94
rect 2786 -61 2884 -27
rect 2918 -60 2952 -27
rect 2518 -214 2552 -183
rect 2618 -133 2652 -95
rect 2618 -214 2652 -183
rect 2718 -132 2752 -94
rect 2986 -61 3084 -27
rect 3118 -60 3152 -27
rect 2718 -214 2752 -183
rect 2818 -133 2852 -95
rect 2818 -214 2852 -183
rect 2918 -132 2952 -94
rect 3186 -61 3284 -27
rect 3318 -60 3352 -27
rect 2918 -214 2952 -183
rect 3018 -133 3052 -95
rect 3018 -214 3052 -183
rect 3118 -132 3152 -94
rect 3386 -61 3484 -27
rect 3518 -60 3552 -27
rect 3118 -214 3152 -183
rect 3218 -133 3252 -95
rect 3218 -214 3252 -183
rect 3318 -132 3352 -94
rect 3586 -61 3684 -27
rect 3718 -60 3752 -27
rect 3318 -214 3352 -183
rect 3418 -133 3452 -95
rect 3418 -214 3452 -183
rect 3518 -132 3552 -94
rect 3786 -61 3884 -27
rect 3918 -60 3952 -27
rect 3518 -214 3552 -183
rect 3618 -133 3652 -95
rect 3618 -214 3652 -183
rect 3718 -132 3752 -94
rect 3986 -61 4084 -27
rect 4118 -60 4152 -27
rect 3718 -214 3752 -183
rect 3818 -133 3852 -95
rect 3818 -214 3852 -183
rect 3918 -132 3952 -94
rect 4186 -61 4284 -27
rect 4318 -60 4352 -27
rect 3918 -214 3952 -183
rect 4018 -133 4052 -95
rect 4018 -214 4052 -183
rect 4118 -132 4152 -94
rect 4386 -61 4484 -27
rect 4518 -60 4552 -27
rect 4118 -214 4152 -183
rect 4218 -133 4252 -95
rect 4218 -214 4252 -183
rect 4318 -132 4352 -94
rect 4586 -61 4684 -27
rect 4718 -60 4752 -27
rect 4318 -214 4352 -183
rect 4418 -133 4452 -95
rect 4418 -214 4452 -183
rect 4518 -132 4552 -94
rect 4786 -61 4884 -27
rect 4918 -60 4952 -27
rect 4518 -214 4552 -183
rect 4618 -133 4652 -95
rect 4618 -214 4652 -183
rect 4718 -132 4752 -94
rect 4986 -61 5084 -27
rect 5118 -60 5152 -27
rect 4718 -214 4752 -183
rect 4818 -133 4852 -95
rect 4818 -214 4852 -183
rect 4918 -132 4952 -94
rect 5186 -61 5284 -27
rect 5318 -60 5352 -27
rect 4918 -214 4952 -183
rect 5018 -133 5052 -95
rect 5018 -214 5052 -183
rect 5118 -132 5152 -94
rect 5386 -61 5484 -27
rect 5518 -60 5552 -27
rect 5118 -214 5152 -183
rect 5218 -133 5252 -95
rect 5218 -214 5252 -183
rect 5318 -132 5352 -94
rect 5586 -61 5684 -27
rect 5718 -60 5752 -27
rect 5318 -214 5352 -183
rect 5418 -133 5452 -95
rect 5418 -214 5452 -183
rect 5518 -132 5552 -94
rect 5786 -61 5884 -27
rect 5918 -60 5952 -27
rect 5518 -214 5552 -183
rect 5618 -133 5652 -95
rect 5618 -214 5652 -183
rect 5718 -132 5752 -94
rect 5986 -61 6084 -27
rect 6118 -60 6152 -27
rect 5718 -214 5752 -183
rect 5818 -133 5852 -95
rect 5818 -214 5852 -183
rect 5918 -132 5952 -94
rect 6186 -61 6284 -27
rect 6318 -60 6352 -27
rect 5918 -214 5952 -183
rect 6018 -133 6052 -95
rect 6018 -214 6052 -183
rect 6118 -132 6152 -94
rect 6386 -61 6484 -27
rect 6518 -60 6552 -27
rect 6118 -214 6152 -183
rect 6218 -133 6252 -95
rect 6218 -214 6252 -183
rect 6318 -132 6352 -94
rect 6586 -61 6684 -27
rect 6718 -60 6752 -27
rect 6318 -214 6352 -183
rect 6418 -133 6452 -95
rect 6418 -214 6452 -183
rect 6518 -132 6552 -94
rect 6786 -61 6884 -27
rect 6918 -60 6952 -27
rect 6518 -214 6552 -183
rect 6618 -133 6652 -95
rect 6618 -214 6652 -183
rect 6718 -132 6752 -94
rect 6986 -61 7084 -27
rect 7118 -60 7152 -27
rect 6718 -214 6752 -183
rect 6818 -133 6852 -95
rect 6818 -214 6852 -183
rect 6918 -132 6952 -94
rect 7186 -61 7284 -27
rect 7318 -60 7352 -27
rect 6918 -214 6952 -183
rect 7018 -133 7052 -95
rect 7018 -214 7052 -183
rect 7118 -132 7152 -94
rect 7386 -61 7484 -27
rect 7518 -60 7552 -27
rect 7118 -214 7152 -183
rect 7218 -133 7252 -95
rect 7218 -214 7252 -183
rect 7318 -132 7352 -94
rect 7586 -61 7684 -27
rect 7718 -60 7752 -27
rect 7318 -214 7352 -183
rect 7418 -133 7452 -95
rect 7418 -214 7452 -183
rect 7518 -132 7552 -94
rect 7786 -61 7884 -27
rect 7918 -60 7952 -27
rect 7518 -214 7552 -183
rect 7618 -133 7652 -95
rect 7618 -214 7652 -183
rect 7718 -132 7752 -94
rect 7986 -61 8084 -27
rect 8118 -60 8152 -27
rect 7718 -214 7752 -183
rect 7818 -133 7852 -95
rect 7818 -214 7852 -183
rect 7918 -132 7952 -94
rect 8186 -61 8284 -27
rect 8318 -60 8352 -27
rect 7918 -214 7952 -183
rect 8018 -133 8052 -95
rect 8018 -214 8052 -183
rect 8118 -132 8152 -94
rect 8386 -61 8484 -27
rect 8518 -60 8552 -27
rect 8118 -214 8152 -183
rect 8218 -133 8252 -95
rect 8218 -214 8252 -183
rect 8318 -132 8352 -94
rect 8586 -61 8684 -27
rect 8718 -60 8752 -27
rect 8318 -214 8352 -183
rect 8418 -133 8452 -95
rect 8418 -214 8452 -183
rect 8518 -132 8552 -94
rect 8786 -61 8884 -27
rect 8918 -60 8952 -27
rect 8518 -214 8552 -183
rect 8618 -133 8652 -95
rect 8618 -214 8652 -183
rect 8718 -132 8752 -94
rect 8986 -61 9084 -27
rect 9118 -60 9152 -27
rect 8718 -214 8752 -183
rect 8818 -133 8852 -95
rect 8818 -214 8852 -183
rect 8918 -132 8952 -94
rect 9186 -61 9284 -27
rect 9318 -60 9352 -27
rect 8918 -214 8952 -183
rect 9018 -133 9052 -95
rect 9018 -214 9052 -183
rect 9118 -132 9152 -94
rect 9386 -61 9484 -27
rect 9518 -60 9552 -27
rect 9118 -214 9152 -183
rect 9218 -133 9252 -95
rect 9218 -214 9252 -183
rect 9318 -132 9352 -94
rect 9586 -61 9684 -27
rect 9718 -60 9752 -27
rect 9318 -214 9352 -183
rect 9418 -133 9452 -95
rect 9418 -214 9452 -183
rect 9518 -132 9552 -94
rect 9786 -61 9884 -27
rect 9918 -60 9952 -27
rect 9518 -214 9552 -183
rect 9618 -133 9652 -95
rect 9618 -214 9652 -183
rect 9718 -132 9752 -94
rect 9986 -61 10084 -27
rect 10118 -60 10152 -27
rect 9718 -214 9752 -183
rect 9818 -133 9852 -95
rect 9818 -214 9852 -183
rect 9918 -132 9952 -94
rect 10186 -61 10284 -27
rect 10318 -60 10352 -27
rect 9918 -214 9952 -183
rect 10018 -133 10052 -95
rect 10018 -214 10052 -183
rect 10118 -132 10152 -94
rect 10386 -61 10484 -27
rect 10518 -60 10552 -27
rect 10118 -214 10152 -183
rect 10218 -133 10252 -95
rect 10218 -214 10252 -183
rect 10318 -132 10352 -94
rect 10586 -61 10684 -27
rect 10718 -60 10752 -27
rect 10318 -214 10352 -183
rect 10418 -133 10452 -95
rect 10418 -214 10452 -183
rect 10518 -132 10552 -94
rect 10786 -61 10884 -27
rect 10918 -60 10952 -27
rect 10518 -214 10552 -183
rect 10618 -133 10652 -95
rect 10618 -214 10652 -183
rect 10718 -132 10752 -94
rect 10986 -61 11084 -27
rect 11118 -60 11152 -27
rect 10718 -214 10752 -183
rect 10818 -133 10852 -95
rect 10818 -214 10852 -183
rect 10918 -132 10952 -94
rect 11186 -61 11284 -27
rect 11318 -60 11352 -27
rect 10918 -214 10952 -183
rect 11018 -133 11052 -95
rect 11018 -214 11052 -183
rect 11118 -132 11152 -94
rect 11386 -61 11484 -27
rect 11518 -60 11552 -27
rect 11118 -214 11152 -183
rect 11218 -133 11252 -95
rect 11218 -214 11252 -183
rect 11318 -132 11352 -94
rect 11586 -61 11684 -27
rect 11718 -60 11752 -27
rect 11318 -214 11352 -183
rect 11418 -133 11452 -95
rect 11418 -214 11452 -183
rect 11518 -132 11552 -94
rect 11786 -61 11884 -27
rect 11918 -60 11952 -27
rect 11518 -214 11552 -183
rect 11618 -133 11652 -95
rect 11618 -214 11652 -183
rect 11718 -132 11752 -94
rect 11986 -61 12084 -27
rect 12118 -60 12152 -27
rect 11718 -214 11752 -183
rect 11818 -133 11852 -95
rect 11818 -214 11852 -183
rect 11918 -132 11952 -94
rect 12186 -61 12284 -27
rect 12318 -60 12352 -27
rect 11918 -214 11952 -183
rect 12018 -133 12052 -95
rect 12018 -214 12052 -183
rect 12118 -132 12152 -94
rect 12386 -61 12484 -27
rect 12518 -60 12552 -27
rect 12118 -214 12152 -183
rect 12218 -133 12252 -95
rect 12218 -214 12252 -183
rect 12318 -132 12352 -94
rect 12586 -61 12684 -27
rect 12718 -60 12752 -27
rect 12318 -214 12352 -183
rect 12418 -133 12452 -95
rect 12418 -214 12452 -183
rect 12518 -132 12552 -94
rect 12786 -61 12802 -27
rect 12518 -214 12552 -183
rect 12618 -133 12652 -95
rect 12618 -214 12652 -183
rect 12718 -132 12752 -94
rect 12718 -214 12752 -183
rect 14548 -149 14564 -115
rect 14598 -149 14632 -115
rect 14666 -149 14682 -115
rect 14548 -208 14682 -149
rect 14824 -149 14847 -115
rect 14881 -149 14915 -115
rect 14949 -149 14983 -115
rect 15017 -149 15051 -115
rect 15085 -149 15108 -115
rect 14824 -208 15108 -149
rect 15234 -149 15257 -115
rect 15291 -149 15325 -115
rect 15359 -149 15393 -115
rect 15427 -149 15461 -115
rect 15495 -149 15518 -115
rect 15234 -208 15518 -149
rect 15660 -149 15676 -115
rect 15710 -149 15744 -115
rect 15778 -149 15794 -115
rect 15660 -208 15794 -149
rect 14532 -242 14558 -208
rect 14596 -242 14630 -208
rect 14664 -242 14694 -208
rect 14808 -242 14842 -208
rect 14881 -242 14914 -208
rect 14949 -242 14983 -208
rect 15020 -242 15051 -208
rect 15092 -242 15124 -208
rect 15218 -242 15249 -208
rect 15291 -242 15321 -208
rect 15359 -242 15393 -208
rect 15427 -242 15461 -208
rect 15499 -242 15534 -208
rect 15648 -242 15677 -208
rect 15712 -242 15746 -208
rect 15783 -242 15810 -208
rect -32 -282 18 -248
rect 52 -282 68 -248
rect 168 -282 218 -248
rect 252 -282 268 -248
rect 368 -282 418 -248
rect 452 -282 468 -248
rect 568 -282 618 -248
rect 652 -282 668 -248
rect 768 -282 818 -248
rect 852 -282 868 -248
rect 968 -282 1018 -248
rect 1052 -282 1068 -248
rect 1168 -282 1218 -248
rect 1252 -282 1268 -248
rect 1368 -282 1418 -248
rect 1452 -282 1468 -248
rect 1568 -282 1618 -248
rect 1652 -282 1668 -248
rect 1768 -282 1818 -248
rect 1852 -282 1868 -248
rect 1968 -282 2018 -248
rect 2052 -282 2068 -248
rect 2168 -282 2218 -248
rect 2252 -282 2268 -248
rect 2368 -282 2418 -248
rect 2452 -282 2468 -248
rect 2568 -282 2618 -248
rect 2652 -282 2668 -248
rect 2768 -282 2818 -248
rect 2852 -282 2868 -248
rect 2968 -282 3018 -248
rect 3052 -282 3068 -248
rect 3168 -282 3218 -248
rect 3252 -282 3268 -248
rect 3368 -282 3418 -248
rect 3452 -282 3468 -248
rect 3568 -282 3618 -248
rect 3652 -282 3668 -248
rect 3768 -282 3818 -248
rect 3852 -282 3868 -248
rect 3968 -282 4018 -248
rect 4052 -282 4068 -248
rect 4168 -282 4218 -248
rect 4252 -282 4268 -248
rect 4368 -282 4418 -248
rect 4452 -282 4468 -248
rect 4568 -282 4618 -248
rect 4652 -282 4668 -248
rect 4768 -282 4818 -248
rect 4852 -282 4868 -248
rect 4968 -282 5018 -248
rect 5052 -282 5068 -248
rect 5168 -282 5218 -248
rect 5252 -282 5268 -248
rect 5368 -282 5418 -248
rect 5452 -282 5468 -248
rect 5568 -282 5618 -248
rect 5652 -282 5668 -248
rect 5768 -282 5818 -248
rect 5852 -282 5868 -248
rect 5968 -282 6018 -248
rect 6052 -282 6068 -248
rect 6168 -282 6218 -248
rect 6252 -282 6268 -248
rect 6368 -282 6418 -248
rect 6452 -282 6468 -248
rect 6568 -282 6618 -248
rect 6652 -282 6668 -248
rect 6768 -282 6818 -248
rect 6852 -282 6868 -248
rect 6968 -282 7018 -248
rect 7052 -282 7068 -248
rect 7168 -282 7218 -248
rect 7252 -282 7268 -248
rect 7368 -282 7418 -248
rect 7452 -282 7468 -248
rect 7568 -282 7618 -248
rect 7652 -282 7668 -248
rect 7768 -282 7818 -248
rect 7852 -282 7868 -248
rect 7968 -282 8018 -248
rect 8052 -282 8068 -248
rect 8168 -282 8218 -248
rect 8252 -282 8268 -248
rect 8368 -282 8418 -248
rect 8452 -282 8468 -248
rect 8568 -282 8618 -248
rect 8652 -282 8668 -248
rect 8768 -282 8818 -248
rect 8852 -282 8868 -248
rect 8968 -282 9018 -248
rect 9052 -282 9068 -248
rect 9168 -282 9218 -248
rect 9252 -282 9268 -248
rect 9368 -282 9418 -248
rect 9452 -282 9468 -248
rect 9568 -282 9618 -248
rect 9652 -282 9668 -248
rect 9768 -282 9818 -248
rect 9852 -282 9868 -248
rect 9968 -282 10018 -248
rect 10052 -282 10068 -248
rect 10168 -282 10218 -248
rect 10252 -282 10268 -248
rect 10368 -282 10418 -248
rect 10452 -282 10468 -248
rect 10568 -282 10618 -248
rect 10652 -282 10668 -248
rect 10768 -282 10818 -248
rect 10852 -282 10868 -248
rect 10968 -282 11018 -248
rect 11052 -282 11068 -248
rect 11168 -282 11218 -248
rect 11252 -282 11268 -248
rect 11368 -282 11418 -248
rect 11452 -282 11468 -248
rect 11568 -282 11618 -248
rect 11652 -282 11668 -248
rect 11768 -282 11818 -248
rect 11852 -282 11868 -248
rect 11968 -282 12018 -248
rect 12052 -282 12068 -248
rect 12168 -282 12218 -248
rect 12252 -282 12268 -248
rect 12368 -282 12418 -248
rect 12452 -282 12468 -248
rect 12568 -282 12618 -248
rect 12652 -282 12668 -248
rect -82 -363 -48 -322
rect -82 -431 -48 -397
rect -82 -561 -48 -469
rect 18 -363 52 -322
rect 18 -431 52 -397
rect 18 -506 52 -469
rect 118 -363 152 -322
rect 118 -431 152 -397
rect -125 -595 -118 -561
rect -84 -595 -82 -561
rect -48 -595 -46 -561
rect -12 -595 -5 -561
rect 44 -577 78 -561
rect 44 -630 78 -611
rect -30 -683 4 -667
rect -30 -803 4 -717
rect 118 -683 152 -469
rect 218 -363 252 -322
rect 218 -431 252 -397
rect 218 -506 252 -469
rect 318 -363 352 -322
rect 318 -431 352 -397
rect 318 -561 352 -469
rect 418 -363 452 -322
rect 418 -431 452 -397
rect 418 -506 452 -469
rect 518 -363 552 -322
rect 518 -431 552 -397
rect 192 -577 226 -561
rect 275 -595 282 -561
rect 316 -595 318 -561
rect 352 -595 354 -561
rect 388 -595 395 -561
rect 444 -577 478 -561
rect 192 -630 226 -611
rect 444 -630 478 -611
rect 118 -733 152 -717
rect 266 -683 300 -667
rect 266 -803 300 -717
rect -30 -837 24 -803
rect 246 -837 300 -803
rect 370 -683 404 -667
rect 370 -803 404 -717
rect 518 -683 552 -469
rect 618 -363 652 -322
rect 618 -431 652 -397
rect 618 -506 652 -469
rect 718 -363 752 -322
rect 718 -431 752 -397
rect 718 -561 752 -469
rect 818 -363 852 -322
rect 818 -431 852 -397
rect 818 -506 852 -469
rect 918 -363 952 -322
rect 918 -431 952 -397
rect 592 -577 626 -561
rect 675 -595 682 -561
rect 716 -595 718 -561
rect 752 -595 754 -561
rect 788 -595 795 -561
rect 844 -577 878 -561
rect 592 -630 626 -611
rect 844 -630 878 -611
rect 518 -733 552 -717
rect 666 -683 700 -667
rect 666 -803 700 -717
rect 370 -837 424 -803
rect 646 -837 700 -803
rect 770 -683 804 -667
rect 770 -803 804 -717
rect 918 -683 952 -469
rect 1018 -363 1052 -322
rect 1018 -431 1052 -397
rect 1018 -506 1052 -469
rect 1118 -363 1152 -322
rect 1118 -431 1152 -397
rect 1118 -561 1152 -469
rect 1218 -363 1252 -322
rect 1218 -431 1252 -397
rect 1218 -506 1252 -469
rect 1318 -363 1352 -322
rect 1318 -431 1352 -397
rect 992 -577 1026 -561
rect 1075 -595 1082 -561
rect 1116 -595 1118 -561
rect 1152 -595 1154 -561
rect 1188 -595 1195 -561
rect 1244 -577 1278 -561
rect 992 -630 1026 -611
rect 1244 -630 1278 -611
rect 918 -733 952 -717
rect 1066 -683 1100 -667
rect 1066 -803 1100 -717
rect 770 -837 824 -803
rect 1046 -837 1100 -803
rect 1170 -683 1204 -667
rect 1170 -803 1204 -717
rect 1318 -683 1352 -469
rect 1418 -363 1452 -322
rect 1418 -431 1452 -397
rect 1418 -506 1452 -469
rect 1518 -363 1552 -322
rect 1518 -431 1552 -397
rect 1518 -561 1552 -469
rect 1618 -363 1652 -322
rect 1618 -431 1652 -397
rect 1618 -506 1652 -469
rect 1718 -363 1752 -322
rect 1718 -431 1752 -397
rect 1392 -577 1426 -561
rect 1475 -595 1482 -561
rect 1516 -595 1518 -561
rect 1552 -595 1554 -561
rect 1588 -595 1595 -561
rect 1644 -577 1678 -561
rect 1392 -630 1426 -611
rect 1644 -630 1678 -611
rect 1318 -733 1352 -717
rect 1466 -683 1500 -667
rect 1466 -803 1500 -717
rect 1170 -837 1224 -803
rect 1446 -837 1500 -803
rect 1570 -683 1604 -667
rect 1570 -803 1604 -717
rect 1718 -683 1752 -469
rect 1818 -363 1852 -322
rect 1818 -431 1852 -397
rect 1818 -506 1852 -469
rect 1918 -363 1952 -322
rect 1918 -431 1952 -397
rect 1918 -561 1952 -469
rect 2018 -363 2052 -322
rect 2018 -431 2052 -397
rect 2018 -506 2052 -469
rect 2118 -363 2152 -322
rect 2118 -431 2152 -397
rect 1792 -577 1826 -561
rect 1875 -595 1882 -561
rect 1916 -595 1918 -561
rect 1952 -595 1954 -561
rect 1988 -595 1995 -561
rect 2044 -577 2078 -561
rect 1792 -630 1826 -611
rect 2044 -630 2078 -611
rect 1718 -733 1752 -717
rect 1866 -683 1900 -667
rect 1866 -803 1900 -717
rect 1570 -837 1624 -803
rect 1846 -837 1900 -803
rect 1970 -683 2004 -667
rect 1970 -803 2004 -717
rect 2118 -683 2152 -469
rect 2218 -363 2252 -322
rect 2218 -431 2252 -397
rect 2218 -506 2252 -469
rect 2318 -363 2352 -322
rect 2318 -431 2352 -397
rect 2318 -561 2352 -469
rect 2418 -363 2452 -322
rect 2418 -431 2452 -397
rect 2418 -506 2452 -469
rect 2518 -363 2552 -322
rect 2518 -431 2552 -397
rect 2192 -577 2226 -561
rect 2275 -595 2282 -561
rect 2316 -595 2318 -561
rect 2352 -595 2354 -561
rect 2388 -595 2395 -561
rect 2444 -577 2478 -561
rect 2192 -630 2226 -611
rect 2444 -630 2478 -611
rect 2118 -733 2152 -717
rect 2266 -683 2300 -667
rect 2266 -803 2300 -717
rect 1970 -837 2024 -803
rect 2246 -837 2300 -803
rect 2370 -683 2404 -667
rect 2370 -803 2404 -717
rect 2518 -683 2552 -469
rect 2618 -363 2652 -322
rect 2618 -431 2652 -397
rect 2618 -506 2652 -469
rect 2718 -363 2752 -322
rect 2718 -431 2752 -397
rect 2718 -561 2752 -469
rect 2818 -363 2852 -322
rect 2818 -431 2852 -397
rect 2818 -506 2852 -469
rect 2918 -363 2952 -322
rect 2918 -431 2952 -397
rect 2592 -577 2626 -561
rect 2675 -595 2682 -561
rect 2716 -595 2718 -561
rect 2752 -595 2754 -561
rect 2788 -595 2795 -561
rect 2844 -577 2878 -561
rect 2592 -630 2626 -611
rect 2844 -630 2878 -611
rect 2518 -733 2552 -717
rect 2666 -683 2700 -667
rect 2666 -803 2700 -717
rect 2370 -837 2424 -803
rect 2646 -837 2700 -803
rect 2770 -683 2804 -667
rect 2770 -803 2804 -717
rect 2918 -683 2952 -469
rect 3018 -363 3052 -322
rect 3018 -431 3052 -397
rect 3018 -506 3052 -469
rect 3118 -363 3152 -322
rect 3118 -431 3152 -397
rect 3118 -561 3152 -469
rect 3218 -363 3252 -322
rect 3218 -431 3252 -397
rect 3218 -506 3252 -469
rect 3318 -363 3352 -322
rect 3318 -431 3352 -397
rect 2992 -577 3026 -561
rect 3075 -595 3082 -561
rect 3116 -595 3118 -561
rect 3152 -595 3154 -561
rect 3188 -595 3195 -561
rect 3244 -577 3278 -561
rect 2992 -630 3026 -611
rect 3244 -630 3278 -611
rect 2918 -733 2952 -717
rect 3066 -683 3100 -667
rect 3066 -803 3100 -717
rect 2770 -837 2824 -803
rect 3046 -837 3100 -803
rect 3170 -683 3204 -667
rect 3170 -803 3204 -717
rect 3318 -683 3352 -469
rect 3418 -363 3452 -322
rect 3418 -431 3452 -397
rect 3418 -506 3452 -469
rect 3518 -363 3552 -322
rect 3518 -431 3552 -397
rect 3518 -561 3552 -469
rect 3618 -363 3652 -322
rect 3618 -431 3652 -397
rect 3618 -506 3652 -469
rect 3718 -363 3752 -322
rect 3718 -431 3752 -397
rect 3392 -577 3426 -561
rect 3475 -595 3482 -561
rect 3516 -595 3518 -561
rect 3552 -595 3554 -561
rect 3588 -595 3595 -561
rect 3644 -577 3678 -561
rect 3392 -630 3426 -611
rect 3644 -630 3678 -611
rect 3318 -733 3352 -717
rect 3466 -683 3500 -667
rect 3466 -803 3500 -717
rect 3170 -837 3224 -803
rect 3446 -837 3500 -803
rect 3570 -683 3604 -667
rect 3570 -803 3604 -717
rect 3718 -683 3752 -469
rect 3818 -363 3852 -322
rect 3818 -431 3852 -397
rect 3818 -506 3852 -469
rect 3918 -363 3952 -322
rect 3918 -431 3952 -397
rect 3918 -561 3952 -469
rect 4018 -363 4052 -322
rect 4018 -431 4052 -397
rect 4018 -506 4052 -469
rect 4118 -363 4152 -322
rect 4118 -431 4152 -397
rect 3792 -577 3826 -561
rect 3875 -595 3882 -561
rect 3916 -595 3918 -561
rect 3952 -595 3954 -561
rect 3988 -595 3995 -561
rect 4044 -577 4078 -561
rect 3792 -630 3826 -611
rect 4044 -630 4078 -611
rect 3718 -733 3752 -717
rect 3866 -683 3900 -667
rect 3866 -803 3900 -717
rect 3570 -837 3624 -803
rect 3846 -837 3900 -803
rect 3970 -683 4004 -667
rect 3970 -803 4004 -717
rect 4118 -683 4152 -469
rect 4218 -363 4252 -322
rect 4218 -431 4252 -397
rect 4218 -506 4252 -469
rect 4318 -363 4352 -322
rect 4318 -431 4352 -397
rect 4318 -561 4352 -469
rect 4418 -363 4452 -322
rect 4418 -431 4452 -397
rect 4418 -506 4452 -469
rect 4518 -363 4552 -322
rect 4518 -431 4552 -397
rect 4192 -577 4226 -561
rect 4275 -595 4282 -561
rect 4316 -595 4318 -561
rect 4352 -595 4354 -561
rect 4388 -595 4395 -561
rect 4444 -577 4478 -561
rect 4192 -630 4226 -611
rect 4444 -630 4478 -611
rect 4118 -733 4152 -717
rect 4266 -683 4300 -667
rect 4266 -803 4300 -717
rect 3970 -837 4024 -803
rect 4246 -837 4300 -803
rect 4370 -683 4404 -667
rect 4370 -803 4404 -717
rect 4518 -683 4552 -469
rect 4618 -363 4652 -322
rect 4618 -431 4652 -397
rect 4618 -506 4652 -469
rect 4718 -363 4752 -322
rect 4718 -431 4752 -397
rect 4718 -561 4752 -469
rect 4818 -363 4852 -322
rect 4818 -431 4852 -397
rect 4818 -506 4852 -469
rect 4918 -363 4952 -322
rect 4918 -431 4952 -397
rect 4592 -577 4626 -561
rect 4675 -595 4682 -561
rect 4716 -595 4718 -561
rect 4752 -595 4754 -561
rect 4788 -595 4795 -561
rect 4844 -577 4878 -561
rect 4592 -630 4626 -611
rect 4844 -630 4878 -611
rect 4518 -733 4552 -717
rect 4666 -683 4700 -667
rect 4666 -803 4700 -717
rect 4370 -837 4424 -803
rect 4646 -837 4700 -803
rect 4770 -683 4804 -667
rect 4770 -803 4804 -717
rect 4918 -683 4952 -469
rect 5018 -363 5052 -322
rect 5018 -431 5052 -397
rect 5018 -506 5052 -469
rect 5118 -363 5152 -322
rect 5118 -431 5152 -397
rect 5118 -561 5152 -469
rect 5218 -363 5252 -322
rect 5218 -431 5252 -397
rect 5218 -506 5252 -469
rect 5318 -363 5352 -322
rect 5318 -431 5352 -397
rect 4992 -577 5026 -561
rect 5075 -595 5082 -561
rect 5116 -595 5118 -561
rect 5152 -595 5154 -561
rect 5188 -595 5195 -561
rect 5244 -577 5278 -561
rect 4992 -630 5026 -611
rect 5244 -630 5278 -611
rect 4918 -733 4952 -717
rect 5066 -683 5100 -667
rect 5066 -803 5100 -717
rect 4770 -837 4824 -803
rect 5046 -837 5100 -803
rect 5170 -683 5204 -667
rect 5170 -803 5204 -717
rect 5318 -683 5352 -469
rect 5418 -363 5452 -322
rect 5418 -431 5452 -397
rect 5418 -506 5452 -469
rect 5518 -363 5552 -322
rect 5518 -431 5552 -397
rect 5518 -561 5552 -469
rect 5618 -363 5652 -322
rect 5618 -431 5652 -397
rect 5618 -506 5652 -469
rect 5718 -363 5752 -322
rect 5718 -431 5752 -397
rect 5392 -577 5426 -561
rect 5475 -595 5482 -561
rect 5516 -595 5518 -561
rect 5552 -595 5554 -561
rect 5588 -595 5595 -561
rect 5644 -577 5678 -561
rect 5392 -630 5426 -611
rect 5644 -630 5678 -611
rect 5318 -733 5352 -717
rect 5466 -683 5500 -667
rect 5466 -803 5500 -717
rect 5170 -837 5224 -803
rect 5446 -837 5500 -803
rect 5570 -683 5604 -667
rect 5570 -803 5604 -717
rect 5718 -683 5752 -469
rect 5818 -363 5852 -322
rect 5818 -431 5852 -397
rect 5818 -506 5852 -469
rect 5918 -363 5952 -322
rect 5918 -431 5952 -397
rect 5918 -561 5952 -469
rect 6018 -363 6052 -322
rect 6018 -431 6052 -397
rect 6018 -506 6052 -469
rect 6118 -363 6152 -322
rect 6118 -431 6152 -397
rect 5792 -577 5826 -561
rect 5875 -595 5882 -561
rect 5916 -595 5918 -561
rect 5952 -595 5954 -561
rect 5988 -595 5995 -561
rect 6044 -577 6078 -561
rect 5792 -630 5826 -611
rect 6044 -630 6078 -611
rect 5718 -733 5752 -717
rect 5866 -683 5900 -667
rect 5866 -803 5900 -717
rect 5570 -837 5624 -803
rect 5846 -837 5900 -803
rect 5970 -683 6004 -667
rect 5970 -803 6004 -717
rect 6118 -683 6152 -469
rect 6218 -363 6252 -322
rect 6218 -431 6252 -397
rect 6218 -506 6252 -469
rect 6318 -363 6352 -322
rect 6318 -431 6352 -397
rect 6318 -561 6352 -469
rect 6418 -363 6452 -322
rect 6418 -431 6452 -397
rect 6418 -506 6452 -469
rect 6518 -363 6552 -322
rect 6518 -431 6552 -397
rect 6192 -577 6226 -561
rect 6275 -595 6282 -561
rect 6316 -595 6318 -561
rect 6352 -595 6354 -561
rect 6388 -595 6395 -561
rect 6444 -577 6478 -561
rect 6192 -630 6226 -611
rect 6444 -630 6478 -611
rect 6118 -733 6152 -717
rect 6266 -683 6300 -667
rect 6266 -803 6300 -717
rect 5970 -837 6024 -803
rect 6246 -837 6300 -803
rect 6370 -683 6404 -667
rect 6370 -803 6404 -717
rect 6518 -683 6552 -469
rect 6618 -363 6652 -322
rect 6618 -431 6652 -397
rect 6618 -506 6652 -469
rect 6718 -363 6752 -322
rect 6718 -431 6752 -397
rect 6718 -561 6752 -469
rect 6818 -363 6852 -322
rect 6818 -431 6852 -397
rect 6818 -506 6852 -469
rect 6918 -363 6952 -322
rect 6918 -431 6952 -397
rect 6592 -577 6626 -561
rect 6675 -595 6682 -561
rect 6716 -595 6718 -561
rect 6752 -595 6754 -561
rect 6788 -595 6795 -561
rect 6844 -577 6878 -561
rect 6592 -630 6626 -611
rect 6844 -630 6878 -611
rect 6518 -733 6552 -717
rect 6666 -683 6700 -667
rect 6666 -803 6700 -717
rect 6370 -837 6424 -803
rect 6646 -837 6700 -803
rect 6770 -683 6804 -667
rect 6770 -803 6804 -717
rect 6918 -683 6952 -469
rect 7018 -363 7052 -322
rect 7018 -431 7052 -397
rect 7018 -506 7052 -469
rect 7118 -363 7152 -322
rect 7118 -431 7152 -397
rect 7118 -561 7152 -469
rect 7218 -363 7252 -322
rect 7218 -431 7252 -397
rect 7218 -506 7252 -469
rect 7318 -363 7352 -322
rect 7318 -431 7352 -397
rect 6992 -577 7026 -561
rect 7075 -595 7082 -561
rect 7116 -595 7118 -561
rect 7152 -595 7154 -561
rect 7188 -595 7195 -561
rect 7244 -577 7278 -561
rect 6992 -630 7026 -611
rect 7244 -630 7278 -611
rect 6918 -733 6952 -717
rect 7066 -683 7100 -667
rect 7066 -803 7100 -717
rect 6770 -837 6824 -803
rect 7046 -837 7100 -803
rect 7170 -683 7204 -667
rect 7170 -803 7204 -717
rect 7318 -683 7352 -469
rect 7418 -363 7452 -322
rect 7418 -431 7452 -397
rect 7418 -506 7452 -469
rect 7518 -363 7552 -322
rect 7518 -431 7552 -397
rect 7518 -561 7552 -469
rect 7618 -363 7652 -322
rect 7618 -431 7652 -397
rect 7618 -506 7652 -469
rect 7718 -363 7752 -322
rect 7718 -431 7752 -397
rect 7392 -577 7426 -561
rect 7475 -595 7482 -561
rect 7516 -595 7518 -561
rect 7552 -595 7554 -561
rect 7588 -595 7595 -561
rect 7644 -577 7678 -561
rect 7392 -630 7426 -611
rect 7644 -630 7678 -611
rect 7318 -733 7352 -717
rect 7466 -683 7500 -667
rect 7466 -803 7500 -717
rect 7170 -837 7224 -803
rect 7446 -837 7500 -803
rect 7570 -683 7604 -667
rect 7570 -803 7604 -717
rect 7718 -683 7752 -469
rect 7818 -363 7852 -322
rect 7818 -431 7852 -397
rect 7818 -506 7852 -469
rect 7918 -363 7952 -322
rect 7918 -431 7952 -397
rect 7918 -561 7952 -469
rect 8018 -363 8052 -322
rect 8018 -431 8052 -397
rect 8018 -506 8052 -469
rect 8118 -363 8152 -322
rect 8118 -431 8152 -397
rect 7792 -577 7826 -561
rect 7875 -595 7882 -561
rect 7916 -595 7918 -561
rect 7952 -595 7954 -561
rect 7988 -595 7995 -561
rect 8044 -577 8078 -561
rect 7792 -630 7826 -611
rect 8044 -630 8078 -611
rect 7718 -733 7752 -717
rect 7866 -683 7900 -667
rect 7866 -803 7900 -717
rect 7570 -837 7624 -803
rect 7846 -837 7900 -803
rect 7970 -683 8004 -667
rect 7970 -803 8004 -717
rect 8118 -683 8152 -469
rect 8218 -363 8252 -322
rect 8218 -431 8252 -397
rect 8218 -506 8252 -469
rect 8318 -363 8352 -322
rect 8318 -431 8352 -397
rect 8318 -561 8352 -469
rect 8418 -363 8452 -322
rect 8418 -431 8452 -397
rect 8418 -506 8452 -469
rect 8518 -363 8552 -322
rect 8518 -431 8552 -397
rect 8192 -577 8226 -561
rect 8275 -595 8282 -561
rect 8316 -595 8318 -561
rect 8352 -595 8354 -561
rect 8388 -595 8395 -561
rect 8444 -577 8478 -561
rect 8192 -630 8226 -611
rect 8444 -630 8478 -611
rect 8118 -733 8152 -717
rect 8266 -683 8300 -667
rect 8266 -803 8300 -717
rect 7970 -837 8024 -803
rect 8246 -837 8300 -803
rect 8370 -683 8404 -667
rect 8370 -803 8404 -717
rect 8518 -683 8552 -469
rect 8618 -363 8652 -322
rect 8618 -431 8652 -397
rect 8618 -506 8652 -469
rect 8718 -363 8752 -322
rect 8718 -431 8752 -397
rect 8718 -561 8752 -469
rect 8818 -363 8852 -322
rect 8818 -431 8852 -397
rect 8818 -506 8852 -469
rect 8918 -363 8952 -322
rect 8918 -431 8952 -397
rect 8592 -577 8626 -561
rect 8675 -595 8682 -561
rect 8716 -595 8718 -561
rect 8752 -595 8754 -561
rect 8788 -595 8795 -561
rect 8844 -577 8878 -561
rect 8592 -630 8626 -611
rect 8844 -630 8878 -611
rect 8518 -733 8552 -717
rect 8666 -683 8700 -667
rect 8666 -803 8700 -717
rect 8370 -837 8424 -803
rect 8646 -837 8700 -803
rect 8770 -683 8804 -667
rect 8770 -803 8804 -717
rect 8918 -683 8952 -469
rect 9018 -363 9052 -322
rect 9018 -431 9052 -397
rect 9018 -506 9052 -469
rect 9118 -363 9152 -322
rect 9118 -431 9152 -397
rect 9118 -561 9152 -469
rect 9218 -363 9252 -322
rect 9218 -431 9252 -397
rect 9218 -506 9252 -469
rect 9318 -363 9352 -322
rect 9318 -431 9352 -397
rect 8992 -577 9026 -561
rect 9075 -595 9082 -561
rect 9116 -595 9118 -561
rect 9152 -595 9154 -561
rect 9188 -595 9195 -561
rect 9244 -577 9278 -561
rect 8992 -630 9026 -611
rect 9244 -630 9278 -611
rect 8918 -733 8952 -717
rect 9066 -683 9100 -667
rect 9066 -803 9100 -717
rect 8770 -837 8824 -803
rect 9046 -837 9100 -803
rect 9170 -683 9204 -667
rect 9170 -803 9204 -717
rect 9318 -683 9352 -469
rect 9418 -363 9452 -322
rect 9418 -431 9452 -397
rect 9418 -506 9452 -469
rect 9518 -363 9552 -322
rect 9518 -431 9552 -397
rect 9518 -561 9552 -469
rect 9618 -363 9652 -322
rect 9618 -431 9652 -397
rect 9618 -506 9652 -469
rect 9718 -363 9752 -322
rect 9718 -431 9752 -397
rect 9392 -577 9426 -561
rect 9475 -595 9482 -561
rect 9516 -595 9518 -561
rect 9552 -595 9554 -561
rect 9588 -595 9595 -561
rect 9644 -577 9678 -561
rect 9392 -630 9426 -611
rect 9644 -630 9678 -611
rect 9318 -733 9352 -717
rect 9466 -683 9500 -667
rect 9466 -803 9500 -717
rect 9170 -837 9224 -803
rect 9446 -837 9500 -803
rect 9570 -683 9604 -667
rect 9570 -803 9604 -717
rect 9718 -683 9752 -469
rect 9818 -363 9852 -322
rect 9818 -431 9852 -397
rect 9818 -506 9852 -469
rect 9918 -363 9952 -322
rect 9918 -431 9952 -397
rect 9918 -561 9952 -469
rect 10018 -363 10052 -322
rect 10018 -431 10052 -397
rect 10018 -506 10052 -469
rect 10118 -363 10152 -322
rect 10118 -431 10152 -397
rect 9792 -577 9826 -561
rect 9875 -595 9882 -561
rect 9916 -595 9918 -561
rect 9952 -595 9954 -561
rect 9988 -595 9995 -561
rect 10044 -577 10078 -561
rect 9792 -630 9826 -611
rect 10044 -630 10078 -611
rect 9718 -733 9752 -717
rect 9866 -683 9900 -667
rect 9866 -803 9900 -717
rect 9570 -837 9624 -803
rect 9846 -837 9900 -803
rect 9970 -683 10004 -667
rect 9970 -803 10004 -717
rect 10118 -683 10152 -469
rect 10218 -363 10252 -322
rect 10218 -431 10252 -397
rect 10218 -506 10252 -469
rect 10318 -363 10352 -322
rect 10318 -431 10352 -397
rect 10318 -561 10352 -469
rect 10418 -363 10452 -322
rect 10418 -431 10452 -397
rect 10418 -506 10452 -469
rect 10518 -363 10552 -322
rect 10518 -431 10552 -397
rect 10192 -577 10226 -561
rect 10275 -595 10282 -561
rect 10316 -595 10318 -561
rect 10352 -595 10354 -561
rect 10388 -595 10395 -561
rect 10444 -577 10478 -561
rect 10192 -630 10226 -611
rect 10444 -630 10478 -611
rect 10118 -733 10152 -717
rect 10266 -683 10300 -667
rect 10266 -803 10300 -717
rect 9970 -837 10024 -803
rect 10246 -837 10300 -803
rect 10370 -683 10404 -667
rect 10370 -803 10404 -717
rect 10518 -683 10552 -469
rect 10618 -363 10652 -322
rect 10618 -431 10652 -397
rect 10618 -506 10652 -469
rect 10718 -363 10752 -322
rect 10718 -431 10752 -397
rect 10718 -561 10752 -469
rect 10818 -363 10852 -322
rect 10818 -431 10852 -397
rect 10818 -506 10852 -469
rect 10918 -363 10952 -322
rect 10918 -431 10952 -397
rect 10592 -577 10626 -561
rect 10675 -595 10682 -561
rect 10716 -595 10718 -561
rect 10752 -595 10754 -561
rect 10788 -595 10795 -561
rect 10844 -577 10878 -561
rect 10592 -630 10626 -611
rect 10844 -630 10878 -611
rect 10518 -733 10552 -717
rect 10666 -683 10700 -667
rect 10666 -803 10700 -717
rect 10370 -837 10424 -803
rect 10646 -837 10700 -803
rect 10770 -683 10804 -667
rect 10770 -803 10804 -717
rect 10918 -683 10952 -469
rect 11018 -363 11052 -322
rect 11018 -431 11052 -397
rect 11018 -506 11052 -469
rect 11118 -363 11152 -322
rect 11118 -431 11152 -397
rect 11118 -561 11152 -469
rect 11218 -363 11252 -322
rect 11218 -431 11252 -397
rect 11218 -506 11252 -469
rect 11318 -363 11352 -322
rect 11318 -431 11352 -397
rect 10992 -577 11026 -561
rect 11075 -595 11082 -561
rect 11116 -595 11118 -561
rect 11152 -595 11154 -561
rect 11188 -595 11195 -561
rect 11244 -577 11278 -561
rect 10992 -630 11026 -611
rect 11244 -630 11278 -611
rect 10918 -733 10952 -717
rect 11066 -683 11100 -667
rect 11066 -803 11100 -717
rect 10770 -837 10824 -803
rect 11046 -837 11100 -803
rect 11170 -683 11204 -667
rect 11170 -803 11204 -717
rect 11318 -683 11352 -469
rect 11418 -363 11452 -322
rect 11418 -431 11452 -397
rect 11418 -506 11452 -469
rect 11518 -363 11552 -322
rect 11518 -431 11552 -397
rect 11518 -561 11552 -469
rect 11618 -363 11652 -322
rect 11618 -431 11652 -397
rect 11618 -506 11652 -469
rect 11718 -363 11752 -322
rect 11718 -431 11752 -397
rect 11392 -577 11426 -561
rect 11475 -595 11482 -561
rect 11516 -595 11518 -561
rect 11552 -595 11554 -561
rect 11588 -595 11595 -561
rect 11644 -577 11678 -561
rect 11392 -630 11426 -611
rect 11644 -630 11678 -611
rect 11318 -733 11352 -717
rect 11466 -683 11500 -667
rect 11466 -803 11500 -717
rect 11170 -837 11224 -803
rect 11446 -837 11500 -803
rect 11570 -683 11604 -667
rect 11570 -803 11604 -717
rect 11718 -683 11752 -469
rect 11818 -363 11852 -322
rect 11818 -431 11852 -397
rect 11818 -506 11852 -469
rect 11918 -363 11952 -322
rect 11918 -431 11952 -397
rect 11918 -561 11952 -469
rect 12018 -363 12052 -322
rect 12018 -431 12052 -397
rect 12018 -506 12052 -469
rect 12118 -363 12152 -322
rect 12118 -431 12152 -397
rect 11792 -577 11826 -561
rect 11875 -595 11882 -561
rect 11916 -595 11918 -561
rect 11952 -595 11954 -561
rect 11988 -595 11995 -561
rect 12044 -577 12078 -561
rect 11792 -630 11826 -611
rect 12044 -630 12078 -611
rect 11718 -733 11752 -717
rect 11866 -683 11900 -667
rect 11866 -803 11900 -717
rect 11570 -837 11624 -803
rect 11846 -837 11900 -803
rect 11970 -683 12004 -667
rect 11970 -803 12004 -717
rect 12118 -683 12152 -469
rect 12218 -363 12252 -322
rect 12218 -431 12252 -397
rect 12218 -506 12252 -469
rect 12318 -363 12352 -322
rect 12318 -431 12352 -397
rect 12318 -561 12352 -469
rect 12418 -363 12452 -322
rect 12418 -431 12452 -397
rect 12418 -506 12452 -469
rect 12518 -363 12552 -322
rect 12518 -431 12552 -397
rect 12192 -577 12226 -561
rect 12275 -595 12282 -561
rect 12316 -595 12318 -561
rect 12352 -595 12354 -561
rect 12388 -595 12395 -561
rect 12444 -577 12478 -561
rect 12192 -630 12226 -611
rect 12444 -630 12478 -611
rect 12118 -733 12152 -717
rect 12266 -683 12300 -667
rect 12266 -803 12300 -717
rect 11970 -837 12024 -803
rect 12246 -837 12300 -803
rect 12370 -683 12404 -667
rect 12370 -803 12404 -717
rect 12518 -683 12552 -469
rect 12618 -363 12652 -322
rect 12618 -431 12652 -397
rect 12618 -506 12652 -469
rect 12718 -363 12752 -322
rect 14532 -342 14560 -308
rect 14596 -342 14630 -308
rect 14666 -342 14694 -308
rect 14734 -309 14768 -292
rect 12718 -431 12752 -397
rect 14808 -342 14841 -308
rect 14881 -342 14913 -308
rect 14949 -342 14983 -308
rect 15019 -342 15051 -308
rect 15091 -342 15124 -308
rect 15218 -342 15251 -308
rect 15291 -342 15323 -308
rect 15359 -342 15393 -308
rect 15429 -342 15461 -308
rect 15501 -342 15534 -308
rect 15574 -309 15608 -292
rect 14734 -408 14768 -343
rect 15648 -342 15676 -308
rect 15712 -342 15746 -308
rect 15782 -342 15810 -308
rect 15574 -408 15608 -343
rect 14532 -442 14558 -408
rect 14596 -442 14630 -408
rect 14664 -442 14694 -408
rect 14808 -442 14842 -408
rect 14881 -442 14914 -408
rect 14949 -442 14983 -408
rect 15020 -442 15051 -408
rect 15092 -442 15124 -408
rect 15218 -442 15249 -408
rect 15291 -442 15321 -408
rect 15359 -442 15393 -408
rect 15427 -442 15461 -408
rect 15499 -442 15534 -408
rect 15648 -442 15677 -408
rect 15712 -442 15746 -408
rect 15783 -442 15810 -408
rect 12718 -561 12752 -469
rect 14532 -542 14560 -508
rect 14596 -542 14630 -508
rect 14666 -542 14694 -508
rect 14734 -509 14768 -492
rect 14808 -542 14841 -508
rect 14881 -542 14913 -508
rect 14949 -542 14983 -508
rect 15019 -542 15051 -508
rect 15091 -542 15124 -508
rect 15218 -542 15251 -508
rect 15291 -542 15323 -508
rect 15359 -542 15393 -508
rect 15429 -542 15461 -508
rect 15501 -542 15534 -508
rect 15574 -509 15608 -492
rect 12592 -577 12626 -561
rect 12675 -595 12682 -561
rect 12716 -595 12718 -561
rect 12752 -595 12754 -561
rect 12788 -595 12795 -561
rect 14734 -608 14768 -543
rect 15648 -542 15676 -508
rect 15712 -542 15746 -508
rect 15782 -542 15810 -508
rect 15574 -608 15608 -543
rect 12592 -630 12626 -611
rect 14532 -642 14558 -608
rect 14596 -642 14630 -608
rect 14664 -642 14694 -608
rect 14808 -642 14842 -608
rect 14881 -642 14914 -608
rect 14949 -642 14983 -608
rect 15020 -642 15051 -608
rect 15092 -642 15124 -608
rect 15218 -642 15249 -608
rect 15291 -642 15321 -608
rect 15359 -642 15393 -608
rect 15427 -642 15461 -608
rect 15499 -642 15534 -608
rect 15648 -642 15677 -608
rect 15712 -642 15746 -608
rect 15783 -642 15810 -608
rect 12518 -733 12552 -717
rect 12666 -683 12700 -667
rect 12666 -803 12700 -717
rect 14532 -742 14560 -708
rect 14596 -742 14630 -708
rect 14666 -742 14694 -708
rect 14734 -709 14768 -692
rect 12370 -837 12424 -803
rect 12646 -837 12700 -803
rect 14808 -742 14841 -708
rect 14881 -742 14913 -708
rect 14949 -742 14983 -708
rect 15019 -742 15051 -708
rect 15091 -742 15124 -708
rect 15218 -742 15251 -708
rect 15291 -742 15323 -708
rect 15359 -742 15393 -708
rect 15429 -742 15461 -708
rect 15501 -742 15534 -708
rect 15574 -709 15608 -692
rect 14734 -808 14768 -743
rect 15648 -742 15676 -708
rect 15712 -742 15746 -708
rect 15782 -742 15810 -708
rect 15574 -808 15608 -743
rect -10 -871 -4 -837
rect 30 -858 68 -837
rect -10 -892 -2 -871
rect 32 -892 66 -858
rect 102 -871 108 -837
rect 100 -892 108 -871
rect -82 -908 -48 -892
rect -82 -958 -48 -942
rect -10 -958 108 -892
rect 162 -871 168 -837
rect 202 -858 240 -837
rect 162 -892 170 -871
rect 204 -892 238 -858
rect 274 -871 280 -837
rect 272 -892 280 -871
rect 162 -908 280 -892
rect 390 -871 396 -837
rect 430 -858 468 -837
rect 390 -892 398 -871
rect 432 -892 466 -858
rect 502 -871 508 -837
rect 500 -892 508 -871
rect -10 -992 -2 -958
rect 32 -992 66 -958
rect 100 -992 108 -958
rect -82 -1008 -48 -992
rect -10 -1008 108 -992
rect 162 -958 280 -942
rect 162 -992 170 -958
rect 204 -992 238 -958
rect 272 -992 280 -958
rect -82 -1058 -48 -1042
rect -10 -1058 108 -1042
rect -10 -1092 -2 -1058
rect 32 -1092 66 -1058
rect 100 -1092 108 -1058
rect -82 -1108 -48 -1092
rect -82 -1158 -48 -1142
rect -10 -1158 108 -1092
rect -10 -1192 -2 -1158
rect 32 -1192 66 -1158
rect 100 -1192 108 -1158
rect -82 -1208 -48 -1192
rect -10 -1208 108 -1192
rect 162 -1058 280 -992
rect 390 -958 508 -892
rect 562 -871 568 -837
rect 602 -858 640 -837
rect 562 -892 570 -871
rect 604 -892 638 -858
rect 674 -871 680 -837
rect 672 -892 680 -871
rect 790 -871 796 -837
rect 830 -858 868 -837
rect 790 -892 798 -871
rect 832 -892 866 -858
rect 902 -871 908 -837
rect 900 -892 908 -871
rect 562 -908 680 -892
rect 718 -908 752 -892
rect 390 -992 398 -958
rect 432 -992 466 -958
rect 500 -992 508 -958
rect 390 -1008 508 -992
rect 562 -958 680 -942
rect 718 -958 752 -942
rect 790 -958 908 -892
rect 962 -871 968 -837
rect 1002 -858 1040 -837
rect 962 -892 970 -871
rect 1004 -892 1038 -858
rect 1074 -871 1080 -837
rect 1072 -892 1080 -871
rect 962 -908 1080 -892
rect 1190 -871 1196 -837
rect 1230 -858 1268 -837
rect 1190 -892 1198 -871
rect 1232 -892 1266 -858
rect 1302 -871 1308 -837
rect 1300 -892 1308 -871
rect 562 -992 570 -958
rect 604 -992 638 -958
rect 672 -992 680 -958
rect 790 -992 798 -958
rect 832 -992 866 -958
rect 900 -992 908 -958
rect 162 -1092 170 -1058
rect 204 -1092 238 -1058
rect 272 -1092 280 -1058
rect 162 -1158 280 -1092
rect 390 -1058 508 -1042
rect 390 -1092 398 -1058
rect 432 -1092 466 -1058
rect 500 -1092 508 -1058
rect 390 -1108 508 -1092
rect 562 -1058 680 -992
rect 718 -1008 752 -992
rect 790 -1008 908 -992
rect 962 -958 1080 -942
rect 962 -992 970 -958
rect 1004 -992 1038 -958
rect 1072 -992 1080 -958
rect 718 -1058 752 -1042
rect 790 -1058 908 -1042
rect 562 -1092 570 -1058
rect 604 -1092 638 -1058
rect 672 -1092 680 -1058
rect 790 -1092 798 -1058
rect 832 -1092 866 -1058
rect 900 -1092 908 -1058
rect 562 -1108 680 -1092
rect 718 -1108 752 -1092
rect 162 -1192 170 -1158
rect 204 -1192 238 -1158
rect 272 -1192 280 -1158
rect 162 -1208 280 -1192
rect 390 -1158 508 -1142
rect 390 -1192 398 -1158
rect 432 -1192 466 -1158
rect 500 -1192 508 -1158
rect -82 -1258 -48 -1242
rect -10 -1258 108 -1242
rect -10 -1292 -2 -1258
rect 32 -1292 66 -1258
rect 100 -1292 108 -1258
rect -82 -1308 -48 -1292
rect -82 -1358 -48 -1342
rect -10 -1358 108 -1292
rect -10 -1392 -2 -1358
rect 32 -1392 66 -1358
rect 100 -1392 108 -1358
rect -82 -1408 -48 -1392
rect -10 -1408 108 -1392
rect 162 -1258 280 -1242
rect 162 -1292 170 -1258
rect 204 -1292 238 -1258
rect 272 -1292 280 -1258
rect 162 -1358 280 -1292
rect 162 -1392 170 -1358
rect 204 -1392 238 -1358
rect 272 -1392 280 -1358
rect 162 -1408 280 -1392
rect 390 -1258 508 -1192
rect 390 -1292 398 -1258
rect 432 -1292 466 -1258
rect 500 -1292 508 -1258
rect 390 -1358 508 -1292
rect 390 -1392 398 -1358
rect 432 -1392 466 -1358
rect 500 -1392 508 -1358
rect 390 -1408 508 -1392
rect 562 -1158 680 -1142
rect 718 -1158 752 -1142
rect 790 -1158 908 -1092
rect 562 -1192 570 -1158
rect 604 -1192 638 -1158
rect 672 -1192 680 -1158
rect 790 -1192 798 -1158
rect 832 -1192 866 -1158
rect 900 -1192 908 -1158
rect 562 -1258 680 -1192
rect 718 -1208 752 -1192
rect 790 -1208 908 -1192
rect 962 -1058 1080 -992
rect 1190 -958 1308 -892
rect 1362 -871 1368 -837
rect 1402 -858 1440 -837
rect 1362 -892 1370 -871
rect 1404 -892 1438 -858
rect 1474 -871 1480 -837
rect 1472 -892 1480 -871
rect 1590 -871 1596 -837
rect 1630 -858 1668 -837
rect 1590 -892 1598 -871
rect 1632 -892 1666 -858
rect 1702 -871 1708 -837
rect 1700 -892 1708 -871
rect 1362 -908 1480 -892
rect 1518 -908 1552 -892
rect 1190 -992 1198 -958
rect 1232 -992 1266 -958
rect 1300 -992 1308 -958
rect 1190 -1008 1308 -992
rect 1362 -958 1480 -942
rect 1518 -958 1552 -942
rect 1590 -958 1708 -892
rect 1762 -871 1768 -837
rect 1802 -858 1840 -837
rect 1762 -892 1770 -871
rect 1804 -892 1838 -858
rect 1874 -871 1880 -837
rect 1872 -892 1880 -871
rect 1762 -908 1880 -892
rect 1990 -871 1996 -837
rect 2030 -858 2068 -837
rect 1990 -892 1998 -871
rect 2032 -892 2066 -858
rect 2102 -871 2108 -837
rect 2100 -892 2108 -871
rect 1362 -992 1370 -958
rect 1404 -992 1438 -958
rect 1472 -992 1480 -958
rect 1590 -992 1598 -958
rect 1632 -992 1666 -958
rect 1700 -992 1708 -958
rect 962 -1092 970 -1058
rect 1004 -1092 1038 -1058
rect 1072 -1092 1080 -1058
rect 962 -1158 1080 -1092
rect 1190 -1058 1308 -1042
rect 1190 -1092 1198 -1058
rect 1232 -1092 1266 -1058
rect 1300 -1092 1308 -1058
rect 1190 -1108 1308 -1092
rect 1362 -1058 1480 -992
rect 1518 -1008 1552 -992
rect 1590 -1008 1708 -992
rect 1762 -958 1880 -942
rect 1762 -992 1770 -958
rect 1804 -992 1838 -958
rect 1872 -992 1880 -958
rect 1518 -1058 1552 -1042
rect 1590 -1058 1708 -1042
rect 1362 -1092 1370 -1058
rect 1404 -1092 1438 -1058
rect 1472 -1092 1480 -1058
rect 1590 -1092 1598 -1058
rect 1632 -1092 1666 -1058
rect 1700 -1092 1708 -1058
rect 1362 -1108 1480 -1092
rect 1518 -1108 1552 -1092
rect 962 -1192 970 -1158
rect 1004 -1192 1038 -1158
rect 1072 -1192 1080 -1158
rect 962 -1208 1080 -1192
rect 1190 -1158 1308 -1142
rect 1190 -1192 1198 -1158
rect 1232 -1192 1266 -1158
rect 1300 -1192 1308 -1158
rect 718 -1258 752 -1242
rect 790 -1258 908 -1242
rect 562 -1292 570 -1258
rect 604 -1292 638 -1258
rect 672 -1292 680 -1258
rect 790 -1292 798 -1258
rect 832 -1292 866 -1258
rect 900 -1292 908 -1258
rect 562 -1358 680 -1292
rect 718 -1308 752 -1292
rect 790 -1308 908 -1292
rect 962 -1258 1080 -1242
rect 962 -1292 970 -1258
rect 1004 -1292 1038 -1258
rect 1072 -1292 1080 -1258
rect 962 -1308 1080 -1292
rect 1190 -1258 1308 -1192
rect 1190 -1292 1198 -1258
rect 1232 -1292 1266 -1258
rect 1300 -1292 1308 -1258
rect 1190 -1308 1308 -1292
rect 1362 -1158 1480 -1142
rect 1518 -1158 1552 -1142
rect 1590 -1158 1708 -1092
rect 1362 -1192 1370 -1158
rect 1404 -1192 1438 -1158
rect 1472 -1192 1480 -1158
rect 1590 -1192 1598 -1158
rect 1632 -1192 1666 -1158
rect 1700 -1192 1708 -1158
rect 1362 -1258 1480 -1192
rect 1518 -1208 1552 -1192
rect 1590 -1208 1708 -1192
rect 1762 -1058 1880 -992
rect 1990 -958 2108 -892
rect 2162 -871 2168 -837
rect 2202 -858 2240 -837
rect 2162 -892 2170 -871
rect 2204 -892 2238 -858
rect 2274 -871 2280 -837
rect 2272 -892 2280 -871
rect 2390 -871 2396 -837
rect 2430 -858 2468 -837
rect 2390 -892 2398 -871
rect 2432 -892 2466 -858
rect 2502 -871 2508 -837
rect 2500 -892 2508 -871
rect 2162 -908 2280 -892
rect 2318 -908 2352 -892
rect 1990 -992 1998 -958
rect 2032 -992 2066 -958
rect 2100 -992 2108 -958
rect 1990 -1008 2108 -992
rect 2162 -958 2280 -942
rect 2318 -958 2352 -942
rect 2390 -958 2508 -892
rect 2562 -871 2568 -837
rect 2602 -858 2640 -837
rect 2562 -892 2570 -871
rect 2604 -892 2638 -858
rect 2674 -871 2680 -837
rect 2672 -892 2680 -871
rect 2562 -908 2680 -892
rect 2790 -871 2796 -837
rect 2830 -858 2868 -837
rect 2790 -892 2798 -871
rect 2832 -892 2866 -858
rect 2902 -871 2908 -837
rect 2900 -892 2908 -871
rect 2162 -992 2170 -958
rect 2204 -992 2238 -958
rect 2272 -992 2280 -958
rect 2390 -992 2398 -958
rect 2432 -992 2466 -958
rect 2500 -992 2508 -958
rect 1762 -1092 1770 -1058
rect 1804 -1092 1838 -1058
rect 1872 -1092 1880 -1058
rect 1762 -1158 1880 -1092
rect 1990 -1058 2108 -1042
rect 1990 -1092 1998 -1058
rect 2032 -1092 2066 -1058
rect 2100 -1092 2108 -1058
rect 1990 -1108 2108 -1092
rect 2162 -1058 2280 -992
rect 2318 -1008 2352 -992
rect 2390 -1008 2508 -992
rect 2562 -958 2680 -942
rect 2562 -992 2570 -958
rect 2604 -992 2638 -958
rect 2672 -992 2680 -958
rect 2318 -1058 2352 -1042
rect 2390 -1058 2508 -1042
rect 2162 -1092 2170 -1058
rect 2204 -1092 2238 -1058
rect 2272 -1092 2280 -1058
rect 2390 -1092 2398 -1058
rect 2432 -1092 2466 -1058
rect 2500 -1092 2508 -1058
rect 2162 -1108 2280 -1092
rect 2318 -1108 2352 -1092
rect 1762 -1192 1770 -1158
rect 1804 -1192 1838 -1158
rect 1872 -1192 1880 -1158
rect 1762 -1208 1880 -1192
rect 1990 -1158 2108 -1142
rect 1990 -1192 1998 -1158
rect 2032 -1192 2066 -1158
rect 2100 -1192 2108 -1158
rect 1518 -1258 1552 -1242
rect 1590 -1258 1708 -1242
rect 1362 -1292 1370 -1258
rect 1404 -1292 1438 -1258
rect 1472 -1292 1480 -1258
rect 1590 -1292 1598 -1258
rect 1632 -1292 1666 -1258
rect 1700 -1292 1708 -1258
rect 1362 -1308 1480 -1292
rect 1518 -1308 1552 -1292
rect 718 -1358 752 -1342
rect 790 -1358 908 -1342
rect 562 -1392 570 -1358
rect 604 -1392 638 -1358
rect 672 -1392 680 -1358
rect 790 -1392 798 -1358
rect 832 -1392 866 -1358
rect 900 -1392 908 -1358
rect 562 -1408 680 -1392
rect 718 -1408 752 -1392
rect -82 -1458 -48 -1442
rect -10 -1458 108 -1442
rect -10 -1492 -2 -1458
rect 32 -1492 66 -1458
rect 100 -1492 108 -1458
rect -82 -1508 -48 -1492
rect -82 -1558 -48 -1542
rect -10 -1558 108 -1492
rect -10 -1592 -2 -1558
rect 32 -1592 66 -1558
rect 100 -1592 108 -1558
rect -82 -1608 -48 -1592
rect -10 -1608 108 -1592
rect 162 -1458 280 -1442
rect 162 -1492 170 -1458
rect 204 -1492 238 -1458
rect 272 -1492 280 -1458
rect 162 -1558 280 -1492
rect 162 -1592 170 -1558
rect 204 -1592 238 -1558
rect 272 -1592 280 -1558
rect 162 -1608 280 -1592
rect 390 -1458 508 -1442
rect 390 -1492 398 -1458
rect 432 -1492 466 -1458
rect 500 -1492 508 -1458
rect 390 -1558 508 -1492
rect 390 -1592 398 -1558
rect 432 -1592 466 -1558
rect 500 -1592 508 -1558
rect 390 -1608 508 -1592
rect 562 -1458 680 -1442
rect 718 -1458 752 -1442
rect 790 -1458 908 -1392
rect 562 -1492 570 -1458
rect 604 -1492 638 -1458
rect 672 -1492 680 -1458
rect 790 -1492 798 -1458
rect 832 -1492 866 -1458
rect 900 -1492 908 -1458
rect 562 -1558 680 -1492
rect 718 -1508 752 -1492
rect 718 -1558 752 -1542
rect 790 -1558 908 -1492
rect 562 -1592 570 -1558
rect 604 -1592 638 -1558
rect 672 -1592 680 -1558
rect 790 -1592 798 -1558
rect 832 -1592 866 -1558
rect 900 -1592 908 -1558
rect 562 -1608 680 -1592
rect 718 -1608 752 -1592
rect 790 -1608 908 -1592
rect 962 -1358 1080 -1342
rect 962 -1392 970 -1358
rect 1004 -1392 1038 -1358
rect 1072 -1392 1080 -1358
rect 962 -1458 1080 -1392
rect 962 -1492 970 -1458
rect 1004 -1492 1038 -1458
rect 1072 -1492 1080 -1458
rect 962 -1558 1080 -1492
rect 962 -1592 970 -1558
rect 1004 -1592 1038 -1558
rect 1072 -1592 1080 -1558
rect 962 -1608 1080 -1592
rect 1190 -1358 1308 -1342
rect 1190 -1392 1198 -1358
rect 1232 -1392 1266 -1358
rect 1300 -1392 1308 -1358
rect 1190 -1458 1308 -1392
rect 1190 -1492 1198 -1458
rect 1232 -1492 1266 -1458
rect 1300 -1492 1308 -1458
rect 1190 -1558 1308 -1492
rect 1190 -1592 1198 -1558
rect 1232 -1592 1266 -1558
rect 1300 -1592 1308 -1558
rect 1190 -1608 1308 -1592
rect 1362 -1358 1480 -1342
rect 1518 -1358 1552 -1342
rect 1590 -1358 1708 -1292
rect 1362 -1392 1370 -1358
rect 1404 -1392 1438 -1358
rect 1472 -1392 1480 -1358
rect 1590 -1392 1598 -1358
rect 1632 -1392 1666 -1358
rect 1700 -1392 1708 -1358
rect 1362 -1458 1480 -1392
rect 1518 -1408 1552 -1392
rect 1590 -1408 1708 -1392
rect 1762 -1258 1880 -1242
rect 1762 -1292 1770 -1258
rect 1804 -1292 1838 -1258
rect 1872 -1292 1880 -1258
rect 1762 -1358 1880 -1292
rect 1762 -1392 1770 -1358
rect 1804 -1392 1838 -1358
rect 1872 -1392 1880 -1358
rect 1762 -1408 1880 -1392
rect 1990 -1258 2108 -1192
rect 1990 -1292 1998 -1258
rect 2032 -1292 2066 -1258
rect 2100 -1292 2108 -1258
rect 1990 -1358 2108 -1292
rect 1990 -1392 1998 -1358
rect 2032 -1392 2066 -1358
rect 2100 -1392 2108 -1358
rect 1990 -1408 2108 -1392
rect 2162 -1158 2280 -1142
rect 2318 -1158 2352 -1142
rect 2390 -1158 2508 -1092
rect 2162 -1192 2170 -1158
rect 2204 -1192 2238 -1158
rect 2272 -1192 2280 -1158
rect 2390 -1192 2398 -1158
rect 2432 -1192 2466 -1158
rect 2500 -1192 2508 -1158
rect 2162 -1258 2280 -1192
rect 2318 -1208 2352 -1192
rect 2390 -1208 2508 -1192
rect 2562 -1058 2680 -992
rect 2790 -958 2908 -892
rect 2962 -871 2968 -837
rect 3002 -858 3040 -837
rect 2962 -892 2970 -871
rect 3004 -892 3038 -858
rect 3074 -871 3080 -837
rect 3072 -892 3080 -871
rect 3190 -871 3196 -837
rect 3230 -858 3268 -837
rect 3190 -892 3198 -871
rect 3232 -892 3266 -858
rect 3302 -871 3308 -837
rect 3300 -892 3308 -871
rect 2962 -908 3080 -892
rect 3118 -908 3152 -892
rect 2790 -992 2798 -958
rect 2832 -992 2866 -958
rect 2900 -992 2908 -958
rect 2790 -1008 2908 -992
rect 2962 -958 3080 -942
rect 3118 -958 3152 -942
rect 3190 -958 3308 -892
rect 3362 -871 3368 -837
rect 3402 -858 3440 -837
rect 3362 -892 3370 -871
rect 3404 -892 3438 -858
rect 3474 -871 3480 -837
rect 3472 -892 3480 -871
rect 3362 -908 3480 -892
rect 3590 -871 3596 -837
rect 3630 -858 3668 -837
rect 3590 -892 3598 -871
rect 3632 -892 3666 -858
rect 3702 -871 3708 -837
rect 3700 -892 3708 -871
rect 2962 -992 2970 -958
rect 3004 -992 3038 -958
rect 3072 -992 3080 -958
rect 3190 -992 3198 -958
rect 3232 -992 3266 -958
rect 3300 -992 3308 -958
rect 2562 -1092 2570 -1058
rect 2604 -1092 2638 -1058
rect 2672 -1092 2680 -1058
rect 2562 -1158 2680 -1092
rect 2790 -1058 2908 -1042
rect 2790 -1092 2798 -1058
rect 2832 -1092 2866 -1058
rect 2900 -1092 2908 -1058
rect 2790 -1108 2908 -1092
rect 2962 -1058 3080 -992
rect 3118 -1008 3152 -992
rect 3190 -1008 3308 -992
rect 3362 -958 3480 -942
rect 3362 -992 3370 -958
rect 3404 -992 3438 -958
rect 3472 -992 3480 -958
rect 3118 -1058 3152 -1042
rect 3190 -1058 3308 -1042
rect 2962 -1092 2970 -1058
rect 3004 -1092 3038 -1058
rect 3072 -1092 3080 -1058
rect 3190 -1092 3198 -1058
rect 3232 -1092 3266 -1058
rect 3300 -1092 3308 -1058
rect 2962 -1108 3080 -1092
rect 3118 -1108 3152 -1092
rect 2562 -1192 2570 -1158
rect 2604 -1192 2638 -1158
rect 2672 -1192 2680 -1158
rect 2562 -1208 2680 -1192
rect 2790 -1158 2908 -1142
rect 2790 -1192 2798 -1158
rect 2832 -1192 2866 -1158
rect 2900 -1192 2908 -1158
rect 2318 -1258 2352 -1242
rect 2390 -1258 2508 -1242
rect 2162 -1292 2170 -1258
rect 2204 -1292 2238 -1258
rect 2272 -1292 2280 -1258
rect 2390 -1292 2398 -1258
rect 2432 -1292 2466 -1258
rect 2500 -1292 2508 -1258
rect 2162 -1358 2280 -1292
rect 2318 -1308 2352 -1292
rect 2390 -1308 2508 -1292
rect 2562 -1258 2680 -1242
rect 2562 -1292 2570 -1258
rect 2604 -1292 2638 -1258
rect 2672 -1292 2680 -1258
rect 2562 -1308 2680 -1292
rect 2790 -1258 2908 -1192
rect 2790 -1292 2798 -1258
rect 2832 -1292 2866 -1258
rect 2900 -1292 2908 -1258
rect 2790 -1308 2908 -1292
rect 2962 -1158 3080 -1142
rect 3118 -1158 3152 -1142
rect 3190 -1158 3308 -1092
rect 2962 -1192 2970 -1158
rect 3004 -1192 3038 -1158
rect 3072 -1192 3080 -1158
rect 3190 -1192 3198 -1158
rect 3232 -1192 3266 -1158
rect 3300 -1192 3308 -1158
rect 2962 -1258 3080 -1192
rect 3118 -1208 3152 -1192
rect 3190 -1208 3308 -1192
rect 3362 -1058 3480 -992
rect 3590 -958 3708 -892
rect 3762 -871 3768 -837
rect 3802 -858 3840 -837
rect 3762 -892 3770 -871
rect 3804 -892 3838 -858
rect 3874 -871 3880 -837
rect 3872 -892 3880 -871
rect 3990 -871 3996 -837
rect 4030 -858 4068 -837
rect 3990 -892 3998 -871
rect 4032 -892 4066 -858
rect 4102 -871 4108 -837
rect 4100 -892 4108 -871
rect 3762 -908 3880 -892
rect 3918 -908 3952 -892
rect 3590 -992 3598 -958
rect 3632 -992 3666 -958
rect 3700 -992 3708 -958
rect 3590 -1008 3708 -992
rect 3762 -958 3880 -942
rect 3918 -958 3952 -942
rect 3990 -958 4108 -892
rect 4162 -871 4168 -837
rect 4202 -858 4240 -837
rect 4162 -892 4170 -871
rect 4204 -892 4238 -858
rect 4274 -871 4280 -837
rect 4272 -892 4280 -871
rect 4162 -908 4280 -892
rect 4390 -871 4396 -837
rect 4430 -858 4468 -837
rect 4390 -892 4398 -871
rect 4432 -892 4466 -858
rect 4502 -871 4508 -837
rect 4500 -892 4508 -871
rect 3762 -992 3770 -958
rect 3804 -992 3838 -958
rect 3872 -992 3880 -958
rect 3990 -992 3998 -958
rect 4032 -992 4066 -958
rect 4100 -992 4108 -958
rect 3362 -1092 3370 -1058
rect 3404 -1092 3438 -1058
rect 3472 -1092 3480 -1058
rect 3362 -1158 3480 -1092
rect 3590 -1058 3708 -1042
rect 3590 -1092 3598 -1058
rect 3632 -1092 3666 -1058
rect 3700 -1092 3708 -1058
rect 3590 -1108 3708 -1092
rect 3762 -1058 3880 -992
rect 3918 -1008 3952 -992
rect 3990 -1008 4108 -992
rect 4162 -958 4280 -942
rect 4162 -992 4170 -958
rect 4204 -992 4238 -958
rect 4272 -992 4280 -958
rect 3918 -1058 3952 -1042
rect 3990 -1058 4108 -1042
rect 3762 -1092 3770 -1058
rect 3804 -1092 3838 -1058
rect 3872 -1092 3880 -1058
rect 3990 -1092 3998 -1058
rect 4032 -1092 4066 -1058
rect 4100 -1092 4108 -1058
rect 3762 -1108 3880 -1092
rect 3918 -1108 3952 -1092
rect 3362 -1192 3370 -1158
rect 3404 -1192 3438 -1158
rect 3472 -1192 3480 -1158
rect 3362 -1208 3480 -1192
rect 3590 -1158 3708 -1142
rect 3590 -1192 3598 -1158
rect 3632 -1192 3666 -1158
rect 3700 -1192 3708 -1158
rect 3118 -1258 3152 -1242
rect 3190 -1258 3308 -1242
rect 2962 -1292 2970 -1258
rect 3004 -1292 3038 -1258
rect 3072 -1292 3080 -1258
rect 3190 -1292 3198 -1258
rect 3232 -1292 3266 -1258
rect 3300 -1292 3308 -1258
rect 2962 -1308 3080 -1292
rect 3118 -1308 3152 -1292
rect 2318 -1358 2352 -1342
rect 2390 -1358 2508 -1342
rect 2162 -1392 2170 -1358
rect 2204 -1392 2238 -1358
rect 2272 -1392 2280 -1358
rect 2390 -1392 2398 -1358
rect 2432 -1392 2466 -1358
rect 2500 -1392 2508 -1358
rect 2162 -1408 2280 -1392
rect 2318 -1408 2352 -1392
rect 1518 -1458 1552 -1442
rect 1590 -1458 1708 -1442
rect 1362 -1492 1370 -1458
rect 1404 -1492 1438 -1458
rect 1472 -1492 1480 -1458
rect 1590 -1492 1598 -1458
rect 1632 -1492 1666 -1458
rect 1700 -1492 1708 -1458
rect 1362 -1558 1480 -1492
rect 1518 -1508 1552 -1492
rect 1590 -1508 1708 -1492
rect 1762 -1458 1880 -1442
rect 1762 -1492 1770 -1458
rect 1804 -1492 1838 -1458
rect 1872 -1492 1880 -1458
rect 1762 -1508 1880 -1492
rect 1990 -1458 2108 -1442
rect 1990 -1492 1998 -1458
rect 2032 -1492 2066 -1458
rect 2100 -1492 2108 -1458
rect 1990 -1508 2108 -1492
rect 2162 -1458 2280 -1442
rect 2318 -1458 2352 -1442
rect 2390 -1458 2508 -1392
rect 2162 -1492 2170 -1458
rect 2204 -1492 2238 -1458
rect 2272 -1492 2280 -1458
rect 2390 -1492 2398 -1458
rect 2432 -1492 2466 -1458
rect 2500 -1492 2508 -1458
rect 2162 -1508 2280 -1492
rect 2318 -1508 2352 -1492
rect 2390 -1508 2508 -1492
rect 2562 -1358 2680 -1342
rect 2562 -1392 2570 -1358
rect 2604 -1392 2638 -1358
rect 2672 -1392 2680 -1358
rect 2562 -1458 2680 -1392
rect 2562 -1492 2570 -1458
rect 2604 -1492 2638 -1458
rect 2672 -1492 2680 -1458
rect 2562 -1508 2680 -1492
rect 2790 -1358 2908 -1342
rect 2790 -1392 2798 -1358
rect 2832 -1392 2866 -1358
rect 2900 -1392 2908 -1358
rect 2790 -1458 2908 -1392
rect 2790 -1492 2798 -1458
rect 2832 -1492 2866 -1458
rect 2900 -1492 2908 -1458
rect 2790 -1508 2908 -1492
rect 2962 -1358 3080 -1342
rect 3118 -1358 3152 -1342
rect 3190 -1358 3308 -1292
rect 2962 -1392 2970 -1358
rect 3004 -1392 3038 -1358
rect 3072 -1392 3080 -1358
rect 3190 -1392 3198 -1358
rect 3232 -1392 3266 -1358
rect 3300 -1392 3308 -1358
rect 2962 -1458 3080 -1392
rect 3118 -1408 3152 -1392
rect 3190 -1408 3308 -1392
rect 3362 -1258 3480 -1242
rect 3362 -1292 3370 -1258
rect 3404 -1292 3438 -1258
rect 3472 -1292 3480 -1258
rect 3362 -1358 3480 -1292
rect 3362 -1392 3370 -1358
rect 3404 -1392 3438 -1358
rect 3472 -1392 3480 -1358
rect 3362 -1408 3480 -1392
rect 3590 -1258 3708 -1192
rect 3590 -1292 3598 -1258
rect 3632 -1292 3666 -1258
rect 3700 -1292 3708 -1258
rect 3590 -1358 3708 -1292
rect 3590 -1392 3598 -1358
rect 3632 -1392 3666 -1358
rect 3700 -1392 3708 -1358
rect 3590 -1408 3708 -1392
rect 3762 -1158 3880 -1142
rect 3918 -1158 3952 -1142
rect 3990 -1158 4108 -1092
rect 3762 -1192 3770 -1158
rect 3804 -1192 3838 -1158
rect 3872 -1192 3880 -1158
rect 3990 -1192 3998 -1158
rect 4032 -1192 4066 -1158
rect 4100 -1192 4108 -1158
rect 3762 -1258 3880 -1192
rect 3918 -1208 3952 -1192
rect 3990 -1208 4108 -1192
rect 4162 -1058 4280 -992
rect 4390 -958 4508 -892
rect 4562 -871 4568 -837
rect 4602 -858 4640 -837
rect 4562 -892 4570 -871
rect 4604 -892 4638 -858
rect 4674 -871 4680 -837
rect 4672 -892 4680 -871
rect 4790 -871 4796 -837
rect 4830 -858 4868 -837
rect 4790 -892 4798 -871
rect 4832 -892 4866 -858
rect 4902 -871 4908 -837
rect 4900 -892 4908 -871
rect 4562 -908 4680 -892
rect 4718 -908 4752 -892
rect 4390 -992 4398 -958
rect 4432 -992 4466 -958
rect 4500 -992 4508 -958
rect 4390 -1008 4508 -992
rect 4562 -958 4680 -942
rect 4718 -958 4752 -942
rect 4790 -958 4908 -892
rect 4962 -871 4968 -837
rect 5002 -858 5040 -837
rect 4962 -892 4970 -871
rect 5004 -892 5038 -858
rect 5074 -871 5080 -837
rect 5072 -892 5080 -871
rect 4962 -908 5080 -892
rect 5190 -871 5196 -837
rect 5230 -858 5268 -837
rect 5190 -892 5198 -871
rect 5232 -892 5266 -858
rect 5302 -871 5308 -837
rect 5300 -892 5308 -871
rect 4562 -992 4570 -958
rect 4604 -992 4638 -958
rect 4672 -992 4680 -958
rect 4790 -992 4798 -958
rect 4832 -992 4866 -958
rect 4900 -992 4908 -958
rect 4162 -1092 4170 -1058
rect 4204 -1092 4238 -1058
rect 4272 -1092 4280 -1058
rect 4162 -1158 4280 -1092
rect 4390 -1058 4508 -1042
rect 4390 -1092 4398 -1058
rect 4432 -1092 4466 -1058
rect 4500 -1092 4508 -1058
rect 4390 -1108 4508 -1092
rect 4562 -1058 4680 -992
rect 4718 -1008 4752 -992
rect 4790 -1008 4908 -992
rect 4962 -958 5080 -942
rect 4962 -992 4970 -958
rect 5004 -992 5038 -958
rect 5072 -992 5080 -958
rect 4718 -1058 4752 -1042
rect 4790 -1058 4908 -1042
rect 4562 -1092 4570 -1058
rect 4604 -1092 4638 -1058
rect 4672 -1092 4680 -1058
rect 4790 -1092 4798 -1058
rect 4832 -1092 4866 -1058
rect 4900 -1092 4908 -1058
rect 4562 -1108 4680 -1092
rect 4718 -1108 4752 -1092
rect 4162 -1192 4170 -1158
rect 4204 -1192 4238 -1158
rect 4272 -1192 4280 -1158
rect 4162 -1208 4280 -1192
rect 4390 -1158 4508 -1142
rect 4390 -1192 4398 -1158
rect 4432 -1192 4466 -1158
rect 4500 -1192 4508 -1158
rect 3918 -1258 3952 -1242
rect 3990 -1258 4108 -1242
rect 3762 -1292 3770 -1258
rect 3804 -1292 3838 -1258
rect 3872 -1292 3880 -1258
rect 3990 -1292 3998 -1258
rect 4032 -1292 4066 -1258
rect 4100 -1292 4108 -1258
rect 3762 -1358 3880 -1292
rect 3918 -1308 3952 -1292
rect 3990 -1308 4108 -1292
rect 4162 -1258 4280 -1242
rect 4162 -1292 4170 -1258
rect 4204 -1292 4238 -1258
rect 4272 -1292 4280 -1258
rect 4162 -1308 4280 -1292
rect 4390 -1258 4508 -1192
rect 4390 -1292 4398 -1258
rect 4432 -1292 4466 -1258
rect 4500 -1292 4508 -1258
rect 4390 -1308 4508 -1292
rect 4562 -1158 4680 -1142
rect 4718 -1158 4752 -1142
rect 4790 -1158 4908 -1092
rect 4562 -1192 4570 -1158
rect 4604 -1192 4638 -1158
rect 4672 -1192 4680 -1158
rect 4790 -1192 4798 -1158
rect 4832 -1192 4866 -1158
rect 4900 -1192 4908 -1158
rect 4562 -1258 4680 -1192
rect 4718 -1208 4752 -1192
rect 4790 -1208 4908 -1192
rect 4962 -1058 5080 -992
rect 5190 -958 5308 -892
rect 5362 -871 5368 -837
rect 5402 -858 5440 -837
rect 5362 -892 5370 -871
rect 5404 -892 5438 -858
rect 5474 -871 5480 -837
rect 5472 -892 5480 -871
rect 5590 -871 5596 -837
rect 5630 -858 5668 -837
rect 5590 -892 5598 -871
rect 5632 -892 5666 -858
rect 5702 -871 5708 -837
rect 5700 -892 5708 -871
rect 5362 -908 5480 -892
rect 5518 -908 5552 -892
rect 5190 -992 5198 -958
rect 5232 -992 5266 -958
rect 5300 -992 5308 -958
rect 5190 -1008 5308 -992
rect 5362 -958 5480 -942
rect 5518 -958 5552 -942
rect 5590 -958 5708 -892
rect 5762 -871 5768 -837
rect 5802 -858 5840 -837
rect 5762 -892 5770 -871
rect 5804 -892 5838 -858
rect 5874 -871 5880 -837
rect 5872 -892 5880 -871
rect 5762 -908 5880 -892
rect 5990 -871 5996 -837
rect 6030 -858 6068 -837
rect 5990 -892 5998 -871
rect 6032 -892 6066 -858
rect 6102 -871 6108 -837
rect 6100 -892 6108 -871
rect 5362 -992 5370 -958
rect 5404 -992 5438 -958
rect 5472 -992 5480 -958
rect 5590 -992 5598 -958
rect 5632 -992 5666 -958
rect 5700 -992 5708 -958
rect 4962 -1092 4970 -1058
rect 5004 -1092 5038 -1058
rect 5072 -1092 5080 -1058
rect 4962 -1158 5080 -1092
rect 5190 -1058 5308 -1042
rect 5190 -1092 5198 -1058
rect 5232 -1092 5266 -1058
rect 5300 -1092 5308 -1058
rect 5190 -1108 5308 -1092
rect 5362 -1058 5480 -992
rect 5518 -1008 5552 -992
rect 5590 -1008 5708 -992
rect 5762 -958 5880 -942
rect 5762 -992 5770 -958
rect 5804 -992 5838 -958
rect 5872 -992 5880 -958
rect 5518 -1058 5552 -1042
rect 5590 -1058 5708 -1042
rect 5362 -1092 5370 -1058
rect 5404 -1092 5438 -1058
rect 5472 -1092 5480 -1058
rect 5590 -1092 5598 -1058
rect 5632 -1092 5666 -1058
rect 5700 -1092 5708 -1058
rect 5362 -1108 5480 -1092
rect 5518 -1108 5552 -1092
rect 4962 -1192 4970 -1158
rect 5004 -1192 5038 -1158
rect 5072 -1192 5080 -1158
rect 4962 -1208 5080 -1192
rect 5190 -1158 5308 -1142
rect 5190 -1192 5198 -1158
rect 5232 -1192 5266 -1158
rect 5300 -1192 5308 -1158
rect 4718 -1258 4752 -1242
rect 4790 -1258 4908 -1242
rect 4562 -1292 4570 -1258
rect 4604 -1292 4638 -1258
rect 4672 -1292 4680 -1258
rect 4790 -1292 4798 -1258
rect 4832 -1292 4866 -1258
rect 4900 -1292 4908 -1258
rect 4562 -1308 4680 -1292
rect 4718 -1308 4752 -1292
rect 3918 -1358 3952 -1342
rect 3990 -1358 4108 -1342
rect 3762 -1392 3770 -1358
rect 3804 -1392 3838 -1358
rect 3872 -1392 3880 -1358
rect 3990 -1392 3998 -1358
rect 4032 -1392 4066 -1358
rect 4100 -1392 4108 -1358
rect 3762 -1408 3880 -1392
rect 3918 -1408 3952 -1392
rect 3118 -1458 3152 -1442
rect 3190 -1458 3308 -1442
rect 2962 -1492 2970 -1458
rect 3004 -1492 3038 -1458
rect 3072 -1492 3080 -1458
rect 3190 -1492 3198 -1458
rect 3232 -1492 3266 -1458
rect 3300 -1492 3308 -1458
rect 2962 -1508 3080 -1492
rect 3118 -1508 3152 -1492
rect 1518 -1558 1552 -1542
rect 1590 -1558 1708 -1542
rect 1362 -1592 1370 -1558
rect 1404 -1592 1438 -1558
rect 1472 -1592 1480 -1558
rect 1590 -1592 1598 -1558
rect 1632 -1592 1666 -1558
rect 1700 -1592 1708 -1558
rect 1362 -1608 1480 -1592
rect 1518 -1608 1552 -1592
rect -82 -1658 -48 -1642
rect -10 -1658 108 -1642
rect -10 -1692 -2 -1658
rect 32 -1692 66 -1658
rect 100 -1692 108 -1658
rect -82 -1708 -48 -1692
rect -82 -1758 -48 -1742
rect -10 -1758 108 -1692
rect -10 -1792 -2 -1758
rect 32 -1792 66 -1758
rect 100 -1792 108 -1758
rect -82 -1808 -48 -1792
rect -10 -1808 108 -1792
rect 162 -1658 280 -1642
rect 162 -1692 170 -1658
rect 204 -1692 238 -1658
rect 272 -1692 280 -1658
rect 162 -1758 280 -1692
rect 162 -1792 170 -1758
rect 204 -1792 238 -1758
rect 272 -1792 280 -1758
rect 162 -1808 280 -1792
rect 390 -1658 508 -1642
rect 390 -1692 398 -1658
rect 432 -1692 466 -1658
rect 500 -1692 508 -1658
rect 390 -1758 508 -1692
rect 390 -1792 398 -1758
rect 432 -1792 466 -1758
rect 500 -1792 508 -1758
rect 390 -1808 508 -1792
rect 562 -1658 680 -1642
rect 718 -1658 752 -1642
rect 790 -1658 908 -1642
rect 562 -1692 570 -1658
rect 604 -1692 638 -1658
rect 672 -1692 680 -1658
rect 790 -1692 798 -1658
rect 832 -1692 866 -1658
rect 900 -1692 908 -1658
rect 562 -1758 680 -1692
rect 718 -1708 752 -1692
rect 718 -1758 752 -1742
rect 790 -1758 908 -1692
rect 562 -1792 570 -1758
rect 604 -1792 638 -1758
rect 672 -1792 680 -1758
rect 790 -1792 798 -1758
rect 832 -1792 866 -1758
rect 900 -1792 908 -1758
rect 562 -1808 680 -1792
rect 718 -1808 752 -1792
rect 790 -1808 908 -1792
rect 962 -1658 1080 -1642
rect 962 -1692 970 -1658
rect 1004 -1692 1038 -1658
rect 1072 -1692 1080 -1658
rect 962 -1758 1080 -1692
rect 962 -1792 970 -1758
rect 1004 -1792 1038 -1758
rect 1072 -1792 1080 -1758
rect 962 -1808 1080 -1792
rect 1190 -1658 1308 -1642
rect 1190 -1692 1198 -1658
rect 1232 -1692 1266 -1658
rect 1300 -1692 1308 -1658
rect 1190 -1758 1308 -1692
rect 1190 -1792 1198 -1758
rect 1232 -1792 1266 -1758
rect 1300 -1792 1308 -1758
rect 1190 -1808 1308 -1792
rect 1362 -1658 1480 -1642
rect 1518 -1658 1552 -1642
rect 1590 -1658 1708 -1592
rect 1362 -1692 1370 -1658
rect 1404 -1692 1438 -1658
rect 1472 -1692 1480 -1658
rect 1590 -1692 1598 -1658
rect 1632 -1692 1666 -1658
rect 1700 -1692 1708 -1658
rect 1362 -1758 1480 -1692
rect 1518 -1708 1552 -1692
rect 1518 -1758 1552 -1742
rect 1590 -1758 1708 -1692
rect 1362 -1792 1370 -1758
rect 1404 -1792 1438 -1758
rect 1472 -1792 1480 -1758
rect 1590 -1792 1598 -1758
rect 1632 -1792 1666 -1758
rect 1700 -1792 1708 -1758
rect 1362 -1808 1480 -1792
rect 1518 -1808 1552 -1792
rect 1590 -1808 1708 -1792
rect 1762 -1558 1880 -1542
rect 1762 -1592 1770 -1558
rect 1804 -1592 1838 -1558
rect 1872 -1592 1880 -1558
rect 1762 -1658 1880 -1592
rect 1762 -1692 1770 -1658
rect 1804 -1692 1838 -1658
rect 1872 -1692 1880 -1658
rect 1762 -1758 1880 -1692
rect 1762 -1792 1770 -1758
rect 1804 -1792 1838 -1758
rect 1872 -1792 1880 -1758
rect 1762 -1808 1880 -1792
rect 1990 -1558 2108 -1542
rect 1990 -1592 1998 -1558
rect 2032 -1592 2066 -1558
rect 2100 -1592 2108 -1558
rect 1990 -1658 2108 -1592
rect 1990 -1692 1998 -1658
rect 2032 -1692 2066 -1658
rect 2100 -1692 2108 -1658
rect 1990 -1758 2108 -1692
rect 1990 -1792 1998 -1758
rect 2032 -1792 2066 -1758
rect 2100 -1792 2108 -1758
rect 1990 -1808 2108 -1792
rect 2162 -1558 2280 -1542
rect 2318 -1558 2352 -1542
rect 2390 -1558 2508 -1542
rect 2162 -1592 2170 -1558
rect 2204 -1592 2238 -1558
rect 2272 -1592 2280 -1558
rect 2390 -1592 2398 -1558
rect 2432 -1592 2466 -1558
rect 2500 -1592 2508 -1558
rect 2162 -1658 2280 -1592
rect 2318 -1608 2352 -1592
rect 2318 -1658 2352 -1642
rect 2390 -1658 2508 -1592
rect 2162 -1692 2170 -1658
rect 2204 -1692 2238 -1658
rect 2272 -1692 2280 -1658
rect 2390 -1692 2398 -1658
rect 2432 -1692 2466 -1658
rect 2500 -1692 2508 -1658
rect 2162 -1758 2280 -1692
rect 2318 -1708 2352 -1692
rect 2318 -1758 2352 -1742
rect 2390 -1758 2508 -1692
rect 2162 -1792 2170 -1758
rect 2204 -1792 2238 -1758
rect 2272 -1792 2280 -1758
rect 2390 -1792 2398 -1758
rect 2432 -1792 2466 -1758
rect 2500 -1792 2508 -1758
rect 2162 -1808 2280 -1792
rect 2318 -1808 2352 -1792
rect 2390 -1808 2508 -1792
rect 2562 -1558 2680 -1542
rect 2562 -1592 2570 -1558
rect 2604 -1592 2638 -1558
rect 2672 -1592 2680 -1558
rect 2562 -1658 2680 -1592
rect 2562 -1692 2570 -1658
rect 2604 -1692 2638 -1658
rect 2672 -1692 2680 -1658
rect 2562 -1758 2680 -1692
rect 2562 -1792 2570 -1758
rect 2604 -1792 2638 -1758
rect 2672 -1792 2680 -1758
rect 2562 -1808 2680 -1792
rect 2790 -1558 2908 -1542
rect 2790 -1592 2798 -1558
rect 2832 -1592 2866 -1558
rect 2900 -1592 2908 -1558
rect 2790 -1658 2908 -1592
rect 2790 -1692 2798 -1658
rect 2832 -1692 2866 -1658
rect 2900 -1692 2908 -1658
rect 2790 -1758 2908 -1692
rect 2790 -1792 2798 -1758
rect 2832 -1792 2866 -1758
rect 2900 -1792 2908 -1758
rect 2790 -1808 2908 -1792
rect 2962 -1558 3080 -1542
rect 3118 -1558 3152 -1542
rect 3190 -1558 3308 -1492
rect 2962 -1592 2970 -1558
rect 3004 -1592 3038 -1558
rect 3072 -1592 3080 -1558
rect 3190 -1592 3198 -1558
rect 3232 -1592 3266 -1558
rect 3300 -1592 3308 -1558
rect 2962 -1658 3080 -1592
rect 3118 -1608 3152 -1592
rect 3190 -1608 3308 -1592
rect 3362 -1458 3480 -1442
rect 3362 -1492 3370 -1458
rect 3404 -1492 3438 -1458
rect 3472 -1492 3480 -1458
rect 3362 -1558 3480 -1492
rect 3362 -1592 3370 -1558
rect 3404 -1592 3438 -1558
rect 3472 -1592 3480 -1558
rect 3362 -1608 3480 -1592
rect 3590 -1458 3708 -1442
rect 3590 -1492 3598 -1458
rect 3632 -1492 3666 -1458
rect 3700 -1492 3708 -1458
rect 3590 -1558 3708 -1492
rect 3590 -1592 3598 -1558
rect 3632 -1592 3666 -1558
rect 3700 -1592 3708 -1558
rect 3590 -1608 3708 -1592
rect 3762 -1458 3880 -1442
rect 3918 -1458 3952 -1442
rect 3990 -1458 4108 -1392
rect 3762 -1492 3770 -1458
rect 3804 -1492 3838 -1458
rect 3872 -1492 3880 -1458
rect 3990 -1492 3998 -1458
rect 4032 -1492 4066 -1458
rect 4100 -1492 4108 -1458
rect 3762 -1558 3880 -1492
rect 3918 -1508 3952 -1492
rect 3918 -1558 3952 -1542
rect 3990 -1558 4108 -1492
rect 3762 -1592 3770 -1558
rect 3804 -1592 3838 -1558
rect 3872 -1592 3880 -1558
rect 3990 -1592 3998 -1558
rect 4032 -1592 4066 -1558
rect 4100 -1592 4108 -1558
rect 3762 -1608 3880 -1592
rect 3918 -1608 3952 -1592
rect 3990 -1608 4108 -1592
rect 4162 -1358 4280 -1342
rect 4162 -1392 4170 -1358
rect 4204 -1392 4238 -1358
rect 4272 -1392 4280 -1358
rect 4162 -1458 4280 -1392
rect 4162 -1492 4170 -1458
rect 4204 -1492 4238 -1458
rect 4272 -1492 4280 -1458
rect 4162 -1558 4280 -1492
rect 4162 -1592 4170 -1558
rect 4204 -1592 4238 -1558
rect 4272 -1592 4280 -1558
rect 4162 -1608 4280 -1592
rect 4390 -1358 4508 -1342
rect 4390 -1392 4398 -1358
rect 4432 -1392 4466 -1358
rect 4500 -1392 4508 -1358
rect 4390 -1458 4508 -1392
rect 4390 -1492 4398 -1458
rect 4432 -1492 4466 -1458
rect 4500 -1492 4508 -1458
rect 4390 -1558 4508 -1492
rect 4390 -1592 4398 -1558
rect 4432 -1592 4466 -1558
rect 4500 -1592 4508 -1558
rect 4390 -1608 4508 -1592
rect 4562 -1358 4680 -1342
rect 4718 -1358 4752 -1342
rect 4790 -1358 4908 -1292
rect 4562 -1392 4570 -1358
rect 4604 -1392 4638 -1358
rect 4672 -1392 4680 -1358
rect 4790 -1392 4798 -1358
rect 4832 -1392 4866 -1358
rect 4900 -1392 4908 -1358
rect 4562 -1458 4680 -1392
rect 4718 -1408 4752 -1392
rect 4790 -1408 4908 -1392
rect 4962 -1258 5080 -1242
rect 4962 -1292 4970 -1258
rect 5004 -1292 5038 -1258
rect 5072 -1292 5080 -1258
rect 4962 -1358 5080 -1292
rect 4962 -1392 4970 -1358
rect 5004 -1392 5038 -1358
rect 5072 -1392 5080 -1358
rect 4962 -1408 5080 -1392
rect 5190 -1258 5308 -1192
rect 5190 -1292 5198 -1258
rect 5232 -1292 5266 -1258
rect 5300 -1292 5308 -1258
rect 5190 -1358 5308 -1292
rect 5190 -1392 5198 -1358
rect 5232 -1392 5266 -1358
rect 5300 -1392 5308 -1358
rect 5190 -1408 5308 -1392
rect 5362 -1158 5480 -1142
rect 5518 -1158 5552 -1142
rect 5590 -1158 5708 -1092
rect 5362 -1192 5370 -1158
rect 5404 -1192 5438 -1158
rect 5472 -1192 5480 -1158
rect 5590 -1192 5598 -1158
rect 5632 -1192 5666 -1158
rect 5700 -1192 5708 -1158
rect 5362 -1258 5480 -1192
rect 5518 -1208 5552 -1192
rect 5590 -1208 5708 -1192
rect 5762 -1058 5880 -992
rect 5990 -958 6108 -892
rect 6162 -871 6168 -837
rect 6202 -858 6240 -837
rect 6162 -892 6170 -871
rect 6204 -892 6238 -858
rect 6274 -871 6280 -837
rect 6272 -892 6280 -871
rect 6390 -871 6396 -837
rect 6430 -858 6468 -837
rect 6390 -892 6398 -871
rect 6432 -892 6466 -858
rect 6502 -871 6508 -837
rect 6500 -892 6508 -871
rect 6162 -908 6280 -892
rect 6318 -908 6352 -892
rect 5990 -992 5998 -958
rect 6032 -992 6066 -958
rect 6100 -992 6108 -958
rect 5990 -1008 6108 -992
rect 6162 -958 6280 -942
rect 6318 -958 6352 -942
rect 6390 -958 6508 -892
rect 6562 -871 6568 -837
rect 6602 -858 6640 -837
rect 6562 -892 6570 -871
rect 6604 -892 6638 -858
rect 6674 -871 6680 -837
rect 6672 -892 6680 -871
rect 6562 -908 6680 -892
rect 6790 -871 6796 -837
rect 6830 -858 6868 -837
rect 6790 -892 6798 -871
rect 6832 -892 6866 -858
rect 6902 -871 6908 -837
rect 6900 -892 6908 -871
rect 6162 -992 6170 -958
rect 6204 -992 6238 -958
rect 6272 -992 6280 -958
rect 6390 -992 6398 -958
rect 6432 -992 6466 -958
rect 6500 -992 6508 -958
rect 5762 -1092 5770 -1058
rect 5804 -1092 5838 -1058
rect 5872 -1092 5880 -1058
rect 5762 -1158 5880 -1092
rect 5990 -1058 6108 -1042
rect 5990 -1092 5998 -1058
rect 6032 -1092 6066 -1058
rect 6100 -1092 6108 -1058
rect 5990 -1108 6108 -1092
rect 6162 -1058 6280 -992
rect 6318 -1008 6352 -992
rect 6390 -1008 6508 -992
rect 6562 -958 6680 -942
rect 6562 -992 6570 -958
rect 6604 -992 6638 -958
rect 6672 -992 6680 -958
rect 6318 -1058 6352 -1042
rect 6390 -1058 6508 -1042
rect 6162 -1092 6170 -1058
rect 6204 -1092 6238 -1058
rect 6272 -1092 6280 -1058
rect 6390 -1092 6398 -1058
rect 6432 -1092 6466 -1058
rect 6500 -1092 6508 -1058
rect 6162 -1108 6280 -1092
rect 6318 -1108 6352 -1092
rect 5762 -1192 5770 -1158
rect 5804 -1192 5838 -1158
rect 5872 -1192 5880 -1158
rect 5762 -1208 5880 -1192
rect 5990 -1158 6108 -1142
rect 5990 -1192 5998 -1158
rect 6032 -1192 6066 -1158
rect 6100 -1192 6108 -1158
rect 5518 -1258 5552 -1242
rect 5590 -1258 5708 -1242
rect 5362 -1292 5370 -1258
rect 5404 -1292 5438 -1258
rect 5472 -1292 5480 -1258
rect 5590 -1292 5598 -1258
rect 5632 -1292 5666 -1258
rect 5700 -1292 5708 -1258
rect 5362 -1358 5480 -1292
rect 5518 -1308 5552 -1292
rect 5590 -1308 5708 -1292
rect 5762 -1258 5880 -1242
rect 5762 -1292 5770 -1258
rect 5804 -1292 5838 -1258
rect 5872 -1292 5880 -1258
rect 5762 -1308 5880 -1292
rect 5990 -1258 6108 -1192
rect 5990 -1292 5998 -1258
rect 6032 -1292 6066 -1258
rect 6100 -1292 6108 -1258
rect 5990 -1308 6108 -1292
rect 6162 -1158 6280 -1142
rect 6318 -1158 6352 -1142
rect 6390 -1158 6508 -1092
rect 6162 -1192 6170 -1158
rect 6204 -1192 6238 -1158
rect 6272 -1192 6280 -1158
rect 6390 -1192 6398 -1158
rect 6432 -1192 6466 -1158
rect 6500 -1192 6508 -1158
rect 6162 -1258 6280 -1192
rect 6318 -1208 6352 -1192
rect 6390 -1208 6508 -1192
rect 6562 -1058 6680 -992
rect 6790 -958 6908 -892
rect 6962 -871 6968 -837
rect 7002 -858 7040 -837
rect 6962 -892 6970 -871
rect 7004 -892 7038 -858
rect 7074 -871 7080 -837
rect 7072 -892 7080 -871
rect 7190 -871 7196 -837
rect 7230 -858 7268 -837
rect 7190 -892 7198 -871
rect 7232 -892 7266 -858
rect 7302 -871 7308 -837
rect 7300 -892 7308 -871
rect 6962 -908 7080 -892
rect 7118 -908 7152 -892
rect 6790 -992 6798 -958
rect 6832 -992 6866 -958
rect 6900 -992 6908 -958
rect 6790 -1008 6908 -992
rect 6962 -958 7080 -942
rect 7118 -958 7152 -942
rect 7190 -958 7308 -892
rect 7362 -871 7368 -837
rect 7402 -858 7440 -837
rect 7362 -892 7370 -871
rect 7404 -892 7438 -858
rect 7474 -871 7480 -837
rect 7472 -892 7480 -871
rect 7362 -908 7480 -892
rect 7590 -871 7596 -837
rect 7630 -858 7668 -837
rect 7590 -892 7598 -871
rect 7632 -892 7666 -858
rect 7702 -871 7708 -837
rect 7700 -892 7708 -871
rect 6962 -992 6970 -958
rect 7004 -992 7038 -958
rect 7072 -992 7080 -958
rect 7190 -992 7198 -958
rect 7232 -992 7266 -958
rect 7300 -992 7308 -958
rect 6562 -1092 6570 -1058
rect 6604 -1092 6638 -1058
rect 6672 -1092 6680 -1058
rect 6562 -1158 6680 -1092
rect 6790 -1058 6908 -1042
rect 6790 -1092 6798 -1058
rect 6832 -1092 6866 -1058
rect 6900 -1092 6908 -1058
rect 6790 -1108 6908 -1092
rect 6962 -1058 7080 -992
rect 7118 -1008 7152 -992
rect 7190 -1008 7308 -992
rect 7362 -958 7480 -942
rect 7362 -992 7370 -958
rect 7404 -992 7438 -958
rect 7472 -992 7480 -958
rect 7118 -1058 7152 -1042
rect 7190 -1058 7308 -1042
rect 6962 -1092 6970 -1058
rect 7004 -1092 7038 -1058
rect 7072 -1092 7080 -1058
rect 7190 -1092 7198 -1058
rect 7232 -1092 7266 -1058
rect 7300 -1092 7308 -1058
rect 6962 -1108 7080 -1092
rect 7118 -1108 7152 -1092
rect 6562 -1192 6570 -1158
rect 6604 -1192 6638 -1158
rect 6672 -1192 6680 -1158
rect 6562 -1208 6680 -1192
rect 6790 -1158 6908 -1142
rect 6790 -1192 6798 -1158
rect 6832 -1192 6866 -1158
rect 6900 -1192 6908 -1158
rect 6318 -1258 6352 -1242
rect 6390 -1258 6508 -1242
rect 6162 -1292 6170 -1258
rect 6204 -1292 6238 -1258
rect 6272 -1292 6280 -1258
rect 6390 -1292 6398 -1258
rect 6432 -1292 6466 -1258
rect 6500 -1292 6508 -1258
rect 6162 -1308 6280 -1292
rect 6318 -1308 6352 -1292
rect 5518 -1358 5552 -1342
rect 5590 -1358 5708 -1342
rect 5362 -1392 5370 -1358
rect 5404 -1392 5438 -1358
rect 5472 -1392 5480 -1358
rect 5590 -1392 5598 -1358
rect 5632 -1392 5666 -1358
rect 5700 -1392 5708 -1358
rect 5362 -1408 5480 -1392
rect 5518 -1408 5552 -1392
rect 4718 -1458 4752 -1442
rect 4790 -1458 4908 -1442
rect 4562 -1492 4570 -1458
rect 4604 -1492 4638 -1458
rect 4672 -1492 4680 -1458
rect 4790 -1492 4798 -1458
rect 4832 -1492 4866 -1458
rect 4900 -1492 4908 -1458
rect 4562 -1558 4680 -1492
rect 4718 -1508 4752 -1492
rect 4790 -1508 4908 -1492
rect 4962 -1458 5080 -1442
rect 4962 -1492 4970 -1458
rect 5004 -1492 5038 -1458
rect 5072 -1492 5080 -1458
rect 4962 -1508 5080 -1492
rect 5190 -1458 5308 -1442
rect 5190 -1492 5198 -1458
rect 5232 -1492 5266 -1458
rect 5300 -1492 5308 -1458
rect 5190 -1508 5308 -1492
rect 5362 -1458 5480 -1442
rect 5518 -1458 5552 -1442
rect 5590 -1458 5708 -1392
rect 5362 -1492 5370 -1458
rect 5404 -1492 5438 -1458
rect 5472 -1492 5480 -1458
rect 5590 -1492 5598 -1458
rect 5632 -1492 5666 -1458
rect 5700 -1492 5708 -1458
rect 5362 -1508 5480 -1492
rect 5518 -1508 5552 -1492
rect 5590 -1508 5708 -1492
rect 5762 -1358 5880 -1342
rect 5762 -1392 5770 -1358
rect 5804 -1392 5838 -1358
rect 5872 -1392 5880 -1358
rect 5762 -1458 5880 -1392
rect 5762 -1492 5770 -1458
rect 5804 -1492 5838 -1458
rect 5872 -1492 5880 -1458
rect 5762 -1508 5880 -1492
rect 5990 -1358 6108 -1342
rect 5990 -1392 5998 -1358
rect 6032 -1392 6066 -1358
rect 6100 -1392 6108 -1358
rect 5990 -1458 6108 -1392
rect 5990 -1492 5998 -1458
rect 6032 -1492 6066 -1458
rect 6100 -1492 6108 -1458
rect 5990 -1508 6108 -1492
rect 6162 -1358 6280 -1342
rect 6318 -1358 6352 -1342
rect 6390 -1358 6508 -1292
rect 6162 -1392 6170 -1358
rect 6204 -1392 6238 -1358
rect 6272 -1392 6280 -1358
rect 6390 -1392 6398 -1358
rect 6432 -1392 6466 -1358
rect 6500 -1392 6508 -1358
rect 6162 -1458 6280 -1392
rect 6318 -1408 6352 -1392
rect 6390 -1408 6508 -1392
rect 6562 -1258 6680 -1242
rect 6562 -1292 6570 -1258
rect 6604 -1292 6638 -1258
rect 6672 -1292 6680 -1258
rect 6562 -1358 6680 -1292
rect 6562 -1392 6570 -1358
rect 6604 -1392 6638 -1358
rect 6672 -1392 6680 -1358
rect 6562 -1408 6680 -1392
rect 6790 -1258 6908 -1192
rect 6790 -1292 6798 -1258
rect 6832 -1292 6866 -1258
rect 6900 -1292 6908 -1258
rect 6790 -1358 6908 -1292
rect 6790 -1392 6798 -1358
rect 6832 -1392 6866 -1358
rect 6900 -1392 6908 -1358
rect 6790 -1408 6908 -1392
rect 6962 -1158 7080 -1142
rect 7118 -1158 7152 -1142
rect 7190 -1158 7308 -1092
rect 6962 -1192 6970 -1158
rect 7004 -1192 7038 -1158
rect 7072 -1192 7080 -1158
rect 7190 -1192 7198 -1158
rect 7232 -1192 7266 -1158
rect 7300 -1192 7308 -1158
rect 6962 -1258 7080 -1192
rect 7118 -1208 7152 -1192
rect 7190 -1208 7308 -1192
rect 7362 -1058 7480 -992
rect 7590 -958 7708 -892
rect 7762 -871 7768 -837
rect 7802 -858 7840 -837
rect 7762 -892 7770 -871
rect 7804 -892 7838 -858
rect 7874 -871 7880 -837
rect 7872 -892 7880 -871
rect 7990 -871 7996 -837
rect 8030 -858 8068 -837
rect 7990 -892 7998 -871
rect 8032 -892 8066 -858
rect 8102 -871 8108 -837
rect 8100 -892 8108 -871
rect 7762 -908 7880 -892
rect 7918 -908 7952 -892
rect 7590 -992 7598 -958
rect 7632 -992 7666 -958
rect 7700 -992 7708 -958
rect 7590 -1008 7708 -992
rect 7762 -958 7880 -942
rect 7918 -958 7952 -942
rect 7990 -958 8108 -892
rect 8162 -871 8168 -837
rect 8202 -858 8240 -837
rect 8162 -892 8170 -871
rect 8204 -892 8238 -858
rect 8274 -871 8280 -837
rect 8272 -892 8280 -871
rect 8162 -908 8280 -892
rect 8390 -871 8396 -837
rect 8430 -858 8468 -837
rect 8390 -892 8398 -871
rect 8432 -892 8466 -858
rect 8502 -871 8508 -837
rect 8500 -892 8508 -871
rect 7762 -992 7770 -958
rect 7804 -992 7838 -958
rect 7872 -992 7880 -958
rect 7990 -992 7998 -958
rect 8032 -992 8066 -958
rect 8100 -992 8108 -958
rect 7362 -1092 7370 -1058
rect 7404 -1092 7438 -1058
rect 7472 -1092 7480 -1058
rect 7362 -1158 7480 -1092
rect 7590 -1058 7708 -1042
rect 7590 -1092 7598 -1058
rect 7632 -1092 7666 -1058
rect 7700 -1092 7708 -1058
rect 7590 -1108 7708 -1092
rect 7762 -1058 7880 -992
rect 7918 -1008 7952 -992
rect 7990 -1008 8108 -992
rect 8162 -958 8280 -942
rect 8162 -992 8170 -958
rect 8204 -992 8238 -958
rect 8272 -992 8280 -958
rect 7918 -1058 7952 -1042
rect 7990 -1058 8108 -1042
rect 7762 -1092 7770 -1058
rect 7804 -1092 7838 -1058
rect 7872 -1092 7880 -1058
rect 7990 -1092 7998 -1058
rect 8032 -1092 8066 -1058
rect 8100 -1092 8108 -1058
rect 7762 -1108 7880 -1092
rect 7918 -1108 7952 -1092
rect 7362 -1192 7370 -1158
rect 7404 -1192 7438 -1158
rect 7472 -1192 7480 -1158
rect 7362 -1208 7480 -1192
rect 7590 -1158 7708 -1142
rect 7590 -1192 7598 -1158
rect 7632 -1192 7666 -1158
rect 7700 -1192 7708 -1158
rect 7118 -1258 7152 -1242
rect 7190 -1258 7308 -1242
rect 6962 -1292 6970 -1258
rect 7004 -1292 7038 -1258
rect 7072 -1292 7080 -1258
rect 7190 -1292 7198 -1258
rect 7232 -1292 7266 -1258
rect 7300 -1292 7308 -1258
rect 6962 -1358 7080 -1292
rect 7118 -1308 7152 -1292
rect 7190 -1308 7308 -1292
rect 7362 -1258 7480 -1242
rect 7362 -1292 7370 -1258
rect 7404 -1292 7438 -1258
rect 7472 -1292 7480 -1258
rect 7362 -1308 7480 -1292
rect 7590 -1258 7708 -1192
rect 7590 -1292 7598 -1258
rect 7632 -1292 7666 -1258
rect 7700 -1292 7708 -1258
rect 7590 -1308 7708 -1292
rect 7762 -1158 7880 -1142
rect 7918 -1158 7952 -1142
rect 7990 -1158 8108 -1092
rect 7762 -1192 7770 -1158
rect 7804 -1192 7838 -1158
rect 7872 -1192 7880 -1158
rect 7990 -1192 7998 -1158
rect 8032 -1192 8066 -1158
rect 8100 -1192 8108 -1158
rect 7762 -1258 7880 -1192
rect 7918 -1208 7952 -1192
rect 7990 -1208 8108 -1192
rect 8162 -1058 8280 -992
rect 8390 -958 8508 -892
rect 8562 -871 8568 -837
rect 8602 -858 8640 -837
rect 8562 -892 8570 -871
rect 8604 -892 8638 -858
rect 8674 -871 8680 -837
rect 8672 -892 8680 -871
rect 8790 -871 8796 -837
rect 8830 -858 8868 -837
rect 8790 -892 8798 -871
rect 8832 -892 8866 -858
rect 8902 -871 8908 -837
rect 8900 -892 8908 -871
rect 8562 -908 8680 -892
rect 8718 -908 8752 -892
rect 8390 -992 8398 -958
rect 8432 -992 8466 -958
rect 8500 -992 8508 -958
rect 8390 -1008 8508 -992
rect 8562 -958 8680 -942
rect 8718 -958 8752 -942
rect 8790 -958 8908 -892
rect 8962 -871 8968 -837
rect 9002 -858 9040 -837
rect 8962 -892 8970 -871
rect 9004 -892 9038 -858
rect 9074 -871 9080 -837
rect 9072 -892 9080 -871
rect 8962 -908 9080 -892
rect 9190 -871 9196 -837
rect 9230 -858 9268 -837
rect 9190 -892 9198 -871
rect 9232 -892 9266 -858
rect 9302 -871 9308 -837
rect 9300 -892 9308 -871
rect 8562 -992 8570 -958
rect 8604 -992 8638 -958
rect 8672 -992 8680 -958
rect 8790 -992 8798 -958
rect 8832 -992 8866 -958
rect 8900 -992 8908 -958
rect 8162 -1092 8170 -1058
rect 8204 -1092 8238 -1058
rect 8272 -1092 8280 -1058
rect 8162 -1158 8280 -1092
rect 8390 -1058 8508 -1042
rect 8390 -1092 8398 -1058
rect 8432 -1092 8466 -1058
rect 8500 -1092 8508 -1058
rect 8390 -1108 8508 -1092
rect 8562 -1058 8680 -992
rect 8718 -1008 8752 -992
rect 8790 -1008 8908 -992
rect 8962 -958 9080 -942
rect 8962 -992 8970 -958
rect 9004 -992 9038 -958
rect 9072 -992 9080 -958
rect 8718 -1058 8752 -1042
rect 8790 -1058 8908 -1042
rect 8562 -1092 8570 -1058
rect 8604 -1092 8638 -1058
rect 8672 -1092 8680 -1058
rect 8790 -1092 8798 -1058
rect 8832 -1092 8866 -1058
rect 8900 -1092 8908 -1058
rect 8562 -1108 8680 -1092
rect 8718 -1108 8752 -1092
rect 8162 -1192 8170 -1158
rect 8204 -1192 8238 -1158
rect 8272 -1192 8280 -1158
rect 8162 -1208 8280 -1192
rect 8390 -1158 8508 -1142
rect 8390 -1192 8398 -1158
rect 8432 -1192 8466 -1158
rect 8500 -1192 8508 -1158
rect 7918 -1258 7952 -1242
rect 7990 -1258 8108 -1242
rect 7762 -1292 7770 -1258
rect 7804 -1292 7838 -1258
rect 7872 -1292 7880 -1258
rect 7990 -1292 7998 -1258
rect 8032 -1292 8066 -1258
rect 8100 -1292 8108 -1258
rect 7762 -1308 7880 -1292
rect 7918 -1308 7952 -1292
rect 7118 -1358 7152 -1342
rect 7190 -1358 7308 -1342
rect 6962 -1392 6970 -1358
rect 7004 -1392 7038 -1358
rect 7072 -1392 7080 -1358
rect 7190 -1392 7198 -1358
rect 7232 -1392 7266 -1358
rect 7300 -1392 7308 -1358
rect 6962 -1408 7080 -1392
rect 7118 -1408 7152 -1392
rect 6318 -1458 6352 -1442
rect 6390 -1458 6508 -1442
rect 6162 -1492 6170 -1458
rect 6204 -1492 6238 -1458
rect 6272 -1492 6280 -1458
rect 6390 -1492 6398 -1458
rect 6432 -1492 6466 -1458
rect 6500 -1492 6508 -1458
rect 6162 -1508 6280 -1492
rect 6318 -1508 6352 -1492
rect 4718 -1558 4752 -1542
rect 4790 -1558 4908 -1542
rect 4562 -1592 4570 -1558
rect 4604 -1592 4638 -1558
rect 4672 -1592 4680 -1558
rect 4790 -1592 4798 -1558
rect 4832 -1592 4866 -1558
rect 4900 -1592 4908 -1558
rect 4562 -1608 4680 -1592
rect 4718 -1608 4752 -1592
rect 3118 -1658 3152 -1642
rect 3190 -1658 3308 -1642
rect 2962 -1692 2970 -1658
rect 3004 -1692 3038 -1658
rect 3072 -1692 3080 -1658
rect 3190 -1692 3198 -1658
rect 3232 -1692 3266 -1658
rect 3300 -1692 3308 -1658
rect 2962 -1758 3080 -1692
rect 3118 -1708 3152 -1692
rect 3190 -1708 3308 -1692
rect 3362 -1658 3480 -1642
rect 3362 -1692 3370 -1658
rect 3404 -1692 3438 -1658
rect 3472 -1692 3480 -1658
rect 3362 -1708 3480 -1692
rect 3590 -1658 3708 -1642
rect 3590 -1692 3598 -1658
rect 3632 -1692 3666 -1658
rect 3700 -1692 3708 -1658
rect 3590 -1708 3708 -1692
rect 3762 -1658 3880 -1642
rect 3918 -1658 3952 -1642
rect 3990 -1658 4108 -1642
rect 3762 -1692 3770 -1658
rect 3804 -1692 3838 -1658
rect 3872 -1692 3880 -1658
rect 3990 -1692 3998 -1658
rect 4032 -1692 4066 -1658
rect 4100 -1692 4108 -1658
rect 3762 -1708 3880 -1692
rect 3918 -1708 3952 -1692
rect 3990 -1708 4108 -1692
rect 4162 -1658 4280 -1642
rect 4162 -1692 4170 -1658
rect 4204 -1692 4238 -1658
rect 4272 -1692 4280 -1658
rect 4162 -1708 4280 -1692
rect 4390 -1658 4508 -1642
rect 4390 -1692 4398 -1658
rect 4432 -1692 4466 -1658
rect 4500 -1692 4508 -1658
rect 4390 -1708 4508 -1692
rect 4562 -1658 4680 -1642
rect 4718 -1658 4752 -1642
rect 4790 -1658 4908 -1592
rect 4562 -1692 4570 -1658
rect 4604 -1692 4638 -1658
rect 4672 -1692 4680 -1658
rect 4790 -1692 4798 -1658
rect 4832 -1692 4866 -1658
rect 4900 -1692 4908 -1658
rect 4562 -1708 4680 -1692
rect 4718 -1708 4752 -1692
rect 4790 -1708 4908 -1692
rect 4962 -1558 5080 -1542
rect 4962 -1592 4970 -1558
rect 5004 -1592 5038 -1558
rect 5072 -1592 5080 -1558
rect 4962 -1658 5080 -1592
rect 4962 -1692 4970 -1658
rect 5004 -1692 5038 -1658
rect 5072 -1692 5080 -1658
rect 4962 -1708 5080 -1692
rect 5190 -1558 5308 -1542
rect 5190 -1592 5198 -1558
rect 5232 -1592 5266 -1558
rect 5300 -1592 5308 -1558
rect 5190 -1658 5308 -1592
rect 5190 -1692 5198 -1658
rect 5232 -1692 5266 -1658
rect 5300 -1692 5308 -1658
rect 5190 -1708 5308 -1692
rect 5362 -1558 5480 -1542
rect 5518 -1558 5552 -1542
rect 5590 -1558 5708 -1542
rect 5362 -1592 5370 -1558
rect 5404 -1592 5438 -1558
rect 5472 -1592 5480 -1558
rect 5590 -1592 5598 -1558
rect 5632 -1592 5666 -1558
rect 5700 -1592 5708 -1558
rect 5362 -1658 5480 -1592
rect 5518 -1608 5552 -1592
rect 5518 -1658 5552 -1642
rect 5590 -1658 5708 -1592
rect 5362 -1692 5370 -1658
rect 5404 -1692 5438 -1658
rect 5472 -1692 5480 -1658
rect 5590 -1692 5598 -1658
rect 5632 -1692 5666 -1658
rect 5700 -1692 5708 -1658
rect 5362 -1708 5480 -1692
rect 5518 -1708 5552 -1692
rect 5590 -1708 5708 -1692
rect 5762 -1558 5880 -1542
rect 5762 -1592 5770 -1558
rect 5804 -1592 5838 -1558
rect 5872 -1592 5880 -1558
rect 5762 -1658 5880 -1592
rect 5762 -1692 5770 -1658
rect 5804 -1692 5838 -1658
rect 5872 -1692 5880 -1658
rect 5762 -1708 5880 -1692
rect 5990 -1558 6108 -1542
rect 5990 -1592 5998 -1558
rect 6032 -1592 6066 -1558
rect 6100 -1592 6108 -1558
rect 5990 -1658 6108 -1592
rect 5990 -1692 5998 -1658
rect 6032 -1692 6066 -1658
rect 6100 -1692 6108 -1658
rect 5990 -1708 6108 -1692
rect 6162 -1558 6280 -1542
rect 6318 -1558 6352 -1542
rect 6390 -1558 6508 -1492
rect 6162 -1592 6170 -1558
rect 6204 -1592 6238 -1558
rect 6272 -1592 6280 -1558
rect 6390 -1592 6398 -1558
rect 6432 -1592 6466 -1558
rect 6500 -1592 6508 -1558
rect 6162 -1658 6280 -1592
rect 6318 -1608 6352 -1592
rect 6390 -1608 6508 -1592
rect 6562 -1458 6680 -1442
rect 6562 -1492 6570 -1458
rect 6604 -1492 6638 -1458
rect 6672 -1492 6680 -1458
rect 6562 -1558 6680 -1492
rect 6562 -1592 6570 -1558
rect 6604 -1592 6638 -1558
rect 6672 -1592 6680 -1558
rect 6562 -1608 6680 -1592
rect 6790 -1458 6908 -1442
rect 6790 -1492 6798 -1458
rect 6832 -1492 6866 -1458
rect 6900 -1492 6908 -1458
rect 6790 -1558 6908 -1492
rect 6790 -1592 6798 -1558
rect 6832 -1592 6866 -1558
rect 6900 -1592 6908 -1558
rect 6790 -1608 6908 -1592
rect 6962 -1458 7080 -1442
rect 7118 -1458 7152 -1442
rect 7190 -1458 7308 -1392
rect 6962 -1492 6970 -1458
rect 7004 -1492 7038 -1458
rect 7072 -1492 7080 -1458
rect 7190 -1492 7198 -1458
rect 7232 -1492 7266 -1458
rect 7300 -1492 7308 -1458
rect 6962 -1558 7080 -1492
rect 7118 -1508 7152 -1492
rect 7118 -1558 7152 -1542
rect 7190 -1558 7308 -1492
rect 6962 -1592 6970 -1558
rect 7004 -1592 7038 -1558
rect 7072 -1592 7080 -1558
rect 7190 -1592 7198 -1558
rect 7232 -1592 7266 -1558
rect 7300 -1592 7308 -1558
rect 6962 -1608 7080 -1592
rect 7118 -1608 7152 -1592
rect 7190 -1608 7308 -1592
rect 7362 -1358 7480 -1342
rect 7362 -1392 7370 -1358
rect 7404 -1392 7438 -1358
rect 7472 -1392 7480 -1358
rect 7362 -1458 7480 -1392
rect 7362 -1492 7370 -1458
rect 7404 -1492 7438 -1458
rect 7472 -1492 7480 -1458
rect 7362 -1558 7480 -1492
rect 7362 -1592 7370 -1558
rect 7404 -1592 7438 -1558
rect 7472 -1592 7480 -1558
rect 7362 -1608 7480 -1592
rect 7590 -1358 7708 -1342
rect 7590 -1392 7598 -1358
rect 7632 -1392 7666 -1358
rect 7700 -1392 7708 -1358
rect 7590 -1458 7708 -1392
rect 7590 -1492 7598 -1458
rect 7632 -1492 7666 -1458
rect 7700 -1492 7708 -1458
rect 7590 -1558 7708 -1492
rect 7590 -1592 7598 -1558
rect 7632 -1592 7666 -1558
rect 7700 -1592 7708 -1558
rect 7590 -1608 7708 -1592
rect 7762 -1358 7880 -1342
rect 7918 -1358 7952 -1342
rect 7990 -1358 8108 -1292
rect 7762 -1392 7770 -1358
rect 7804 -1392 7838 -1358
rect 7872 -1392 7880 -1358
rect 7990 -1392 7998 -1358
rect 8032 -1392 8066 -1358
rect 8100 -1392 8108 -1358
rect 7762 -1458 7880 -1392
rect 7918 -1408 7952 -1392
rect 7990 -1408 8108 -1392
rect 8162 -1258 8280 -1242
rect 8162 -1292 8170 -1258
rect 8204 -1292 8238 -1258
rect 8272 -1292 8280 -1258
rect 8162 -1358 8280 -1292
rect 8162 -1392 8170 -1358
rect 8204 -1392 8238 -1358
rect 8272 -1392 8280 -1358
rect 8162 -1408 8280 -1392
rect 8390 -1258 8508 -1192
rect 8390 -1292 8398 -1258
rect 8432 -1292 8466 -1258
rect 8500 -1292 8508 -1258
rect 8390 -1358 8508 -1292
rect 8390 -1392 8398 -1358
rect 8432 -1392 8466 -1358
rect 8500 -1392 8508 -1358
rect 8390 -1408 8508 -1392
rect 8562 -1158 8680 -1142
rect 8718 -1158 8752 -1142
rect 8790 -1158 8908 -1092
rect 8562 -1192 8570 -1158
rect 8604 -1192 8638 -1158
rect 8672 -1192 8680 -1158
rect 8790 -1192 8798 -1158
rect 8832 -1192 8866 -1158
rect 8900 -1192 8908 -1158
rect 8562 -1258 8680 -1192
rect 8718 -1208 8752 -1192
rect 8790 -1208 8908 -1192
rect 8962 -1058 9080 -992
rect 9190 -958 9308 -892
rect 9362 -871 9368 -837
rect 9402 -858 9440 -837
rect 9362 -892 9370 -871
rect 9404 -892 9438 -858
rect 9474 -871 9480 -837
rect 9472 -892 9480 -871
rect 9590 -871 9596 -837
rect 9630 -858 9668 -837
rect 9590 -892 9598 -871
rect 9632 -892 9666 -858
rect 9702 -871 9708 -837
rect 9700 -892 9708 -871
rect 9362 -908 9480 -892
rect 9518 -908 9552 -892
rect 9190 -992 9198 -958
rect 9232 -992 9266 -958
rect 9300 -992 9308 -958
rect 9190 -1008 9308 -992
rect 9362 -958 9480 -942
rect 9518 -958 9552 -942
rect 9590 -958 9708 -892
rect 9762 -871 9768 -837
rect 9802 -858 9840 -837
rect 9762 -892 9770 -871
rect 9804 -892 9838 -858
rect 9874 -871 9880 -837
rect 9872 -892 9880 -871
rect 9762 -908 9880 -892
rect 9990 -871 9996 -837
rect 10030 -858 10068 -837
rect 9990 -892 9998 -871
rect 10032 -892 10066 -858
rect 10102 -871 10108 -837
rect 10100 -892 10108 -871
rect 9362 -992 9370 -958
rect 9404 -992 9438 -958
rect 9472 -992 9480 -958
rect 9590 -992 9598 -958
rect 9632 -992 9666 -958
rect 9700 -992 9708 -958
rect 8962 -1092 8970 -1058
rect 9004 -1092 9038 -1058
rect 9072 -1092 9080 -1058
rect 8962 -1158 9080 -1092
rect 9190 -1058 9308 -1042
rect 9190 -1092 9198 -1058
rect 9232 -1092 9266 -1058
rect 9300 -1092 9308 -1058
rect 9190 -1108 9308 -1092
rect 9362 -1058 9480 -992
rect 9518 -1008 9552 -992
rect 9590 -1008 9708 -992
rect 9762 -958 9880 -942
rect 9762 -992 9770 -958
rect 9804 -992 9838 -958
rect 9872 -992 9880 -958
rect 9518 -1058 9552 -1042
rect 9590 -1058 9708 -1042
rect 9362 -1092 9370 -1058
rect 9404 -1092 9438 -1058
rect 9472 -1092 9480 -1058
rect 9590 -1092 9598 -1058
rect 9632 -1092 9666 -1058
rect 9700 -1092 9708 -1058
rect 9362 -1108 9480 -1092
rect 9518 -1108 9552 -1092
rect 8962 -1192 8970 -1158
rect 9004 -1192 9038 -1158
rect 9072 -1192 9080 -1158
rect 8962 -1208 9080 -1192
rect 9190 -1158 9308 -1142
rect 9190 -1192 9198 -1158
rect 9232 -1192 9266 -1158
rect 9300 -1192 9308 -1158
rect 8718 -1258 8752 -1242
rect 8790 -1258 8908 -1242
rect 8562 -1292 8570 -1258
rect 8604 -1292 8638 -1258
rect 8672 -1292 8680 -1258
rect 8790 -1292 8798 -1258
rect 8832 -1292 8866 -1258
rect 8900 -1292 8908 -1258
rect 8562 -1358 8680 -1292
rect 8718 -1308 8752 -1292
rect 8790 -1308 8908 -1292
rect 8962 -1258 9080 -1242
rect 8962 -1292 8970 -1258
rect 9004 -1292 9038 -1258
rect 9072 -1292 9080 -1258
rect 8962 -1308 9080 -1292
rect 9190 -1258 9308 -1192
rect 9190 -1292 9198 -1258
rect 9232 -1292 9266 -1258
rect 9300 -1292 9308 -1258
rect 9190 -1308 9308 -1292
rect 9362 -1158 9480 -1142
rect 9518 -1158 9552 -1142
rect 9590 -1158 9708 -1092
rect 9362 -1192 9370 -1158
rect 9404 -1192 9438 -1158
rect 9472 -1192 9480 -1158
rect 9590 -1192 9598 -1158
rect 9632 -1192 9666 -1158
rect 9700 -1192 9708 -1158
rect 9362 -1258 9480 -1192
rect 9518 -1208 9552 -1192
rect 9590 -1208 9708 -1192
rect 9762 -1058 9880 -992
rect 9990 -958 10108 -892
rect 10162 -871 10168 -837
rect 10202 -858 10240 -837
rect 10162 -892 10170 -871
rect 10204 -892 10238 -858
rect 10274 -871 10280 -837
rect 10272 -892 10280 -871
rect 10390 -871 10396 -837
rect 10430 -858 10468 -837
rect 10390 -892 10398 -871
rect 10432 -892 10466 -858
rect 10502 -871 10508 -837
rect 10500 -892 10508 -871
rect 10162 -908 10280 -892
rect 10318 -908 10352 -892
rect 9990 -992 9998 -958
rect 10032 -992 10066 -958
rect 10100 -992 10108 -958
rect 9990 -1008 10108 -992
rect 10162 -958 10280 -942
rect 10318 -958 10352 -942
rect 10390 -958 10508 -892
rect 10562 -871 10568 -837
rect 10602 -858 10640 -837
rect 10562 -892 10570 -871
rect 10604 -892 10638 -858
rect 10674 -871 10680 -837
rect 10672 -892 10680 -871
rect 10562 -908 10680 -892
rect 10790 -871 10796 -837
rect 10830 -858 10868 -837
rect 10790 -892 10798 -871
rect 10832 -892 10866 -858
rect 10902 -871 10908 -837
rect 10900 -892 10908 -871
rect 10162 -992 10170 -958
rect 10204 -992 10238 -958
rect 10272 -992 10280 -958
rect 10390 -992 10398 -958
rect 10432 -992 10466 -958
rect 10500 -992 10508 -958
rect 9762 -1092 9770 -1058
rect 9804 -1092 9838 -1058
rect 9872 -1092 9880 -1058
rect 9762 -1158 9880 -1092
rect 9990 -1058 10108 -1042
rect 9990 -1092 9998 -1058
rect 10032 -1092 10066 -1058
rect 10100 -1092 10108 -1058
rect 9990 -1108 10108 -1092
rect 10162 -1058 10280 -992
rect 10318 -1008 10352 -992
rect 10390 -1008 10508 -992
rect 10562 -958 10680 -942
rect 10562 -992 10570 -958
rect 10604 -992 10638 -958
rect 10672 -992 10680 -958
rect 10318 -1058 10352 -1042
rect 10390 -1058 10508 -1042
rect 10162 -1092 10170 -1058
rect 10204 -1092 10238 -1058
rect 10272 -1092 10280 -1058
rect 10390 -1092 10398 -1058
rect 10432 -1092 10466 -1058
rect 10500 -1092 10508 -1058
rect 10162 -1108 10280 -1092
rect 10318 -1108 10352 -1092
rect 9762 -1192 9770 -1158
rect 9804 -1192 9838 -1158
rect 9872 -1192 9880 -1158
rect 9762 -1208 9880 -1192
rect 9990 -1158 10108 -1142
rect 9990 -1192 9998 -1158
rect 10032 -1192 10066 -1158
rect 10100 -1192 10108 -1158
rect 9518 -1258 9552 -1242
rect 9590 -1258 9708 -1242
rect 9362 -1292 9370 -1258
rect 9404 -1292 9438 -1258
rect 9472 -1292 9480 -1258
rect 9590 -1292 9598 -1258
rect 9632 -1292 9666 -1258
rect 9700 -1292 9708 -1258
rect 9362 -1308 9480 -1292
rect 9518 -1308 9552 -1292
rect 8718 -1358 8752 -1342
rect 8790 -1358 8908 -1342
rect 8562 -1392 8570 -1358
rect 8604 -1392 8638 -1358
rect 8672 -1392 8680 -1358
rect 8790 -1392 8798 -1358
rect 8832 -1392 8866 -1358
rect 8900 -1392 8908 -1358
rect 8562 -1408 8680 -1392
rect 8718 -1408 8752 -1392
rect 7918 -1458 7952 -1442
rect 7990 -1458 8108 -1442
rect 7762 -1492 7770 -1458
rect 7804 -1492 7838 -1458
rect 7872 -1492 7880 -1458
rect 7990 -1492 7998 -1458
rect 8032 -1492 8066 -1458
rect 8100 -1492 8108 -1458
rect 7762 -1558 7880 -1492
rect 7918 -1508 7952 -1492
rect 7990 -1508 8108 -1492
rect 8162 -1458 8280 -1442
rect 8162 -1492 8170 -1458
rect 8204 -1492 8238 -1458
rect 8272 -1492 8280 -1458
rect 8162 -1508 8280 -1492
rect 8390 -1458 8508 -1442
rect 8390 -1492 8398 -1458
rect 8432 -1492 8466 -1458
rect 8500 -1492 8508 -1458
rect 8390 -1508 8508 -1492
rect 8562 -1458 8680 -1442
rect 8718 -1458 8752 -1442
rect 8790 -1458 8908 -1392
rect 8562 -1492 8570 -1458
rect 8604 -1492 8638 -1458
rect 8672 -1492 8680 -1458
rect 8790 -1492 8798 -1458
rect 8832 -1492 8866 -1458
rect 8900 -1492 8908 -1458
rect 8562 -1508 8680 -1492
rect 8718 -1508 8752 -1492
rect 8790 -1508 8908 -1492
rect 8962 -1358 9080 -1342
rect 8962 -1392 8970 -1358
rect 9004 -1392 9038 -1358
rect 9072 -1392 9080 -1358
rect 8962 -1458 9080 -1392
rect 8962 -1492 8970 -1458
rect 9004 -1492 9038 -1458
rect 9072 -1492 9080 -1458
rect 8962 -1508 9080 -1492
rect 9190 -1358 9308 -1342
rect 9190 -1392 9198 -1358
rect 9232 -1392 9266 -1358
rect 9300 -1392 9308 -1358
rect 9190 -1458 9308 -1392
rect 9190 -1492 9198 -1458
rect 9232 -1492 9266 -1458
rect 9300 -1492 9308 -1458
rect 9190 -1508 9308 -1492
rect 9362 -1358 9480 -1342
rect 9518 -1358 9552 -1342
rect 9590 -1358 9708 -1292
rect 9362 -1392 9370 -1358
rect 9404 -1392 9438 -1358
rect 9472 -1392 9480 -1358
rect 9590 -1392 9598 -1358
rect 9632 -1392 9666 -1358
rect 9700 -1392 9708 -1358
rect 9362 -1458 9480 -1392
rect 9518 -1408 9552 -1392
rect 9590 -1408 9708 -1392
rect 9762 -1258 9880 -1242
rect 9762 -1292 9770 -1258
rect 9804 -1292 9838 -1258
rect 9872 -1292 9880 -1258
rect 9762 -1358 9880 -1292
rect 9762 -1392 9770 -1358
rect 9804 -1392 9838 -1358
rect 9872 -1392 9880 -1358
rect 9762 -1408 9880 -1392
rect 9990 -1258 10108 -1192
rect 9990 -1292 9998 -1258
rect 10032 -1292 10066 -1258
rect 10100 -1292 10108 -1258
rect 9990 -1358 10108 -1292
rect 9990 -1392 9998 -1358
rect 10032 -1392 10066 -1358
rect 10100 -1392 10108 -1358
rect 9990 -1408 10108 -1392
rect 10162 -1158 10280 -1142
rect 10318 -1158 10352 -1142
rect 10390 -1158 10508 -1092
rect 10162 -1192 10170 -1158
rect 10204 -1192 10238 -1158
rect 10272 -1192 10280 -1158
rect 10390 -1192 10398 -1158
rect 10432 -1192 10466 -1158
rect 10500 -1192 10508 -1158
rect 10162 -1258 10280 -1192
rect 10318 -1208 10352 -1192
rect 10390 -1208 10508 -1192
rect 10562 -1058 10680 -992
rect 10790 -958 10908 -892
rect 10962 -871 10968 -837
rect 11002 -858 11040 -837
rect 10962 -892 10970 -871
rect 11004 -892 11038 -858
rect 11074 -871 11080 -837
rect 11072 -892 11080 -871
rect 11190 -871 11196 -837
rect 11230 -858 11268 -837
rect 11190 -892 11198 -871
rect 11232 -892 11266 -858
rect 11302 -871 11308 -837
rect 11300 -892 11308 -871
rect 10962 -908 11080 -892
rect 11118 -908 11152 -892
rect 10790 -992 10798 -958
rect 10832 -992 10866 -958
rect 10900 -992 10908 -958
rect 10790 -1008 10908 -992
rect 10962 -958 11080 -942
rect 11118 -958 11152 -942
rect 11190 -958 11308 -892
rect 11362 -871 11368 -837
rect 11402 -858 11440 -837
rect 11362 -892 11370 -871
rect 11404 -892 11438 -858
rect 11474 -871 11480 -837
rect 11472 -892 11480 -871
rect 11362 -908 11480 -892
rect 11590 -871 11596 -837
rect 11630 -858 11668 -837
rect 11590 -892 11598 -871
rect 11632 -892 11666 -858
rect 11702 -871 11708 -837
rect 11700 -892 11708 -871
rect 10962 -992 10970 -958
rect 11004 -992 11038 -958
rect 11072 -992 11080 -958
rect 11190 -992 11198 -958
rect 11232 -992 11266 -958
rect 11300 -992 11308 -958
rect 10562 -1092 10570 -1058
rect 10604 -1092 10638 -1058
rect 10672 -1092 10680 -1058
rect 10562 -1158 10680 -1092
rect 10790 -1058 10908 -1042
rect 10790 -1092 10798 -1058
rect 10832 -1092 10866 -1058
rect 10900 -1092 10908 -1058
rect 10790 -1108 10908 -1092
rect 10962 -1058 11080 -992
rect 11118 -1008 11152 -992
rect 11190 -1008 11308 -992
rect 11362 -958 11480 -942
rect 11362 -992 11370 -958
rect 11404 -992 11438 -958
rect 11472 -992 11480 -958
rect 11118 -1058 11152 -1042
rect 11190 -1058 11308 -1042
rect 10962 -1092 10970 -1058
rect 11004 -1092 11038 -1058
rect 11072 -1092 11080 -1058
rect 11190 -1092 11198 -1058
rect 11232 -1092 11266 -1058
rect 11300 -1092 11308 -1058
rect 10962 -1108 11080 -1092
rect 11118 -1108 11152 -1092
rect 10562 -1192 10570 -1158
rect 10604 -1192 10638 -1158
rect 10672 -1192 10680 -1158
rect 10562 -1208 10680 -1192
rect 10790 -1158 10908 -1142
rect 10790 -1192 10798 -1158
rect 10832 -1192 10866 -1158
rect 10900 -1192 10908 -1158
rect 10318 -1258 10352 -1242
rect 10390 -1258 10508 -1242
rect 10162 -1292 10170 -1258
rect 10204 -1292 10238 -1258
rect 10272 -1292 10280 -1258
rect 10390 -1292 10398 -1258
rect 10432 -1292 10466 -1258
rect 10500 -1292 10508 -1258
rect 10162 -1358 10280 -1292
rect 10318 -1308 10352 -1292
rect 10390 -1308 10508 -1292
rect 10562 -1258 10680 -1242
rect 10562 -1292 10570 -1258
rect 10604 -1292 10638 -1258
rect 10672 -1292 10680 -1258
rect 10562 -1308 10680 -1292
rect 10790 -1258 10908 -1192
rect 10790 -1292 10798 -1258
rect 10832 -1292 10866 -1258
rect 10900 -1292 10908 -1258
rect 10790 -1308 10908 -1292
rect 10962 -1158 11080 -1142
rect 11118 -1158 11152 -1142
rect 11190 -1158 11308 -1092
rect 10962 -1192 10970 -1158
rect 11004 -1192 11038 -1158
rect 11072 -1192 11080 -1158
rect 11190 -1192 11198 -1158
rect 11232 -1192 11266 -1158
rect 11300 -1192 11308 -1158
rect 10962 -1258 11080 -1192
rect 11118 -1208 11152 -1192
rect 11190 -1208 11308 -1192
rect 11362 -1058 11480 -992
rect 11590 -958 11708 -892
rect 11762 -871 11768 -837
rect 11802 -858 11840 -837
rect 11762 -892 11770 -871
rect 11804 -892 11838 -858
rect 11874 -871 11880 -837
rect 11872 -892 11880 -871
rect 11990 -871 11996 -837
rect 12030 -858 12068 -837
rect 11990 -892 11998 -871
rect 12032 -892 12066 -858
rect 12102 -871 12108 -837
rect 12100 -892 12108 -871
rect 11762 -908 11880 -892
rect 11918 -908 11952 -892
rect 11590 -992 11598 -958
rect 11632 -992 11666 -958
rect 11700 -992 11708 -958
rect 11590 -1008 11708 -992
rect 11762 -958 11880 -942
rect 11918 -958 11952 -942
rect 11990 -958 12108 -892
rect 12162 -871 12168 -837
rect 12202 -858 12240 -837
rect 12162 -892 12170 -871
rect 12204 -892 12238 -858
rect 12274 -871 12280 -837
rect 12272 -892 12280 -871
rect 12162 -908 12280 -892
rect 12390 -871 12396 -837
rect 12430 -858 12468 -837
rect 12390 -892 12398 -871
rect 12432 -892 12466 -858
rect 12502 -871 12508 -837
rect 12500 -892 12508 -871
rect 11762 -992 11770 -958
rect 11804 -992 11838 -958
rect 11872 -992 11880 -958
rect 11990 -992 11998 -958
rect 12032 -992 12066 -958
rect 12100 -992 12108 -958
rect 11362 -1092 11370 -1058
rect 11404 -1092 11438 -1058
rect 11472 -1092 11480 -1058
rect 11362 -1158 11480 -1092
rect 11590 -1058 11708 -1042
rect 11590 -1092 11598 -1058
rect 11632 -1092 11666 -1058
rect 11700 -1092 11708 -1058
rect 11590 -1108 11708 -1092
rect 11762 -1058 11880 -992
rect 11918 -1008 11952 -992
rect 11990 -1008 12108 -992
rect 12162 -958 12280 -942
rect 12162 -992 12170 -958
rect 12204 -992 12238 -958
rect 12272 -992 12280 -958
rect 11918 -1058 11952 -1042
rect 11990 -1058 12108 -1042
rect 11762 -1092 11770 -1058
rect 11804 -1092 11838 -1058
rect 11872 -1092 11880 -1058
rect 11990 -1092 11998 -1058
rect 12032 -1092 12066 -1058
rect 12100 -1092 12108 -1058
rect 11762 -1108 11880 -1092
rect 11918 -1108 11952 -1092
rect 11362 -1192 11370 -1158
rect 11404 -1192 11438 -1158
rect 11472 -1192 11480 -1158
rect 11362 -1208 11480 -1192
rect 11590 -1158 11708 -1142
rect 11590 -1192 11598 -1158
rect 11632 -1192 11666 -1158
rect 11700 -1192 11708 -1158
rect 11118 -1258 11152 -1242
rect 11190 -1258 11308 -1242
rect 10962 -1292 10970 -1258
rect 11004 -1292 11038 -1258
rect 11072 -1292 11080 -1258
rect 11190 -1292 11198 -1258
rect 11232 -1292 11266 -1258
rect 11300 -1292 11308 -1258
rect 10962 -1308 11080 -1292
rect 11118 -1308 11152 -1292
rect 10318 -1358 10352 -1342
rect 10390 -1358 10508 -1342
rect 10162 -1392 10170 -1358
rect 10204 -1392 10238 -1358
rect 10272 -1392 10280 -1358
rect 10390 -1392 10398 -1358
rect 10432 -1392 10466 -1358
rect 10500 -1392 10508 -1358
rect 10162 -1408 10280 -1392
rect 10318 -1408 10352 -1392
rect 9518 -1458 9552 -1442
rect 9590 -1458 9708 -1442
rect 9362 -1492 9370 -1458
rect 9404 -1492 9438 -1458
rect 9472 -1492 9480 -1458
rect 9590 -1492 9598 -1458
rect 9632 -1492 9666 -1458
rect 9700 -1492 9708 -1458
rect 9362 -1508 9480 -1492
rect 9518 -1508 9552 -1492
rect 7918 -1558 7952 -1542
rect 7990 -1558 8108 -1542
rect 7762 -1592 7770 -1558
rect 7804 -1592 7838 -1558
rect 7872 -1592 7880 -1558
rect 7990 -1592 7998 -1558
rect 8032 -1592 8066 -1558
rect 8100 -1592 8108 -1558
rect 7762 -1608 7880 -1592
rect 7918 -1608 7952 -1592
rect 6318 -1658 6352 -1642
rect 6390 -1658 6508 -1642
rect 6162 -1692 6170 -1658
rect 6204 -1692 6238 -1658
rect 6272 -1692 6280 -1658
rect 6390 -1692 6398 -1658
rect 6432 -1692 6466 -1658
rect 6500 -1692 6508 -1658
rect 6162 -1708 6280 -1692
rect 6318 -1708 6352 -1692
rect 3118 -1758 3152 -1742
rect 3190 -1758 3308 -1742
rect 2962 -1792 2970 -1758
rect 3004 -1792 3038 -1758
rect 3072 -1792 3080 -1758
rect 3190 -1792 3198 -1758
rect 3232 -1792 3266 -1758
rect 3300 -1792 3308 -1758
rect 2962 -1808 3080 -1792
rect 3118 -1808 3152 -1792
rect -82 -1858 -48 -1842
rect -10 -1858 108 -1842
rect -10 -1892 -2 -1858
rect 32 -1892 66 -1858
rect 100 -1892 108 -1858
rect -82 -1908 -48 -1892
rect -82 -1958 -48 -1942
rect -10 -1958 108 -1892
rect -10 -1992 -2 -1958
rect 32 -1992 66 -1958
rect 100 -1992 108 -1958
rect -82 -2008 -48 -1992
rect -10 -2008 108 -1992
rect 162 -1858 280 -1842
rect 162 -1892 170 -1858
rect 204 -1892 238 -1858
rect 272 -1892 280 -1858
rect 162 -1958 280 -1892
rect 162 -1992 170 -1958
rect 204 -1992 238 -1958
rect 272 -1992 280 -1958
rect 162 -2008 280 -1992
rect 390 -1858 508 -1842
rect 390 -1892 398 -1858
rect 432 -1892 466 -1858
rect 500 -1892 508 -1858
rect 390 -1958 508 -1892
rect 390 -1992 398 -1958
rect 432 -1992 466 -1958
rect 500 -1992 508 -1958
rect 390 -2008 508 -1992
rect 562 -1858 680 -1842
rect 718 -1858 752 -1842
rect 790 -1858 908 -1842
rect 562 -1892 570 -1858
rect 604 -1892 638 -1858
rect 672 -1892 680 -1858
rect 790 -1892 798 -1858
rect 832 -1892 866 -1858
rect 900 -1892 908 -1858
rect 562 -1958 680 -1892
rect 718 -1908 752 -1892
rect 718 -1958 752 -1942
rect 790 -1958 908 -1892
rect 562 -1992 570 -1958
rect 604 -1992 638 -1958
rect 672 -1992 680 -1958
rect 790 -1992 798 -1958
rect 832 -1992 866 -1958
rect 900 -1992 908 -1958
rect 562 -2008 680 -1992
rect 718 -2008 752 -1992
rect 790 -2008 908 -1992
rect 962 -1858 1080 -1842
rect 962 -1892 970 -1858
rect 1004 -1892 1038 -1858
rect 1072 -1892 1080 -1858
rect 962 -1958 1080 -1892
rect 962 -1992 970 -1958
rect 1004 -1992 1038 -1958
rect 1072 -1992 1080 -1958
rect 962 -2008 1080 -1992
rect 1190 -1858 1308 -1842
rect 1190 -1892 1198 -1858
rect 1232 -1892 1266 -1858
rect 1300 -1892 1308 -1858
rect 1190 -1958 1308 -1892
rect 1190 -1992 1198 -1958
rect 1232 -1992 1266 -1958
rect 1300 -1992 1308 -1958
rect 1190 -2008 1308 -1992
rect 1362 -1858 1480 -1842
rect 1518 -1858 1552 -1842
rect 1590 -1858 1708 -1842
rect 1362 -1892 1370 -1858
rect 1404 -1892 1438 -1858
rect 1472 -1892 1480 -1858
rect 1590 -1892 1598 -1858
rect 1632 -1892 1666 -1858
rect 1700 -1892 1708 -1858
rect 1362 -1958 1480 -1892
rect 1518 -1908 1552 -1892
rect 1518 -1958 1552 -1942
rect 1590 -1958 1708 -1892
rect 1362 -1992 1370 -1958
rect 1404 -1992 1438 -1958
rect 1472 -1992 1480 -1958
rect 1590 -1992 1598 -1958
rect 1632 -1992 1666 -1958
rect 1700 -1992 1708 -1958
rect 1362 -2008 1480 -1992
rect 1518 -2008 1552 -1992
rect 1590 -2008 1708 -1992
rect 1762 -1858 1880 -1842
rect 1762 -1892 1770 -1858
rect 1804 -1892 1838 -1858
rect 1872 -1892 1880 -1858
rect 1762 -1958 1880 -1892
rect 1762 -1992 1770 -1958
rect 1804 -1992 1838 -1958
rect 1872 -1992 1880 -1958
rect 1762 -2008 1880 -1992
rect 1990 -1858 2108 -1842
rect 1990 -1892 1998 -1858
rect 2032 -1892 2066 -1858
rect 2100 -1892 2108 -1858
rect 1990 -1958 2108 -1892
rect 1990 -1992 1998 -1958
rect 2032 -1992 2066 -1958
rect 2100 -1992 2108 -1958
rect 1990 -2008 2108 -1992
rect 2162 -1858 2280 -1842
rect 2318 -1858 2352 -1842
rect 2390 -1858 2508 -1842
rect 2162 -1892 2170 -1858
rect 2204 -1892 2238 -1858
rect 2272 -1892 2280 -1858
rect 2390 -1892 2398 -1858
rect 2432 -1892 2466 -1858
rect 2500 -1892 2508 -1858
rect 2162 -1958 2280 -1892
rect 2318 -1908 2352 -1892
rect 2318 -1958 2352 -1942
rect 2390 -1958 2508 -1892
rect 2162 -1992 2170 -1958
rect 2204 -1992 2238 -1958
rect 2272 -1992 2280 -1958
rect 2390 -1992 2398 -1958
rect 2432 -1992 2466 -1958
rect 2500 -1992 2508 -1958
rect 2162 -2008 2280 -1992
rect 2318 -2008 2352 -1992
rect 2390 -2008 2508 -1992
rect 2562 -1858 2680 -1842
rect 2562 -1892 2570 -1858
rect 2604 -1892 2638 -1858
rect 2672 -1892 2680 -1858
rect 2562 -1958 2680 -1892
rect 2562 -1992 2570 -1958
rect 2604 -1992 2638 -1958
rect 2672 -1992 2680 -1958
rect 2562 -2008 2680 -1992
rect 2790 -1858 2908 -1842
rect 2790 -1892 2798 -1858
rect 2832 -1892 2866 -1858
rect 2900 -1892 2908 -1858
rect 2790 -1958 2908 -1892
rect 2790 -1992 2798 -1958
rect 2832 -1992 2866 -1958
rect 2900 -1992 2908 -1958
rect 2790 -2008 2908 -1992
rect 2962 -1858 3080 -1842
rect 3118 -1858 3152 -1842
rect 3190 -1858 3308 -1792
rect 2962 -1892 2970 -1858
rect 3004 -1892 3038 -1858
rect 3072 -1892 3080 -1858
rect 3190 -1892 3198 -1858
rect 3232 -1892 3266 -1858
rect 3300 -1892 3308 -1858
rect 2962 -1958 3080 -1892
rect 3118 -1908 3152 -1892
rect 3118 -1958 3152 -1942
rect 3190 -1958 3308 -1892
rect 2962 -1992 2970 -1958
rect 3004 -1992 3038 -1958
rect 3072 -1992 3080 -1958
rect 3190 -1992 3198 -1958
rect 3232 -1992 3266 -1958
rect 3300 -1992 3308 -1958
rect 2962 -2008 3080 -1992
rect 3118 -2008 3152 -1992
rect 3190 -2008 3308 -1992
rect 3362 -1758 3480 -1742
rect 3362 -1792 3370 -1758
rect 3404 -1792 3438 -1758
rect 3472 -1792 3480 -1758
rect 3362 -1858 3480 -1792
rect 3362 -1892 3370 -1858
rect 3404 -1892 3438 -1858
rect 3472 -1892 3480 -1858
rect 3362 -1958 3480 -1892
rect 3362 -1992 3370 -1958
rect 3404 -1992 3438 -1958
rect 3472 -1992 3480 -1958
rect 3362 -2008 3480 -1992
rect 3590 -1758 3708 -1742
rect 3590 -1792 3598 -1758
rect 3632 -1792 3666 -1758
rect 3700 -1792 3708 -1758
rect 3590 -1858 3708 -1792
rect 3590 -1892 3598 -1858
rect 3632 -1892 3666 -1858
rect 3700 -1892 3708 -1858
rect 3590 -1958 3708 -1892
rect 3590 -1992 3598 -1958
rect 3632 -1992 3666 -1958
rect 3700 -1992 3708 -1958
rect 3590 -2008 3708 -1992
rect 3762 -1758 3880 -1742
rect 3918 -1758 3952 -1742
rect 3990 -1758 4108 -1742
rect 3762 -1792 3770 -1758
rect 3804 -1792 3838 -1758
rect 3872 -1792 3880 -1758
rect 3990 -1792 3998 -1758
rect 4032 -1792 4066 -1758
rect 4100 -1792 4108 -1758
rect 3762 -1858 3880 -1792
rect 3918 -1808 3952 -1792
rect 3918 -1858 3952 -1842
rect 3990 -1858 4108 -1792
rect 3762 -1892 3770 -1858
rect 3804 -1892 3838 -1858
rect 3872 -1892 3880 -1858
rect 3990 -1892 3998 -1858
rect 4032 -1892 4066 -1858
rect 4100 -1892 4108 -1858
rect 3762 -1958 3880 -1892
rect 3918 -1908 3952 -1892
rect 3918 -1958 3952 -1942
rect 3990 -1958 4108 -1892
rect 3762 -1992 3770 -1958
rect 3804 -1992 3838 -1958
rect 3872 -1992 3880 -1958
rect 3990 -1992 3998 -1958
rect 4032 -1992 4066 -1958
rect 4100 -1992 4108 -1958
rect 3762 -2008 3880 -1992
rect 3918 -2008 3952 -1992
rect 3990 -2008 4108 -1992
rect 4162 -1758 4280 -1742
rect 4162 -1792 4170 -1758
rect 4204 -1792 4238 -1758
rect 4272 -1792 4280 -1758
rect 4162 -1858 4280 -1792
rect 4162 -1892 4170 -1858
rect 4204 -1892 4238 -1858
rect 4272 -1892 4280 -1858
rect 4162 -1958 4280 -1892
rect 4162 -1992 4170 -1958
rect 4204 -1992 4238 -1958
rect 4272 -1992 4280 -1958
rect 4162 -2008 4280 -1992
rect 4390 -1758 4508 -1742
rect 4390 -1792 4398 -1758
rect 4432 -1792 4466 -1758
rect 4500 -1792 4508 -1758
rect 4390 -1858 4508 -1792
rect 4390 -1892 4398 -1858
rect 4432 -1892 4466 -1858
rect 4500 -1892 4508 -1858
rect 4390 -1958 4508 -1892
rect 4390 -1992 4398 -1958
rect 4432 -1992 4466 -1958
rect 4500 -1992 4508 -1958
rect 4390 -2008 4508 -1992
rect 4562 -1758 4680 -1742
rect 4718 -1758 4752 -1742
rect 4790 -1758 4908 -1742
rect 4562 -1792 4570 -1758
rect 4604 -1792 4638 -1758
rect 4672 -1792 4680 -1758
rect 4790 -1792 4798 -1758
rect 4832 -1792 4866 -1758
rect 4900 -1792 4908 -1758
rect 4562 -1858 4680 -1792
rect 4718 -1808 4752 -1792
rect 4718 -1858 4752 -1842
rect 4790 -1858 4908 -1792
rect 4562 -1892 4570 -1858
rect 4604 -1892 4638 -1858
rect 4672 -1892 4680 -1858
rect 4790 -1892 4798 -1858
rect 4832 -1892 4866 -1858
rect 4900 -1892 4908 -1858
rect 4562 -1958 4680 -1892
rect 4718 -1908 4752 -1892
rect 4718 -1958 4752 -1942
rect 4790 -1958 4908 -1892
rect 4562 -1992 4570 -1958
rect 4604 -1992 4638 -1958
rect 4672 -1992 4680 -1958
rect 4790 -1992 4798 -1958
rect 4832 -1992 4866 -1958
rect 4900 -1992 4908 -1958
rect 4562 -2008 4680 -1992
rect 4718 -2008 4752 -1992
rect 4790 -2008 4908 -1992
rect 4962 -1758 5080 -1742
rect 4962 -1792 4970 -1758
rect 5004 -1792 5038 -1758
rect 5072 -1792 5080 -1758
rect 4962 -1858 5080 -1792
rect 4962 -1892 4970 -1858
rect 5004 -1892 5038 -1858
rect 5072 -1892 5080 -1858
rect 4962 -1958 5080 -1892
rect 4962 -1992 4970 -1958
rect 5004 -1992 5038 -1958
rect 5072 -1992 5080 -1958
rect 4962 -2008 5080 -1992
rect 5190 -1758 5308 -1742
rect 5190 -1792 5198 -1758
rect 5232 -1792 5266 -1758
rect 5300 -1792 5308 -1758
rect 5190 -1858 5308 -1792
rect 5190 -1892 5198 -1858
rect 5232 -1892 5266 -1858
rect 5300 -1892 5308 -1858
rect 5190 -1958 5308 -1892
rect 5190 -1992 5198 -1958
rect 5232 -1992 5266 -1958
rect 5300 -1992 5308 -1958
rect 5190 -2008 5308 -1992
rect 5362 -1758 5480 -1742
rect 5518 -1758 5552 -1742
rect 5590 -1758 5708 -1742
rect 5362 -1792 5370 -1758
rect 5404 -1792 5438 -1758
rect 5472 -1792 5480 -1758
rect 5590 -1792 5598 -1758
rect 5632 -1792 5666 -1758
rect 5700 -1792 5708 -1758
rect 5362 -1858 5480 -1792
rect 5518 -1808 5552 -1792
rect 5518 -1858 5552 -1842
rect 5590 -1858 5708 -1792
rect 5362 -1892 5370 -1858
rect 5404 -1892 5438 -1858
rect 5472 -1892 5480 -1858
rect 5590 -1892 5598 -1858
rect 5632 -1892 5666 -1858
rect 5700 -1892 5708 -1858
rect 5362 -1958 5480 -1892
rect 5518 -1908 5552 -1892
rect 5518 -1958 5552 -1942
rect 5590 -1958 5708 -1892
rect 5362 -1992 5370 -1958
rect 5404 -1992 5438 -1958
rect 5472 -1992 5480 -1958
rect 5590 -1992 5598 -1958
rect 5632 -1992 5666 -1958
rect 5700 -1992 5708 -1958
rect 5362 -2008 5480 -1992
rect 5518 -2008 5552 -1992
rect 5590 -2008 5708 -1992
rect 5762 -1758 5880 -1742
rect 5762 -1792 5770 -1758
rect 5804 -1792 5838 -1758
rect 5872 -1792 5880 -1758
rect 5762 -1858 5880 -1792
rect 5762 -1892 5770 -1858
rect 5804 -1892 5838 -1858
rect 5872 -1892 5880 -1858
rect 5762 -1958 5880 -1892
rect 5762 -1992 5770 -1958
rect 5804 -1992 5838 -1958
rect 5872 -1992 5880 -1958
rect 5762 -2008 5880 -1992
rect 5990 -1758 6108 -1742
rect 5990 -1792 5998 -1758
rect 6032 -1792 6066 -1758
rect 6100 -1792 6108 -1758
rect 5990 -1858 6108 -1792
rect 5990 -1892 5998 -1858
rect 6032 -1892 6066 -1858
rect 6100 -1892 6108 -1858
rect 5990 -1958 6108 -1892
rect 5990 -1992 5998 -1958
rect 6032 -1992 6066 -1958
rect 6100 -1992 6108 -1958
rect 5990 -2008 6108 -1992
rect 6162 -1758 6280 -1742
rect 6318 -1758 6352 -1742
rect 6390 -1758 6508 -1692
rect 6162 -1792 6170 -1758
rect 6204 -1792 6238 -1758
rect 6272 -1792 6280 -1758
rect 6390 -1792 6398 -1758
rect 6432 -1792 6466 -1758
rect 6500 -1792 6508 -1758
rect 6162 -1858 6280 -1792
rect 6318 -1808 6352 -1792
rect 6390 -1808 6508 -1792
rect 6562 -1658 6680 -1642
rect 6562 -1692 6570 -1658
rect 6604 -1692 6638 -1658
rect 6672 -1692 6680 -1658
rect 6562 -1758 6680 -1692
rect 6562 -1792 6570 -1758
rect 6604 -1792 6638 -1758
rect 6672 -1792 6680 -1758
rect 6562 -1808 6680 -1792
rect 6790 -1658 6908 -1642
rect 6790 -1692 6798 -1658
rect 6832 -1692 6866 -1658
rect 6900 -1692 6908 -1658
rect 6790 -1758 6908 -1692
rect 6790 -1792 6798 -1758
rect 6832 -1792 6866 -1758
rect 6900 -1792 6908 -1758
rect 6790 -1808 6908 -1792
rect 6962 -1658 7080 -1642
rect 7118 -1658 7152 -1642
rect 7190 -1658 7308 -1642
rect 6962 -1692 6970 -1658
rect 7004 -1692 7038 -1658
rect 7072 -1692 7080 -1658
rect 7190 -1692 7198 -1658
rect 7232 -1692 7266 -1658
rect 7300 -1692 7308 -1658
rect 6962 -1758 7080 -1692
rect 7118 -1708 7152 -1692
rect 7118 -1758 7152 -1742
rect 7190 -1758 7308 -1692
rect 6962 -1792 6970 -1758
rect 7004 -1792 7038 -1758
rect 7072 -1792 7080 -1758
rect 7190 -1792 7198 -1758
rect 7232 -1792 7266 -1758
rect 7300 -1792 7308 -1758
rect 6962 -1808 7080 -1792
rect 7118 -1808 7152 -1792
rect 7190 -1808 7308 -1792
rect 7362 -1658 7480 -1642
rect 7362 -1692 7370 -1658
rect 7404 -1692 7438 -1658
rect 7472 -1692 7480 -1658
rect 7362 -1758 7480 -1692
rect 7362 -1792 7370 -1758
rect 7404 -1792 7438 -1758
rect 7472 -1792 7480 -1758
rect 7362 -1808 7480 -1792
rect 7590 -1658 7708 -1642
rect 7590 -1692 7598 -1658
rect 7632 -1692 7666 -1658
rect 7700 -1692 7708 -1658
rect 7590 -1758 7708 -1692
rect 7590 -1792 7598 -1758
rect 7632 -1792 7666 -1758
rect 7700 -1792 7708 -1758
rect 7590 -1808 7708 -1792
rect 7762 -1658 7880 -1642
rect 7918 -1658 7952 -1642
rect 7990 -1658 8108 -1592
rect 7762 -1692 7770 -1658
rect 7804 -1692 7838 -1658
rect 7872 -1692 7880 -1658
rect 7990 -1692 7998 -1658
rect 8032 -1692 8066 -1658
rect 8100 -1692 8108 -1658
rect 7762 -1758 7880 -1692
rect 7918 -1708 7952 -1692
rect 7918 -1758 7952 -1742
rect 7990 -1758 8108 -1692
rect 7762 -1792 7770 -1758
rect 7804 -1792 7838 -1758
rect 7872 -1792 7880 -1758
rect 7990 -1792 7998 -1758
rect 8032 -1792 8066 -1758
rect 8100 -1792 8108 -1758
rect 7762 -1808 7880 -1792
rect 7918 -1808 7952 -1792
rect 7990 -1808 8108 -1792
rect 8162 -1558 8280 -1542
rect 8162 -1592 8170 -1558
rect 8204 -1592 8238 -1558
rect 8272 -1592 8280 -1558
rect 8162 -1658 8280 -1592
rect 8162 -1692 8170 -1658
rect 8204 -1692 8238 -1658
rect 8272 -1692 8280 -1658
rect 8162 -1758 8280 -1692
rect 8162 -1792 8170 -1758
rect 8204 -1792 8238 -1758
rect 8272 -1792 8280 -1758
rect 8162 -1808 8280 -1792
rect 8390 -1558 8508 -1542
rect 8390 -1592 8398 -1558
rect 8432 -1592 8466 -1558
rect 8500 -1592 8508 -1558
rect 8390 -1658 8508 -1592
rect 8390 -1692 8398 -1658
rect 8432 -1692 8466 -1658
rect 8500 -1692 8508 -1658
rect 8390 -1758 8508 -1692
rect 8390 -1792 8398 -1758
rect 8432 -1792 8466 -1758
rect 8500 -1792 8508 -1758
rect 8390 -1808 8508 -1792
rect 8562 -1558 8680 -1542
rect 8718 -1558 8752 -1542
rect 8790 -1558 8908 -1542
rect 8562 -1592 8570 -1558
rect 8604 -1592 8638 -1558
rect 8672 -1592 8680 -1558
rect 8790 -1592 8798 -1558
rect 8832 -1592 8866 -1558
rect 8900 -1592 8908 -1558
rect 8562 -1658 8680 -1592
rect 8718 -1608 8752 -1592
rect 8718 -1658 8752 -1642
rect 8790 -1658 8908 -1592
rect 8562 -1692 8570 -1658
rect 8604 -1692 8638 -1658
rect 8672 -1692 8680 -1658
rect 8790 -1692 8798 -1658
rect 8832 -1692 8866 -1658
rect 8900 -1692 8908 -1658
rect 8562 -1758 8680 -1692
rect 8718 -1708 8752 -1692
rect 8718 -1758 8752 -1742
rect 8790 -1758 8908 -1692
rect 8562 -1792 8570 -1758
rect 8604 -1792 8638 -1758
rect 8672 -1792 8680 -1758
rect 8790 -1792 8798 -1758
rect 8832 -1792 8866 -1758
rect 8900 -1792 8908 -1758
rect 8562 -1808 8680 -1792
rect 8718 -1808 8752 -1792
rect 8790 -1808 8908 -1792
rect 8962 -1558 9080 -1542
rect 8962 -1592 8970 -1558
rect 9004 -1592 9038 -1558
rect 9072 -1592 9080 -1558
rect 8962 -1658 9080 -1592
rect 8962 -1692 8970 -1658
rect 9004 -1692 9038 -1658
rect 9072 -1692 9080 -1658
rect 8962 -1758 9080 -1692
rect 8962 -1792 8970 -1758
rect 9004 -1792 9038 -1758
rect 9072 -1792 9080 -1758
rect 8962 -1808 9080 -1792
rect 9190 -1558 9308 -1542
rect 9190 -1592 9198 -1558
rect 9232 -1592 9266 -1558
rect 9300 -1592 9308 -1558
rect 9190 -1658 9308 -1592
rect 9190 -1692 9198 -1658
rect 9232 -1692 9266 -1658
rect 9300 -1692 9308 -1658
rect 9190 -1758 9308 -1692
rect 9190 -1792 9198 -1758
rect 9232 -1792 9266 -1758
rect 9300 -1792 9308 -1758
rect 9190 -1808 9308 -1792
rect 9362 -1558 9480 -1542
rect 9518 -1558 9552 -1542
rect 9590 -1558 9708 -1492
rect 9362 -1592 9370 -1558
rect 9404 -1592 9438 -1558
rect 9472 -1592 9480 -1558
rect 9590 -1592 9598 -1558
rect 9632 -1592 9666 -1558
rect 9700 -1592 9708 -1558
rect 9362 -1658 9480 -1592
rect 9518 -1608 9552 -1592
rect 9590 -1608 9708 -1592
rect 9762 -1458 9880 -1442
rect 9762 -1492 9770 -1458
rect 9804 -1492 9838 -1458
rect 9872 -1492 9880 -1458
rect 9762 -1558 9880 -1492
rect 9762 -1592 9770 -1558
rect 9804 -1592 9838 -1558
rect 9872 -1592 9880 -1558
rect 9762 -1608 9880 -1592
rect 9990 -1458 10108 -1442
rect 9990 -1492 9998 -1458
rect 10032 -1492 10066 -1458
rect 10100 -1492 10108 -1458
rect 9990 -1558 10108 -1492
rect 9990 -1592 9998 -1558
rect 10032 -1592 10066 -1558
rect 10100 -1592 10108 -1558
rect 9990 -1608 10108 -1592
rect 10162 -1458 10280 -1442
rect 10318 -1458 10352 -1442
rect 10390 -1458 10508 -1392
rect 10162 -1492 10170 -1458
rect 10204 -1492 10238 -1458
rect 10272 -1492 10280 -1458
rect 10390 -1492 10398 -1458
rect 10432 -1492 10466 -1458
rect 10500 -1492 10508 -1458
rect 10162 -1558 10280 -1492
rect 10318 -1508 10352 -1492
rect 10318 -1558 10352 -1542
rect 10390 -1558 10508 -1492
rect 10162 -1592 10170 -1558
rect 10204 -1592 10238 -1558
rect 10272 -1592 10280 -1558
rect 10390 -1592 10398 -1558
rect 10432 -1592 10466 -1558
rect 10500 -1592 10508 -1558
rect 10162 -1608 10280 -1592
rect 10318 -1608 10352 -1592
rect 10390 -1608 10508 -1592
rect 10562 -1358 10680 -1342
rect 10562 -1392 10570 -1358
rect 10604 -1392 10638 -1358
rect 10672 -1392 10680 -1358
rect 10562 -1458 10680 -1392
rect 10562 -1492 10570 -1458
rect 10604 -1492 10638 -1458
rect 10672 -1492 10680 -1458
rect 10562 -1558 10680 -1492
rect 10562 -1592 10570 -1558
rect 10604 -1592 10638 -1558
rect 10672 -1592 10680 -1558
rect 10562 -1608 10680 -1592
rect 10790 -1358 10908 -1342
rect 10790 -1392 10798 -1358
rect 10832 -1392 10866 -1358
rect 10900 -1392 10908 -1358
rect 10790 -1458 10908 -1392
rect 10790 -1492 10798 -1458
rect 10832 -1492 10866 -1458
rect 10900 -1492 10908 -1458
rect 10790 -1558 10908 -1492
rect 10790 -1592 10798 -1558
rect 10832 -1592 10866 -1558
rect 10900 -1592 10908 -1558
rect 10790 -1608 10908 -1592
rect 10962 -1358 11080 -1342
rect 11118 -1358 11152 -1342
rect 11190 -1358 11308 -1292
rect 10962 -1392 10970 -1358
rect 11004 -1392 11038 -1358
rect 11072 -1392 11080 -1358
rect 11190 -1392 11198 -1358
rect 11232 -1392 11266 -1358
rect 11300 -1392 11308 -1358
rect 10962 -1458 11080 -1392
rect 11118 -1408 11152 -1392
rect 11190 -1408 11308 -1392
rect 11362 -1258 11480 -1242
rect 11362 -1292 11370 -1258
rect 11404 -1292 11438 -1258
rect 11472 -1292 11480 -1258
rect 11362 -1358 11480 -1292
rect 11362 -1392 11370 -1358
rect 11404 -1392 11438 -1358
rect 11472 -1392 11480 -1358
rect 11362 -1408 11480 -1392
rect 11590 -1258 11708 -1192
rect 11590 -1292 11598 -1258
rect 11632 -1292 11666 -1258
rect 11700 -1292 11708 -1258
rect 11590 -1358 11708 -1292
rect 11590 -1392 11598 -1358
rect 11632 -1392 11666 -1358
rect 11700 -1392 11708 -1358
rect 11590 -1408 11708 -1392
rect 11762 -1158 11880 -1142
rect 11918 -1158 11952 -1142
rect 11990 -1158 12108 -1092
rect 11762 -1192 11770 -1158
rect 11804 -1192 11838 -1158
rect 11872 -1192 11880 -1158
rect 11990 -1192 11998 -1158
rect 12032 -1192 12066 -1158
rect 12100 -1192 12108 -1158
rect 11762 -1258 11880 -1192
rect 11918 -1208 11952 -1192
rect 11990 -1208 12108 -1192
rect 12162 -1058 12280 -992
rect 12390 -958 12508 -892
rect 12562 -871 12568 -837
rect 12602 -858 12640 -837
rect 12562 -892 12570 -871
rect 12604 -892 12638 -858
rect 12674 -871 12680 -837
rect 14532 -842 14558 -808
rect 14596 -842 14630 -808
rect 14664 -842 14694 -808
rect 14808 -842 14842 -808
rect 14881 -842 14914 -808
rect 14949 -842 14983 -808
rect 15020 -842 15051 -808
rect 15092 -842 15124 -808
rect 15218 -842 15249 -808
rect 15291 -842 15321 -808
rect 15359 -842 15393 -808
rect 15427 -842 15461 -808
rect 15499 -842 15534 -808
rect 15648 -842 15677 -808
rect 15712 -842 15746 -808
rect 15783 -842 15810 -808
rect 12672 -892 12680 -871
rect 12562 -908 12680 -892
rect 12718 -908 12752 -892
rect 14532 -942 14560 -908
rect 14596 -942 14630 -908
rect 14666 -942 14694 -908
rect 14734 -909 14768 -892
rect 12390 -992 12398 -958
rect 12432 -992 12466 -958
rect 12500 -992 12508 -958
rect 12390 -1008 12508 -992
rect 12562 -958 12680 -942
rect 12718 -958 12752 -942
rect 14808 -942 14841 -908
rect 14881 -942 14913 -908
rect 14949 -942 14983 -908
rect 15019 -942 15051 -908
rect 15091 -942 15124 -908
rect 15218 -942 15251 -908
rect 15291 -942 15323 -908
rect 15359 -942 15393 -908
rect 15429 -942 15461 -908
rect 15501 -942 15534 -908
rect 15574 -909 15608 -892
rect 12562 -992 12570 -958
rect 12604 -992 12638 -958
rect 12672 -992 12680 -958
rect 12162 -1092 12170 -1058
rect 12204 -1092 12238 -1058
rect 12272 -1092 12280 -1058
rect 12162 -1158 12280 -1092
rect 12390 -1058 12508 -1042
rect 12390 -1092 12398 -1058
rect 12432 -1092 12466 -1058
rect 12500 -1092 12508 -1058
rect 12390 -1108 12508 -1092
rect 12562 -1058 12680 -992
rect 12718 -1008 12752 -992
rect 14734 -1008 14768 -943
rect 15648 -942 15676 -908
rect 15712 -942 15746 -908
rect 15782 -942 15810 -908
rect 15574 -1008 15608 -943
rect 14532 -1042 14558 -1008
rect 14596 -1042 14630 -1008
rect 14664 -1042 14694 -1008
rect 14808 -1042 14842 -1008
rect 14881 -1042 14914 -1008
rect 14949 -1042 14983 -1008
rect 15020 -1042 15051 -1008
rect 15092 -1042 15124 -1008
rect 15218 -1042 15249 -1008
rect 15291 -1042 15321 -1008
rect 15359 -1042 15393 -1008
rect 15427 -1042 15461 -1008
rect 15499 -1042 15534 -1008
rect 15648 -1042 15677 -1008
rect 15712 -1042 15746 -1008
rect 15783 -1042 15810 -1008
rect 12718 -1058 12752 -1042
rect 12562 -1092 12570 -1058
rect 12604 -1092 12638 -1058
rect 12672 -1092 12680 -1058
rect 12562 -1108 12680 -1092
rect 12718 -1108 12752 -1092
rect 14532 -1142 14560 -1108
rect 14596 -1142 14630 -1108
rect 14666 -1142 14694 -1108
rect 14734 -1109 14768 -1092
rect 12162 -1192 12170 -1158
rect 12204 -1192 12238 -1158
rect 12272 -1192 12280 -1158
rect 12162 -1208 12280 -1192
rect 12390 -1158 12508 -1142
rect 12390 -1192 12398 -1158
rect 12432 -1192 12466 -1158
rect 12500 -1192 12508 -1158
rect 11918 -1258 11952 -1242
rect 11990 -1258 12108 -1242
rect 11762 -1292 11770 -1258
rect 11804 -1292 11838 -1258
rect 11872 -1292 11880 -1258
rect 11990 -1292 11998 -1258
rect 12032 -1292 12066 -1258
rect 12100 -1292 12108 -1258
rect 11762 -1358 11880 -1292
rect 11918 -1308 11952 -1292
rect 11990 -1308 12108 -1292
rect 12162 -1258 12280 -1242
rect 12162 -1292 12170 -1258
rect 12204 -1292 12238 -1258
rect 12272 -1292 12280 -1258
rect 12162 -1308 12280 -1292
rect 12390 -1258 12508 -1192
rect 12390 -1292 12398 -1258
rect 12432 -1292 12466 -1258
rect 12500 -1292 12508 -1258
rect 12390 -1308 12508 -1292
rect 12562 -1158 12680 -1142
rect 12718 -1158 12752 -1142
rect 14808 -1142 14841 -1108
rect 14881 -1142 14913 -1108
rect 14949 -1142 14983 -1108
rect 15019 -1142 15051 -1108
rect 15091 -1142 15124 -1108
rect 15218 -1142 15251 -1108
rect 15291 -1142 15323 -1108
rect 15359 -1142 15393 -1108
rect 15429 -1142 15461 -1108
rect 15501 -1142 15534 -1108
rect 15574 -1109 15608 -1092
rect 12562 -1192 12570 -1158
rect 12604 -1192 12638 -1158
rect 12672 -1192 12680 -1158
rect 12562 -1258 12680 -1192
rect 12718 -1208 12752 -1192
rect 14734 -1208 14768 -1143
rect 15648 -1142 15676 -1108
rect 15712 -1142 15746 -1108
rect 15782 -1142 15810 -1108
rect 15574 -1208 15608 -1143
rect 14532 -1242 14558 -1208
rect 14596 -1242 14630 -1208
rect 14664 -1242 14694 -1208
rect 14808 -1242 14842 -1208
rect 14881 -1242 14914 -1208
rect 14949 -1242 14983 -1208
rect 15020 -1242 15051 -1208
rect 15092 -1242 15124 -1208
rect 15218 -1242 15249 -1208
rect 15291 -1242 15321 -1208
rect 15359 -1242 15393 -1208
rect 15427 -1242 15461 -1208
rect 15499 -1242 15534 -1208
rect 15648 -1242 15677 -1208
rect 15712 -1242 15746 -1208
rect 15783 -1242 15810 -1208
rect 12718 -1258 12752 -1242
rect 12562 -1292 12570 -1258
rect 12604 -1292 12638 -1258
rect 12672 -1292 12680 -1258
rect 12562 -1308 12680 -1292
rect 12718 -1308 12752 -1292
rect 14532 -1342 14560 -1308
rect 14596 -1342 14630 -1308
rect 14666 -1342 14694 -1308
rect 14734 -1309 14768 -1292
rect 11918 -1358 11952 -1342
rect 11990 -1358 12108 -1342
rect 11762 -1392 11770 -1358
rect 11804 -1392 11838 -1358
rect 11872 -1392 11880 -1358
rect 11990 -1392 11998 -1358
rect 12032 -1392 12066 -1358
rect 12100 -1392 12108 -1358
rect 11762 -1408 11880 -1392
rect 11918 -1408 11952 -1392
rect 11118 -1458 11152 -1442
rect 11190 -1458 11308 -1442
rect 10962 -1492 10970 -1458
rect 11004 -1492 11038 -1458
rect 11072 -1492 11080 -1458
rect 11190 -1492 11198 -1458
rect 11232 -1492 11266 -1458
rect 11300 -1492 11308 -1458
rect 10962 -1558 11080 -1492
rect 11118 -1508 11152 -1492
rect 11190 -1508 11308 -1492
rect 11362 -1458 11480 -1442
rect 11362 -1492 11370 -1458
rect 11404 -1492 11438 -1458
rect 11472 -1492 11480 -1458
rect 11362 -1508 11480 -1492
rect 11590 -1458 11708 -1442
rect 11590 -1492 11598 -1458
rect 11632 -1492 11666 -1458
rect 11700 -1492 11708 -1458
rect 11590 -1508 11708 -1492
rect 11762 -1458 11880 -1442
rect 11918 -1458 11952 -1442
rect 11990 -1458 12108 -1392
rect 11762 -1492 11770 -1458
rect 11804 -1492 11838 -1458
rect 11872 -1492 11880 -1458
rect 11990 -1492 11998 -1458
rect 12032 -1492 12066 -1458
rect 12100 -1492 12108 -1458
rect 11762 -1508 11880 -1492
rect 11918 -1508 11952 -1492
rect 11990 -1508 12108 -1492
rect 12162 -1358 12280 -1342
rect 12162 -1392 12170 -1358
rect 12204 -1392 12238 -1358
rect 12272 -1392 12280 -1358
rect 12162 -1458 12280 -1392
rect 12162 -1492 12170 -1458
rect 12204 -1492 12238 -1458
rect 12272 -1492 12280 -1458
rect 12162 -1508 12280 -1492
rect 12390 -1358 12508 -1342
rect 12390 -1392 12398 -1358
rect 12432 -1392 12466 -1358
rect 12500 -1392 12508 -1358
rect 12390 -1458 12508 -1392
rect 12390 -1492 12398 -1458
rect 12432 -1492 12466 -1458
rect 12500 -1492 12508 -1458
rect 12390 -1508 12508 -1492
rect 12562 -1358 12680 -1342
rect 12718 -1358 12752 -1342
rect 14808 -1342 14841 -1308
rect 14881 -1342 14913 -1308
rect 14949 -1342 14983 -1308
rect 15019 -1342 15051 -1308
rect 15091 -1342 15124 -1308
rect 15218 -1342 15251 -1308
rect 15291 -1342 15323 -1308
rect 15359 -1342 15393 -1308
rect 15429 -1342 15461 -1308
rect 15501 -1342 15534 -1308
rect 15574 -1309 15608 -1292
rect 12562 -1392 12570 -1358
rect 12604 -1392 12638 -1358
rect 12672 -1392 12680 -1358
rect 12562 -1458 12680 -1392
rect 12718 -1408 12752 -1392
rect 14734 -1408 14768 -1343
rect 15648 -1342 15676 -1308
rect 15712 -1342 15746 -1308
rect 15782 -1342 15810 -1308
rect 15574 -1408 15608 -1343
rect 14532 -1442 14558 -1408
rect 14596 -1442 14630 -1408
rect 14664 -1442 14694 -1408
rect 14808 -1442 14842 -1408
rect 14881 -1442 14914 -1408
rect 14949 -1442 14983 -1408
rect 15020 -1442 15051 -1408
rect 15092 -1442 15124 -1408
rect 15218 -1442 15249 -1408
rect 15291 -1442 15321 -1408
rect 15359 -1442 15393 -1408
rect 15427 -1442 15461 -1408
rect 15499 -1442 15534 -1408
rect 15648 -1442 15677 -1408
rect 15712 -1442 15746 -1408
rect 15783 -1442 15810 -1408
rect 12718 -1458 12752 -1442
rect 12562 -1492 12570 -1458
rect 12604 -1492 12638 -1458
rect 12672 -1492 12680 -1458
rect 12562 -1508 12680 -1492
rect 12718 -1508 12752 -1492
rect 14532 -1542 14560 -1508
rect 14596 -1542 14630 -1508
rect 14666 -1542 14694 -1508
rect 14734 -1509 14768 -1492
rect 11118 -1558 11152 -1542
rect 11190 -1558 11308 -1542
rect 10962 -1592 10970 -1558
rect 11004 -1592 11038 -1558
rect 11072 -1592 11080 -1558
rect 11190 -1592 11198 -1558
rect 11232 -1592 11266 -1558
rect 11300 -1592 11308 -1558
rect 10962 -1608 11080 -1592
rect 11118 -1608 11152 -1592
rect 9518 -1658 9552 -1642
rect 9590 -1658 9708 -1642
rect 9362 -1692 9370 -1658
rect 9404 -1692 9438 -1658
rect 9472 -1692 9480 -1658
rect 9590 -1692 9598 -1658
rect 9632 -1692 9666 -1658
rect 9700 -1692 9708 -1658
rect 9362 -1758 9480 -1692
rect 9518 -1708 9552 -1692
rect 9590 -1708 9708 -1692
rect 9762 -1658 9880 -1642
rect 9762 -1692 9770 -1658
rect 9804 -1692 9838 -1658
rect 9872 -1692 9880 -1658
rect 9762 -1708 9880 -1692
rect 9990 -1658 10108 -1642
rect 9990 -1692 9998 -1658
rect 10032 -1692 10066 -1658
rect 10100 -1692 10108 -1658
rect 9990 -1708 10108 -1692
rect 10162 -1658 10280 -1642
rect 10318 -1658 10352 -1642
rect 10390 -1658 10508 -1642
rect 10162 -1692 10170 -1658
rect 10204 -1692 10238 -1658
rect 10272 -1692 10280 -1658
rect 10390 -1692 10398 -1658
rect 10432 -1692 10466 -1658
rect 10500 -1692 10508 -1658
rect 10162 -1708 10280 -1692
rect 10318 -1708 10352 -1692
rect 10390 -1708 10508 -1692
rect 10562 -1658 10680 -1642
rect 10562 -1692 10570 -1658
rect 10604 -1692 10638 -1658
rect 10672 -1692 10680 -1658
rect 10562 -1708 10680 -1692
rect 10790 -1658 10908 -1642
rect 10790 -1692 10798 -1658
rect 10832 -1692 10866 -1658
rect 10900 -1692 10908 -1658
rect 10790 -1708 10908 -1692
rect 10962 -1658 11080 -1642
rect 11118 -1658 11152 -1642
rect 11190 -1658 11308 -1592
rect 10962 -1692 10970 -1658
rect 11004 -1692 11038 -1658
rect 11072 -1692 11080 -1658
rect 11190 -1692 11198 -1658
rect 11232 -1692 11266 -1658
rect 11300 -1692 11308 -1658
rect 10962 -1708 11080 -1692
rect 11118 -1708 11152 -1692
rect 11190 -1708 11308 -1692
rect 11362 -1558 11480 -1542
rect 11362 -1592 11370 -1558
rect 11404 -1592 11438 -1558
rect 11472 -1592 11480 -1558
rect 11362 -1658 11480 -1592
rect 11362 -1692 11370 -1658
rect 11404 -1692 11438 -1658
rect 11472 -1692 11480 -1658
rect 11362 -1708 11480 -1692
rect 11590 -1558 11708 -1542
rect 11590 -1592 11598 -1558
rect 11632 -1592 11666 -1558
rect 11700 -1592 11708 -1558
rect 11590 -1658 11708 -1592
rect 11590 -1692 11598 -1658
rect 11632 -1692 11666 -1658
rect 11700 -1692 11708 -1658
rect 11590 -1708 11708 -1692
rect 11762 -1558 11880 -1542
rect 11918 -1558 11952 -1542
rect 11990 -1558 12108 -1542
rect 11762 -1592 11770 -1558
rect 11804 -1592 11838 -1558
rect 11872 -1592 11880 -1558
rect 11990 -1592 11998 -1558
rect 12032 -1592 12066 -1558
rect 12100 -1592 12108 -1558
rect 11762 -1658 11880 -1592
rect 11918 -1608 11952 -1592
rect 11918 -1658 11952 -1642
rect 11990 -1658 12108 -1592
rect 11762 -1692 11770 -1658
rect 11804 -1692 11838 -1658
rect 11872 -1692 11880 -1658
rect 11990 -1692 11998 -1658
rect 12032 -1692 12066 -1658
rect 12100 -1692 12108 -1658
rect 11762 -1708 11880 -1692
rect 11918 -1708 11952 -1692
rect 11990 -1708 12108 -1692
rect 12162 -1558 12280 -1542
rect 12162 -1592 12170 -1558
rect 12204 -1592 12238 -1558
rect 12272 -1592 12280 -1558
rect 12162 -1658 12280 -1592
rect 12162 -1692 12170 -1658
rect 12204 -1692 12238 -1658
rect 12272 -1692 12280 -1658
rect 12162 -1708 12280 -1692
rect 12390 -1558 12508 -1542
rect 12390 -1592 12398 -1558
rect 12432 -1592 12466 -1558
rect 12500 -1592 12508 -1558
rect 12390 -1658 12508 -1592
rect 12390 -1692 12398 -1658
rect 12432 -1692 12466 -1658
rect 12500 -1692 12508 -1658
rect 12390 -1708 12508 -1692
rect 12562 -1558 12680 -1542
rect 12718 -1558 12752 -1542
rect 14808 -1542 14841 -1508
rect 14881 -1542 14913 -1508
rect 14949 -1542 14983 -1508
rect 15019 -1542 15051 -1508
rect 15091 -1542 15124 -1508
rect 15218 -1542 15251 -1508
rect 15291 -1542 15323 -1508
rect 15359 -1542 15393 -1508
rect 15429 -1542 15461 -1508
rect 15501 -1542 15534 -1508
rect 15574 -1509 15608 -1492
rect 12562 -1592 12570 -1558
rect 12604 -1592 12638 -1558
rect 12672 -1592 12680 -1558
rect 12562 -1658 12680 -1592
rect 12718 -1608 12752 -1592
rect 14734 -1608 14768 -1543
rect 15648 -1542 15676 -1508
rect 15712 -1542 15746 -1508
rect 15782 -1542 15810 -1508
rect 15574 -1608 15608 -1543
rect 14532 -1642 14558 -1608
rect 14596 -1642 14630 -1608
rect 14664 -1642 14694 -1608
rect 14808 -1642 14842 -1608
rect 14881 -1642 14914 -1608
rect 14949 -1642 14983 -1608
rect 15020 -1642 15051 -1608
rect 15092 -1642 15124 -1608
rect 15218 -1642 15249 -1608
rect 15291 -1642 15321 -1608
rect 15359 -1642 15393 -1608
rect 15427 -1642 15461 -1608
rect 15499 -1642 15534 -1608
rect 15648 -1642 15677 -1608
rect 15712 -1642 15746 -1608
rect 15783 -1642 15810 -1608
rect 12718 -1658 12752 -1642
rect 12562 -1692 12570 -1658
rect 12604 -1692 12638 -1658
rect 12672 -1692 12680 -1658
rect 12562 -1708 12680 -1692
rect 12718 -1708 12752 -1692
rect 14532 -1742 14560 -1708
rect 14596 -1742 14630 -1708
rect 14666 -1742 14694 -1708
rect 14734 -1709 14768 -1692
rect 9518 -1758 9552 -1742
rect 9590 -1758 9708 -1742
rect 9362 -1792 9370 -1758
rect 9404 -1792 9438 -1758
rect 9472 -1792 9480 -1758
rect 9590 -1792 9598 -1758
rect 9632 -1792 9666 -1758
rect 9700 -1792 9708 -1758
rect 9362 -1808 9480 -1792
rect 9518 -1808 9552 -1792
rect 6318 -1858 6352 -1842
rect 6390 -1858 6508 -1842
rect 6162 -1892 6170 -1858
rect 6204 -1892 6238 -1858
rect 6272 -1892 6280 -1858
rect 6390 -1892 6398 -1858
rect 6432 -1892 6466 -1858
rect 6500 -1892 6508 -1858
rect 6162 -1958 6280 -1892
rect 6318 -1908 6352 -1892
rect 6390 -1908 6508 -1892
rect 6562 -1858 6680 -1842
rect 6562 -1892 6570 -1858
rect 6604 -1892 6638 -1858
rect 6672 -1892 6680 -1858
rect 6562 -1908 6680 -1892
rect 6790 -1858 6908 -1842
rect 6790 -1892 6798 -1858
rect 6832 -1892 6866 -1858
rect 6900 -1892 6908 -1858
rect 6790 -1908 6908 -1892
rect 6962 -1858 7080 -1842
rect 7118 -1858 7152 -1842
rect 7190 -1858 7308 -1842
rect 6962 -1892 6970 -1858
rect 7004 -1892 7038 -1858
rect 7072 -1892 7080 -1858
rect 7190 -1892 7198 -1858
rect 7232 -1892 7266 -1858
rect 7300 -1892 7308 -1858
rect 6962 -1908 7080 -1892
rect 7118 -1908 7152 -1892
rect 7190 -1908 7308 -1892
rect 7362 -1858 7480 -1842
rect 7362 -1892 7370 -1858
rect 7404 -1892 7438 -1858
rect 7472 -1892 7480 -1858
rect 7362 -1908 7480 -1892
rect 7590 -1858 7708 -1842
rect 7590 -1892 7598 -1858
rect 7632 -1892 7666 -1858
rect 7700 -1892 7708 -1858
rect 7590 -1908 7708 -1892
rect 7762 -1858 7880 -1842
rect 7918 -1858 7952 -1842
rect 7990 -1858 8108 -1842
rect 7762 -1892 7770 -1858
rect 7804 -1892 7838 -1858
rect 7872 -1892 7880 -1858
rect 7990 -1892 7998 -1858
rect 8032 -1892 8066 -1858
rect 8100 -1892 8108 -1858
rect 7762 -1908 7880 -1892
rect 7918 -1908 7952 -1892
rect 7990 -1908 8108 -1892
rect 8162 -1858 8280 -1842
rect 8162 -1892 8170 -1858
rect 8204 -1892 8238 -1858
rect 8272 -1892 8280 -1858
rect 8162 -1908 8280 -1892
rect 8390 -1858 8508 -1842
rect 8390 -1892 8398 -1858
rect 8432 -1892 8466 -1858
rect 8500 -1892 8508 -1858
rect 8390 -1908 8508 -1892
rect 8562 -1858 8680 -1842
rect 8718 -1858 8752 -1842
rect 8790 -1858 8908 -1842
rect 8562 -1892 8570 -1858
rect 8604 -1892 8638 -1858
rect 8672 -1892 8680 -1858
rect 8790 -1892 8798 -1858
rect 8832 -1892 8866 -1858
rect 8900 -1892 8908 -1858
rect 8562 -1908 8680 -1892
rect 8718 -1908 8752 -1892
rect 8790 -1908 8908 -1892
rect 8962 -1858 9080 -1842
rect 8962 -1892 8970 -1858
rect 9004 -1892 9038 -1858
rect 9072 -1892 9080 -1858
rect 8962 -1908 9080 -1892
rect 9190 -1858 9308 -1842
rect 9190 -1892 9198 -1858
rect 9232 -1892 9266 -1858
rect 9300 -1892 9308 -1858
rect 9190 -1908 9308 -1892
rect 9362 -1858 9480 -1842
rect 9518 -1858 9552 -1842
rect 9590 -1858 9708 -1792
rect 9362 -1892 9370 -1858
rect 9404 -1892 9438 -1858
rect 9472 -1892 9480 -1858
rect 9590 -1892 9598 -1858
rect 9632 -1892 9666 -1858
rect 9700 -1892 9708 -1858
rect 9362 -1908 9480 -1892
rect 9518 -1908 9552 -1892
rect 9590 -1908 9708 -1892
rect 9762 -1758 9880 -1742
rect 9762 -1792 9770 -1758
rect 9804 -1792 9838 -1758
rect 9872 -1792 9880 -1758
rect 9762 -1858 9880 -1792
rect 9762 -1892 9770 -1858
rect 9804 -1892 9838 -1858
rect 9872 -1892 9880 -1858
rect 9762 -1908 9880 -1892
rect 9990 -1758 10108 -1742
rect 9990 -1792 9998 -1758
rect 10032 -1792 10066 -1758
rect 10100 -1792 10108 -1758
rect 9990 -1858 10108 -1792
rect 9990 -1892 9998 -1858
rect 10032 -1892 10066 -1858
rect 10100 -1892 10108 -1858
rect 9990 -1908 10108 -1892
rect 10162 -1758 10280 -1742
rect 10318 -1758 10352 -1742
rect 10390 -1758 10508 -1742
rect 10162 -1792 10170 -1758
rect 10204 -1792 10238 -1758
rect 10272 -1792 10280 -1758
rect 10390 -1792 10398 -1758
rect 10432 -1792 10466 -1758
rect 10500 -1792 10508 -1758
rect 10162 -1858 10280 -1792
rect 10318 -1808 10352 -1792
rect 10318 -1858 10352 -1842
rect 10390 -1858 10508 -1792
rect 10162 -1892 10170 -1858
rect 10204 -1892 10238 -1858
rect 10272 -1892 10280 -1858
rect 10390 -1892 10398 -1858
rect 10432 -1892 10466 -1858
rect 10500 -1892 10508 -1858
rect 10162 -1908 10280 -1892
rect 10318 -1908 10352 -1892
rect 10390 -1908 10508 -1892
rect 10562 -1758 10680 -1742
rect 10562 -1792 10570 -1758
rect 10604 -1792 10638 -1758
rect 10672 -1792 10680 -1758
rect 10562 -1858 10680 -1792
rect 10562 -1892 10570 -1858
rect 10604 -1892 10638 -1858
rect 10672 -1892 10680 -1858
rect 10562 -1908 10680 -1892
rect 10790 -1758 10908 -1742
rect 10790 -1792 10798 -1758
rect 10832 -1792 10866 -1758
rect 10900 -1792 10908 -1758
rect 10790 -1858 10908 -1792
rect 10790 -1892 10798 -1858
rect 10832 -1892 10866 -1858
rect 10900 -1892 10908 -1858
rect 10790 -1908 10908 -1892
rect 10962 -1758 11080 -1742
rect 11118 -1758 11152 -1742
rect 11190 -1758 11308 -1742
rect 10962 -1792 10970 -1758
rect 11004 -1792 11038 -1758
rect 11072 -1792 11080 -1758
rect 11190 -1792 11198 -1758
rect 11232 -1792 11266 -1758
rect 11300 -1792 11308 -1758
rect 10962 -1858 11080 -1792
rect 11118 -1808 11152 -1792
rect 11118 -1858 11152 -1842
rect 11190 -1858 11308 -1792
rect 10962 -1892 10970 -1858
rect 11004 -1892 11038 -1858
rect 11072 -1892 11080 -1858
rect 11190 -1892 11198 -1858
rect 11232 -1892 11266 -1858
rect 11300 -1892 11308 -1858
rect 10962 -1908 11080 -1892
rect 11118 -1908 11152 -1892
rect 11190 -1908 11308 -1892
rect 11362 -1758 11480 -1742
rect 11362 -1792 11370 -1758
rect 11404 -1792 11438 -1758
rect 11472 -1792 11480 -1758
rect 11362 -1858 11480 -1792
rect 11362 -1892 11370 -1858
rect 11404 -1892 11438 -1858
rect 11472 -1892 11480 -1858
rect 11362 -1908 11480 -1892
rect 11590 -1758 11708 -1742
rect 11590 -1792 11598 -1758
rect 11632 -1792 11666 -1758
rect 11700 -1792 11708 -1758
rect 11590 -1858 11708 -1792
rect 11590 -1892 11598 -1858
rect 11632 -1892 11666 -1858
rect 11700 -1892 11708 -1858
rect 11590 -1908 11708 -1892
rect 11762 -1758 11880 -1742
rect 11918 -1758 11952 -1742
rect 11990 -1758 12108 -1742
rect 11762 -1792 11770 -1758
rect 11804 -1792 11838 -1758
rect 11872 -1792 11880 -1758
rect 11990 -1792 11998 -1758
rect 12032 -1792 12066 -1758
rect 12100 -1792 12108 -1758
rect 11762 -1858 11880 -1792
rect 11918 -1808 11952 -1792
rect 11918 -1858 11952 -1842
rect 11990 -1858 12108 -1792
rect 11762 -1892 11770 -1858
rect 11804 -1892 11838 -1858
rect 11872 -1892 11880 -1858
rect 11990 -1892 11998 -1858
rect 12032 -1892 12066 -1858
rect 12100 -1892 12108 -1858
rect 11762 -1908 11880 -1892
rect 11918 -1908 11952 -1892
rect 11990 -1908 12108 -1892
rect 12162 -1758 12280 -1742
rect 12162 -1792 12170 -1758
rect 12204 -1792 12238 -1758
rect 12272 -1792 12280 -1758
rect 12162 -1858 12280 -1792
rect 12162 -1892 12170 -1858
rect 12204 -1892 12238 -1858
rect 12272 -1892 12280 -1858
rect 12162 -1908 12280 -1892
rect 12390 -1758 12508 -1742
rect 12390 -1792 12398 -1758
rect 12432 -1792 12466 -1758
rect 12500 -1792 12508 -1758
rect 12390 -1858 12508 -1792
rect 12390 -1892 12398 -1858
rect 12432 -1892 12466 -1858
rect 12500 -1892 12508 -1858
rect 12390 -1908 12508 -1892
rect 12562 -1758 12680 -1742
rect 12718 -1758 12752 -1742
rect 14808 -1742 14841 -1708
rect 14881 -1742 14913 -1708
rect 14949 -1742 14983 -1708
rect 15019 -1742 15051 -1708
rect 15091 -1742 15124 -1708
rect 15218 -1742 15251 -1708
rect 15291 -1742 15323 -1708
rect 15359 -1742 15393 -1708
rect 15429 -1742 15461 -1708
rect 15501 -1742 15534 -1708
rect 15574 -1709 15608 -1692
rect 12562 -1792 12570 -1758
rect 12604 -1792 12638 -1758
rect 12672 -1792 12680 -1758
rect 12562 -1858 12680 -1792
rect 12718 -1808 12752 -1792
rect 14734 -1808 14768 -1743
rect 15648 -1742 15676 -1708
rect 15712 -1742 15746 -1708
rect 15782 -1742 15810 -1708
rect 15574 -1808 15608 -1743
rect 14532 -1842 14558 -1808
rect 14596 -1842 14630 -1808
rect 14664 -1842 14694 -1808
rect 14808 -1842 14842 -1808
rect 14881 -1842 14914 -1808
rect 14949 -1842 14983 -1808
rect 15020 -1842 15051 -1808
rect 15092 -1842 15124 -1808
rect 15218 -1842 15249 -1808
rect 15291 -1842 15321 -1808
rect 15359 -1842 15393 -1808
rect 15427 -1842 15461 -1808
rect 15499 -1842 15534 -1808
rect 15648 -1842 15677 -1808
rect 15712 -1842 15746 -1808
rect 15783 -1842 15810 -1808
rect 12718 -1858 12752 -1842
rect 12562 -1892 12570 -1858
rect 12604 -1892 12638 -1858
rect 12672 -1892 12680 -1858
rect 12562 -1908 12680 -1892
rect 12718 -1908 12752 -1892
rect 14532 -1942 14560 -1908
rect 14596 -1942 14630 -1908
rect 14666 -1942 14694 -1908
rect 14734 -1909 14768 -1892
rect 6318 -1958 6352 -1942
rect 6390 -1958 6508 -1942
rect 6162 -1992 6170 -1958
rect 6204 -1992 6238 -1958
rect 6272 -1992 6280 -1958
rect 6390 -1992 6398 -1958
rect 6432 -1992 6466 -1958
rect 6500 -1992 6508 -1958
rect 6162 -2008 6280 -1992
rect 6318 -2008 6352 -1992
rect -82 -2058 -48 -2042
rect -10 -2058 108 -2042
rect -10 -2092 -2 -2058
rect 32 -2092 66 -2058
rect 100 -2092 108 -2058
rect -10 -2117 108 -2092
rect 162 -2058 280 -2042
rect 162 -2092 170 -2058
rect 204 -2092 238 -2058
rect 272 -2092 280 -2058
rect 162 -2117 280 -2092
rect 390 -2058 508 -2042
rect 390 -2092 398 -2058
rect 432 -2092 466 -2058
rect 500 -2092 508 -2058
rect 390 -2117 508 -2092
rect 562 -2058 680 -2042
rect 718 -2058 752 -2042
rect 790 -2058 908 -2042
rect 562 -2092 570 -2058
rect 604 -2092 638 -2058
rect 672 -2092 680 -2058
rect 562 -2117 680 -2092
rect 790 -2092 798 -2058
rect 832 -2092 866 -2058
rect 900 -2092 908 -2058
rect 790 -2117 908 -2092
rect 962 -2058 1080 -2042
rect 962 -2092 970 -2058
rect 1004 -2092 1038 -2058
rect 1072 -2092 1080 -2058
rect 962 -2117 1080 -2092
rect 1190 -2058 1308 -2042
rect 1190 -2092 1198 -2058
rect 1232 -2092 1266 -2058
rect 1300 -2092 1308 -2058
rect 1190 -2117 1308 -2092
rect 1362 -2058 1480 -2042
rect 1518 -2058 1552 -2042
rect 1590 -2058 1708 -2042
rect 1362 -2092 1370 -2058
rect 1404 -2092 1438 -2058
rect 1472 -2092 1480 -2058
rect 1362 -2117 1480 -2092
rect 1590 -2092 1598 -2058
rect 1632 -2092 1666 -2058
rect 1700 -2092 1708 -2058
rect 1590 -2117 1708 -2092
rect 1762 -2058 1880 -2042
rect 1762 -2092 1770 -2058
rect 1804 -2092 1838 -2058
rect 1872 -2092 1880 -2058
rect 1762 -2117 1880 -2092
rect 1990 -2058 2108 -2042
rect 1990 -2092 1998 -2058
rect 2032 -2092 2066 -2058
rect 2100 -2092 2108 -2058
rect 1990 -2117 2108 -2092
rect 2162 -2058 2280 -2042
rect 2318 -2058 2352 -2042
rect 2390 -2058 2508 -2042
rect 2162 -2092 2170 -2058
rect 2204 -2092 2238 -2058
rect 2272 -2092 2280 -2058
rect 2162 -2117 2280 -2092
rect 2390 -2092 2398 -2058
rect 2432 -2092 2466 -2058
rect 2500 -2092 2508 -2058
rect 2390 -2117 2508 -2092
rect 2562 -2058 2680 -2042
rect 2562 -2092 2570 -2058
rect 2604 -2092 2638 -2058
rect 2672 -2092 2680 -2058
rect 2562 -2117 2680 -2092
rect 2790 -2058 2908 -2042
rect 2790 -2092 2798 -2058
rect 2832 -2092 2866 -2058
rect 2900 -2092 2908 -2058
rect 2790 -2117 2908 -2092
rect 2962 -2058 3080 -2042
rect 3118 -2058 3152 -2042
rect 3190 -2058 3308 -2042
rect 2962 -2092 2970 -2058
rect 3004 -2092 3038 -2058
rect 3072 -2092 3080 -2058
rect 2962 -2117 3080 -2092
rect 3190 -2092 3198 -2058
rect 3232 -2092 3266 -2058
rect 3300 -2092 3308 -2058
rect 3190 -2117 3308 -2092
rect 3362 -2058 3480 -2042
rect 3362 -2092 3370 -2058
rect 3404 -2092 3438 -2058
rect 3472 -2092 3480 -2058
rect 3362 -2117 3480 -2092
rect 3590 -2058 3708 -2042
rect 3590 -2092 3598 -2058
rect 3632 -2092 3666 -2058
rect 3700 -2092 3708 -2058
rect 3590 -2117 3708 -2092
rect 3762 -2058 3880 -2042
rect 3918 -2058 3952 -2042
rect 3990 -2058 4108 -2042
rect 3762 -2092 3770 -2058
rect 3804 -2092 3838 -2058
rect 3872 -2092 3880 -2058
rect 3762 -2117 3880 -2092
rect 3990 -2092 3998 -2058
rect 4032 -2092 4066 -2058
rect 4100 -2092 4108 -2058
rect 3990 -2117 4108 -2092
rect 4162 -2058 4280 -2042
rect 4162 -2092 4170 -2058
rect 4204 -2092 4238 -2058
rect 4272 -2092 4280 -2058
rect 4162 -2117 4280 -2092
rect 4390 -2058 4508 -2042
rect 4390 -2092 4398 -2058
rect 4432 -2092 4466 -2058
rect 4500 -2092 4508 -2058
rect 4390 -2117 4508 -2092
rect 4562 -2058 4680 -2042
rect 4718 -2058 4752 -2042
rect 4790 -2058 4908 -2042
rect 4562 -2092 4570 -2058
rect 4604 -2092 4638 -2058
rect 4672 -2092 4680 -2058
rect 4562 -2117 4680 -2092
rect 4790 -2092 4798 -2058
rect 4832 -2092 4866 -2058
rect 4900 -2092 4908 -2058
rect 4790 -2117 4908 -2092
rect 4962 -2058 5080 -2042
rect 4962 -2092 4970 -2058
rect 5004 -2092 5038 -2058
rect 5072 -2092 5080 -2058
rect 4962 -2117 5080 -2092
rect 5190 -2058 5308 -2042
rect 5190 -2092 5198 -2058
rect 5232 -2092 5266 -2058
rect 5300 -2092 5308 -2058
rect 5190 -2117 5308 -2092
rect 5362 -2058 5480 -2042
rect 5518 -2058 5552 -2042
rect 5590 -2058 5708 -2042
rect 5362 -2092 5370 -2058
rect 5404 -2092 5438 -2058
rect 5472 -2092 5480 -2058
rect 5362 -2117 5480 -2092
rect 5590 -2092 5598 -2058
rect 5632 -2092 5666 -2058
rect 5700 -2092 5708 -2058
rect 5590 -2117 5708 -2092
rect 5762 -2058 5880 -2042
rect 5762 -2092 5770 -2058
rect 5804 -2092 5838 -2058
rect 5872 -2092 5880 -2058
rect 5762 -2117 5880 -2092
rect 5990 -2058 6108 -2042
rect 5990 -2092 5998 -2058
rect 6032 -2092 6066 -2058
rect 6100 -2092 6108 -2058
rect 5990 -2117 6108 -2092
rect 6162 -2058 6280 -2042
rect 6318 -2058 6352 -2042
rect 6390 -2058 6508 -1992
rect 6162 -2092 6170 -2058
rect 6204 -2092 6238 -2058
rect 6272 -2092 6280 -2058
rect 6162 -2117 6280 -2092
rect 6390 -2092 6398 -2058
rect 6432 -2092 6466 -2058
rect 6500 -2092 6508 -2058
rect 6390 -2117 6508 -2092
rect 6562 -1958 6680 -1942
rect 6562 -1992 6570 -1958
rect 6604 -1992 6638 -1958
rect 6672 -1992 6680 -1958
rect 6562 -2058 6680 -1992
rect 6562 -2092 6570 -2058
rect 6604 -2092 6638 -2058
rect 6672 -2092 6680 -2058
rect 6562 -2117 6680 -2092
rect 6790 -1958 6908 -1942
rect 6790 -1992 6798 -1958
rect 6832 -1992 6866 -1958
rect 6900 -1992 6908 -1958
rect 6790 -2058 6908 -1992
rect 6790 -2092 6798 -2058
rect 6832 -2092 6866 -2058
rect 6900 -2092 6908 -2058
rect 6790 -2117 6908 -2092
rect 6962 -1958 7080 -1942
rect 7118 -1958 7152 -1942
rect 7190 -1958 7308 -1942
rect 6962 -1992 6970 -1958
rect 7004 -1992 7038 -1958
rect 7072 -1992 7080 -1958
rect 7190 -1992 7198 -1958
rect 7232 -1992 7266 -1958
rect 7300 -1992 7308 -1958
rect 6962 -2058 7080 -1992
rect 7118 -2008 7152 -1992
rect 7118 -2058 7152 -2042
rect 7190 -2058 7308 -1992
rect 6962 -2092 6970 -2058
rect 7004 -2092 7038 -2058
rect 7072 -2092 7080 -2058
rect 6962 -2117 7080 -2092
rect 7190 -2092 7198 -2058
rect 7232 -2092 7266 -2058
rect 7300 -2092 7308 -2058
rect 7190 -2117 7308 -2092
rect 7362 -1958 7480 -1942
rect 7362 -1992 7370 -1958
rect 7404 -1992 7438 -1958
rect 7472 -1992 7480 -1958
rect 7362 -2058 7480 -1992
rect 7362 -2092 7370 -2058
rect 7404 -2092 7438 -2058
rect 7472 -2092 7480 -2058
rect 7362 -2117 7480 -2092
rect 7590 -1958 7708 -1942
rect 7590 -1992 7598 -1958
rect 7632 -1992 7666 -1958
rect 7700 -1992 7708 -1958
rect 7590 -2058 7708 -1992
rect 7590 -2092 7598 -2058
rect 7632 -2092 7666 -2058
rect 7700 -2092 7708 -2058
rect 7590 -2117 7708 -2092
rect 7762 -1958 7880 -1942
rect 7918 -1958 7952 -1942
rect 7990 -1958 8108 -1942
rect 7762 -1992 7770 -1958
rect 7804 -1992 7838 -1958
rect 7872 -1992 7880 -1958
rect 7990 -1992 7998 -1958
rect 8032 -1992 8066 -1958
rect 8100 -1992 8108 -1958
rect 7762 -2058 7880 -1992
rect 7918 -2008 7952 -1992
rect 7918 -2058 7952 -2042
rect 7990 -2058 8108 -1992
rect 7762 -2092 7770 -2058
rect 7804 -2092 7838 -2058
rect 7872 -2092 7880 -2058
rect 7762 -2117 7880 -2092
rect 7990 -2092 7998 -2058
rect 8032 -2092 8066 -2058
rect 8100 -2092 8108 -2058
rect 7990 -2117 8108 -2092
rect 8162 -1958 8280 -1942
rect 8162 -1992 8170 -1958
rect 8204 -1992 8238 -1958
rect 8272 -1992 8280 -1958
rect 8162 -2058 8280 -1992
rect 8162 -2092 8170 -2058
rect 8204 -2092 8238 -2058
rect 8272 -2092 8280 -2058
rect 8162 -2117 8280 -2092
rect 8390 -1958 8508 -1942
rect 8390 -1992 8398 -1958
rect 8432 -1992 8466 -1958
rect 8500 -1992 8508 -1958
rect 8390 -2058 8508 -1992
rect 8390 -2092 8398 -2058
rect 8432 -2092 8466 -2058
rect 8500 -2092 8508 -2058
rect 8390 -2117 8508 -2092
rect 8562 -1958 8680 -1942
rect 8718 -1958 8752 -1942
rect 8790 -1958 8908 -1942
rect 8562 -1992 8570 -1958
rect 8604 -1992 8638 -1958
rect 8672 -1992 8680 -1958
rect 8790 -1992 8798 -1958
rect 8832 -1992 8866 -1958
rect 8900 -1992 8908 -1958
rect 8562 -2058 8680 -1992
rect 8718 -2008 8752 -1992
rect 8718 -2058 8752 -2042
rect 8790 -2058 8908 -1992
rect 8562 -2092 8570 -2058
rect 8604 -2092 8638 -2058
rect 8672 -2092 8680 -2058
rect 8562 -2117 8680 -2092
rect 8790 -2092 8798 -2058
rect 8832 -2092 8866 -2058
rect 8900 -2092 8908 -2058
rect 8790 -2117 8908 -2092
rect 8962 -1958 9080 -1942
rect 8962 -1992 8970 -1958
rect 9004 -1992 9038 -1958
rect 9072 -1992 9080 -1958
rect 8962 -2058 9080 -1992
rect 8962 -2092 8970 -2058
rect 9004 -2092 9038 -2058
rect 9072 -2092 9080 -2058
rect 8962 -2117 9080 -2092
rect 9190 -1958 9308 -1942
rect 9190 -1992 9198 -1958
rect 9232 -1992 9266 -1958
rect 9300 -1992 9308 -1958
rect 9190 -2058 9308 -1992
rect 9190 -2092 9198 -2058
rect 9232 -2092 9266 -2058
rect 9300 -2092 9308 -2058
rect 9190 -2117 9308 -2092
rect 9362 -1958 9480 -1942
rect 9518 -1958 9552 -1942
rect 9590 -1958 9708 -1942
rect 9362 -1992 9370 -1958
rect 9404 -1992 9438 -1958
rect 9472 -1992 9480 -1958
rect 9590 -1992 9598 -1958
rect 9632 -1992 9666 -1958
rect 9700 -1992 9708 -1958
rect 9362 -2058 9480 -1992
rect 9518 -2008 9552 -1992
rect 9518 -2058 9552 -2042
rect 9590 -2058 9708 -1992
rect 9362 -2092 9370 -2058
rect 9404 -2092 9438 -2058
rect 9472 -2092 9480 -2058
rect 9362 -2117 9480 -2092
rect 9590 -2092 9598 -2058
rect 9632 -2092 9666 -2058
rect 9700 -2092 9708 -2058
rect 9590 -2117 9708 -2092
rect 9762 -1958 9880 -1942
rect 9762 -1992 9770 -1958
rect 9804 -1992 9838 -1958
rect 9872 -1992 9880 -1958
rect 9762 -2058 9880 -1992
rect 9762 -2092 9770 -2058
rect 9804 -2092 9838 -2058
rect 9872 -2092 9880 -2058
rect 9762 -2117 9880 -2092
rect 9990 -1958 10108 -1942
rect 9990 -1992 9998 -1958
rect 10032 -1992 10066 -1958
rect 10100 -1992 10108 -1958
rect 9990 -2058 10108 -1992
rect 9990 -2092 9998 -2058
rect 10032 -2092 10066 -2058
rect 10100 -2092 10108 -2058
rect 9990 -2117 10108 -2092
rect 10162 -1958 10280 -1942
rect 10318 -1958 10352 -1942
rect 10390 -1958 10508 -1942
rect 10162 -1992 10170 -1958
rect 10204 -1992 10238 -1958
rect 10272 -1992 10280 -1958
rect 10390 -1992 10398 -1958
rect 10432 -1992 10466 -1958
rect 10500 -1992 10508 -1958
rect 10162 -2058 10280 -1992
rect 10318 -2008 10352 -1992
rect 10318 -2058 10352 -2042
rect 10390 -2058 10508 -1992
rect 10162 -2092 10170 -2058
rect 10204 -2092 10238 -2058
rect 10272 -2092 10280 -2058
rect 10162 -2117 10280 -2092
rect 10390 -2092 10398 -2058
rect 10432 -2092 10466 -2058
rect 10500 -2092 10508 -2058
rect 10390 -2117 10508 -2092
rect 10562 -1958 10680 -1942
rect 10562 -1992 10570 -1958
rect 10604 -1992 10638 -1958
rect 10672 -1992 10680 -1958
rect 10562 -2058 10680 -1992
rect 10562 -2092 10570 -2058
rect 10604 -2092 10638 -2058
rect 10672 -2092 10680 -2058
rect 10562 -2117 10680 -2092
rect 10790 -1958 10908 -1942
rect 10790 -1992 10798 -1958
rect 10832 -1992 10866 -1958
rect 10900 -1992 10908 -1958
rect 10790 -2058 10908 -1992
rect 10790 -2092 10798 -2058
rect 10832 -2092 10866 -2058
rect 10900 -2092 10908 -2058
rect 10790 -2117 10908 -2092
rect 10962 -1958 11080 -1942
rect 11118 -1958 11152 -1942
rect 11190 -1958 11308 -1942
rect 10962 -1992 10970 -1958
rect 11004 -1992 11038 -1958
rect 11072 -1992 11080 -1958
rect 11190 -1992 11198 -1958
rect 11232 -1992 11266 -1958
rect 11300 -1992 11308 -1958
rect 10962 -2058 11080 -1992
rect 11118 -2008 11152 -1992
rect 11118 -2058 11152 -2042
rect 11190 -2058 11308 -1992
rect 10962 -2092 10970 -2058
rect 11004 -2092 11038 -2058
rect 11072 -2092 11080 -2058
rect 10962 -2117 11080 -2092
rect 11190 -2092 11198 -2058
rect 11232 -2092 11266 -2058
rect 11300 -2092 11308 -2058
rect 11190 -2117 11308 -2092
rect 11362 -1958 11480 -1942
rect 11362 -1992 11370 -1958
rect 11404 -1992 11438 -1958
rect 11472 -1992 11480 -1958
rect 11362 -2058 11480 -1992
rect 11362 -2092 11370 -2058
rect 11404 -2092 11438 -2058
rect 11472 -2092 11480 -2058
rect 11362 -2117 11480 -2092
rect 11590 -1958 11708 -1942
rect 11590 -1992 11598 -1958
rect 11632 -1992 11666 -1958
rect 11700 -1992 11708 -1958
rect 11590 -2058 11708 -1992
rect 11590 -2092 11598 -2058
rect 11632 -2092 11666 -2058
rect 11700 -2092 11708 -2058
rect 11590 -2117 11708 -2092
rect 11762 -1958 11880 -1942
rect 11918 -1958 11952 -1942
rect 11990 -1958 12108 -1942
rect 11762 -1992 11770 -1958
rect 11804 -1992 11838 -1958
rect 11872 -1992 11880 -1958
rect 11990 -1992 11998 -1958
rect 12032 -1992 12066 -1958
rect 12100 -1992 12108 -1958
rect 11762 -2058 11880 -1992
rect 11918 -2008 11952 -1992
rect 11918 -2058 11952 -2042
rect 11990 -2058 12108 -1992
rect 11762 -2092 11770 -2058
rect 11804 -2092 11838 -2058
rect 11872 -2092 11880 -2058
rect 11762 -2117 11880 -2092
rect 11990 -2092 11998 -2058
rect 12032 -2092 12066 -2058
rect 12100 -2092 12108 -2058
rect 11990 -2117 12108 -2092
rect 12162 -1958 12280 -1942
rect 12162 -1992 12170 -1958
rect 12204 -1992 12238 -1958
rect 12272 -1992 12280 -1958
rect 12162 -2058 12280 -1992
rect 12162 -2092 12170 -2058
rect 12204 -2092 12238 -2058
rect 12272 -2092 12280 -2058
rect 12162 -2117 12280 -2092
rect 12390 -1958 12508 -1942
rect 12390 -1992 12398 -1958
rect 12432 -1992 12466 -1958
rect 12500 -1992 12508 -1958
rect 12390 -2058 12508 -1992
rect 12390 -2092 12398 -2058
rect 12432 -2092 12466 -2058
rect 12500 -2092 12508 -2058
rect 12390 -2117 12508 -2092
rect 12562 -1958 12680 -1942
rect 12718 -1958 12752 -1942
rect 14808 -1942 14841 -1908
rect 14881 -1942 14913 -1908
rect 14949 -1942 14983 -1908
rect 15019 -1942 15051 -1908
rect 15091 -1942 15124 -1908
rect 15218 -1942 15251 -1908
rect 15291 -1942 15323 -1908
rect 15359 -1942 15393 -1908
rect 15429 -1942 15461 -1908
rect 15501 -1942 15534 -1908
rect 15574 -1909 15608 -1892
rect 12562 -1992 12570 -1958
rect 12604 -1992 12638 -1958
rect 12672 -1992 12680 -1958
rect 12562 -2058 12680 -1992
rect 12718 -2008 12752 -1992
rect 14734 -2008 14768 -1943
rect 15648 -1942 15676 -1908
rect 15712 -1942 15746 -1908
rect 15782 -1942 15810 -1908
rect 15574 -2008 15608 -1943
rect 14532 -2042 14558 -2008
rect 14596 -2042 14630 -2008
rect 14664 -2042 14694 -2008
rect 14808 -2042 14842 -2008
rect 14881 -2042 14914 -2008
rect 14949 -2042 14983 -2008
rect 15020 -2042 15051 -2008
rect 15092 -2042 15124 -2008
rect 15218 -2042 15249 -2008
rect 15291 -2042 15321 -2008
rect 15359 -2042 15393 -2008
rect 15427 -2042 15461 -2008
rect 15499 -2042 15534 -2008
rect 15648 -2042 15677 -2008
rect 15712 -2042 15746 -2008
rect 15783 -2042 15810 -2008
rect 12718 -2058 12752 -2042
rect 12562 -2092 12570 -2058
rect 12604 -2092 12638 -2058
rect 12672 -2092 12680 -2058
rect 12562 -2117 12680 -2092
rect 14548 -2101 14682 -2042
rect -65 -2135 12735 -2117
rect 14548 -2135 14564 -2101
rect 14598 -2135 14632 -2101
rect 14666 -2135 14682 -2101
rect 14824 -2101 15108 -2042
rect 14824 -2135 14847 -2101
rect 14881 -2135 14915 -2101
rect 14949 -2135 14983 -2101
rect 15017 -2135 15051 -2101
rect 15085 -2135 15108 -2101
rect 15234 -2101 15518 -2042
rect 15234 -2135 15257 -2101
rect 15291 -2135 15325 -2101
rect 15359 -2135 15393 -2101
rect 15427 -2135 15461 -2101
rect 15495 -2135 15518 -2101
rect 15660 -2101 15794 -2042
rect 15660 -2135 15676 -2101
rect 15710 -2135 15744 -2101
rect 15778 -2135 15794 -2101
rect -65 -2169 -4 -2135
rect 30 -2151 68 -2135
rect 30 -2169 32 -2151
rect -65 -2185 32 -2169
rect 66 -2169 68 -2151
rect 102 -2169 168 -2135
rect 202 -2151 240 -2135
rect 202 -2169 204 -2151
rect 66 -2185 204 -2169
rect 238 -2169 240 -2151
rect 274 -2169 396 -2135
rect 430 -2151 468 -2135
rect 430 -2169 432 -2151
rect 238 -2185 432 -2169
rect 466 -2169 468 -2151
rect 502 -2169 568 -2135
rect 602 -2151 640 -2135
rect 602 -2169 604 -2151
rect 466 -2185 604 -2169
rect 638 -2169 640 -2151
rect 674 -2169 796 -2135
rect 830 -2151 868 -2135
rect 830 -2169 832 -2151
rect 638 -2185 832 -2169
rect 866 -2169 868 -2151
rect 902 -2169 968 -2135
rect 1002 -2151 1040 -2135
rect 1002 -2169 1004 -2151
rect 866 -2185 1004 -2169
rect 1038 -2169 1040 -2151
rect 1074 -2169 1196 -2135
rect 1230 -2151 1268 -2135
rect 1230 -2169 1232 -2151
rect 1038 -2185 1232 -2169
rect 1266 -2169 1268 -2151
rect 1302 -2169 1368 -2135
rect 1402 -2151 1440 -2135
rect 1402 -2169 1404 -2151
rect 1266 -2185 1404 -2169
rect 1438 -2169 1440 -2151
rect 1474 -2169 1596 -2135
rect 1630 -2151 1668 -2135
rect 1630 -2169 1632 -2151
rect 1438 -2185 1632 -2169
rect 1666 -2169 1668 -2151
rect 1702 -2169 1768 -2135
rect 1802 -2151 1840 -2135
rect 1802 -2169 1804 -2151
rect 1666 -2185 1804 -2169
rect 1838 -2169 1840 -2151
rect 1874 -2169 1996 -2135
rect 2030 -2151 2068 -2135
rect 2030 -2169 2032 -2151
rect 1838 -2185 2032 -2169
rect 2066 -2169 2068 -2151
rect 2102 -2169 2168 -2135
rect 2202 -2151 2240 -2135
rect 2202 -2169 2204 -2151
rect 2066 -2185 2204 -2169
rect 2238 -2169 2240 -2151
rect 2274 -2169 2396 -2135
rect 2430 -2151 2468 -2135
rect 2430 -2169 2432 -2151
rect 2238 -2185 2432 -2169
rect 2466 -2169 2468 -2151
rect 2502 -2169 2568 -2135
rect 2602 -2151 2640 -2135
rect 2602 -2169 2604 -2151
rect 2466 -2185 2604 -2169
rect 2638 -2169 2640 -2151
rect 2674 -2169 2796 -2135
rect 2830 -2151 2868 -2135
rect 2830 -2169 2832 -2151
rect 2638 -2185 2832 -2169
rect 2866 -2169 2868 -2151
rect 2902 -2169 2968 -2135
rect 3002 -2151 3040 -2135
rect 3002 -2169 3004 -2151
rect 2866 -2185 3004 -2169
rect 3038 -2169 3040 -2151
rect 3074 -2169 3196 -2135
rect 3230 -2151 3268 -2135
rect 3230 -2169 3232 -2151
rect 3038 -2185 3232 -2169
rect 3266 -2169 3268 -2151
rect 3302 -2169 3368 -2135
rect 3402 -2151 3440 -2135
rect 3402 -2169 3404 -2151
rect 3266 -2185 3404 -2169
rect 3438 -2169 3440 -2151
rect 3474 -2169 3596 -2135
rect 3630 -2151 3668 -2135
rect 3630 -2169 3632 -2151
rect 3438 -2185 3632 -2169
rect 3666 -2169 3668 -2151
rect 3702 -2169 3768 -2135
rect 3802 -2151 3840 -2135
rect 3802 -2169 3804 -2151
rect 3666 -2185 3804 -2169
rect 3838 -2169 3840 -2151
rect 3874 -2169 3996 -2135
rect 4030 -2151 4068 -2135
rect 4030 -2169 4032 -2151
rect 3838 -2185 4032 -2169
rect 4066 -2169 4068 -2151
rect 4102 -2169 4168 -2135
rect 4202 -2151 4240 -2135
rect 4202 -2169 4204 -2151
rect 4066 -2185 4204 -2169
rect 4238 -2169 4240 -2151
rect 4274 -2169 4396 -2135
rect 4430 -2151 4468 -2135
rect 4430 -2169 4432 -2151
rect 4238 -2185 4432 -2169
rect 4466 -2169 4468 -2151
rect 4502 -2169 4568 -2135
rect 4602 -2151 4640 -2135
rect 4602 -2169 4604 -2151
rect 4466 -2185 4604 -2169
rect 4638 -2169 4640 -2151
rect 4674 -2169 4796 -2135
rect 4830 -2151 4868 -2135
rect 4830 -2169 4832 -2151
rect 4638 -2185 4832 -2169
rect 4866 -2169 4868 -2151
rect 4902 -2169 4968 -2135
rect 5002 -2151 5040 -2135
rect 5002 -2169 5004 -2151
rect 4866 -2185 5004 -2169
rect 5038 -2169 5040 -2151
rect 5074 -2169 5196 -2135
rect 5230 -2151 5268 -2135
rect 5230 -2169 5232 -2151
rect 5038 -2185 5232 -2169
rect 5266 -2169 5268 -2151
rect 5302 -2169 5368 -2135
rect 5402 -2151 5440 -2135
rect 5402 -2169 5404 -2151
rect 5266 -2185 5404 -2169
rect 5438 -2169 5440 -2151
rect 5474 -2169 5596 -2135
rect 5630 -2151 5668 -2135
rect 5630 -2169 5632 -2151
rect 5438 -2185 5632 -2169
rect 5666 -2169 5668 -2151
rect 5702 -2169 5768 -2135
rect 5802 -2151 5840 -2135
rect 5802 -2169 5804 -2151
rect 5666 -2185 5804 -2169
rect 5838 -2169 5840 -2151
rect 5874 -2169 5996 -2135
rect 6030 -2151 6068 -2135
rect 6030 -2169 6032 -2151
rect 5838 -2185 6032 -2169
rect 6066 -2169 6068 -2151
rect 6102 -2169 6168 -2135
rect 6202 -2151 6240 -2135
rect 6202 -2169 6204 -2151
rect 6066 -2185 6204 -2169
rect 6238 -2169 6240 -2151
rect 6274 -2169 6396 -2135
rect 6430 -2151 6468 -2135
rect 6430 -2169 6432 -2151
rect 6238 -2185 6432 -2169
rect 6466 -2169 6468 -2151
rect 6502 -2169 6568 -2135
rect 6602 -2151 6640 -2135
rect 6602 -2169 6604 -2151
rect 6466 -2185 6604 -2169
rect 6638 -2169 6640 -2151
rect 6674 -2169 6796 -2135
rect 6830 -2151 6868 -2135
rect 6830 -2169 6832 -2151
rect 6638 -2185 6832 -2169
rect 6866 -2169 6868 -2151
rect 6902 -2169 6968 -2135
rect 7002 -2151 7040 -2135
rect 7002 -2169 7004 -2151
rect 6866 -2185 7004 -2169
rect 7038 -2169 7040 -2151
rect 7074 -2169 7196 -2135
rect 7230 -2151 7268 -2135
rect 7230 -2169 7232 -2151
rect 7038 -2185 7232 -2169
rect 7266 -2169 7268 -2151
rect 7302 -2169 7368 -2135
rect 7402 -2151 7440 -2135
rect 7402 -2169 7404 -2151
rect 7266 -2185 7404 -2169
rect 7438 -2169 7440 -2151
rect 7474 -2169 7596 -2135
rect 7630 -2151 7668 -2135
rect 7630 -2169 7632 -2151
rect 7438 -2185 7632 -2169
rect 7666 -2169 7668 -2151
rect 7702 -2169 7768 -2135
rect 7802 -2151 7840 -2135
rect 7802 -2169 7804 -2151
rect 7666 -2185 7804 -2169
rect 7838 -2169 7840 -2151
rect 7874 -2169 7996 -2135
rect 8030 -2151 8068 -2135
rect 8030 -2169 8032 -2151
rect 7838 -2185 8032 -2169
rect 8066 -2169 8068 -2151
rect 8102 -2169 8168 -2135
rect 8202 -2151 8240 -2135
rect 8202 -2169 8204 -2151
rect 8066 -2185 8204 -2169
rect 8238 -2169 8240 -2151
rect 8274 -2169 8396 -2135
rect 8430 -2151 8468 -2135
rect 8430 -2169 8432 -2151
rect 8238 -2185 8432 -2169
rect 8466 -2169 8468 -2151
rect 8502 -2169 8568 -2135
rect 8602 -2151 8640 -2135
rect 8602 -2169 8604 -2151
rect 8466 -2185 8604 -2169
rect 8638 -2169 8640 -2151
rect 8674 -2169 8796 -2135
rect 8830 -2151 8868 -2135
rect 8830 -2169 8832 -2151
rect 8638 -2185 8832 -2169
rect 8866 -2169 8868 -2151
rect 8902 -2169 8968 -2135
rect 9002 -2151 9040 -2135
rect 9002 -2169 9004 -2151
rect 8866 -2185 9004 -2169
rect 9038 -2169 9040 -2151
rect 9074 -2169 9196 -2135
rect 9230 -2151 9268 -2135
rect 9230 -2169 9232 -2151
rect 9038 -2185 9232 -2169
rect 9266 -2169 9268 -2151
rect 9302 -2169 9368 -2135
rect 9402 -2151 9440 -2135
rect 9402 -2169 9404 -2151
rect 9266 -2185 9404 -2169
rect 9438 -2169 9440 -2151
rect 9474 -2169 9596 -2135
rect 9630 -2151 9668 -2135
rect 9630 -2169 9632 -2151
rect 9438 -2185 9632 -2169
rect 9666 -2169 9668 -2151
rect 9702 -2169 9768 -2135
rect 9802 -2151 9840 -2135
rect 9802 -2169 9804 -2151
rect 9666 -2185 9804 -2169
rect 9838 -2169 9840 -2151
rect 9874 -2169 9996 -2135
rect 10030 -2151 10068 -2135
rect 10030 -2169 10032 -2151
rect 9838 -2185 10032 -2169
rect 10066 -2169 10068 -2151
rect 10102 -2169 10168 -2135
rect 10202 -2151 10240 -2135
rect 10202 -2169 10204 -2151
rect 10066 -2185 10204 -2169
rect 10238 -2169 10240 -2151
rect 10274 -2169 10396 -2135
rect 10430 -2151 10468 -2135
rect 10430 -2169 10432 -2151
rect 10238 -2185 10432 -2169
rect 10466 -2169 10468 -2151
rect 10502 -2169 10568 -2135
rect 10602 -2151 10640 -2135
rect 10602 -2169 10604 -2151
rect 10466 -2185 10604 -2169
rect 10638 -2169 10640 -2151
rect 10674 -2169 10796 -2135
rect 10830 -2151 10868 -2135
rect 10830 -2169 10832 -2151
rect 10638 -2185 10832 -2169
rect 10866 -2169 10868 -2151
rect 10902 -2169 10968 -2135
rect 11002 -2151 11040 -2135
rect 11002 -2169 11004 -2151
rect 10866 -2185 11004 -2169
rect 11038 -2169 11040 -2151
rect 11074 -2169 11196 -2135
rect 11230 -2151 11268 -2135
rect 11230 -2169 11232 -2151
rect 11038 -2185 11232 -2169
rect 11266 -2169 11268 -2151
rect 11302 -2169 11368 -2135
rect 11402 -2151 11440 -2135
rect 11402 -2169 11404 -2151
rect 11266 -2185 11404 -2169
rect 11438 -2169 11440 -2151
rect 11474 -2169 11596 -2135
rect 11630 -2151 11668 -2135
rect 11630 -2169 11632 -2151
rect 11438 -2185 11632 -2169
rect 11666 -2169 11668 -2151
rect 11702 -2169 11768 -2135
rect 11802 -2151 11840 -2135
rect 11802 -2169 11804 -2151
rect 11666 -2185 11804 -2169
rect 11838 -2169 11840 -2151
rect 11874 -2169 11996 -2135
rect 12030 -2151 12068 -2135
rect 12030 -2169 12032 -2151
rect 11838 -2185 12032 -2169
rect 12066 -2169 12068 -2151
rect 12102 -2169 12168 -2135
rect 12202 -2151 12240 -2135
rect 12202 -2169 12204 -2151
rect 12066 -2185 12204 -2169
rect 12238 -2169 12240 -2151
rect 12274 -2169 12396 -2135
rect 12430 -2151 12468 -2135
rect 12430 -2169 12432 -2151
rect 12238 -2185 12432 -2169
rect 12466 -2169 12468 -2151
rect 12502 -2169 12568 -2135
rect 12602 -2151 12640 -2135
rect 12602 -2169 12604 -2151
rect 12466 -2185 12604 -2169
rect 12638 -2169 12640 -2151
rect 12674 -2169 12735 -2135
rect 12638 -2185 12735 -2169
rect -65 -2187 12735 -2185
<< viali >>
rect 118 4983 152 5017
rect 318 4983 352 5017
rect 518 4983 552 5017
rect 718 4983 752 5017
rect 918 4983 952 5017
rect 1118 4983 1152 5017
rect 1318 4983 1352 5017
rect 1518 4983 1552 5017
rect 1718 4983 1752 5017
rect 1918 4983 1952 5017
rect 2118 4983 2152 5017
rect 2318 4983 2352 5017
rect 2518 4983 2552 5017
rect 2718 4983 2752 5017
rect 2918 4983 2952 5017
rect 3118 4983 3152 5017
rect 3318 4983 3352 5017
rect 3518 4983 3552 5017
rect 3718 4983 3752 5017
rect 3918 4983 3952 5017
rect 4118 4983 4152 5017
rect 4318 4983 4352 5017
rect 4518 4983 4552 5017
rect 4718 4983 4752 5017
rect 4918 4983 4952 5017
rect 5118 4983 5152 5017
rect 5318 4983 5352 5017
rect 5518 4983 5552 5017
rect 5718 4983 5752 5017
rect 5918 4983 5952 5017
rect 6118 4983 6152 5017
rect 6318 4983 6352 5017
rect 6518 4983 6552 5017
rect 6718 4983 6752 5017
rect 6918 4983 6952 5017
rect 7118 4983 7152 5017
rect 7318 4983 7352 5017
rect 7518 4983 7552 5017
rect 7718 4983 7752 5017
rect 7918 4983 7952 5017
rect 8118 4983 8152 5017
rect 8318 4983 8352 5017
rect 8518 4983 8552 5017
rect 8718 4983 8752 5017
rect 8918 4983 8952 5017
rect 9118 4983 9152 5017
rect 9318 4983 9352 5017
rect 9518 4983 9552 5017
rect 9718 4983 9752 5017
rect 9918 4983 9952 5017
rect 10118 4983 10152 5017
rect 10318 4983 10352 5017
rect 10518 4983 10552 5017
rect 10718 4983 10752 5017
rect 10918 4983 10952 5017
rect 11118 4983 11152 5017
rect 11318 4983 11352 5017
rect 11518 4983 11552 5017
rect 11718 4983 11752 5017
rect 11918 4983 11952 5017
rect 12118 4983 12152 5017
rect 12318 4983 12352 5017
rect 12518 4983 12552 5017
rect 12718 4983 12752 5017
rect 18 4860 52 4894
rect 218 4876 252 4910
rect 418 4860 452 4894
rect 618 4876 652 4910
rect 818 4860 852 4894
rect 1018 4876 1052 4910
rect 1218 4860 1252 4894
rect 1418 4876 1452 4910
rect 1618 4860 1652 4894
rect 1818 4876 1852 4910
rect 2018 4860 2052 4894
rect 2218 4876 2252 4910
rect 2418 4860 2452 4894
rect 2618 4876 2652 4910
rect 2818 4860 2852 4894
rect 3018 4876 3052 4910
rect 3218 4860 3252 4894
rect 3418 4876 3452 4910
rect 3618 4860 3652 4894
rect 3818 4876 3852 4910
rect 4018 4860 4052 4894
rect 4218 4876 4252 4910
rect 4418 4860 4452 4894
rect 4618 4876 4652 4910
rect 4818 4860 4852 4894
rect 5018 4876 5052 4910
rect 5218 4860 5252 4894
rect 5418 4876 5452 4910
rect 5618 4860 5652 4894
rect 5818 4876 5852 4910
rect 6018 4860 6052 4894
rect 6218 4876 6252 4910
rect 6418 4860 6452 4894
rect 6618 4876 6652 4910
rect 6818 4860 6852 4894
rect 7018 4876 7052 4910
rect 7218 4860 7252 4894
rect 7418 4876 7452 4910
rect 7618 4860 7652 4894
rect 7818 4876 7852 4910
rect 8018 4860 8052 4894
rect 8218 4876 8252 4910
rect 8418 4860 8452 4894
rect 8618 4876 8652 4910
rect 8818 4860 8852 4894
rect 9018 4876 9052 4910
rect 9218 4860 9252 4894
rect 9418 4876 9452 4910
rect 9618 4860 9652 4894
rect 9818 4876 9852 4910
rect 10018 4860 10052 4894
rect 10218 4876 10252 4910
rect 10418 4860 10452 4894
rect 10618 4876 10652 4910
rect 10818 4860 10852 4894
rect 11018 4876 11052 4910
rect 11218 4860 11252 4894
rect 11418 4876 11452 4910
rect 11618 4860 11652 4894
rect 11818 4876 11852 4910
rect 12018 4860 12052 4894
rect 12218 4876 12252 4910
rect 12418 4860 12452 4894
rect 12618 4876 12652 4910
rect 12916 4857 12950 4891
rect 13120 4879 13154 4913
rect 13278 4874 13312 4908
rect 13378 4874 13412 4908
rect 13478 4874 13512 4908
rect 13578 4874 13612 4908
rect 18 4753 24 4787
rect 24 4753 52 4787
rect 118 4753 152 4787
rect 218 4753 252 4787
rect 318 4753 346 4787
rect 346 4753 352 4787
rect 418 4753 424 4787
rect 424 4753 452 4787
rect 518 4753 552 4787
rect 618 4753 652 4787
rect 718 4753 752 4787
rect 818 4753 852 4787
rect 918 4753 952 4787
rect 1018 4753 1052 4787
rect 1118 4753 1146 4787
rect 1146 4753 1152 4787
rect 1218 4753 1224 4787
rect 1224 4753 1252 4787
rect 1318 4753 1352 4787
rect 1418 4753 1452 4787
rect 1518 4753 1552 4787
rect 1618 4753 1652 4787
rect 1718 4753 1752 4787
rect 1818 4753 1852 4787
rect 1918 4753 1952 4787
rect 2018 4753 2052 4787
rect 2118 4753 2152 4787
rect 2218 4753 2252 4787
rect 2318 4753 2346 4787
rect 2346 4753 2352 4787
rect 2418 4753 2424 4787
rect 2424 4753 2452 4787
rect 2518 4753 2552 4787
rect 2618 4753 2652 4787
rect 2718 4753 2752 4787
rect 2818 4753 2852 4787
rect 2918 4753 2952 4787
rect 3018 4753 3052 4787
rect 3118 4753 3146 4787
rect 3146 4753 3152 4787
rect 3218 4753 3224 4787
rect 3224 4753 3252 4787
rect 3318 4753 3352 4787
rect 3418 4753 3446 4787
rect 3446 4753 3452 4787
rect 3518 4753 3524 4787
rect 3524 4753 3552 4787
rect 3618 4753 3652 4787
rect 3718 4753 3752 4787
rect 3818 4753 3852 4787
rect 3918 4753 3952 4787
rect 4018 4753 4052 4787
rect 4118 4753 4152 4787
rect 4218 4753 4246 4787
rect 4246 4753 4252 4787
rect 4318 4753 4324 4787
rect 4324 4753 4352 4787
rect 4418 4753 4452 4787
rect 4518 4753 4552 4787
rect 4618 4753 4652 4787
rect 4718 4753 4752 4787
rect 4818 4753 4852 4787
rect 4918 4753 4952 4787
rect 5018 4753 5052 4787
rect 5118 4753 5152 4787
rect 5218 4753 5252 4787
rect 5318 4753 5352 4787
rect 5418 4753 5452 4787
rect 5518 4753 5552 4787
rect 5618 4753 5652 4787
rect 5718 4753 5752 4787
rect 5818 4753 5852 4787
rect 5918 4753 5952 4787
rect 6018 4753 6052 4787
rect 6118 4753 6152 4787
rect 6218 4753 6252 4787
rect 6318 4753 6352 4787
rect 6418 4753 6446 4787
rect 6446 4753 6452 4787
rect 6518 4753 6524 4787
rect 6524 4753 6552 4787
rect 6618 4753 6652 4787
rect 6718 4753 6752 4787
rect 6818 4753 6852 4787
rect 6918 4753 6952 4787
rect 7018 4753 7052 4787
rect 7118 4753 7152 4787
rect 7218 4753 7252 4787
rect 7318 4753 7352 4787
rect 7418 4753 7452 4787
rect 7518 4753 7552 4787
rect 7618 4753 7652 4787
rect 7718 4753 7752 4787
rect 7818 4753 7852 4787
rect 7918 4753 7952 4787
rect 8018 4753 8052 4787
rect 8118 4753 8152 4787
rect 8218 4753 8252 4787
rect 8318 4753 8352 4787
rect 8418 4753 8452 4787
rect 8518 4753 8552 4787
rect 8618 4753 8652 4787
rect 8718 4753 8752 4787
rect 8818 4753 8852 4787
rect 8918 4753 8952 4787
rect 9018 4753 9052 4787
rect 9118 4753 9152 4787
rect 9218 4753 9252 4787
rect 9318 4753 9352 4787
rect 9418 4753 9452 4787
rect 9518 4753 9552 4787
rect 9618 4753 9652 4787
rect 9718 4753 9752 4787
rect 9818 4753 9846 4787
rect 9846 4753 9852 4787
rect 9918 4753 9924 4787
rect 9924 4753 9952 4787
rect 10018 4753 10052 4787
rect 10118 4753 10152 4787
rect 10218 4753 10252 4787
rect 10318 4753 10352 4787
rect 10418 4753 10452 4787
rect 10518 4753 10552 4787
rect 10618 4753 10652 4787
rect 10718 4753 10746 4787
rect 10746 4753 10752 4787
rect 10818 4753 10824 4787
rect 10824 4753 10852 4787
rect 10918 4753 10952 4787
rect 11018 4753 11052 4787
rect 11118 4753 11152 4787
rect 11218 4753 11252 4787
rect 11318 4753 11352 4787
rect 11418 4753 11452 4787
rect 11518 4753 11552 4787
rect 11618 4753 11646 4787
rect 11646 4753 11652 4787
rect 11718 4753 11724 4787
rect 11724 4753 11752 4787
rect 11818 4753 11852 4787
rect 11918 4753 11952 4787
rect 12018 4753 12052 4787
rect 12118 4753 12152 4787
rect 12218 4753 12252 4787
rect 12318 4753 12352 4787
rect 12418 4753 12446 4787
rect 12446 4753 12452 4787
rect 12518 4753 12524 4787
rect 12524 4753 12552 4787
rect 12618 4753 12652 4787
rect 12718 4753 12752 4787
rect 12818 4753 12846 4787
rect 12846 4753 12852 4787
rect 12916 4768 12924 4802
rect 12924 4768 12950 4802
rect 13120 4738 13146 4772
rect 13146 4738 13154 4772
rect 18 4613 52 4647
rect 118 4613 152 4647
rect 218 4613 252 4647
rect 318 4613 352 4647
rect 418 4613 452 4647
rect 518 4613 552 4647
rect 618 4613 652 4647
rect 718 4613 752 4647
rect 818 4613 852 4647
rect 918 4613 952 4647
rect 1018 4613 1052 4647
rect 1118 4613 1146 4647
rect 1146 4613 1152 4647
rect 1218 4613 1224 4647
rect 1224 4613 1252 4647
rect 1318 4613 1352 4647
rect 1418 4613 1452 4647
rect 1518 4613 1552 4647
rect 1618 4613 1652 4647
rect 1718 4613 1752 4647
rect 1818 4613 1852 4647
rect 1918 4613 1952 4647
rect 2018 4613 2052 4647
rect 2118 4613 2152 4647
rect 2218 4613 2252 4647
rect 2318 4613 2352 4647
rect 2418 4613 2452 4647
rect 2518 4613 2552 4647
rect 2618 4613 2652 4647
rect 2718 4613 2752 4647
rect 2818 4613 2852 4647
rect 2918 4613 2946 4647
rect 2946 4613 2952 4647
rect 3018 4613 3024 4647
rect 3024 4613 3052 4647
rect 3118 4613 3152 4647
rect 3218 4613 3252 4647
rect 3318 4613 3352 4647
rect 3418 4613 3452 4647
rect 3518 4613 3552 4647
rect 3618 4613 3646 4647
rect 3646 4613 3652 4647
rect 3718 4613 3724 4647
rect 3724 4613 3752 4647
rect 3818 4613 3852 4647
rect 3918 4613 3952 4647
rect 4018 4613 4052 4647
rect 4118 4613 4152 4647
rect 4218 4613 4252 4647
rect 4318 4613 4352 4647
rect 4418 4613 4452 4647
rect 4518 4613 4552 4647
rect 4618 4613 4652 4647
rect 4718 4613 4746 4647
rect 4746 4613 4752 4647
rect 4818 4613 4824 4647
rect 4824 4613 4852 4647
rect 4918 4613 4952 4647
rect 5018 4613 5046 4647
rect 5046 4613 5052 4647
rect 5118 4613 5124 4647
rect 5124 4613 5152 4647
rect 5218 4613 5252 4647
rect 5318 4613 5352 4647
rect 5418 4613 5452 4647
rect 5518 4613 5552 4647
rect 5618 4613 5652 4647
rect 5718 4613 5752 4647
rect 5818 4613 5846 4647
rect 5846 4613 5852 4647
rect 5918 4613 5924 4647
rect 5924 4613 5952 4647
rect 6018 4613 6052 4647
rect 6118 4613 6152 4647
rect 6218 4613 6252 4647
rect 6318 4613 6352 4647
rect 6418 4613 6446 4647
rect 6446 4613 6452 4647
rect 6518 4613 6524 4647
rect 6524 4613 6552 4647
rect 6618 4613 6652 4647
rect 6718 4613 6752 4647
rect 6818 4613 6852 4647
rect 6918 4613 6952 4647
rect 7018 4613 7052 4647
rect 7118 4613 7152 4647
rect 7218 4613 7252 4647
rect 7318 4613 7352 4647
rect 7418 4613 7452 4647
rect 7518 4613 7552 4647
rect 7618 4613 7652 4647
rect 7718 4613 7752 4647
rect 7818 4613 7852 4647
rect 7918 4613 7952 4647
rect 8018 4613 8052 4647
rect 8118 4613 8152 4647
rect 8218 4613 8252 4647
rect 8318 4613 8352 4647
rect 8418 4613 8452 4647
rect 8518 4613 8552 4647
rect 8618 4613 8652 4647
rect 8718 4613 8746 4647
rect 8746 4613 8752 4647
rect 8818 4613 8824 4647
rect 8824 4613 8852 4647
rect 8918 4613 8952 4647
rect 9018 4613 9052 4647
rect 9118 4613 9152 4647
rect 9218 4613 9252 4647
rect 9318 4613 9352 4647
rect 9418 4613 9452 4647
rect 9518 4613 9552 4647
rect 9618 4613 9652 4647
rect 9718 4613 9752 4647
rect 9818 4613 9852 4647
rect 9918 4613 9952 4647
rect 10018 4613 10052 4647
rect 10118 4613 10152 4647
rect 10218 4613 10252 4647
rect 10318 4613 10352 4647
rect 10418 4613 10452 4647
rect 10518 4613 10552 4647
rect 10618 4613 10652 4647
rect 10718 4613 10752 4647
rect 10818 4613 10852 4647
rect 10918 4613 10952 4647
rect 11018 4613 11052 4647
rect 11118 4613 11152 4647
rect 11218 4613 11252 4647
rect 11318 4613 11352 4647
rect 11418 4613 11452 4647
rect 11518 4613 11552 4647
rect 11618 4613 11652 4647
rect 11718 4613 11752 4647
rect 11818 4613 11852 4647
rect 11918 4613 11952 4647
rect 12018 4613 12052 4647
rect 12118 4613 12152 4647
rect 12218 4613 12252 4647
rect 12318 4613 12352 4647
rect 12418 4613 12452 4647
rect 12518 4613 12552 4647
rect 12618 4613 12646 4647
rect 12646 4613 12652 4647
rect 12718 4613 12724 4647
rect 12724 4613 12752 4647
rect 12818 4613 12846 4647
rect 12846 4613 12852 4647
rect 12916 4628 12924 4662
rect 12924 4628 12950 4662
rect 13120 4598 13146 4632
rect 13146 4598 13154 4632
rect 18 4473 52 4507
rect 118 4473 152 4507
rect 218 4473 252 4507
rect 318 4473 346 4507
rect 346 4473 352 4507
rect 418 4473 424 4507
rect 424 4473 452 4507
rect 518 4473 552 4507
rect 618 4473 652 4507
rect 718 4473 752 4507
rect 818 4473 852 4507
rect 918 4473 952 4507
rect 1018 4473 1052 4507
rect 1118 4473 1152 4507
rect 1218 4473 1252 4507
rect 1318 4473 1352 4507
rect 1418 4473 1452 4507
rect 1518 4473 1552 4507
rect 1618 4473 1646 4507
rect 1646 4473 1652 4507
rect 1718 4473 1724 4507
rect 1724 4473 1752 4507
rect 1818 4473 1846 4507
rect 1846 4473 1852 4507
rect 1918 4473 1924 4507
rect 1924 4473 1952 4507
rect 2018 4473 2052 4507
rect 2118 4473 2152 4507
rect 2218 4473 2252 4507
rect 2318 4473 2346 4507
rect 2346 4473 2352 4507
rect 2418 4473 2424 4507
rect 2424 4473 2452 4507
rect 2518 4473 2552 4507
rect 2618 4473 2646 4507
rect 2646 4473 2652 4507
rect 2718 4473 2724 4507
rect 2724 4473 2752 4507
rect 2818 4473 2846 4507
rect 2846 4473 2852 4507
rect 2918 4473 2924 4507
rect 2924 4473 2952 4507
rect 3018 4473 3052 4507
rect 3118 4473 3152 4507
rect 3218 4473 3252 4507
rect 3318 4473 3352 4507
rect 3418 4473 3452 4507
rect 3518 4473 3552 4507
rect 3618 4473 3652 4507
rect 3718 4473 3746 4507
rect 3746 4473 3752 4507
rect 3818 4473 3824 4507
rect 3824 4473 3852 4507
rect 3918 4473 3952 4507
rect 4018 4473 4052 4507
rect 4118 4473 4152 4507
rect 4218 4473 4252 4507
rect 4318 4473 4352 4507
rect 4418 4473 4452 4507
rect 4518 4473 4552 4507
rect 4618 4473 4652 4507
rect 4718 4473 4752 4507
rect 4818 4473 4852 4507
rect 4918 4473 4952 4507
rect 5018 4473 5046 4507
rect 5046 4473 5052 4507
rect 5118 4473 5124 4507
rect 5124 4473 5152 4507
rect 5218 4473 5252 4507
rect 5318 4473 5346 4507
rect 5346 4473 5352 4507
rect 5418 4473 5424 4507
rect 5424 4473 5452 4507
rect 5518 4473 5552 4507
rect 5618 4473 5652 4507
rect 5718 4473 5752 4507
rect 5818 4473 5852 4507
rect 5918 4473 5952 4507
rect 6018 4473 6046 4507
rect 6046 4473 6052 4507
rect 6118 4473 6124 4507
rect 6124 4473 6152 4507
rect 6218 4473 6252 4507
rect 6318 4473 6352 4507
rect 6418 4473 6452 4507
rect 6518 4473 6552 4507
rect 6618 4473 6652 4507
rect 6718 4473 6752 4507
rect 6818 4473 6852 4507
rect 6918 4473 6952 4507
rect 7018 4473 7052 4507
rect 7118 4473 7152 4507
rect 7218 4473 7252 4507
rect 7318 4473 7352 4507
rect 7418 4473 7452 4507
rect 7518 4473 7552 4507
rect 7618 4473 7652 4507
rect 7718 4473 7752 4507
rect 7818 4473 7852 4507
rect 7918 4473 7952 4507
rect 8018 4473 8046 4507
rect 8046 4473 8052 4507
rect 8118 4473 8124 4507
rect 8124 4473 8152 4507
rect 8218 4473 8252 4507
rect 8318 4473 8346 4507
rect 8346 4473 8352 4507
rect 8418 4473 8424 4507
rect 8424 4473 8452 4507
rect 8518 4473 8552 4507
rect 8618 4473 8652 4507
rect 8718 4473 8752 4507
rect 8818 4473 8846 4507
rect 8846 4473 8852 4507
rect 8918 4473 8924 4507
rect 8924 4473 8952 4507
rect 9018 4473 9046 4507
rect 9046 4473 9052 4507
rect 9118 4473 9124 4507
rect 9124 4473 9152 4507
rect 9218 4473 9252 4507
rect 9318 4473 9346 4507
rect 9346 4473 9352 4507
rect 9418 4473 9424 4507
rect 9424 4473 9452 4507
rect 9518 4473 9552 4507
rect 9618 4473 9646 4507
rect 9646 4473 9652 4507
rect 9718 4473 9724 4507
rect 9724 4473 9752 4507
rect 9818 4473 9852 4507
rect 9918 4473 9946 4507
rect 9946 4473 9952 4507
rect 10018 4473 10024 4507
rect 10024 4473 10052 4507
rect 10118 4473 10152 4507
rect 10218 4473 10246 4507
rect 10246 4473 10252 4507
rect 10318 4473 10324 4507
rect 10324 4473 10352 4507
rect 10418 4473 10452 4507
rect 10518 4473 10546 4507
rect 10546 4473 10552 4507
rect 10618 4473 10624 4507
rect 10624 4473 10652 4507
rect 10718 4473 10746 4507
rect 10746 4473 10752 4507
rect 10818 4473 10824 4507
rect 10824 4473 10852 4507
rect 10918 4473 10946 4507
rect 10946 4473 10952 4507
rect 11018 4473 11024 4507
rect 11024 4473 11052 4507
rect 11118 4473 11152 4507
rect 11218 4473 11246 4507
rect 11246 4473 11252 4507
rect 11318 4473 11324 4507
rect 11324 4473 11352 4507
rect 11418 4473 11452 4507
rect 11518 4473 11552 4507
rect 11618 4473 11652 4507
rect 11718 4473 11752 4507
rect 11818 4473 11852 4507
rect 11918 4473 11952 4507
rect 12018 4473 12052 4507
rect 12118 4473 12152 4507
rect 12218 4473 12252 4507
rect 12318 4473 12352 4507
rect 12418 4473 12446 4507
rect 12446 4473 12452 4507
rect 12518 4473 12524 4507
rect 12524 4473 12552 4507
rect 12618 4473 12652 4507
rect 12718 4473 12752 4507
rect 12818 4473 12846 4507
rect 12846 4473 12852 4507
rect 12916 4488 12924 4522
rect 12924 4488 12950 4522
rect 13120 4458 13146 4492
rect 13146 4458 13154 4492
rect 18 4333 24 4367
rect 24 4333 52 4367
rect 118 4333 152 4367
rect 218 4333 252 4367
rect 318 4333 352 4367
rect 418 4333 452 4367
rect 518 4333 552 4367
rect 618 4333 652 4367
rect 718 4333 752 4367
rect 818 4333 852 4367
rect 918 4333 952 4367
rect 1018 4333 1052 4367
rect 1118 4333 1152 4367
rect 1218 4333 1246 4367
rect 1246 4333 1252 4367
rect 1318 4333 1324 4367
rect 1324 4333 1352 4367
rect 1418 4333 1452 4367
rect 1518 4333 1552 4367
rect 1618 4333 1652 4367
rect 1718 4333 1752 4367
rect 1818 4333 1852 4367
rect 1918 4333 1946 4367
rect 1946 4333 1952 4367
rect 2018 4333 2024 4367
rect 2024 4333 2052 4367
rect 2118 4333 2152 4367
rect 2218 4333 2252 4367
rect 2318 4333 2352 4367
rect 2418 4333 2452 4367
rect 2518 4333 2552 4367
rect 2618 4333 2652 4367
rect 2718 4333 2752 4367
rect 2818 4333 2852 4367
rect 2918 4333 2952 4367
rect 3018 4333 3052 4367
rect 3118 4333 3152 4367
rect 3218 4333 3252 4367
rect 3318 4333 3352 4367
rect 3418 4333 3452 4367
rect 3518 4333 3552 4367
rect 3618 4333 3652 4367
rect 3718 4333 3746 4367
rect 3746 4333 3752 4367
rect 3818 4333 3824 4367
rect 3824 4333 3852 4367
rect 3918 4333 3952 4367
rect 4018 4333 4052 4367
rect 4118 4333 4152 4367
rect 4218 4333 4252 4367
rect 4318 4333 4352 4367
rect 4418 4333 4452 4367
rect 4518 4333 4552 4367
rect 4618 4333 4652 4367
rect 4718 4333 4752 4367
rect 4818 4333 4852 4367
rect 4918 4333 4952 4367
rect 5018 4333 5052 4367
rect 5118 4333 5152 4367
rect 5218 4333 5252 4367
rect 5318 4333 5352 4367
rect 5418 4333 5452 4367
rect 5518 4333 5552 4367
rect 5618 4333 5652 4367
rect 5718 4333 5752 4367
rect 5818 4333 5852 4367
rect 5918 4333 5952 4367
rect 6018 4333 6046 4367
rect 6046 4333 6052 4367
rect 6118 4333 6124 4367
rect 6124 4333 6152 4367
rect 6218 4333 6252 4367
rect 6318 4333 6352 4367
rect 6418 4333 6452 4367
rect 6518 4333 6552 4367
rect 6618 4333 6646 4367
rect 6646 4333 6652 4367
rect 6718 4333 6724 4367
rect 6724 4333 6752 4367
rect 6818 4333 6852 4367
rect 6918 4333 6952 4367
rect 7018 4333 7052 4367
rect 7118 4333 7152 4367
rect 7218 4333 7252 4367
rect 7318 4333 7346 4367
rect 7346 4333 7352 4367
rect 7418 4333 7424 4367
rect 7424 4333 7452 4367
rect 7518 4333 7552 4367
rect 7618 4333 7652 4367
rect 7718 4333 7752 4367
rect 7818 4333 7852 4367
rect 7918 4333 7952 4367
rect 8018 4333 8052 4367
rect 8118 4333 8152 4367
rect 8218 4333 8252 4367
rect 8318 4333 8352 4367
rect 8418 4333 8452 4367
rect 8518 4333 8552 4367
rect 8618 4333 8652 4367
rect 8718 4333 8752 4367
rect 8818 4333 8852 4367
rect 8918 4333 8952 4367
rect 9018 4333 9052 4367
rect 9118 4333 9152 4367
rect 9218 4333 9252 4367
rect 9318 4333 9352 4367
rect 9418 4333 9452 4367
rect 9518 4333 9552 4367
rect 9618 4333 9652 4367
rect 9718 4333 9752 4367
rect 9818 4333 9852 4367
rect 9918 4333 9952 4367
rect 10018 4333 10052 4367
rect 10118 4333 10152 4367
rect 10218 4333 10252 4367
rect 10318 4333 10352 4367
rect 10418 4333 10452 4367
rect 10518 4333 10552 4367
rect 10618 4333 10652 4367
rect 10718 4333 10752 4367
rect 10818 4333 10846 4367
rect 10846 4333 10852 4367
rect 10918 4333 10924 4367
rect 10924 4333 10952 4367
rect 11018 4333 11052 4367
rect 11118 4333 11146 4367
rect 11146 4333 11152 4367
rect 11218 4333 11224 4367
rect 11224 4333 11252 4367
rect 11318 4333 11352 4367
rect 11418 4333 11452 4367
rect 11518 4333 11552 4367
rect 11618 4333 11652 4367
rect 11718 4333 11752 4367
rect 11818 4333 11852 4367
rect 11918 4333 11946 4367
rect 11946 4333 11952 4367
rect 12018 4333 12024 4367
rect 12024 4333 12052 4367
rect 12118 4333 12152 4367
rect 12218 4333 12252 4367
rect 12318 4333 12352 4367
rect 12418 4333 12452 4367
rect 12518 4333 12552 4367
rect 12618 4333 12652 4367
rect 12718 4333 12752 4367
rect 12818 4333 12846 4367
rect 12846 4333 12852 4367
rect 12916 4348 12924 4382
rect 12924 4348 12950 4382
rect 13120 4318 13146 4352
rect 13146 4318 13154 4352
rect 18 4193 52 4227
rect 118 4193 152 4227
rect 218 4193 252 4227
rect 318 4193 352 4227
rect 418 4193 452 4227
rect 518 4193 546 4227
rect 546 4193 552 4227
rect 618 4193 624 4227
rect 624 4193 652 4227
rect 718 4193 752 4227
rect 818 4193 852 4227
rect 918 4193 952 4227
rect 1018 4193 1052 4227
rect 1118 4193 1146 4227
rect 1146 4193 1152 4227
rect 1218 4193 1224 4227
rect 1224 4193 1252 4227
rect 1318 4193 1352 4227
rect 1418 4193 1452 4227
rect 1518 4193 1552 4227
rect 1618 4193 1652 4227
rect 1718 4193 1752 4227
rect 1818 4193 1852 4227
rect 1918 4193 1946 4227
rect 1946 4193 1952 4227
rect 2018 4193 2024 4227
rect 2024 4193 2052 4227
rect 2118 4193 2152 4227
rect 2218 4193 2252 4227
rect 2318 4193 2352 4227
rect 2418 4193 2452 4227
rect 2518 4193 2552 4227
rect 2618 4193 2652 4227
rect 2718 4193 2752 4227
rect 2818 4193 2852 4227
rect 2918 4193 2952 4227
rect 3018 4193 3052 4227
rect 3118 4193 3152 4227
rect 3218 4193 3252 4227
rect 3318 4193 3352 4227
rect 3418 4193 3452 4227
rect 3518 4193 3552 4227
rect 3618 4193 3652 4227
rect 3718 4193 3752 4227
rect 3818 4193 3852 4227
rect 3918 4193 3952 4227
rect 4018 4193 4046 4227
rect 4046 4193 4052 4227
rect 4118 4193 4124 4227
rect 4124 4193 4152 4227
rect 4218 4193 4246 4227
rect 4246 4193 4252 4227
rect 4318 4193 4324 4227
rect 4324 4193 4352 4227
rect 4418 4193 4446 4227
rect 4446 4193 4452 4227
rect 4518 4193 4524 4227
rect 4524 4193 4552 4227
rect 4618 4193 4646 4227
rect 4646 4193 4652 4227
rect 4718 4193 4724 4227
rect 4724 4193 4752 4227
rect 4818 4193 4846 4227
rect 4846 4193 4852 4227
rect 4918 4193 4924 4227
rect 4924 4193 4952 4227
rect 5018 4193 5052 4227
rect 5118 4193 5152 4227
rect 5218 4193 5252 4227
rect 5318 4193 5352 4227
rect 5418 4193 5452 4227
rect 5518 4193 5546 4227
rect 5546 4193 5552 4227
rect 5618 4193 5624 4227
rect 5624 4193 5652 4227
rect 5718 4193 5752 4227
rect 5818 4193 5852 4227
rect 5918 4193 5952 4227
rect 6018 4193 6046 4227
rect 6046 4193 6052 4227
rect 6118 4193 6124 4227
rect 6124 4193 6152 4227
rect 6218 4193 6246 4227
rect 6246 4193 6252 4227
rect 6318 4193 6324 4227
rect 6324 4193 6352 4227
rect 6418 4193 6446 4227
rect 6446 4193 6452 4227
rect 6518 4193 6524 4227
rect 6524 4193 6552 4227
rect 6618 4193 6646 4227
rect 6646 4193 6652 4227
rect 6718 4193 6724 4227
rect 6724 4193 6752 4227
rect 6818 4193 6852 4227
rect 6918 4193 6952 4227
rect 7018 4193 7052 4227
rect 7118 4193 7146 4227
rect 7146 4193 7152 4227
rect 7218 4193 7224 4227
rect 7224 4193 7252 4227
rect 7318 4193 7352 4227
rect 7418 4193 7452 4227
rect 7518 4193 7552 4227
rect 7618 4193 7652 4227
rect 7718 4193 7752 4227
rect 7818 4193 7852 4227
rect 7918 4193 7952 4227
rect 8018 4193 8052 4227
rect 8118 4193 8146 4227
rect 8146 4193 8152 4227
rect 8218 4193 8224 4227
rect 8224 4193 8252 4227
rect 8318 4193 8346 4227
rect 8346 4193 8352 4227
rect 8418 4193 8424 4227
rect 8424 4193 8452 4227
rect 8518 4193 8546 4227
rect 8546 4193 8552 4227
rect 8618 4193 8624 4227
rect 8624 4193 8652 4227
rect 8718 4193 8746 4227
rect 8746 4193 8752 4227
rect 8818 4193 8824 4227
rect 8824 4193 8852 4227
rect 8918 4193 8946 4227
rect 8946 4193 8952 4227
rect 9018 4193 9024 4227
rect 9024 4193 9052 4227
rect 9118 4193 9152 4227
rect 9218 4193 9252 4227
rect 9318 4193 9346 4227
rect 9346 4193 9352 4227
rect 9418 4193 9424 4227
rect 9424 4193 9452 4227
rect 9518 4193 9546 4227
rect 9546 4193 9552 4227
rect 9618 4193 9624 4227
rect 9624 4193 9652 4227
rect 9718 4193 9746 4227
rect 9746 4193 9752 4227
rect 9818 4193 9824 4227
rect 9824 4193 9852 4227
rect 9918 4193 9952 4227
rect 10018 4193 10046 4227
rect 10046 4193 10052 4227
rect 10118 4193 10124 4227
rect 10124 4193 10152 4227
rect 10218 4193 10252 4227
rect 10318 4193 10352 4227
rect 10418 4193 10452 4227
rect 10518 4193 10552 4227
rect 10618 4193 10652 4227
rect 10718 4193 10752 4227
rect 10818 4193 10852 4227
rect 10918 4193 10946 4227
rect 10946 4193 10952 4227
rect 11018 4193 11024 4227
rect 11024 4193 11052 4227
rect 11118 4193 11152 4227
rect 11218 4193 11252 4227
rect 11318 4193 11346 4227
rect 11346 4193 11352 4227
rect 11418 4193 11424 4227
rect 11424 4193 11452 4227
rect 11518 4193 11546 4227
rect 11546 4193 11552 4227
rect 11618 4193 11624 4227
rect 11624 4193 11652 4227
rect 11718 4193 11752 4227
rect 11818 4193 11852 4227
rect 11918 4193 11952 4227
rect 12018 4193 12052 4227
rect 12118 4193 12152 4227
rect 12218 4193 12252 4227
rect 12318 4193 12352 4227
rect 12418 4193 12452 4227
rect 12518 4193 12552 4227
rect 12618 4193 12652 4227
rect 12718 4193 12752 4227
rect 12818 4193 12852 4227
rect 12916 4208 12924 4242
rect 12924 4208 12950 4242
rect 13120 4178 13146 4212
rect 13146 4178 13154 4212
rect 18 4053 24 4087
rect 24 4053 52 4087
rect 118 4053 152 4087
rect 218 4053 246 4087
rect 246 4053 252 4087
rect 318 4053 324 4087
rect 324 4053 352 4087
rect 418 4053 446 4087
rect 446 4053 452 4087
rect 518 4053 524 4087
rect 524 4053 552 4087
rect 618 4053 652 4087
rect 718 4053 752 4087
rect 818 4053 852 4087
rect 918 4053 952 4087
rect 1018 4053 1052 4087
rect 1118 4053 1152 4087
rect 1218 4053 1252 4087
rect 1318 4053 1346 4087
rect 1346 4053 1352 4087
rect 1418 4053 1424 4087
rect 1424 4053 1452 4087
rect 1518 4053 1552 4087
rect 1618 4053 1646 4087
rect 1646 4053 1652 4087
rect 1718 4053 1724 4087
rect 1724 4053 1752 4087
rect 1818 4053 1852 4087
rect 1918 4053 1952 4087
rect 2018 4053 2052 4087
rect 2118 4053 2152 4087
rect 2218 4053 2246 4087
rect 2246 4053 2252 4087
rect 2318 4053 2324 4087
rect 2324 4053 2352 4087
rect 2418 4053 2452 4087
rect 2518 4053 2552 4087
rect 2618 4053 2646 4087
rect 2646 4053 2652 4087
rect 2718 4053 2724 4087
rect 2724 4053 2752 4087
rect 2818 4053 2852 4087
rect 2918 4053 2946 4087
rect 2946 4053 2952 4087
rect 3018 4053 3024 4087
rect 3024 4053 3052 4087
rect 3118 4053 3152 4087
rect 3218 4053 3246 4087
rect 3246 4053 3252 4087
rect 3318 4053 3324 4087
rect 3324 4053 3352 4087
rect 3418 4053 3452 4087
rect 3518 4053 3552 4087
rect 3618 4053 3652 4087
rect 3718 4053 3752 4087
rect 3818 4053 3852 4087
rect 3918 4053 3952 4087
rect 4018 4053 4052 4087
rect 4118 4053 4146 4087
rect 4146 4053 4152 4087
rect 4218 4053 4224 4087
rect 4224 4053 4252 4087
rect 4318 4053 4346 4087
rect 4346 4053 4352 4087
rect 4418 4053 4424 4087
rect 4424 4053 4452 4087
rect 4518 4053 4546 4087
rect 4546 4053 4552 4087
rect 4618 4053 4624 4087
rect 4624 4053 4652 4087
rect 4718 4053 4746 4087
rect 4746 4053 4752 4087
rect 4818 4053 4824 4087
rect 4824 4053 4852 4087
rect 4918 4053 4946 4087
rect 4946 4053 4952 4087
rect 5018 4053 5024 4087
rect 5024 4053 5052 4087
rect 5118 4053 5152 4087
rect 5218 4053 5246 4087
rect 5246 4053 5252 4087
rect 5318 4053 5324 4087
rect 5324 4053 5352 4087
rect 5418 4053 5452 4087
rect 5518 4053 5552 4087
rect 5618 4053 5646 4087
rect 5646 4053 5652 4087
rect 5718 4053 5724 4087
rect 5724 4053 5752 4087
rect 5818 4053 5852 4087
rect 5918 4053 5952 4087
rect 6018 4053 6052 4087
rect 6118 4053 6152 4087
rect 6218 4053 6252 4087
rect 6318 4053 6352 4087
rect 6418 4053 6452 4087
rect 6518 4053 6552 4087
rect 6618 4053 6652 4087
rect 6718 4053 6752 4087
rect 6818 4053 6852 4087
rect 6918 4053 6952 4087
rect 7018 4053 7052 4087
rect 7118 4053 7152 4087
rect 7218 4053 7252 4087
rect 7318 4053 7346 4087
rect 7346 4053 7352 4087
rect 7418 4053 7424 4087
rect 7424 4053 7452 4087
rect 7518 4053 7552 4087
rect 7618 4053 7646 4087
rect 7646 4053 7652 4087
rect 7718 4053 7724 4087
rect 7724 4053 7752 4087
rect 7818 4053 7846 4087
rect 7846 4053 7852 4087
rect 7918 4053 7924 4087
rect 7924 4053 7952 4087
rect 8018 4053 8052 4087
rect 8118 4053 8152 4087
rect 8218 4053 8252 4087
rect 8318 4053 8352 4087
rect 8418 4053 8452 4087
rect 8518 4053 8552 4087
rect 8618 4053 8652 4087
rect 8718 4053 8746 4087
rect 8746 4053 8752 4087
rect 8818 4053 8824 4087
rect 8824 4053 8852 4087
rect 8918 4053 8946 4087
rect 8946 4053 8952 4087
rect 9018 4053 9024 4087
rect 9024 4053 9052 4087
rect 9118 4053 9152 4087
rect 9218 4053 9252 4087
rect 9318 4053 9352 4087
rect 9418 4053 9452 4087
rect 9518 4053 9546 4087
rect 9546 4053 9552 4087
rect 9618 4053 9624 4087
rect 9624 4053 9652 4087
rect 9718 4053 9752 4087
rect 9818 4053 9852 4087
rect 9918 4053 9952 4087
rect 10018 4053 10052 4087
rect 10118 4053 10152 4087
rect 10218 4053 10252 4087
rect 10318 4053 10352 4087
rect 10418 4053 10452 4087
rect 10518 4053 10552 4087
rect 10618 4053 10646 4087
rect 10646 4053 10652 4087
rect 10718 4053 10724 4087
rect 10724 4053 10752 4087
rect 10818 4053 10846 4087
rect 10846 4053 10852 4087
rect 10918 4053 10924 4087
rect 10924 4053 10952 4087
rect 11018 4053 11052 4087
rect 11118 4053 11152 4087
rect 11218 4053 11252 4087
rect 11318 4053 11346 4087
rect 11346 4053 11352 4087
rect 11418 4053 11424 4087
rect 11424 4053 11452 4087
rect 11518 4053 11546 4087
rect 11546 4053 11552 4087
rect 11618 4053 11624 4087
rect 11624 4053 11652 4087
rect 11718 4053 11752 4087
rect 11818 4053 11846 4087
rect 11846 4053 11852 4087
rect 11918 4053 11924 4087
rect 11924 4053 11952 4087
rect 12018 4053 12052 4087
rect 12118 4053 12152 4087
rect 12218 4053 12252 4087
rect 12318 4053 12352 4087
rect 12418 4053 12452 4087
rect 12518 4053 12552 4087
rect 12618 4053 12646 4087
rect 12646 4053 12652 4087
rect 12718 4053 12724 4087
rect 12724 4053 12752 4087
rect 12818 4053 12846 4087
rect 12846 4053 12852 4087
rect 12916 4068 12924 4102
rect 12924 4068 12950 4102
rect 13120 4038 13146 4072
rect 13146 4038 13154 4072
rect 18 3913 24 3947
rect 24 3913 52 3947
rect 118 3913 152 3947
rect 218 3913 252 3947
rect 318 3913 352 3947
rect 418 3913 452 3947
rect 518 3913 552 3947
rect 618 3913 652 3947
rect 718 3913 752 3947
rect 818 3913 852 3947
rect 918 3913 952 3947
rect 1018 3913 1052 3947
rect 1118 3913 1152 3947
rect 1218 3913 1252 3947
rect 1318 3913 1352 3947
rect 1418 3913 1452 3947
rect 1518 3913 1552 3947
rect 1618 3913 1652 3947
rect 1718 3913 1752 3947
rect 1818 3913 1852 3947
rect 1918 3913 1946 3947
rect 1946 3913 1952 3947
rect 2018 3913 2024 3947
rect 2024 3913 2052 3947
rect 2118 3913 2152 3947
rect 2218 3913 2252 3947
rect 2318 3913 2352 3947
rect 2418 3913 2452 3947
rect 2518 3913 2552 3947
rect 2618 3913 2652 3947
rect 2718 3913 2752 3947
rect 2818 3913 2852 3947
rect 2918 3913 2952 3947
rect 3018 3913 3052 3947
rect 3118 3913 3152 3947
rect 3218 3913 3252 3947
rect 3318 3913 3352 3947
rect 3418 3913 3452 3947
rect 3518 3913 3552 3947
rect 3618 3913 3652 3947
rect 3718 3913 3752 3947
rect 3818 3913 3852 3947
rect 3918 3913 3946 3947
rect 3946 3913 3952 3947
rect 4018 3913 4024 3947
rect 4024 3913 4052 3947
rect 4118 3913 4146 3947
rect 4146 3913 4152 3947
rect 4218 3913 4224 3947
rect 4224 3913 4252 3947
rect 4318 3913 4352 3947
rect 4418 3913 4452 3947
rect 4518 3913 4552 3947
rect 4618 3913 4652 3947
rect 4718 3913 4752 3947
rect 4818 3913 4852 3947
rect 4918 3913 4952 3947
rect 5018 3913 5046 3947
rect 5046 3913 5052 3947
rect 5118 3913 5124 3947
rect 5124 3913 5152 3947
rect 5218 3913 5246 3947
rect 5246 3913 5252 3947
rect 5318 3913 5324 3947
rect 5324 3913 5352 3947
rect 5418 3913 5452 3947
rect 5518 3913 5546 3947
rect 5546 3913 5552 3947
rect 5618 3913 5624 3947
rect 5624 3913 5652 3947
rect 5718 3913 5752 3947
rect 5818 3913 5852 3947
rect 5918 3913 5946 3947
rect 5946 3913 5952 3947
rect 6018 3913 6024 3947
rect 6024 3913 6052 3947
rect 6118 3913 6152 3947
rect 6218 3913 6252 3947
rect 6318 3913 6352 3947
rect 6418 3913 6452 3947
rect 6518 3913 6552 3947
rect 6618 3913 6652 3947
rect 6718 3913 6752 3947
rect 6818 3913 6852 3947
rect 6918 3913 6946 3947
rect 6946 3913 6952 3947
rect 7018 3913 7024 3947
rect 7024 3913 7052 3947
rect 7118 3913 7146 3947
rect 7146 3913 7152 3947
rect 7218 3913 7224 3947
rect 7224 3913 7252 3947
rect 7318 3913 7352 3947
rect 7418 3913 7452 3947
rect 7518 3913 7552 3947
rect 7618 3913 7652 3947
rect 7718 3913 7752 3947
rect 7818 3913 7852 3947
rect 7918 3913 7952 3947
rect 8018 3913 8052 3947
rect 8118 3913 8152 3947
rect 8218 3913 8252 3947
rect 8318 3913 8352 3947
rect 8418 3913 8452 3947
rect 8518 3913 8552 3947
rect 8618 3913 8652 3947
rect 8718 3913 8746 3947
rect 8746 3913 8752 3947
rect 8818 3913 8824 3947
rect 8824 3913 8852 3947
rect 8918 3913 8952 3947
rect 9018 3913 9052 3947
rect 9118 3913 9152 3947
rect 9218 3913 9252 3947
rect 9318 3913 9352 3947
rect 9418 3913 9452 3947
rect 9518 3913 9546 3947
rect 9546 3913 9552 3947
rect 9618 3913 9624 3947
rect 9624 3913 9652 3947
rect 9718 3913 9752 3947
rect 9818 3913 9852 3947
rect 9918 3913 9952 3947
rect 10018 3913 10052 3947
rect 10118 3913 10152 3947
rect 10218 3913 10252 3947
rect 10318 3913 10352 3947
rect 10418 3913 10452 3947
rect 10518 3913 10552 3947
rect 10618 3913 10652 3947
rect 10718 3913 10752 3947
rect 10818 3913 10852 3947
rect 10918 3913 10952 3947
rect 11018 3913 11046 3947
rect 11046 3913 11052 3947
rect 11118 3913 11124 3947
rect 11124 3913 11152 3947
rect 11218 3913 11252 3947
rect 11318 3913 11352 3947
rect 11418 3913 11452 3947
rect 11518 3913 11552 3947
rect 11618 3913 11652 3947
rect 11718 3913 11752 3947
rect 11818 3913 11852 3947
rect 11918 3913 11952 3947
rect 12018 3913 12052 3947
rect 12118 3913 12152 3947
rect 12218 3913 12252 3947
rect 12318 3913 12352 3947
rect 12418 3913 12452 3947
rect 12518 3913 12552 3947
rect 12618 3913 12652 3947
rect 12718 3913 12752 3947
rect 12818 3913 12846 3947
rect 12846 3913 12852 3947
rect 12916 3928 12924 3962
rect 12924 3928 12950 3962
rect 13120 3898 13146 3932
rect 13146 3898 13154 3932
rect 18 3773 24 3807
rect 24 3773 52 3807
rect 118 3773 152 3807
rect 218 3773 252 3807
rect 318 3773 352 3807
rect 418 3773 452 3807
rect 518 3773 552 3807
rect 618 3773 652 3807
rect 718 3773 752 3807
rect 818 3773 852 3807
rect 918 3773 952 3807
rect 1018 3773 1052 3807
rect 1118 3773 1152 3807
rect 1218 3773 1252 3807
rect 1318 3773 1352 3807
rect 1418 3773 1452 3807
rect 1518 3773 1552 3807
rect 1618 3773 1652 3807
rect 1718 3773 1752 3807
rect 1818 3773 1852 3807
rect 1918 3773 1952 3807
rect 2018 3773 2052 3807
rect 2118 3773 2146 3807
rect 2146 3773 2152 3807
rect 2218 3773 2224 3807
rect 2224 3773 2252 3807
rect 2318 3773 2352 3807
rect 2418 3773 2452 3807
rect 2518 3773 2546 3807
rect 2546 3773 2552 3807
rect 2618 3773 2624 3807
rect 2624 3773 2652 3807
rect 2718 3773 2746 3807
rect 2746 3773 2752 3807
rect 2818 3773 2824 3807
rect 2824 3773 2852 3807
rect 2918 3773 2952 3807
rect 3018 3773 3052 3807
rect 3118 3773 3146 3807
rect 3146 3773 3152 3807
rect 3218 3773 3224 3807
rect 3224 3773 3252 3807
rect 3318 3773 3352 3807
rect 3418 3773 3452 3807
rect 3518 3773 3552 3807
rect 3618 3773 3652 3807
rect 3718 3773 3752 3807
rect 3818 3773 3852 3807
rect 3918 3773 3952 3807
rect 4018 3773 4052 3807
rect 4118 3773 4152 3807
rect 4218 3773 4252 3807
rect 4318 3773 4352 3807
rect 4418 3773 4452 3807
rect 4518 3773 4546 3807
rect 4546 3773 4552 3807
rect 4618 3773 4624 3807
rect 4624 3773 4652 3807
rect 4718 3773 4752 3807
rect 4818 3773 4852 3807
rect 4918 3773 4952 3807
rect 5018 3773 5052 3807
rect 5118 3773 5152 3807
rect 5218 3773 5252 3807
rect 5318 3773 5352 3807
rect 5418 3773 5446 3807
rect 5446 3773 5452 3807
rect 5518 3773 5524 3807
rect 5524 3773 5552 3807
rect 5618 3773 5652 3807
rect 5718 3773 5752 3807
rect 5818 3773 5852 3807
rect 5918 3773 5946 3807
rect 5946 3773 5952 3807
rect 6018 3773 6024 3807
rect 6024 3773 6052 3807
rect 6118 3773 6152 3807
rect 6218 3773 6252 3807
rect 6318 3773 6352 3807
rect 6418 3773 6452 3807
rect 6518 3773 6552 3807
rect 6618 3773 6652 3807
rect 6718 3773 6752 3807
rect 6818 3773 6852 3807
rect 6918 3773 6952 3807
rect 7018 3773 7052 3807
rect 7118 3773 7152 3807
rect 7218 3773 7252 3807
rect 7318 3773 7352 3807
rect 7418 3773 7452 3807
rect 7518 3773 7552 3807
rect 7618 3773 7646 3807
rect 7646 3773 7652 3807
rect 7718 3773 7724 3807
rect 7724 3773 7752 3807
rect 7818 3773 7852 3807
rect 7918 3773 7952 3807
rect 8018 3773 8052 3807
rect 8118 3773 8152 3807
rect 8218 3773 8252 3807
rect 8318 3773 8352 3807
rect 8418 3773 8452 3807
rect 8518 3773 8552 3807
rect 8618 3773 8652 3807
rect 8718 3773 8752 3807
rect 8818 3773 8852 3807
rect 8918 3773 8952 3807
rect 9018 3773 9052 3807
rect 9118 3773 9152 3807
rect 9218 3773 9252 3807
rect 9318 3773 9352 3807
rect 9418 3773 9446 3807
rect 9446 3773 9452 3807
rect 9518 3773 9524 3807
rect 9524 3773 9552 3807
rect 9618 3773 9652 3807
rect 9718 3773 9752 3807
rect 9818 3773 9852 3807
rect 9918 3773 9952 3807
rect 10018 3773 10046 3807
rect 10046 3773 10052 3807
rect 10118 3773 10124 3807
rect 10124 3773 10152 3807
rect 10218 3773 10252 3807
rect 10318 3773 10352 3807
rect 10418 3773 10452 3807
rect 10518 3773 10552 3807
rect 10618 3773 10652 3807
rect 10718 3773 10752 3807
rect 10818 3773 10852 3807
rect 10918 3773 10952 3807
rect 11018 3773 11052 3807
rect 11118 3773 11146 3807
rect 11146 3773 11152 3807
rect 11218 3773 11224 3807
rect 11224 3773 11252 3807
rect 11318 3773 11352 3807
rect 11418 3773 11452 3807
rect 11518 3773 11546 3807
rect 11546 3773 11552 3807
rect 11618 3773 11624 3807
rect 11624 3773 11652 3807
rect 11718 3773 11752 3807
rect 11818 3773 11852 3807
rect 11918 3773 11952 3807
rect 12018 3773 12052 3807
rect 12118 3773 12146 3807
rect 12146 3773 12152 3807
rect 12218 3773 12224 3807
rect 12224 3773 12252 3807
rect 12318 3773 12352 3807
rect 12418 3773 12452 3807
rect 12518 3773 12552 3807
rect 12618 3773 12652 3807
rect 12718 3773 12752 3807
rect 12818 3773 12852 3807
rect 12916 3788 12924 3822
rect 12924 3788 12950 3822
rect 13120 3758 13146 3792
rect 13146 3758 13154 3792
rect 18 3650 52 3684
rect 218 3666 252 3700
rect 418 3650 452 3684
rect 618 3666 652 3700
rect 818 3650 852 3684
rect 1018 3666 1052 3700
rect 1218 3650 1252 3684
rect 1418 3666 1452 3700
rect 1618 3650 1652 3684
rect 1818 3666 1852 3700
rect 2018 3650 2052 3684
rect 2218 3666 2252 3700
rect 2418 3650 2452 3684
rect 2618 3666 2652 3700
rect 2818 3650 2852 3684
rect 3018 3666 3052 3700
rect 3218 3650 3252 3684
rect 3418 3666 3452 3700
rect 3618 3650 3652 3684
rect 3818 3666 3852 3700
rect 4018 3650 4052 3684
rect 4218 3666 4252 3700
rect 4418 3650 4452 3684
rect 4618 3666 4652 3700
rect 4818 3650 4852 3684
rect 5018 3666 5052 3700
rect 5218 3650 5252 3684
rect 5418 3666 5452 3700
rect 5618 3650 5652 3684
rect 5818 3666 5852 3700
rect 6018 3650 6052 3684
rect 6218 3666 6252 3700
rect 6418 3650 6452 3684
rect 6618 3666 6652 3700
rect 6818 3650 6852 3684
rect 7018 3666 7052 3700
rect 7218 3650 7252 3684
rect 7418 3666 7452 3700
rect 7618 3650 7652 3684
rect 7818 3666 7852 3700
rect 8018 3650 8052 3684
rect 8218 3666 8252 3700
rect 8418 3650 8452 3684
rect 8618 3666 8652 3700
rect 8818 3650 8852 3684
rect 9018 3666 9052 3700
rect 9218 3650 9252 3684
rect 9418 3666 9452 3700
rect 9618 3650 9652 3684
rect 9818 3666 9852 3700
rect 10018 3650 10052 3684
rect 10218 3666 10252 3700
rect 10418 3650 10452 3684
rect 10618 3666 10652 3700
rect 10818 3650 10852 3684
rect 11018 3666 11052 3700
rect 11218 3650 11252 3684
rect 11418 3666 11452 3700
rect 11618 3650 11652 3684
rect 11818 3666 11852 3700
rect 12018 3650 12052 3684
rect 12218 3666 12252 3700
rect 12418 3650 12452 3684
rect 12618 3666 12652 3700
rect 12916 3647 12950 3681
rect 13120 3669 13154 3703
rect 13278 3664 13312 3698
rect 13378 3664 13412 3698
rect 13478 3664 13512 3698
rect 13578 3664 13612 3698
rect 18 3543 52 3577
rect 118 3543 152 3577
rect 218 3543 252 3577
rect 318 3543 352 3577
rect 418 3543 452 3577
rect 518 3543 552 3577
rect 618 3543 652 3577
rect 718 3543 752 3577
rect 818 3543 846 3577
rect 846 3543 852 3577
rect 918 3543 924 3577
rect 924 3543 952 3577
rect 1018 3543 1046 3577
rect 1046 3543 1052 3577
rect 1118 3543 1124 3577
rect 1124 3543 1152 3577
rect 1218 3543 1252 3577
rect 1318 3543 1352 3577
rect 1418 3543 1452 3577
rect 1518 3543 1552 3577
rect 1618 3543 1652 3577
rect 1718 3543 1752 3577
rect 1818 3543 1852 3577
rect 1918 3543 1952 3577
rect 2018 3543 2052 3577
rect 2118 3543 2152 3577
rect 2218 3543 2252 3577
rect 2318 3543 2352 3577
rect 2418 3543 2452 3577
rect 2518 3543 2546 3577
rect 2546 3543 2552 3577
rect 2618 3543 2624 3577
rect 2624 3543 2652 3577
rect 2718 3543 2752 3577
rect 2818 3543 2852 3577
rect 2918 3543 2952 3577
rect 3018 3543 3052 3577
rect 3118 3543 3146 3577
rect 3146 3543 3152 3577
rect 3218 3543 3224 3577
rect 3224 3543 3252 3577
rect 3318 3543 3352 3577
rect 3418 3543 3452 3577
rect 3518 3543 3552 3577
rect 3618 3543 3652 3577
rect 3718 3543 3752 3577
rect 3818 3543 3852 3577
rect 3918 3543 3952 3577
rect 4018 3543 4052 3577
rect 4118 3543 4152 3577
rect 4218 3543 4252 3577
rect 4318 3543 4352 3577
rect 4418 3543 4446 3577
rect 4446 3543 4452 3577
rect 4518 3543 4524 3577
rect 4524 3543 4552 3577
rect 4618 3543 4652 3577
rect 4718 3543 4752 3577
rect 4818 3543 4852 3577
rect 4918 3543 4952 3577
rect 5018 3543 5052 3577
rect 5118 3543 5152 3577
rect 5218 3543 5252 3577
rect 5318 3543 5352 3577
rect 5418 3543 5452 3577
rect 5518 3543 5552 3577
rect 5618 3543 5652 3577
rect 5718 3543 5746 3577
rect 5746 3543 5752 3577
rect 5818 3543 5824 3577
rect 5824 3543 5852 3577
rect 5918 3543 5952 3577
rect 6018 3543 6052 3577
rect 6118 3543 6152 3577
rect 6218 3543 6252 3577
rect 6318 3543 6352 3577
rect 6418 3543 6452 3577
rect 6518 3543 6552 3577
rect 6618 3543 6652 3577
rect 6718 3543 6752 3577
rect 6818 3543 6852 3577
rect 6918 3543 6952 3577
rect 7018 3543 7052 3577
rect 7118 3543 7152 3577
rect 7218 3543 7252 3577
rect 7318 3543 7352 3577
rect 7418 3543 7452 3577
rect 7518 3543 7552 3577
rect 7618 3543 7652 3577
rect 7718 3543 7752 3577
rect 7818 3543 7852 3577
rect 7918 3543 7952 3577
rect 8018 3543 8052 3577
rect 8118 3543 8152 3577
rect 8218 3543 8252 3577
rect 8318 3543 8352 3577
rect 8418 3543 8452 3577
rect 8518 3543 8552 3577
rect 8618 3543 8652 3577
rect 8718 3543 8752 3577
rect 8818 3543 8852 3577
rect 8918 3543 8946 3577
rect 8946 3543 8952 3577
rect 9018 3543 9024 3577
rect 9024 3543 9052 3577
rect 9118 3543 9146 3577
rect 9146 3543 9152 3577
rect 9218 3543 9224 3577
rect 9224 3543 9252 3577
rect 9318 3543 9346 3577
rect 9346 3543 9352 3577
rect 9418 3543 9424 3577
rect 9424 3543 9452 3577
rect 9518 3543 9552 3577
rect 9618 3543 9652 3577
rect 9718 3543 9752 3577
rect 9818 3543 9852 3577
rect 9918 3543 9952 3577
rect 10018 3543 10046 3577
rect 10046 3543 10052 3577
rect 10118 3543 10124 3577
rect 10124 3543 10152 3577
rect 10218 3543 10252 3577
rect 10318 3543 10352 3577
rect 10418 3543 10452 3577
rect 10518 3543 10552 3577
rect 10618 3543 10646 3577
rect 10646 3543 10652 3577
rect 10718 3543 10724 3577
rect 10724 3543 10752 3577
rect 10818 3543 10852 3577
rect 10918 3543 10952 3577
rect 11018 3543 11052 3577
rect 11118 3543 11152 3577
rect 11218 3543 11252 3577
rect 11318 3543 11352 3577
rect 11418 3543 11446 3577
rect 11446 3543 11452 3577
rect 11518 3543 11524 3577
rect 11524 3543 11552 3577
rect 11618 3543 11652 3577
rect 11718 3543 11752 3577
rect 11818 3543 11852 3577
rect 11918 3543 11952 3577
rect 12018 3543 12052 3577
rect 12118 3543 12152 3577
rect 12218 3543 12252 3577
rect 12318 3543 12352 3577
rect 12418 3543 12452 3577
rect 12518 3543 12552 3577
rect 12618 3543 12652 3577
rect 12718 3543 12752 3577
rect 12818 3543 12852 3577
rect 12916 3558 12924 3592
rect 12924 3558 12950 3592
rect 13120 3528 13146 3562
rect 13146 3528 13154 3562
rect 18 3403 24 3437
rect 24 3403 52 3437
rect 118 3403 152 3437
rect 218 3403 252 3437
rect 318 3403 346 3437
rect 346 3403 352 3437
rect 418 3403 424 3437
rect 424 3403 452 3437
rect 518 3403 546 3437
rect 546 3403 552 3437
rect 618 3403 624 3437
rect 624 3403 652 3437
rect 718 3403 746 3437
rect 746 3403 752 3437
rect 818 3403 824 3437
rect 824 3403 852 3437
rect 918 3403 946 3437
rect 946 3403 952 3437
rect 1018 3403 1024 3437
rect 1024 3403 1052 3437
rect 1118 3403 1152 3437
rect 1218 3403 1252 3437
rect 1318 3403 1352 3437
rect 1418 3403 1452 3437
rect 1518 3403 1552 3437
rect 1618 3403 1652 3437
rect 1718 3403 1752 3437
rect 1818 3403 1852 3437
rect 1918 3403 1952 3437
rect 2018 3403 2052 3437
rect 2118 3403 2152 3437
rect 2218 3403 2252 3437
rect 2318 3403 2352 3437
rect 2418 3403 2452 3437
rect 2518 3403 2552 3437
rect 2618 3403 2652 3437
rect 2718 3403 2752 3437
rect 2818 3403 2852 3437
rect 2918 3403 2952 3437
rect 3018 3403 3052 3437
rect 3118 3403 3152 3437
rect 3218 3403 3252 3437
rect 3318 3403 3352 3437
rect 3418 3403 3452 3437
rect 3518 3403 3552 3437
rect 3618 3403 3652 3437
rect 3718 3403 3752 3437
rect 3818 3403 3846 3437
rect 3846 3403 3852 3437
rect 3918 3403 3924 3437
rect 3924 3403 3952 3437
rect 4018 3403 4052 3437
rect 4118 3403 4152 3437
rect 4218 3403 4252 3437
rect 4318 3403 4352 3437
rect 4418 3403 4446 3437
rect 4446 3403 4452 3437
rect 4518 3403 4524 3437
rect 4524 3403 4552 3437
rect 4618 3403 4652 3437
rect 4718 3403 4752 3437
rect 4818 3403 4846 3437
rect 4846 3403 4852 3437
rect 4918 3403 4924 3437
rect 4924 3403 4952 3437
rect 5018 3403 5046 3437
rect 5046 3403 5052 3437
rect 5118 3403 5124 3437
rect 5124 3403 5152 3437
rect 5218 3403 5252 3437
rect 5318 3403 5352 3437
rect 5418 3403 5452 3437
rect 5518 3403 5552 3437
rect 5618 3403 5652 3437
rect 5718 3403 5752 3437
rect 5818 3403 5852 3437
rect 5918 3403 5952 3437
rect 6018 3403 6046 3437
rect 6046 3403 6052 3437
rect 6118 3403 6124 3437
rect 6124 3403 6152 3437
rect 6218 3403 6252 3437
rect 6318 3403 6352 3437
rect 6418 3403 6446 3437
rect 6446 3403 6452 3437
rect 6518 3403 6524 3437
rect 6524 3403 6552 3437
rect 6618 3403 6652 3437
rect 6718 3403 6746 3437
rect 6746 3403 6752 3437
rect 6818 3403 6824 3437
rect 6824 3403 6852 3437
rect 6918 3403 6952 3437
rect 7018 3403 7052 3437
rect 7118 3403 7152 3437
rect 7218 3403 7252 3437
rect 7318 3403 7352 3437
rect 7418 3403 7452 3437
rect 7518 3403 7552 3437
rect 7618 3403 7652 3437
rect 7718 3403 7752 3437
rect 7818 3403 7852 3437
rect 7918 3403 7952 3437
rect 8018 3403 8052 3437
rect 8118 3403 8152 3437
rect 8218 3403 8252 3437
rect 8318 3403 8352 3437
rect 8418 3403 8452 3437
rect 8518 3403 8552 3437
rect 8618 3403 8652 3437
rect 8718 3403 8752 3437
rect 8818 3403 8852 3437
rect 8918 3403 8952 3437
rect 9018 3403 9052 3437
rect 9118 3403 9152 3437
rect 9218 3403 9252 3437
rect 9318 3403 9352 3437
rect 9418 3403 9446 3437
rect 9446 3403 9452 3437
rect 9518 3403 9524 3437
rect 9524 3403 9552 3437
rect 9618 3403 9652 3437
rect 9718 3403 9746 3437
rect 9746 3403 9752 3437
rect 9818 3403 9824 3437
rect 9824 3403 9852 3437
rect 9918 3403 9952 3437
rect 10018 3403 10052 3437
rect 10118 3403 10152 3437
rect 10218 3403 10252 3437
rect 10318 3403 10352 3437
rect 10418 3403 10452 3437
rect 10518 3403 10552 3437
rect 10618 3403 10652 3437
rect 10718 3403 10752 3437
rect 10818 3403 10852 3437
rect 10918 3403 10952 3437
rect 11018 3403 11052 3437
rect 11118 3403 11152 3437
rect 11218 3403 11252 3437
rect 11318 3403 11352 3437
rect 11418 3403 11446 3437
rect 11446 3403 11452 3437
rect 11518 3403 11524 3437
rect 11524 3403 11552 3437
rect 11618 3403 11652 3437
rect 11718 3403 11752 3437
rect 11818 3403 11852 3437
rect 11918 3403 11952 3437
rect 12018 3403 12052 3437
rect 12118 3403 12146 3437
rect 12146 3403 12152 3437
rect 12218 3403 12224 3437
rect 12224 3403 12252 3437
rect 12318 3403 12352 3437
rect 12418 3403 12452 3437
rect 12518 3403 12552 3437
rect 12618 3403 12652 3437
rect 12718 3403 12752 3437
rect 12818 3403 12846 3437
rect 12846 3403 12852 3437
rect 12916 3418 12924 3452
rect 12924 3418 12950 3452
rect 13120 3388 13146 3422
rect 13146 3388 13154 3422
rect 18 3263 52 3297
rect 118 3263 152 3297
rect 218 3263 252 3297
rect 318 3263 352 3297
rect 418 3263 452 3297
rect 518 3263 552 3297
rect 618 3263 652 3297
rect 718 3263 746 3297
rect 746 3263 752 3297
rect 818 3263 824 3297
rect 824 3263 852 3297
rect 918 3263 946 3297
rect 946 3263 952 3297
rect 1018 3263 1024 3297
rect 1024 3263 1052 3297
rect 1118 3263 1152 3297
rect 1218 3263 1252 3297
rect 1318 3263 1352 3297
rect 1418 3263 1452 3297
rect 1518 3263 1552 3297
rect 1618 3263 1652 3297
rect 1718 3263 1752 3297
rect 1818 3263 1852 3297
rect 1918 3263 1952 3297
rect 2018 3263 2052 3297
rect 2118 3263 2152 3297
rect 2218 3263 2252 3297
rect 2318 3263 2352 3297
rect 2418 3263 2452 3297
rect 2518 3263 2552 3297
rect 2618 3263 2652 3297
rect 2718 3263 2746 3297
rect 2746 3263 2752 3297
rect 2818 3263 2824 3297
rect 2824 3263 2852 3297
rect 2918 3263 2952 3297
rect 3018 3263 3052 3297
rect 3118 3263 3152 3297
rect 3218 3263 3246 3297
rect 3246 3263 3252 3297
rect 3318 3263 3324 3297
rect 3324 3263 3352 3297
rect 3418 3263 3446 3297
rect 3446 3263 3452 3297
rect 3518 3263 3524 3297
rect 3524 3263 3552 3297
rect 3618 3263 3652 3297
rect 3718 3263 3752 3297
rect 3818 3263 3852 3297
rect 3918 3263 3952 3297
rect 4018 3263 4052 3297
rect 4118 3263 4152 3297
rect 4218 3263 4252 3297
rect 4318 3263 4352 3297
rect 4418 3263 4452 3297
rect 4518 3263 4552 3297
rect 4618 3263 4652 3297
rect 4718 3263 4752 3297
rect 4818 3263 4852 3297
rect 4918 3263 4952 3297
rect 5018 3263 5052 3297
rect 5118 3263 5152 3297
rect 5218 3263 5252 3297
rect 5318 3263 5352 3297
rect 5418 3263 5452 3297
rect 5518 3263 5552 3297
rect 5618 3263 5652 3297
rect 5718 3263 5752 3297
rect 5818 3263 5852 3297
rect 5918 3263 5952 3297
rect 6018 3263 6052 3297
rect 6118 3263 6152 3297
rect 6218 3263 6252 3297
rect 6318 3263 6352 3297
rect 6418 3263 6452 3297
rect 6518 3263 6552 3297
rect 6618 3263 6652 3297
rect 6718 3263 6752 3297
rect 6818 3263 6852 3297
rect 6918 3263 6952 3297
rect 7018 3263 7052 3297
rect 7118 3263 7152 3297
rect 7218 3263 7252 3297
rect 7318 3263 7346 3297
rect 7346 3263 7352 3297
rect 7418 3263 7424 3297
rect 7424 3263 7452 3297
rect 7518 3263 7552 3297
rect 7618 3263 7652 3297
rect 7718 3263 7752 3297
rect 7818 3263 7852 3297
rect 7918 3263 7952 3297
rect 8018 3263 8052 3297
rect 8118 3263 8152 3297
rect 8218 3263 8252 3297
rect 8318 3263 8352 3297
rect 8418 3263 8452 3297
rect 8518 3263 8552 3297
rect 8618 3263 8652 3297
rect 8718 3263 8752 3297
rect 8818 3263 8852 3297
rect 8918 3263 8952 3297
rect 9018 3263 9052 3297
rect 9118 3263 9152 3297
rect 9218 3263 9252 3297
rect 9318 3263 9352 3297
rect 9418 3263 9452 3297
rect 9518 3263 9546 3297
rect 9546 3263 9552 3297
rect 9618 3263 9624 3297
rect 9624 3263 9652 3297
rect 9718 3263 9752 3297
rect 9818 3263 9852 3297
rect 9918 3263 9952 3297
rect 10018 3263 10052 3297
rect 10118 3263 10152 3297
rect 10218 3263 10252 3297
rect 10318 3263 10346 3297
rect 10346 3263 10352 3297
rect 10418 3263 10424 3297
rect 10424 3263 10452 3297
rect 10518 3263 10546 3297
rect 10546 3263 10552 3297
rect 10618 3263 10624 3297
rect 10624 3263 10652 3297
rect 10718 3263 10752 3297
rect 10818 3263 10852 3297
rect 10918 3263 10952 3297
rect 11018 3263 11052 3297
rect 11118 3263 11152 3297
rect 11218 3263 11252 3297
rect 11318 3263 11352 3297
rect 11418 3263 11452 3297
rect 11518 3263 11552 3297
rect 11618 3263 11652 3297
rect 11718 3263 11752 3297
rect 11818 3263 11852 3297
rect 11918 3263 11952 3297
rect 12018 3263 12052 3297
rect 12118 3263 12152 3297
rect 12218 3263 12252 3297
rect 12318 3263 12352 3297
rect 12418 3263 12446 3297
rect 12446 3263 12452 3297
rect 12518 3263 12524 3297
rect 12524 3263 12552 3297
rect 12618 3263 12652 3297
rect 12718 3263 12752 3297
rect 12818 3263 12852 3297
rect 12916 3278 12924 3312
rect 12924 3278 12950 3312
rect 13120 3248 13146 3282
rect 13146 3248 13154 3282
rect 18 3123 24 3157
rect 24 3123 52 3157
rect 118 3123 146 3157
rect 146 3123 152 3157
rect 218 3123 224 3157
rect 224 3123 252 3157
rect 318 3123 352 3157
rect 418 3123 452 3157
rect 518 3123 552 3157
rect 618 3123 652 3157
rect 718 3123 752 3157
rect 818 3123 852 3157
rect 918 3123 952 3157
rect 1018 3123 1052 3157
rect 1118 3123 1152 3157
rect 1218 3123 1252 3157
rect 1318 3123 1346 3157
rect 1346 3123 1352 3157
rect 1418 3123 1424 3157
rect 1424 3123 1452 3157
rect 1518 3123 1552 3157
rect 1618 3123 1652 3157
rect 1718 3123 1752 3157
rect 1818 3123 1852 3157
rect 1918 3123 1952 3157
rect 2018 3123 2052 3157
rect 2118 3123 2152 3157
rect 2218 3123 2252 3157
rect 2318 3123 2352 3157
rect 2418 3123 2452 3157
rect 2518 3123 2546 3157
rect 2546 3123 2552 3157
rect 2618 3123 2624 3157
rect 2624 3123 2652 3157
rect 2718 3123 2752 3157
rect 2818 3123 2852 3157
rect 2918 3123 2952 3157
rect 3018 3123 3052 3157
rect 3118 3123 3152 3157
rect 3218 3123 3246 3157
rect 3246 3123 3252 3157
rect 3318 3123 3324 3157
rect 3324 3123 3352 3157
rect 3418 3123 3452 3157
rect 3518 3123 3552 3157
rect 3618 3123 3646 3157
rect 3646 3123 3652 3157
rect 3718 3123 3724 3157
rect 3724 3123 3752 3157
rect 3818 3123 3852 3157
rect 3918 3123 3952 3157
rect 4018 3123 4052 3157
rect 4118 3123 4152 3157
rect 4218 3123 4252 3157
rect 4318 3123 4352 3157
rect 4418 3123 4452 3157
rect 4518 3123 4552 3157
rect 4618 3123 4652 3157
rect 4718 3123 4752 3157
rect 4818 3123 4852 3157
rect 4918 3123 4952 3157
rect 5018 3123 5052 3157
rect 5118 3123 5152 3157
rect 5218 3123 5252 3157
rect 5318 3123 5352 3157
rect 5418 3123 5446 3157
rect 5446 3123 5452 3157
rect 5518 3123 5524 3157
rect 5524 3123 5552 3157
rect 5618 3123 5646 3157
rect 5646 3123 5652 3157
rect 5718 3123 5724 3157
rect 5724 3123 5752 3157
rect 5818 3123 5846 3157
rect 5846 3123 5852 3157
rect 5918 3123 5924 3157
rect 5924 3123 5952 3157
rect 6018 3123 6052 3157
rect 6118 3123 6152 3157
rect 6218 3123 6252 3157
rect 6318 3123 6346 3157
rect 6346 3123 6352 3157
rect 6418 3123 6424 3157
rect 6424 3123 6452 3157
rect 6518 3123 6546 3157
rect 6546 3123 6552 3157
rect 6618 3123 6624 3157
rect 6624 3123 6652 3157
rect 6718 3123 6752 3157
rect 6818 3123 6852 3157
rect 6918 3123 6952 3157
rect 7018 3123 7046 3157
rect 7046 3123 7052 3157
rect 7118 3123 7124 3157
rect 7124 3123 7152 3157
rect 7218 3123 7252 3157
rect 7318 3123 7352 3157
rect 7418 3123 7452 3157
rect 7518 3123 7552 3157
rect 7618 3123 7652 3157
rect 7718 3123 7752 3157
rect 7818 3123 7852 3157
rect 7918 3123 7952 3157
rect 8018 3123 8052 3157
rect 8118 3123 8146 3157
rect 8146 3123 8152 3157
rect 8218 3123 8224 3157
rect 8224 3123 8252 3157
rect 8318 3123 8352 3157
rect 8418 3123 8452 3157
rect 8518 3123 8552 3157
rect 8618 3123 8652 3157
rect 8718 3123 8752 3157
rect 8818 3123 8846 3157
rect 8846 3123 8852 3157
rect 8918 3123 8924 3157
rect 8924 3123 8952 3157
rect 9018 3123 9052 3157
rect 9118 3123 9152 3157
rect 9218 3123 9252 3157
rect 9318 3123 9352 3157
rect 9418 3123 9452 3157
rect 9518 3123 9552 3157
rect 9618 3123 9652 3157
rect 9718 3123 9752 3157
rect 9818 3123 9852 3157
rect 9918 3123 9946 3157
rect 9946 3123 9952 3157
rect 10018 3123 10024 3157
rect 10024 3123 10052 3157
rect 10118 3123 10146 3157
rect 10146 3123 10152 3157
rect 10218 3123 10224 3157
rect 10224 3123 10252 3157
rect 10318 3123 10346 3157
rect 10346 3123 10352 3157
rect 10418 3123 10424 3157
rect 10424 3123 10452 3157
rect 10518 3123 10552 3157
rect 10618 3123 10652 3157
rect 10718 3123 10752 3157
rect 10818 3123 10846 3157
rect 10846 3123 10852 3157
rect 10918 3123 10924 3157
rect 10924 3123 10952 3157
rect 11018 3123 11052 3157
rect 11118 3123 11152 3157
rect 11218 3123 11252 3157
rect 11318 3123 11352 3157
rect 11418 3123 11452 3157
rect 11518 3123 11546 3157
rect 11546 3123 11552 3157
rect 11618 3123 11624 3157
rect 11624 3123 11652 3157
rect 11718 3123 11752 3157
rect 11818 3123 11852 3157
rect 11918 3123 11952 3157
rect 12018 3123 12052 3157
rect 12118 3123 12152 3157
rect 12218 3123 12252 3157
rect 12318 3123 12352 3157
rect 12418 3123 12452 3157
rect 12518 3123 12552 3157
rect 12618 3123 12652 3157
rect 12718 3123 12752 3157
rect 12818 3123 12852 3157
rect 12916 3138 12924 3172
rect 12924 3138 12950 3172
rect 13120 3108 13146 3142
rect 13146 3108 13154 3142
rect 18 2983 52 3017
rect 118 2983 152 3017
rect 218 2983 252 3017
rect 318 2983 352 3017
rect 418 2983 452 3017
rect 518 2983 552 3017
rect 618 2983 646 3017
rect 646 2983 652 3017
rect 718 2983 724 3017
rect 724 2983 752 3017
rect 818 2983 852 3017
rect 918 2983 952 3017
rect 1018 2983 1052 3017
rect 1118 2983 1152 3017
rect 1218 2983 1252 3017
rect 1318 2983 1352 3017
rect 1418 2983 1452 3017
rect 1518 2983 1552 3017
rect 1618 2983 1652 3017
rect 1718 2983 1752 3017
rect 1818 2983 1852 3017
rect 1918 2983 1952 3017
rect 2018 2983 2046 3017
rect 2046 2983 2052 3017
rect 2118 2983 2124 3017
rect 2124 2983 2152 3017
rect 2218 2983 2252 3017
rect 2318 2983 2352 3017
rect 2418 2983 2452 3017
rect 2518 2983 2552 3017
rect 2618 2983 2652 3017
rect 2718 2983 2752 3017
rect 2818 2983 2852 3017
rect 2918 2983 2952 3017
rect 3018 2983 3046 3017
rect 3046 2983 3052 3017
rect 3118 2983 3124 3017
rect 3124 2983 3152 3017
rect 3218 2983 3252 3017
rect 3318 2983 3352 3017
rect 3418 2983 3452 3017
rect 3518 2983 3552 3017
rect 3618 2983 3652 3017
rect 3718 2983 3752 3017
rect 3818 2983 3846 3017
rect 3846 2983 3852 3017
rect 3918 2983 3924 3017
rect 3924 2983 3952 3017
rect 4018 2983 4052 3017
rect 4118 2983 4152 3017
rect 4218 2983 4252 3017
rect 4318 2983 4352 3017
rect 4418 2983 4452 3017
rect 4518 2983 4546 3017
rect 4546 2983 4552 3017
rect 4618 2983 4624 3017
rect 4624 2983 4652 3017
rect 4718 2983 4752 3017
rect 4818 2983 4852 3017
rect 4918 2983 4946 3017
rect 4946 2983 4952 3017
rect 5018 2983 5024 3017
rect 5024 2983 5052 3017
rect 5118 2983 5152 3017
rect 5218 2983 5252 3017
rect 5318 2983 5352 3017
rect 5418 2983 5452 3017
rect 5518 2983 5552 3017
rect 5618 2983 5652 3017
rect 5718 2983 5752 3017
rect 5818 2983 5852 3017
rect 5918 2983 5946 3017
rect 5946 2983 5952 3017
rect 6018 2983 6024 3017
rect 6024 2983 6052 3017
rect 6118 2983 6152 3017
rect 6218 2983 6252 3017
rect 6318 2983 6352 3017
rect 6418 2983 6452 3017
rect 6518 2983 6552 3017
rect 6618 2983 6652 3017
rect 6718 2983 6752 3017
rect 6818 2983 6852 3017
rect 6918 2983 6952 3017
rect 7018 2983 7052 3017
rect 7118 2983 7152 3017
rect 7218 2983 7252 3017
rect 7318 2983 7352 3017
rect 7418 2983 7452 3017
rect 7518 2983 7552 3017
rect 7618 2983 7652 3017
rect 7718 2983 7752 3017
rect 7818 2983 7852 3017
rect 7918 2983 7952 3017
rect 8018 2983 8046 3017
rect 8046 2983 8052 3017
rect 8118 2983 8124 3017
rect 8124 2983 8152 3017
rect 8218 2983 8252 3017
rect 8318 2983 8352 3017
rect 8418 2983 8452 3017
rect 8518 2983 8552 3017
rect 8618 2983 8652 3017
rect 8718 2983 8752 3017
rect 8818 2983 8846 3017
rect 8846 2983 8852 3017
rect 8918 2983 8924 3017
rect 8924 2983 8952 3017
rect 9018 2983 9052 3017
rect 9118 2983 9146 3017
rect 9146 2983 9152 3017
rect 9218 2983 9224 3017
rect 9224 2983 9252 3017
rect 9318 2983 9352 3017
rect 9418 2983 9446 3017
rect 9446 2983 9452 3017
rect 9518 2983 9524 3017
rect 9524 2983 9552 3017
rect 9618 2983 9652 3017
rect 9718 2983 9752 3017
rect 9818 2983 9852 3017
rect 9918 2983 9952 3017
rect 10018 2983 10052 3017
rect 10118 2983 10152 3017
rect 10218 2983 10252 3017
rect 10318 2983 10352 3017
rect 10418 2983 10452 3017
rect 10518 2983 10552 3017
rect 10618 2983 10652 3017
rect 10718 2983 10752 3017
rect 10818 2983 10852 3017
rect 10918 2983 10952 3017
rect 11018 2983 11052 3017
rect 11118 2983 11152 3017
rect 11218 2983 11252 3017
rect 11318 2983 11352 3017
rect 11418 2983 11452 3017
rect 11518 2983 11546 3017
rect 11546 2983 11552 3017
rect 11618 2983 11624 3017
rect 11624 2983 11652 3017
rect 11718 2983 11752 3017
rect 11818 2983 11852 3017
rect 11918 2983 11952 3017
rect 12018 2983 12052 3017
rect 12118 2983 12152 3017
rect 12218 2983 12252 3017
rect 12318 2983 12352 3017
rect 12418 2983 12452 3017
rect 12518 2983 12552 3017
rect 12618 2983 12652 3017
rect 12718 2983 12752 3017
rect 12818 2983 12846 3017
rect 12846 2983 12852 3017
rect 12916 2998 12924 3032
rect 12924 2998 12950 3032
rect 13120 2968 13146 3002
rect 13146 2968 13154 3002
rect 18 2843 24 2877
rect 24 2843 52 2877
rect 118 2843 152 2877
rect 218 2843 252 2877
rect 318 2843 352 2877
rect 418 2843 452 2877
rect 518 2843 552 2877
rect 618 2843 652 2877
rect 718 2843 752 2877
rect 818 2843 846 2877
rect 846 2843 852 2877
rect 918 2843 924 2877
rect 924 2843 952 2877
rect 1018 2843 1052 2877
rect 1118 2843 1152 2877
rect 1218 2843 1252 2877
rect 1318 2843 1352 2877
rect 1418 2843 1452 2877
rect 1518 2843 1552 2877
rect 1618 2843 1652 2877
rect 1718 2843 1752 2877
rect 1818 2843 1852 2877
rect 1918 2843 1952 2877
rect 2018 2843 2052 2877
rect 2118 2843 2152 2877
rect 2218 2843 2252 2877
rect 2318 2843 2352 2877
rect 2418 2843 2452 2877
rect 2518 2843 2552 2877
rect 2618 2843 2646 2877
rect 2646 2843 2652 2877
rect 2718 2843 2724 2877
rect 2724 2843 2752 2877
rect 2818 2843 2852 2877
rect 2918 2843 2946 2877
rect 2946 2843 2952 2877
rect 3018 2843 3024 2877
rect 3024 2843 3052 2877
rect 3118 2843 3152 2877
rect 3218 2843 3252 2877
rect 3318 2843 3346 2877
rect 3346 2843 3352 2877
rect 3418 2843 3424 2877
rect 3424 2843 3452 2877
rect 3518 2843 3552 2877
rect 3618 2843 3652 2877
rect 3718 2843 3752 2877
rect 3818 2843 3852 2877
rect 3918 2843 3946 2877
rect 3946 2843 3952 2877
rect 4018 2843 4024 2877
rect 4024 2843 4052 2877
rect 4118 2843 4152 2877
rect 4218 2843 4252 2877
rect 4318 2843 4352 2877
rect 4418 2843 4452 2877
rect 4518 2843 4552 2877
rect 4618 2843 4652 2877
rect 4718 2843 4752 2877
rect 4818 2843 4852 2877
rect 4918 2843 4952 2877
rect 5018 2843 5052 2877
rect 5118 2843 5152 2877
rect 5218 2843 5252 2877
rect 5318 2843 5346 2877
rect 5346 2843 5352 2877
rect 5418 2843 5424 2877
rect 5424 2843 5452 2877
rect 5518 2843 5552 2877
rect 5618 2843 5652 2877
rect 5718 2843 5752 2877
rect 5818 2843 5852 2877
rect 5918 2843 5952 2877
rect 6018 2843 6046 2877
rect 6046 2843 6052 2877
rect 6118 2843 6124 2877
rect 6124 2843 6152 2877
rect 6218 2843 6252 2877
rect 6318 2843 6352 2877
rect 6418 2843 6452 2877
rect 6518 2843 6552 2877
rect 6618 2843 6652 2877
rect 6718 2843 6752 2877
rect 6818 2843 6852 2877
rect 6918 2843 6946 2877
rect 6946 2843 6952 2877
rect 7018 2843 7024 2877
rect 7024 2843 7052 2877
rect 7118 2843 7152 2877
rect 7218 2843 7252 2877
rect 7318 2843 7346 2877
rect 7346 2843 7352 2877
rect 7418 2843 7424 2877
rect 7424 2843 7452 2877
rect 7518 2843 7552 2877
rect 7618 2843 7652 2877
rect 7718 2843 7752 2877
rect 7818 2843 7852 2877
rect 7918 2843 7946 2877
rect 7946 2843 7952 2877
rect 8018 2843 8024 2877
rect 8024 2843 8052 2877
rect 8118 2843 8152 2877
rect 8218 2843 8252 2877
rect 8318 2843 8352 2877
rect 8418 2843 8452 2877
rect 8518 2843 8552 2877
rect 8618 2843 8652 2877
rect 8718 2843 8746 2877
rect 8746 2843 8752 2877
rect 8818 2843 8824 2877
rect 8824 2843 8852 2877
rect 8918 2843 8952 2877
rect 9018 2843 9052 2877
rect 9118 2843 9152 2877
rect 9218 2843 9252 2877
rect 9318 2843 9352 2877
rect 9418 2843 9452 2877
rect 9518 2843 9552 2877
rect 9618 2843 9652 2877
rect 9718 2843 9752 2877
rect 9818 2843 9852 2877
rect 9918 2843 9952 2877
rect 10018 2843 10052 2877
rect 10118 2843 10152 2877
rect 10218 2843 10252 2877
rect 10318 2843 10352 2877
rect 10418 2843 10452 2877
rect 10518 2843 10546 2877
rect 10546 2843 10552 2877
rect 10618 2843 10624 2877
rect 10624 2843 10652 2877
rect 10718 2843 10752 2877
rect 10818 2843 10852 2877
rect 10918 2843 10952 2877
rect 11018 2843 11052 2877
rect 11118 2843 11152 2877
rect 11218 2843 11252 2877
rect 11318 2843 11346 2877
rect 11346 2843 11352 2877
rect 11418 2843 11424 2877
rect 11424 2843 11452 2877
rect 11518 2843 11552 2877
rect 11618 2843 11652 2877
rect 11718 2843 11752 2877
rect 11818 2843 11846 2877
rect 11846 2843 11852 2877
rect 11918 2843 11924 2877
rect 11924 2843 11952 2877
rect 12018 2843 12052 2877
rect 12118 2843 12152 2877
rect 12218 2843 12252 2877
rect 12318 2843 12352 2877
rect 12418 2843 12452 2877
rect 12518 2843 12552 2877
rect 12618 2843 12652 2877
rect 12718 2843 12752 2877
rect 12818 2843 12846 2877
rect 12846 2843 12852 2877
rect 12916 2858 12924 2892
rect 12924 2858 12950 2892
rect 13120 2828 13146 2862
rect 13146 2828 13154 2862
rect 18 2703 52 2737
rect 118 2703 152 2737
rect 218 2703 252 2737
rect 318 2703 352 2737
rect 418 2703 452 2737
rect 518 2703 552 2737
rect 618 2703 652 2737
rect 718 2703 752 2737
rect 818 2703 852 2737
rect 918 2703 952 2737
rect 1018 2703 1052 2737
rect 1118 2703 1146 2737
rect 1146 2703 1152 2737
rect 1218 2703 1224 2737
rect 1224 2703 1252 2737
rect 1318 2703 1352 2737
rect 1418 2703 1452 2737
rect 1518 2703 1552 2737
rect 1618 2703 1652 2737
rect 1718 2703 1752 2737
rect 1818 2703 1852 2737
rect 1918 2703 1952 2737
rect 2018 2703 2052 2737
rect 2118 2703 2152 2737
rect 2218 2703 2252 2737
rect 2318 2703 2346 2737
rect 2346 2703 2352 2737
rect 2418 2703 2424 2737
rect 2424 2703 2452 2737
rect 2518 2703 2552 2737
rect 2618 2703 2652 2737
rect 2718 2703 2752 2737
rect 2818 2703 2852 2737
rect 2918 2703 2952 2737
rect 3018 2703 3052 2737
rect 3118 2703 3152 2737
rect 3218 2703 3252 2737
rect 3318 2703 3352 2737
rect 3418 2703 3452 2737
rect 3518 2703 3552 2737
rect 3618 2703 3652 2737
rect 3718 2703 3752 2737
rect 3818 2703 3852 2737
rect 3918 2703 3952 2737
rect 4018 2703 4052 2737
rect 4118 2703 4146 2737
rect 4146 2703 4152 2737
rect 4218 2703 4224 2737
rect 4224 2703 4252 2737
rect 4318 2703 4352 2737
rect 4418 2703 4452 2737
rect 4518 2703 4552 2737
rect 4618 2703 4652 2737
rect 4718 2703 4746 2737
rect 4746 2703 4752 2737
rect 4818 2703 4824 2737
rect 4824 2703 4852 2737
rect 4918 2703 4952 2737
rect 5018 2703 5052 2737
rect 5118 2703 5146 2737
rect 5146 2703 5152 2737
rect 5218 2703 5224 2737
rect 5224 2703 5252 2737
rect 5318 2703 5346 2737
rect 5346 2703 5352 2737
rect 5418 2703 5424 2737
rect 5424 2703 5452 2737
rect 5518 2703 5552 2737
rect 5618 2703 5652 2737
rect 5718 2703 5752 2737
rect 5818 2703 5852 2737
rect 5918 2703 5952 2737
rect 6018 2703 6046 2737
rect 6046 2703 6052 2737
rect 6118 2703 6124 2737
rect 6124 2703 6152 2737
rect 6218 2703 6246 2737
rect 6246 2703 6252 2737
rect 6318 2703 6324 2737
rect 6324 2703 6352 2737
rect 6418 2703 6452 2737
rect 6518 2703 6546 2737
rect 6546 2703 6552 2737
rect 6618 2703 6624 2737
rect 6624 2703 6652 2737
rect 6718 2703 6752 2737
rect 6818 2703 6852 2737
rect 6918 2703 6952 2737
rect 7018 2703 7052 2737
rect 7118 2703 7152 2737
rect 7218 2703 7252 2737
rect 7318 2703 7352 2737
rect 7418 2703 7452 2737
rect 7518 2703 7552 2737
rect 7618 2703 7652 2737
rect 7718 2703 7752 2737
rect 7818 2703 7852 2737
rect 7918 2703 7952 2737
rect 8018 2703 8052 2737
rect 8118 2703 8152 2737
rect 8218 2703 8246 2737
rect 8246 2703 8252 2737
rect 8318 2703 8324 2737
rect 8324 2703 8352 2737
rect 8418 2703 8452 2737
rect 8518 2703 8552 2737
rect 8618 2703 8652 2737
rect 8718 2703 8746 2737
rect 8746 2703 8752 2737
rect 8818 2703 8824 2737
rect 8824 2703 8852 2737
rect 8918 2703 8946 2737
rect 8946 2703 8952 2737
rect 9018 2703 9024 2737
rect 9024 2703 9052 2737
rect 9118 2703 9146 2737
rect 9146 2703 9152 2737
rect 9218 2703 9224 2737
rect 9224 2703 9252 2737
rect 9318 2703 9346 2737
rect 9346 2703 9352 2737
rect 9418 2703 9424 2737
rect 9424 2703 9452 2737
rect 9518 2703 9546 2737
rect 9546 2703 9552 2737
rect 9618 2703 9624 2737
rect 9624 2703 9652 2737
rect 9718 2703 9752 2737
rect 9818 2703 9852 2737
rect 9918 2703 9946 2737
rect 9946 2703 9952 2737
rect 10018 2703 10024 2737
rect 10024 2703 10052 2737
rect 10118 2703 10152 2737
rect 10218 2703 10252 2737
rect 10318 2703 10352 2737
rect 10418 2703 10446 2737
rect 10446 2703 10452 2737
rect 10518 2703 10524 2737
rect 10524 2703 10552 2737
rect 10618 2703 10646 2737
rect 10646 2703 10652 2737
rect 10718 2703 10724 2737
rect 10724 2703 10752 2737
rect 10818 2703 10852 2737
rect 10918 2703 10952 2737
rect 11018 2703 11052 2737
rect 11118 2703 11152 2737
rect 11218 2703 11252 2737
rect 11318 2703 11352 2737
rect 11418 2703 11452 2737
rect 11518 2703 11552 2737
rect 11618 2703 11646 2737
rect 11646 2703 11652 2737
rect 11718 2703 11724 2737
rect 11724 2703 11752 2737
rect 11818 2703 11852 2737
rect 11918 2703 11952 2737
rect 12018 2703 12052 2737
rect 12118 2703 12152 2737
rect 12218 2703 12252 2737
rect 12318 2703 12352 2737
rect 12418 2703 12452 2737
rect 12518 2703 12552 2737
rect 12618 2703 12652 2737
rect 12718 2703 12752 2737
rect 12818 2703 12852 2737
rect 12916 2718 12924 2752
rect 12924 2718 12950 2752
rect 13120 2688 13146 2722
rect 13146 2688 13154 2722
rect 18 2563 52 2597
rect 118 2563 152 2597
rect 218 2563 252 2597
rect 318 2563 352 2597
rect 418 2563 452 2597
rect 518 2563 552 2597
rect 618 2563 652 2597
rect 718 2563 752 2597
rect 818 2563 852 2597
rect 918 2563 952 2597
rect 1018 2563 1052 2597
rect 1118 2563 1152 2597
rect 1218 2563 1252 2597
rect 1318 2563 1352 2597
rect 1418 2563 1452 2597
rect 1518 2563 1552 2597
rect 1618 2563 1652 2597
rect 1718 2563 1752 2597
rect 1818 2563 1852 2597
rect 1918 2563 1952 2597
rect 2018 2563 2052 2597
rect 2118 2563 2152 2597
rect 2218 2563 2252 2597
rect 2318 2563 2352 2597
rect 2418 2563 2452 2597
rect 2518 2563 2546 2597
rect 2546 2563 2552 2597
rect 2618 2563 2624 2597
rect 2624 2563 2652 2597
rect 2718 2563 2752 2597
rect 2818 2563 2852 2597
rect 2918 2563 2952 2597
rect 3018 2563 3052 2597
rect 3118 2563 3152 2597
rect 3218 2563 3252 2597
rect 3318 2563 3346 2597
rect 3346 2563 3352 2597
rect 3418 2563 3424 2597
rect 3424 2563 3452 2597
rect 3518 2563 3552 2597
rect 3618 2563 3652 2597
rect 3718 2563 3752 2597
rect 3818 2563 3852 2597
rect 3918 2563 3946 2597
rect 3946 2563 3952 2597
rect 4018 2563 4024 2597
rect 4024 2563 4052 2597
rect 4118 2563 4146 2597
rect 4146 2563 4152 2597
rect 4218 2563 4224 2597
rect 4224 2563 4252 2597
rect 4318 2563 4346 2597
rect 4346 2563 4352 2597
rect 4418 2563 4424 2597
rect 4424 2563 4452 2597
rect 4518 2563 4552 2597
rect 4618 2563 4652 2597
rect 4718 2563 4746 2597
rect 4746 2563 4752 2597
rect 4818 2563 4824 2597
rect 4824 2563 4852 2597
rect 4918 2563 4952 2597
rect 5018 2563 5052 2597
rect 5118 2563 5152 2597
rect 5218 2563 5252 2597
rect 5318 2563 5352 2597
rect 5418 2563 5452 2597
rect 5518 2563 5552 2597
rect 5618 2563 5652 2597
rect 5718 2563 5752 2597
rect 5818 2563 5852 2597
rect 5918 2563 5952 2597
rect 6018 2563 6052 2597
rect 6118 2563 6152 2597
rect 6218 2563 6246 2597
rect 6246 2563 6252 2597
rect 6318 2563 6324 2597
rect 6324 2563 6352 2597
rect 6418 2563 6452 2597
rect 6518 2563 6552 2597
rect 6618 2563 6652 2597
rect 6718 2563 6746 2597
rect 6746 2563 6752 2597
rect 6818 2563 6824 2597
rect 6824 2563 6852 2597
rect 6918 2563 6952 2597
rect 7018 2563 7052 2597
rect 7118 2563 7152 2597
rect 7218 2563 7252 2597
rect 7318 2563 7352 2597
rect 7418 2563 7452 2597
rect 7518 2563 7552 2597
rect 7618 2563 7652 2597
rect 7718 2563 7752 2597
rect 7818 2563 7852 2597
rect 7918 2563 7952 2597
rect 8018 2563 8052 2597
rect 8118 2563 8152 2597
rect 8218 2563 8246 2597
rect 8246 2563 8252 2597
rect 8318 2563 8324 2597
rect 8324 2563 8352 2597
rect 8418 2563 8446 2597
rect 8446 2563 8452 2597
rect 8518 2563 8524 2597
rect 8524 2563 8552 2597
rect 8618 2563 8652 2597
rect 8718 2563 8746 2597
rect 8746 2563 8752 2597
rect 8818 2563 8824 2597
rect 8824 2563 8852 2597
rect 8918 2563 8952 2597
rect 9018 2563 9046 2597
rect 9046 2563 9052 2597
rect 9118 2563 9124 2597
rect 9124 2563 9152 2597
rect 9218 2563 9246 2597
rect 9246 2563 9252 2597
rect 9318 2563 9324 2597
rect 9324 2563 9352 2597
rect 9418 2563 9452 2597
rect 9518 2563 9546 2597
rect 9546 2563 9552 2597
rect 9618 2563 9624 2597
rect 9624 2563 9652 2597
rect 9718 2563 9752 2597
rect 9818 2563 9852 2597
rect 9918 2563 9946 2597
rect 9946 2563 9952 2597
rect 10018 2563 10024 2597
rect 10024 2563 10052 2597
rect 10118 2563 10152 2597
rect 10218 2563 10252 2597
rect 10318 2563 10352 2597
rect 10418 2563 10452 2597
rect 10518 2563 10552 2597
rect 10618 2563 10652 2597
rect 10718 2563 10752 2597
rect 10818 2563 10852 2597
rect 10918 2563 10946 2597
rect 10946 2563 10952 2597
rect 11018 2563 11024 2597
rect 11024 2563 11052 2597
rect 11118 2563 11146 2597
rect 11146 2563 11152 2597
rect 11218 2563 11224 2597
rect 11224 2563 11252 2597
rect 11318 2563 11346 2597
rect 11346 2563 11352 2597
rect 11418 2563 11424 2597
rect 11424 2563 11452 2597
rect 11518 2563 11552 2597
rect 11618 2563 11646 2597
rect 11646 2563 11652 2597
rect 11718 2563 11724 2597
rect 11724 2563 11752 2597
rect 11818 2563 11852 2597
rect 11918 2563 11952 2597
rect 12018 2563 12052 2597
rect 12118 2563 12152 2597
rect 12218 2563 12252 2597
rect 12318 2563 12352 2597
rect 12418 2563 12452 2597
rect 12518 2563 12552 2597
rect 12618 2563 12652 2597
rect 12718 2563 12752 2597
rect 12818 2563 12852 2597
rect 12916 2578 12924 2612
rect 12924 2578 12950 2612
rect 13120 2548 13146 2582
rect 13146 2548 13154 2582
rect 18 2440 52 2474
rect 218 2456 252 2490
rect 418 2440 452 2474
rect 618 2456 652 2490
rect 818 2440 852 2474
rect 1018 2456 1052 2490
rect 1218 2440 1252 2474
rect 1418 2456 1452 2490
rect 1618 2440 1652 2474
rect 1818 2456 1852 2490
rect 2018 2440 2052 2474
rect 2218 2456 2252 2490
rect 2418 2440 2452 2474
rect 2618 2456 2652 2490
rect 2818 2440 2852 2474
rect 3018 2456 3052 2490
rect 3218 2440 3252 2474
rect 3418 2456 3452 2490
rect 3618 2440 3652 2474
rect 3818 2456 3852 2490
rect 4018 2440 4052 2474
rect 4218 2456 4252 2490
rect 4418 2440 4452 2474
rect 4618 2456 4652 2490
rect 4818 2440 4852 2474
rect 5018 2456 5052 2490
rect 5218 2440 5252 2474
rect 5418 2456 5452 2490
rect 5618 2440 5652 2474
rect 5818 2456 5852 2490
rect 6018 2440 6052 2474
rect 6218 2456 6252 2490
rect 6418 2440 6452 2474
rect 6618 2456 6652 2490
rect 6818 2440 6852 2474
rect 7018 2456 7052 2490
rect 7218 2440 7252 2474
rect 7418 2456 7452 2490
rect 7618 2440 7652 2474
rect 7818 2456 7852 2490
rect 8018 2440 8052 2474
rect 8218 2456 8252 2490
rect 8418 2440 8452 2474
rect 8618 2456 8652 2490
rect 8818 2440 8852 2474
rect 9018 2456 9052 2490
rect 9218 2440 9252 2474
rect 9418 2456 9452 2490
rect 9618 2440 9652 2474
rect 9818 2456 9852 2490
rect 10018 2440 10052 2474
rect 10218 2456 10252 2490
rect 10418 2440 10452 2474
rect 10618 2456 10652 2490
rect 10818 2440 10852 2474
rect 11018 2456 11052 2490
rect 11218 2440 11252 2474
rect 11418 2456 11452 2490
rect 11618 2440 11652 2474
rect 11818 2456 11852 2490
rect 12018 2440 12052 2474
rect 12218 2456 12252 2490
rect 12418 2440 12452 2474
rect 12618 2456 12652 2490
rect 12916 2437 12950 2471
rect 13120 2459 13154 2493
rect 13278 2454 13312 2488
rect 13378 2454 13412 2488
rect 13478 2454 13512 2488
rect 13578 2454 13612 2488
rect 18 2333 24 2367
rect 24 2333 52 2367
rect 118 2333 146 2367
rect 146 2333 152 2367
rect 218 2333 224 2367
rect 224 2333 252 2367
rect 318 2333 352 2367
rect 418 2333 446 2367
rect 446 2333 452 2367
rect 518 2333 524 2367
rect 524 2333 552 2367
rect 618 2333 646 2367
rect 646 2333 652 2367
rect 718 2333 724 2367
rect 724 2333 752 2367
rect 818 2333 852 2367
rect 918 2333 952 2367
rect 1018 2333 1052 2367
rect 1118 2333 1152 2367
rect 1218 2333 1252 2367
rect 1318 2333 1352 2367
rect 1418 2333 1452 2367
rect 1518 2333 1552 2367
rect 1618 2333 1652 2367
rect 1718 2333 1752 2367
rect 1818 2333 1852 2367
rect 1918 2333 1952 2367
rect 2018 2333 2052 2367
rect 2118 2333 2152 2367
rect 2218 2333 2252 2367
rect 2318 2333 2346 2367
rect 2346 2333 2352 2367
rect 2418 2333 2424 2367
rect 2424 2333 2452 2367
rect 2518 2333 2552 2367
rect 2618 2333 2646 2367
rect 2646 2333 2652 2367
rect 2718 2333 2724 2367
rect 2724 2333 2752 2367
rect 2818 2333 2852 2367
rect 2918 2333 2952 2367
rect 3018 2333 3052 2367
rect 3118 2333 3152 2367
rect 3218 2333 3252 2367
rect 3318 2333 3352 2367
rect 3418 2333 3452 2367
rect 3518 2333 3552 2367
rect 3618 2333 3652 2367
rect 3718 2333 3752 2367
rect 3818 2333 3852 2367
rect 3918 2333 3952 2367
rect 4018 2333 4052 2367
rect 4118 2333 4152 2367
rect 4218 2333 4252 2367
rect 4318 2333 4352 2367
rect 4418 2333 4452 2367
rect 4518 2333 4552 2367
rect 4618 2333 4652 2367
rect 4718 2333 4752 2367
rect 4818 2333 4852 2367
rect 4918 2333 4952 2367
rect 5018 2333 5052 2367
rect 5118 2333 5152 2367
rect 5218 2333 5252 2367
rect 5318 2333 5352 2367
rect 5418 2333 5452 2367
rect 5518 2333 5552 2367
rect 5618 2333 5652 2367
rect 5718 2333 5752 2367
rect 5818 2333 5852 2367
rect 5918 2333 5952 2367
rect 6018 2333 6052 2367
rect 6118 2333 6152 2367
rect 6218 2333 6252 2367
rect 6318 2333 6352 2367
rect 6418 2333 6452 2367
rect 6518 2333 6552 2367
rect 6618 2333 6652 2367
rect 6718 2333 6752 2367
rect 6818 2333 6852 2367
rect 6918 2333 6946 2367
rect 6946 2333 6952 2367
rect 7018 2333 7024 2367
rect 7024 2333 7052 2367
rect 7118 2333 7152 2367
rect 7218 2333 7246 2367
rect 7246 2333 7252 2367
rect 7318 2333 7324 2367
rect 7324 2333 7352 2367
rect 7418 2333 7452 2367
rect 7518 2333 7552 2367
rect 7618 2333 7652 2367
rect 7718 2333 7752 2367
rect 7818 2333 7852 2367
rect 7918 2333 7952 2367
rect 8018 2333 8052 2367
rect 8118 2333 8152 2367
rect 8218 2333 8252 2367
rect 8318 2333 8352 2367
rect 8418 2333 8452 2367
rect 8518 2333 8546 2367
rect 8546 2333 8552 2367
rect 8618 2333 8624 2367
rect 8624 2333 8652 2367
rect 8718 2333 8752 2367
rect 8818 2333 8852 2367
rect 8918 2333 8952 2367
rect 9018 2333 9052 2367
rect 9118 2333 9152 2367
rect 9218 2333 9252 2367
rect 9318 2333 9352 2367
rect 9418 2333 9452 2367
rect 9518 2333 9552 2367
rect 9618 2333 9646 2367
rect 9646 2333 9652 2367
rect 9718 2333 9724 2367
rect 9724 2333 9752 2367
rect 9818 2333 9852 2367
rect 9918 2333 9952 2367
rect 10018 2333 10052 2367
rect 10118 2333 10152 2367
rect 10218 2333 10252 2367
rect 10318 2333 10352 2367
rect 10418 2333 10452 2367
rect 10518 2333 10552 2367
rect 10618 2333 10652 2367
rect 10718 2333 10752 2367
rect 10818 2333 10852 2367
rect 10918 2333 10952 2367
rect 11018 2333 11052 2367
rect 11118 2333 11152 2367
rect 11218 2333 11252 2367
rect 11318 2333 11352 2367
rect 11418 2333 11452 2367
rect 11518 2333 11552 2367
rect 11618 2333 11652 2367
rect 11718 2333 11746 2367
rect 11746 2333 11752 2367
rect 11818 2333 11824 2367
rect 11824 2333 11852 2367
rect 11918 2333 11946 2367
rect 11946 2333 11952 2367
rect 12018 2333 12024 2367
rect 12024 2333 12052 2367
rect 12118 2333 12152 2367
rect 12218 2333 12252 2367
rect 12318 2333 12352 2367
rect 12418 2333 12452 2367
rect 12518 2333 12546 2367
rect 12546 2333 12552 2367
rect 12618 2333 12624 2367
rect 12624 2333 12652 2367
rect 12718 2333 12752 2367
rect 12818 2333 12852 2367
rect 12916 2348 12924 2382
rect 12924 2348 12950 2382
rect 13120 2318 13146 2352
rect 13146 2318 13154 2352
rect 18 2193 24 2227
rect 24 2193 52 2227
rect 118 2193 152 2227
rect 218 2193 252 2227
rect 318 2193 352 2227
rect 418 2193 452 2227
rect 518 2193 552 2227
rect 618 2193 652 2227
rect 718 2193 752 2227
rect 818 2193 846 2227
rect 846 2193 852 2227
rect 918 2193 924 2227
rect 924 2193 952 2227
rect 1018 2193 1046 2227
rect 1046 2193 1052 2227
rect 1118 2193 1124 2227
rect 1124 2193 1152 2227
rect 1218 2193 1252 2227
rect 1318 2193 1352 2227
rect 1418 2193 1452 2227
rect 1518 2193 1552 2227
rect 1618 2193 1652 2227
rect 1718 2193 1752 2227
rect 1818 2193 1852 2227
rect 1918 2193 1952 2227
rect 2018 2193 2052 2227
rect 2118 2193 2152 2227
rect 2218 2193 2252 2227
rect 2318 2193 2352 2227
rect 2418 2193 2452 2227
rect 2518 2193 2552 2227
rect 2618 2193 2646 2227
rect 2646 2193 2652 2227
rect 2718 2193 2724 2227
rect 2724 2193 2752 2227
rect 2818 2193 2846 2227
rect 2846 2193 2852 2227
rect 2918 2193 2924 2227
rect 2924 2193 2952 2227
rect 3018 2193 3046 2227
rect 3046 2193 3052 2227
rect 3118 2193 3124 2227
rect 3124 2193 3152 2227
rect 3218 2193 3252 2227
rect 3318 2193 3346 2227
rect 3346 2193 3352 2227
rect 3418 2193 3424 2227
rect 3424 2193 3452 2227
rect 3518 2193 3552 2227
rect 3618 2193 3646 2227
rect 3646 2193 3652 2227
rect 3718 2193 3724 2227
rect 3724 2193 3752 2227
rect 3818 2193 3846 2227
rect 3846 2193 3852 2227
rect 3918 2193 3924 2227
rect 3924 2193 3952 2227
rect 4018 2193 4052 2227
rect 4118 2193 4152 2227
rect 4218 2193 4252 2227
rect 4318 2193 4346 2227
rect 4346 2193 4352 2227
rect 4418 2193 4424 2227
rect 4424 2193 4452 2227
rect 4518 2193 4552 2227
rect 4618 2193 4652 2227
rect 4718 2193 4752 2227
rect 4818 2193 4852 2227
rect 4918 2193 4952 2227
rect 5018 2193 5052 2227
rect 5118 2193 5152 2227
rect 5218 2193 5252 2227
rect 5318 2193 5352 2227
rect 5418 2193 5452 2227
rect 5518 2193 5552 2227
rect 5618 2193 5652 2227
rect 5718 2193 5752 2227
rect 5818 2193 5852 2227
rect 5918 2193 5952 2227
rect 6018 2193 6052 2227
rect 6118 2193 6146 2227
rect 6146 2193 6152 2227
rect 6218 2193 6224 2227
rect 6224 2193 6252 2227
rect 6318 2193 6352 2227
rect 6418 2193 6446 2227
rect 6446 2193 6452 2227
rect 6518 2193 6524 2227
rect 6524 2193 6552 2227
rect 6618 2193 6652 2227
rect 6718 2193 6746 2227
rect 6746 2193 6752 2227
rect 6818 2193 6824 2227
rect 6824 2193 6852 2227
rect 6918 2193 6946 2227
rect 6946 2193 6952 2227
rect 7018 2193 7024 2227
rect 7024 2193 7052 2227
rect 7118 2193 7152 2227
rect 7218 2193 7252 2227
rect 7318 2193 7352 2227
rect 7418 2193 7452 2227
rect 7518 2193 7546 2227
rect 7546 2193 7552 2227
rect 7618 2193 7624 2227
rect 7624 2193 7652 2227
rect 7718 2193 7746 2227
rect 7746 2193 7752 2227
rect 7818 2193 7824 2227
rect 7824 2193 7852 2227
rect 7918 2193 7952 2227
rect 8018 2193 8052 2227
rect 8118 2193 8152 2227
rect 8218 2193 8252 2227
rect 8318 2193 8352 2227
rect 8418 2193 8452 2227
rect 8518 2193 8552 2227
rect 8618 2193 8652 2227
rect 8718 2193 8752 2227
rect 8818 2193 8846 2227
rect 8846 2193 8852 2227
rect 8918 2193 8924 2227
rect 8924 2193 8952 2227
rect 9018 2193 9046 2227
rect 9046 2193 9052 2227
rect 9118 2193 9124 2227
rect 9124 2193 9152 2227
rect 9218 2193 9246 2227
rect 9246 2193 9252 2227
rect 9318 2193 9324 2227
rect 9324 2193 9352 2227
rect 9418 2193 9452 2227
rect 9518 2193 9546 2227
rect 9546 2193 9552 2227
rect 9618 2193 9624 2227
rect 9624 2193 9652 2227
rect 9718 2193 9752 2227
rect 9818 2193 9852 2227
rect 9918 2193 9952 2227
rect 10018 2193 10052 2227
rect 10118 2193 10152 2227
rect 10218 2193 10252 2227
rect 10318 2193 10352 2227
rect 10418 2193 10452 2227
rect 10518 2193 10546 2227
rect 10546 2193 10552 2227
rect 10618 2193 10624 2227
rect 10624 2193 10652 2227
rect 10718 2193 10752 2227
rect 10818 2193 10852 2227
rect 10918 2193 10952 2227
rect 11018 2193 11052 2227
rect 11118 2193 11152 2227
rect 11218 2193 11252 2227
rect 11318 2193 11352 2227
rect 11418 2193 11452 2227
rect 11518 2193 11552 2227
rect 11618 2193 11652 2227
rect 11718 2193 11752 2227
rect 11818 2193 11852 2227
rect 11918 2193 11952 2227
rect 12018 2193 12046 2227
rect 12046 2193 12052 2227
rect 12118 2193 12124 2227
rect 12124 2193 12152 2227
rect 12218 2193 12252 2227
rect 12318 2193 12346 2227
rect 12346 2193 12352 2227
rect 12418 2193 12424 2227
rect 12424 2193 12452 2227
rect 12518 2193 12552 2227
rect 12618 2193 12646 2227
rect 12646 2193 12652 2227
rect 12718 2193 12724 2227
rect 12724 2193 12752 2227
rect 12818 2193 12846 2227
rect 12846 2193 12852 2227
rect 12916 2208 12924 2242
rect 12924 2208 12950 2242
rect 13120 2178 13146 2212
rect 13146 2178 13154 2212
rect 18 2053 52 2087
rect 118 2053 152 2087
rect 218 2053 252 2087
rect 318 2053 352 2087
rect 418 2053 452 2087
rect 518 2053 552 2087
rect 618 2053 652 2087
rect 718 2053 746 2087
rect 746 2053 752 2087
rect 818 2053 824 2087
rect 824 2053 852 2087
rect 918 2053 952 2087
rect 1018 2053 1052 2087
rect 1118 2053 1152 2087
rect 1218 2053 1252 2087
rect 1318 2053 1352 2087
rect 1418 2053 1446 2087
rect 1446 2053 1452 2087
rect 1518 2053 1524 2087
rect 1524 2053 1552 2087
rect 1618 2053 1652 2087
rect 1718 2053 1752 2087
rect 1818 2053 1852 2087
rect 1918 2053 1952 2087
rect 2018 2053 2052 2087
rect 2118 2053 2152 2087
rect 2218 2053 2252 2087
rect 2318 2053 2352 2087
rect 2418 2053 2452 2087
rect 2518 2053 2552 2087
rect 2618 2053 2652 2087
rect 2718 2053 2746 2087
rect 2746 2053 2752 2087
rect 2818 2053 2824 2087
rect 2824 2053 2852 2087
rect 2918 2053 2946 2087
rect 2946 2053 2952 2087
rect 3018 2053 3024 2087
rect 3024 2053 3052 2087
rect 3118 2053 3152 2087
rect 3218 2053 3252 2087
rect 3318 2053 3352 2087
rect 3418 2053 3452 2087
rect 3518 2053 3546 2087
rect 3546 2053 3552 2087
rect 3618 2053 3624 2087
rect 3624 2053 3652 2087
rect 3718 2053 3752 2087
rect 3818 2053 3852 2087
rect 3918 2053 3952 2087
rect 4018 2053 4052 2087
rect 4118 2053 4152 2087
rect 4218 2053 4252 2087
rect 4318 2053 4352 2087
rect 4418 2053 4452 2087
rect 4518 2053 4552 2087
rect 4618 2053 4646 2087
rect 4646 2053 4652 2087
rect 4718 2053 4724 2087
rect 4724 2053 4752 2087
rect 4818 2053 4852 2087
rect 4918 2053 4946 2087
rect 4946 2053 4952 2087
rect 5018 2053 5024 2087
rect 5024 2053 5052 2087
rect 5118 2053 5152 2087
rect 5218 2053 5252 2087
rect 5318 2053 5352 2087
rect 5418 2053 5452 2087
rect 5518 2053 5552 2087
rect 5618 2053 5652 2087
rect 5718 2053 5746 2087
rect 5746 2053 5752 2087
rect 5818 2053 5824 2087
rect 5824 2053 5852 2087
rect 5918 2053 5952 2087
rect 6018 2053 6052 2087
rect 6118 2053 6152 2087
rect 6218 2053 6252 2087
rect 6318 2053 6352 2087
rect 6418 2053 6452 2087
rect 6518 2053 6552 2087
rect 6618 2053 6646 2087
rect 6646 2053 6652 2087
rect 6718 2053 6724 2087
rect 6724 2053 6752 2087
rect 6818 2053 6846 2087
rect 6846 2053 6852 2087
rect 6918 2053 6924 2087
rect 6924 2053 6952 2087
rect 7018 2053 7052 2087
rect 7118 2053 7152 2087
rect 7218 2053 7252 2087
rect 7318 2053 7352 2087
rect 7418 2053 7452 2087
rect 7518 2053 7552 2087
rect 7618 2053 7652 2087
rect 7718 2053 7752 2087
rect 7818 2053 7852 2087
rect 7918 2053 7952 2087
rect 8018 2053 8052 2087
rect 8118 2053 8146 2087
rect 8146 2053 8152 2087
rect 8218 2053 8224 2087
rect 8224 2053 8252 2087
rect 8318 2053 8346 2087
rect 8346 2053 8352 2087
rect 8418 2053 8424 2087
rect 8424 2053 8452 2087
rect 8518 2053 8552 2087
rect 8618 2053 8652 2087
rect 8718 2053 8746 2087
rect 8746 2053 8752 2087
rect 8818 2053 8824 2087
rect 8824 2053 8852 2087
rect 8918 2053 8946 2087
rect 8946 2053 8952 2087
rect 9018 2053 9024 2087
rect 9024 2053 9052 2087
rect 9118 2053 9152 2087
rect 9218 2053 9246 2087
rect 9246 2053 9252 2087
rect 9318 2053 9324 2087
rect 9324 2053 9352 2087
rect 9418 2053 9452 2087
rect 9518 2053 9552 2087
rect 9618 2053 9652 2087
rect 9718 2053 9752 2087
rect 9818 2053 9852 2087
rect 9918 2053 9952 2087
rect 10018 2053 10052 2087
rect 10118 2053 10152 2087
rect 10218 2053 10252 2087
rect 10318 2053 10352 2087
rect 10418 2053 10452 2087
rect 10518 2053 10552 2087
rect 10618 2053 10652 2087
rect 10718 2053 10752 2087
rect 10818 2053 10852 2087
rect 10918 2053 10952 2087
rect 11018 2053 11052 2087
rect 11118 2053 11152 2087
rect 11218 2053 11246 2087
rect 11246 2053 11252 2087
rect 11318 2053 11324 2087
rect 11324 2053 11352 2087
rect 11418 2053 11446 2087
rect 11446 2053 11452 2087
rect 11518 2053 11524 2087
rect 11524 2053 11552 2087
rect 11618 2053 11652 2087
rect 11718 2053 11752 2087
rect 11818 2053 11852 2087
rect 11918 2053 11952 2087
rect 12018 2053 12052 2087
rect 12118 2053 12152 2087
rect 12218 2053 12252 2087
rect 12318 2053 12352 2087
rect 12418 2053 12452 2087
rect 12518 2053 12552 2087
rect 12618 2053 12646 2087
rect 12646 2053 12652 2087
rect 12718 2053 12724 2087
rect 12724 2053 12752 2087
rect 12818 2053 12846 2087
rect 12846 2053 12852 2087
rect 12916 2068 12924 2102
rect 12924 2068 12950 2102
rect 13120 2038 13146 2072
rect 13146 2038 13154 2072
rect 18 1913 52 1947
rect 118 1913 152 1947
rect 218 1913 252 1947
rect 318 1913 352 1947
rect 418 1913 452 1947
rect 518 1913 552 1947
rect 618 1913 652 1947
rect 718 1913 752 1947
rect 818 1913 852 1947
rect 918 1913 946 1947
rect 946 1913 952 1947
rect 1018 1913 1024 1947
rect 1024 1913 1052 1947
rect 1118 1913 1152 1947
rect 1218 1913 1252 1947
rect 1318 1913 1352 1947
rect 1418 1913 1452 1947
rect 1518 1913 1546 1947
rect 1546 1913 1552 1947
rect 1618 1913 1624 1947
rect 1624 1913 1652 1947
rect 1718 1913 1752 1947
rect 1818 1913 1852 1947
rect 1918 1913 1952 1947
rect 2018 1913 2052 1947
rect 2118 1913 2152 1947
rect 2218 1913 2252 1947
rect 2318 1913 2352 1947
rect 2418 1913 2452 1947
rect 2518 1913 2552 1947
rect 2618 1913 2652 1947
rect 2718 1913 2752 1947
rect 2818 1913 2852 1947
rect 2918 1913 2952 1947
rect 3018 1913 3052 1947
rect 3118 1913 3152 1947
rect 3218 1913 3252 1947
rect 3318 1913 3352 1947
rect 3418 1913 3452 1947
rect 3518 1913 3552 1947
rect 3618 1913 3646 1947
rect 3646 1913 3652 1947
rect 3718 1913 3724 1947
rect 3724 1913 3752 1947
rect 3818 1913 3852 1947
rect 3918 1913 3952 1947
rect 4018 1913 4052 1947
rect 4118 1913 4152 1947
rect 4218 1913 4246 1947
rect 4246 1913 4252 1947
rect 4318 1913 4324 1947
rect 4324 1913 4352 1947
rect 4418 1913 4446 1947
rect 4446 1913 4452 1947
rect 4518 1913 4524 1947
rect 4524 1913 4552 1947
rect 4618 1913 4646 1947
rect 4646 1913 4652 1947
rect 4718 1913 4724 1947
rect 4724 1913 4752 1947
rect 4818 1913 4852 1947
rect 4918 1913 4952 1947
rect 5018 1913 5052 1947
rect 5118 1913 5146 1947
rect 5146 1913 5152 1947
rect 5218 1913 5224 1947
rect 5224 1913 5252 1947
rect 5318 1913 5352 1947
rect 5418 1913 5452 1947
rect 5518 1913 5552 1947
rect 5618 1913 5652 1947
rect 5718 1913 5746 1947
rect 5746 1913 5752 1947
rect 5818 1913 5824 1947
rect 5824 1913 5852 1947
rect 5918 1913 5952 1947
rect 6018 1913 6052 1947
rect 6118 1913 6152 1947
rect 6218 1913 6252 1947
rect 6318 1913 6352 1947
rect 6418 1913 6452 1947
rect 6518 1913 6552 1947
rect 6618 1913 6652 1947
rect 6718 1913 6746 1947
rect 6746 1913 6752 1947
rect 6818 1913 6824 1947
rect 6824 1913 6852 1947
rect 6918 1913 6946 1947
rect 6946 1913 6952 1947
rect 7018 1913 7024 1947
rect 7024 1913 7052 1947
rect 7118 1913 7152 1947
rect 7218 1913 7252 1947
rect 7318 1913 7352 1947
rect 7418 1913 7452 1947
rect 7518 1913 7552 1947
rect 7618 1913 7652 1947
rect 7718 1913 7752 1947
rect 7818 1913 7852 1947
rect 7918 1913 7952 1947
rect 8018 1913 8052 1947
rect 8118 1913 8152 1947
rect 8218 1913 8252 1947
rect 8318 1913 8352 1947
rect 8418 1913 8452 1947
rect 8518 1913 8552 1947
rect 8618 1913 8652 1947
rect 8718 1913 8752 1947
rect 8818 1913 8852 1947
rect 8918 1913 8952 1947
rect 9018 1913 9052 1947
rect 9118 1913 9152 1947
rect 9218 1913 9252 1947
rect 9318 1913 9352 1947
rect 9418 1913 9452 1947
rect 9518 1913 9552 1947
rect 9618 1913 9652 1947
rect 9718 1913 9752 1947
rect 9818 1913 9852 1947
rect 9918 1913 9952 1947
rect 10018 1913 10052 1947
rect 10118 1913 10152 1947
rect 10218 1913 10252 1947
rect 10318 1913 10352 1947
rect 10418 1913 10452 1947
rect 10518 1913 10552 1947
rect 10618 1913 10652 1947
rect 10718 1913 10752 1947
rect 10818 1913 10852 1947
rect 10918 1913 10952 1947
rect 11018 1913 11046 1947
rect 11046 1913 11052 1947
rect 11118 1913 11124 1947
rect 11124 1913 11152 1947
rect 11218 1913 11246 1947
rect 11246 1913 11252 1947
rect 11318 1913 11324 1947
rect 11324 1913 11352 1947
rect 11418 1913 11452 1947
rect 11518 1913 11552 1947
rect 11618 1913 11652 1947
rect 11718 1913 11752 1947
rect 11818 1913 11852 1947
rect 11918 1913 11952 1947
rect 12018 1913 12052 1947
rect 12118 1913 12152 1947
rect 12218 1913 12252 1947
rect 12318 1913 12352 1947
rect 12418 1913 12452 1947
rect 12518 1913 12552 1947
rect 12618 1913 12646 1947
rect 12646 1913 12652 1947
rect 12718 1913 12724 1947
rect 12724 1913 12752 1947
rect 12818 1913 12846 1947
rect 12846 1913 12852 1947
rect 12916 1928 12924 1962
rect 12924 1928 12950 1962
rect 13120 1898 13146 1932
rect 13146 1898 13154 1932
rect 18 1773 52 1807
rect 118 1773 152 1807
rect 218 1773 252 1807
rect 318 1773 352 1807
rect 418 1773 452 1807
rect 518 1773 552 1807
rect 618 1773 652 1807
rect 718 1773 752 1807
rect 818 1773 852 1807
rect 918 1773 952 1807
rect 1018 1773 1052 1807
rect 1118 1773 1152 1807
rect 1218 1773 1252 1807
rect 1318 1773 1352 1807
rect 1418 1773 1452 1807
rect 1518 1773 1552 1807
rect 1618 1773 1652 1807
rect 1718 1773 1752 1807
rect 1818 1773 1852 1807
rect 1918 1773 1952 1807
rect 2018 1773 2052 1807
rect 2118 1773 2152 1807
rect 2218 1773 2252 1807
rect 2318 1773 2352 1807
rect 2418 1773 2452 1807
rect 2518 1773 2552 1807
rect 2618 1773 2652 1807
rect 2718 1773 2752 1807
rect 2818 1773 2852 1807
rect 2918 1773 2952 1807
rect 3018 1773 3052 1807
rect 3118 1773 3146 1807
rect 3146 1773 3152 1807
rect 3218 1773 3224 1807
rect 3224 1773 3252 1807
rect 3318 1773 3346 1807
rect 3346 1773 3352 1807
rect 3418 1773 3424 1807
rect 3424 1773 3452 1807
rect 3518 1773 3552 1807
rect 3618 1773 3652 1807
rect 3718 1773 3752 1807
rect 3818 1773 3852 1807
rect 3918 1773 3946 1807
rect 3946 1773 3952 1807
rect 4018 1773 4024 1807
rect 4024 1773 4052 1807
rect 4118 1773 4146 1807
rect 4146 1773 4152 1807
rect 4218 1773 4224 1807
rect 4224 1773 4252 1807
rect 4318 1773 4352 1807
rect 4418 1773 4452 1807
rect 4518 1773 4552 1807
rect 4618 1773 4652 1807
rect 4718 1773 4752 1807
rect 4818 1773 4846 1807
rect 4846 1773 4852 1807
rect 4918 1773 4924 1807
rect 4924 1773 4952 1807
rect 5018 1773 5052 1807
rect 5118 1773 5152 1807
rect 5218 1773 5252 1807
rect 5318 1773 5352 1807
rect 5418 1773 5452 1807
rect 5518 1773 5552 1807
rect 5618 1773 5652 1807
rect 5718 1773 5752 1807
rect 5818 1773 5852 1807
rect 5918 1773 5952 1807
rect 6018 1773 6052 1807
rect 6118 1773 6152 1807
rect 6218 1773 6252 1807
rect 6318 1773 6346 1807
rect 6346 1773 6352 1807
rect 6418 1773 6424 1807
rect 6424 1773 6452 1807
rect 6518 1773 6552 1807
rect 6618 1773 6652 1807
rect 6718 1773 6752 1807
rect 6818 1773 6852 1807
rect 6918 1773 6952 1807
rect 7018 1773 7052 1807
rect 7118 1773 7146 1807
rect 7146 1773 7152 1807
rect 7218 1773 7224 1807
rect 7224 1773 7252 1807
rect 7318 1773 7352 1807
rect 7418 1773 7446 1807
rect 7446 1773 7452 1807
rect 7518 1773 7524 1807
rect 7524 1773 7552 1807
rect 7618 1773 7652 1807
rect 7718 1773 7746 1807
rect 7746 1773 7752 1807
rect 7818 1773 7824 1807
rect 7824 1773 7852 1807
rect 7918 1773 7952 1807
rect 8018 1773 8046 1807
rect 8046 1773 8052 1807
rect 8118 1773 8124 1807
rect 8124 1773 8152 1807
rect 8218 1773 8252 1807
rect 8318 1773 8352 1807
rect 8418 1773 8452 1807
rect 8518 1773 8552 1807
rect 8618 1773 8646 1807
rect 8646 1773 8652 1807
rect 8718 1773 8724 1807
rect 8724 1773 8752 1807
rect 8818 1773 8852 1807
rect 8918 1773 8952 1807
rect 9018 1773 9052 1807
rect 9118 1773 9152 1807
rect 9218 1773 9252 1807
rect 9318 1773 9352 1807
rect 9418 1773 9452 1807
rect 9518 1773 9552 1807
rect 9618 1773 9652 1807
rect 9718 1773 9752 1807
rect 9818 1773 9846 1807
rect 9846 1773 9852 1807
rect 9918 1773 9924 1807
rect 9924 1773 9952 1807
rect 10018 1773 10046 1807
rect 10046 1773 10052 1807
rect 10118 1773 10124 1807
rect 10124 1773 10152 1807
rect 10218 1773 10246 1807
rect 10246 1773 10252 1807
rect 10318 1773 10324 1807
rect 10324 1773 10352 1807
rect 10418 1773 10446 1807
rect 10446 1773 10452 1807
rect 10518 1773 10524 1807
rect 10524 1773 10552 1807
rect 10618 1773 10652 1807
rect 10718 1773 10746 1807
rect 10746 1773 10752 1807
rect 10818 1773 10824 1807
rect 10824 1773 10852 1807
rect 10918 1773 10952 1807
rect 11018 1773 11052 1807
rect 11118 1773 11152 1807
rect 11218 1773 11252 1807
rect 11318 1773 11352 1807
rect 11418 1773 11452 1807
rect 11518 1773 11552 1807
rect 11618 1773 11646 1807
rect 11646 1773 11652 1807
rect 11718 1773 11724 1807
rect 11724 1773 11752 1807
rect 11818 1773 11852 1807
rect 11918 1773 11946 1807
rect 11946 1773 11952 1807
rect 12018 1773 12024 1807
rect 12024 1773 12052 1807
rect 12118 1773 12152 1807
rect 12218 1773 12252 1807
rect 12318 1773 12352 1807
rect 12418 1773 12452 1807
rect 12518 1773 12552 1807
rect 12618 1773 12652 1807
rect 12718 1773 12752 1807
rect 12818 1773 12846 1807
rect 12846 1773 12852 1807
rect 12916 1788 12924 1822
rect 12924 1788 12950 1822
rect 13120 1758 13146 1792
rect 13146 1758 13154 1792
rect 18 1633 52 1667
rect 118 1633 152 1667
rect 218 1633 252 1667
rect 318 1633 352 1667
rect 418 1633 452 1667
rect 518 1633 552 1667
rect 618 1633 646 1667
rect 646 1633 652 1667
rect 718 1633 724 1667
rect 724 1633 752 1667
rect 818 1633 852 1667
rect 918 1633 952 1667
rect 1018 1633 1046 1667
rect 1046 1633 1052 1667
rect 1118 1633 1124 1667
rect 1124 1633 1152 1667
rect 1218 1633 1246 1667
rect 1246 1633 1252 1667
rect 1318 1633 1324 1667
rect 1324 1633 1352 1667
rect 1418 1633 1452 1667
rect 1518 1633 1546 1667
rect 1546 1633 1552 1667
rect 1618 1633 1624 1667
rect 1624 1633 1652 1667
rect 1718 1633 1752 1667
rect 1818 1633 1852 1667
rect 1918 1633 1952 1667
rect 2018 1633 2052 1667
rect 2118 1633 2152 1667
rect 2218 1633 2252 1667
rect 2318 1633 2352 1667
rect 2418 1633 2452 1667
rect 2518 1633 2552 1667
rect 2618 1633 2646 1667
rect 2646 1633 2652 1667
rect 2718 1633 2724 1667
rect 2724 1633 2752 1667
rect 2818 1633 2852 1667
rect 2918 1633 2952 1667
rect 3018 1633 3052 1667
rect 3118 1633 3152 1667
rect 3218 1633 3252 1667
rect 3318 1633 3352 1667
rect 3418 1633 3452 1667
rect 3518 1633 3552 1667
rect 3618 1633 3652 1667
rect 3718 1633 3746 1667
rect 3746 1633 3752 1667
rect 3818 1633 3824 1667
rect 3824 1633 3852 1667
rect 3918 1633 3946 1667
rect 3946 1633 3952 1667
rect 4018 1633 4024 1667
rect 4024 1633 4052 1667
rect 4118 1633 4146 1667
rect 4146 1633 4152 1667
rect 4218 1633 4224 1667
rect 4224 1633 4252 1667
rect 4318 1633 4352 1667
rect 4418 1633 4446 1667
rect 4446 1633 4452 1667
rect 4518 1633 4524 1667
rect 4524 1633 4552 1667
rect 4618 1633 4652 1667
rect 4718 1633 4752 1667
rect 4818 1633 4852 1667
rect 4918 1633 4946 1667
rect 4946 1633 4952 1667
rect 5018 1633 5024 1667
rect 5024 1633 5052 1667
rect 5118 1633 5152 1667
rect 5218 1633 5246 1667
rect 5246 1633 5252 1667
rect 5318 1633 5324 1667
rect 5324 1633 5352 1667
rect 5418 1633 5452 1667
rect 5518 1633 5552 1667
rect 5618 1633 5646 1667
rect 5646 1633 5652 1667
rect 5718 1633 5724 1667
rect 5724 1633 5752 1667
rect 5818 1633 5852 1667
rect 5918 1633 5946 1667
rect 5946 1633 5952 1667
rect 6018 1633 6024 1667
rect 6024 1633 6052 1667
rect 6118 1633 6146 1667
rect 6146 1633 6152 1667
rect 6218 1633 6224 1667
rect 6224 1633 6252 1667
rect 6318 1633 6352 1667
rect 6418 1633 6452 1667
rect 6518 1633 6546 1667
rect 6546 1633 6552 1667
rect 6618 1633 6624 1667
rect 6624 1633 6652 1667
rect 6718 1633 6752 1667
rect 6818 1633 6852 1667
rect 6918 1633 6952 1667
rect 7018 1633 7052 1667
rect 7118 1633 7152 1667
rect 7218 1633 7252 1667
rect 7318 1633 7352 1667
rect 7418 1633 7452 1667
rect 7518 1633 7552 1667
rect 7618 1633 7652 1667
rect 7718 1633 7752 1667
rect 7818 1633 7852 1667
rect 7918 1633 7952 1667
rect 8018 1633 8052 1667
rect 8118 1633 8152 1667
rect 8218 1633 8252 1667
rect 8318 1633 8352 1667
rect 8418 1633 8452 1667
rect 8518 1633 8552 1667
rect 8618 1633 8652 1667
rect 8718 1633 8752 1667
rect 8818 1633 8852 1667
rect 8918 1633 8952 1667
rect 9018 1633 9052 1667
rect 9118 1633 9152 1667
rect 9218 1633 9252 1667
rect 9318 1633 9352 1667
rect 9418 1633 9452 1667
rect 9518 1633 9546 1667
rect 9546 1633 9552 1667
rect 9618 1633 9624 1667
rect 9624 1633 9652 1667
rect 9718 1633 9752 1667
rect 9818 1633 9852 1667
rect 9918 1633 9952 1667
rect 10018 1633 10052 1667
rect 10118 1633 10152 1667
rect 10218 1633 10252 1667
rect 10318 1633 10352 1667
rect 10418 1633 10452 1667
rect 10518 1633 10552 1667
rect 10618 1633 10652 1667
rect 10718 1633 10752 1667
rect 10818 1633 10852 1667
rect 10918 1633 10946 1667
rect 10946 1633 10952 1667
rect 11018 1633 11024 1667
rect 11024 1633 11052 1667
rect 11118 1633 11152 1667
rect 11218 1633 11252 1667
rect 11318 1633 11352 1667
rect 11418 1633 11452 1667
rect 11518 1633 11552 1667
rect 11618 1633 11652 1667
rect 11718 1633 11746 1667
rect 11746 1633 11752 1667
rect 11818 1633 11824 1667
rect 11824 1633 11852 1667
rect 11918 1633 11952 1667
rect 12018 1633 12052 1667
rect 12118 1633 12152 1667
rect 12218 1633 12252 1667
rect 12318 1633 12352 1667
rect 12418 1633 12452 1667
rect 12518 1633 12552 1667
rect 12618 1633 12652 1667
rect 12718 1633 12752 1667
rect 12818 1633 12852 1667
rect 12916 1648 12924 1682
rect 12924 1648 12950 1682
rect 13120 1618 13146 1652
rect 13146 1618 13154 1652
rect 18 1493 52 1527
rect 118 1493 152 1527
rect 218 1493 252 1527
rect 318 1493 352 1527
rect 418 1493 446 1527
rect 446 1493 452 1527
rect 518 1493 524 1527
rect 524 1493 552 1527
rect 618 1493 652 1527
rect 718 1493 752 1527
rect 818 1493 852 1527
rect 918 1493 952 1527
rect 1018 1493 1052 1527
rect 1118 1493 1152 1527
rect 1218 1493 1252 1527
rect 1318 1493 1352 1527
rect 1418 1493 1452 1527
rect 1518 1493 1552 1527
rect 1618 1493 1652 1527
rect 1718 1493 1752 1527
rect 1818 1493 1852 1527
rect 1918 1493 1952 1527
rect 2018 1493 2052 1527
rect 2118 1493 2152 1527
rect 2218 1493 2252 1527
rect 2318 1493 2352 1527
rect 2418 1493 2452 1527
rect 2518 1493 2546 1527
rect 2546 1493 2552 1527
rect 2618 1493 2624 1527
rect 2624 1493 2652 1527
rect 2718 1493 2752 1527
rect 2818 1493 2852 1527
rect 2918 1493 2952 1527
rect 3018 1493 3052 1527
rect 3118 1493 3146 1527
rect 3146 1493 3152 1527
rect 3218 1493 3224 1527
rect 3224 1493 3252 1527
rect 3318 1493 3352 1527
rect 3418 1493 3452 1527
rect 3518 1493 3546 1527
rect 3546 1493 3552 1527
rect 3618 1493 3624 1527
rect 3624 1493 3652 1527
rect 3718 1493 3752 1527
rect 3818 1493 3852 1527
rect 3918 1493 3952 1527
rect 4018 1493 4046 1527
rect 4046 1493 4052 1527
rect 4118 1493 4124 1527
rect 4124 1493 4152 1527
rect 4218 1493 4252 1527
rect 4318 1493 4352 1527
rect 4418 1493 4452 1527
rect 4518 1493 4552 1527
rect 4618 1493 4652 1527
rect 4718 1493 4752 1527
rect 4818 1493 4846 1527
rect 4846 1493 4852 1527
rect 4918 1493 4924 1527
rect 4924 1493 4952 1527
rect 5018 1493 5052 1527
rect 5118 1493 5152 1527
rect 5218 1493 5252 1527
rect 5318 1493 5352 1527
rect 5418 1493 5452 1527
rect 5518 1493 5552 1527
rect 5618 1493 5652 1527
rect 5718 1493 5752 1527
rect 5818 1493 5846 1527
rect 5846 1493 5852 1527
rect 5918 1493 5924 1527
rect 5924 1493 5952 1527
rect 6018 1493 6046 1527
rect 6046 1493 6052 1527
rect 6118 1493 6124 1527
rect 6124 1493 6152 1527
rect 6218 1493 6252 1527
rect 6318 1493 6346 1527
rect 6346 1493 6352 1527
rect 6418 1493 6424 1527
rect 6424 1493 6452 1527
rect 6518 1493 6552 1527
rect 6618 1493 6652 1527
rect 6718 1493 6752 1527
rect 6818 1493 6852 1527
rect 6918 1493 6952 1527
rect 7018 1493 7052 1527
rect 7118 1493 7152 1527
rect 7218 1493 7252 1527
rect 7318 1493 7352 1527
rect 7418 1493 7452 1527
rect 7518 1493 7552 1527
rect 7618 1493 7652 1527
rect 7718 1493 7746 1527
rect 7746 1493 7752 1527
rect 7818 1493 7824 1527
rect 7824 1493 7852 1527
rect 7918 1493 7946 1527
rect 7946 1493 7952 1527
rect 8018 1493 8024 1527
rect 8024 1493 8052 1527
rect 8118 1493 8152 1527
rect 8218 1493 8252 1527
rect 8318 1493 8352 1527
rect 8418 1493 8452 1527
rect 8518 1493 8546 1527
rect 8546 1493 8552 1527
rect 8618 1493 8624 1527
rect 8624 1493 8652 1527
rect 8718 1493 8752 1527
rect 8818 1493 8852 1527
rect 8918 1493 8952 1527
rect 9018 1493 9052 1527
rect 9118 1493 9152 1527
rect 9218 1493 9252 1527
rect 9318 1493 9346 1527
rect 9346 1493 9352 1527
rect 9418 1493 9424 1527
rect 9424 1493 9452 1527
rect 9518 1493 9552 1527
rect 9618 1493 9652 1527
rect 9718 1493 9752 1527
rect 9818 1493 9852 1527
rect 9918 1493 9952 1527
rect 10018 1493 10052 1527
rect 10118 1493 10152 1527
rect 10218 1493 10252 1527
rect 10318 1493 10352 1527
rect 10418 1493 10452 1527
rect 10518 1493 10552 1527
rect 10618 1493 10652 1527
rect 10718 1493 10752 1527
rect 10818 1493 10852 1527
rect 10918 1493 10946 1527
rect 10946 1493 10952 1527
rect 11018 1493 11024 1527
rect 11024 1493 11052 1527
rect 11118 1493 11146 1527
rect 11146 1493 11152 1527
rect 11218 1493 11224 1527
rect 11224 1493 11252 1527
rect 11318 1493 11352 1527
rect 11418 1493 11452 1527
rect 11518 1493 11552 1527
rect 11618 1493 11652 1527
rect 11718 1493 11752 1527
rect 11818 1493 11852 1527
rect 11918 1493 11952 1527
rect 12018 1493 12046 1527
rect 12046 1493 12052 1527
rect 12118 1493 12124 1527
rect 12124 1493 12152 1527
rect 12218 1493 12252 1527
rect 12318 1493 12352 1527
rect 12418 1493 12446 1527
rect 12446 1493 12452 1527
rect 12518 1493 12524 1527
rect 12524 1493 12552 1527
rect 12618 1493 12652 1527
rect 12718 1493 12752 1527
rect 12818 1493 12852 1527
rect 12916 1508 12924 1542
rect 12924 1508 12950 1542
rect 13120 1478 13146 1512
rect 13146 1478 13154 1512
rect 18 1353 52 1387
rect 118 1353 152 1387
rect 218 1353 252 1387
rect 318 1353 352 1387
rect 418 1353 452 1387
rect 518 1353 552 1387
rect 618 1353 652 1387
rect 718 1353 752 1387
rect 818 1353 846 1387
rect 846 1353 852 1387
rect 918 1353 924 1387
rect 924 1353 952 1387
rect 1018 1353 1052 1387
rect 1118 1353 1152 1387
rect 1218 1353 1252 1387
rect 1318 1353 1352 1387
rect 1418 1353 1452 1387
rect 1518 1353 1552 1387
rect 1618 1353 1652 1387
rect 1718 1353 1752 1387
rect 1818 1353 1852 1387
rect 1918 1353 1952 1387
rect 2018 1353 2052 1387
rect 2118 1353 2152 1387
rect 2218 1353 2252 1387
rect 2318 1353 2352 1387
rect 2418 1353 2452 1387
rect 2518 1353 2552 1387
rect 2618 1353 2652 1387
rect 2718 1353 2752 1387
rect 2818 1353 2846 1387
rect 2846 1353 2852 1387
rect 2918 1353 2924 1387
rect 2924 1353 2952 1387
rect 3018 1353 3052 1387
rect 3118 1353 3152 1387
rect 3218 1353 3252 1387
rect 3318 1353 3352 1387
rect 3418 1353 3452 1387
rect 3518 1353 3552 1387
rect 3618 1353 3652 1387
rect 3718 1353 3752 1387
rect 3818 1353 3852 1387
rect 3918 1353 3952 1387
rect 4018 1353 4052 1387
rect 4118 1353 4152 1387
rect 4218 1353 4252 1387
rect 4318 1353 4352 1387
rect 4418 1353 4452 1387
rect 4518 1353 4552 1387
rect 4618 1353 4646 1387
rect 4646 1353 4652 1387
rect 4718 1353 4724 1387
rect 4724 1353 4752 1387
rect 4818 1353 4846 1387
rect 4846 1353 4852 1387
rect 4918 1353 4924 1387
rect 4924 1353 4952 1387
rect 5018 1353 5052 1387
rect 5118 1353 5146 1387
rect 5146 1353 5152 1387
rect 5218 1353 5224 1387
rect 5224 1353 5252 1387
rect 5318 1353 5352 1387
rect 5418 1353 5452 1387
rect 5518 1353 5552 1387
rect 5618 1353 5652 1387
rect 5718 1353 5752 1387
rect 5818 1353 5852 1387
rect 5918 1353 5952 1387
rect 6018 1353 6052 1387
rect 6118 1353 6152 1387
rect 6218 1353 6246 1387
rect 6246 1353 6252 1387
rect 6318 1353 6324 1387
rect 6324 1353 6352 1387
rect 6418 1353 6446 1387
rect 6446 1353 6452 1387
rect 6518 1353 6524 1387
rect 6524 1353 6552 1387
rect 6618 1353 6652 1387
rect 6718 1353 6746 1387
rect 6746 1353 6752 1387
rect 6818 1353 6824 1387
rect 6824 1353 6852 1387
rect 6918 1353 6946 1387
rect 6946 1353 6952 1387
rect 7018 1353 7024 1387
rect 7024 1353 7052 1387
rect 7118 1353 7152 1387
rect 7218 1353 7252 1387
rect 7318 1353 7352 1387
rect 7418 1353 7452 1387
rect 7518 1353 7552 1387
rect 7618 1353 7652 1387
rect 7718 1353 7752 1387
rect 7818 1353 7852 1387
rect 7918 1353 7946 1387
rect 7946 1353 7952 1387
rect 8018 1353 8024 1387
rect 8024 1353 8052 1387
rect 8118 1353 8152 1387
rect 8218 1353 8252 1387
rect 8318 1353 8352 1387
rect 8418 1353 8452 1387
rect 8518 1353 8552 1387
rect 8618 1353 8652 1387
rect 8718 1353 8752 1387
rect 8818 1353 8852 1387
rect 8918 1353 8952 1387
rect 9018 1353 9052 1387
rect 9118 1353 9152 1387
rect 9218 1353 9252 1387
rect 9318 1353 9346 1387
rect 9346 1353 9352 1387
rect 9418 1353 9424 1387
rect 9424 1353 9452 1387
rect 9518 1353 9552 1387
rect 9618 1353 9652 1387
rect 9718 1353 9752 1387
rect 9818 1353 9852 1387
rect 9918 1353 9952 1387
rect 10018 1353 10052 1387
rect 10118 1353 10152 1387
rect 10218 1353 10246 1387
rect 10246 1353 10252 1387
rect 10318 1353 10324 1387
rect 10324 1353 10352 1387
rect 10418 1353 10452 1387
rect 10518 1353 10552 1387
rect 10618 1353 10652 1387
rect 10718 1353 10752 1387
rect 10818 1353 10852 1387
rect 10918 1353 10952 1387
rect 11018 1353 11052 1387
rect 11118 1353 11146 1387
rect 11146 1353 11152 1387
rect 11218 1353 11224 1387
rect 11224 1353 11252 1387
rect 11318 1353 11352 1387
rect 11418 1353 11452 1387
rect 11518 1353 11552 1387
rect 11618 1353 11652 1387
rect 11718 1353 11746 1387
rect 11746 1353 11752 1387
rect 11818 1353 11824 1387
rect 11824 1353 11852 1387
rect 11918 1353 11952 1387
rect 12018 1353 12052 1387
rect 12118 1353 12152 1387
rect 12218 1353 12252 1387
rect 12318 1353 12352 1387
rect 12418 1353 12446 1387
rect 12446 1353 12452 1387
rect 12518 1353 12524 1387
rect 12524 1353 12552 1387
rect 12618 1353 12652 1387
rect 12718 1353 12752 1387
rect 12818 1353 12852 1387
rect 12916 1368 12924 1402
rect 12924 1368 12950 1402
rect 13120 1338 13146 1372
rect 13146 1338 13154 1372
rect 18 1230 52 1264
rect 218 1246 252 1280
rect 418 1230 452 1264
rect 618 1246 652 1280
rect 818 1230 852 1264
rect 1018 1246 1052 1280
rect 1218 1230 1252 1264
rect 1418 1246 1452 1280
rect 1618 1230 1652 1264
rect 1818 1246 1852 1280
rect 2018 1230 2052 1264
rect 2218 1246 2252 1280
rect 2418 1230 2452 1264
rect 2618 1246 2652 1280
rect 2818 1230 2852 1264
rect 3018 1246 3052 1280
rect 3218 1230 3252 1264
rect 3418 1246 3452 1280
rect 3618 1230 3652 1264
rect 3818 1246 3852 1280
rect 4018 1230 4052 1264
rect 4218 1246 4252 1280
rect 4418 1230 4452 1264
rect 4618 1246 4652 1280
rect 4818 1230 4852 1264
rect 5018 1246 5052 1280
rect 5218 1230 5252 1264
rect 5418 1246 5452 1280
rect 5618 1230 5652 1264
rect 5818 1246 5852 1280
rect 6018 1230 6052 1264
rect 6218 1246 6252 1280
rect 6418 1230 6452 1264
rect 6618 1246 6652 1280
rect 6818 1230 6852 1264
rect 7018 1246 7052 1280
rect 7218 1230 7252 1264
rect 7418 1246 7452 1280
rect 7618 1230 7652 1264
rect 7818 1246 7852 1280
rect 8018 1230 8052 1264
rect 8218 1246 8252 1280
rect 8418 1230 8452 1264
rect 8618 1246 8652 1280
rect 8818 1230 8852 1264
rect 9018 1246 9052 1280
rect 9218 1230 9252 1264
rect 9418 1246 9452 1280
rect 9618 1230 9652 1264
rect 9818 1246 9852 1280
rect 10018 1230 10052 1264
rect 10218 1246 10252 1280
rect 10418 1230 10452 1264
rect 10618 1246 10652 1280
rect 10818 1230 10852 1264
rect 11018 1246 11052 1280
rect 11218 1230 11252 1264
rect 11418 1246 11452 1280
rect 11618 1230 11652 1264
rect 11818 1246 11852 1280
rect 12018 1230 12052 1264
rect 12218 1246 12252 1280
rect 12418 1230 12452 1264
rect 12618 1246 12652 1280
rect 12916 1227 12950 1261
rect 13120 1249 13154 1283
rect 13278 1244 13312 1278
rect 13378 1244 13412 1278
rect 13478 1244 13512 1278
rect 13578 1244 13612 1278
rect 18 1123 52 1157
rect 118 1123 152 1157
rect 218 1123 252 1157
rect 318 1123 352 1157
rect 418 1123 452 1157
rect 518 1123 552 1157
rect 618 1123 652 1157
rect 718 1123 752 1157
rect 818 1123 852 1157
rect 918 1123 952 1157
rect 1018 1123 1052 1157
rect 1118 1123 1152 1157
rect 1218 1123 1252 1157
rect 1318 1123 1352 1157
rect 1418 1123 1452 1157
rect 1518 1123 1552 1157
rect 1618 1123 1652 1157
rect 1718 1123 1746 1157
rect 1746 1123 1752 1157
rect 1818 1123 1824 1157
rect 1824 1123 1852 1157
rect 1918 1123 1952 1157
rect 2018 1123 2046 1157
rect 2046 1123 2052 1157
rect 2118 1123 2124 1157
rect 2124 1123 2152 1157
rect 2218 1123 2252 1157
rect 2318 1123 2352 1157
rect 2418 1123 2452 1157
rect 2518 1123 2552 1157
rect 2618 1123 2652 1157
rect 2718 1123 2752 1157
rect 2818 1123 2852 1157
rect 2918 1123 2952 1157
rect 3018 1123 3046 1157
rect 3046 1123 3052 1157
rect 3118 1123 3124 1157
rect 3124 1123 3152 1157
rect 3218 1123 3246 1157
rect 3246 1123 3252 1157
rect 3318 1123 3324 1157
rect 3324 1123 3352 1157
rect 3418 1123 3452 1157
rect 3518 1123 3552 1157
rect 3618 1123 3652 1157
rect 3718 1123 3746 1157
rect 3746 1123 3752 1157
rect 3818 1123 3824 1157
rect 3824 1123 3852 1157
rect 3918 1123 3952 1157
rect 4018 1123 4052 1157
rect 4118 1123 4152 1157
rect 4218 1123 4252 1157
rect 4318 1123 4352 1157
rect 4418 1123 4446 1157
rect 4446 1123 4452 1157
rect 4518 1123 4524 1157
rect 4524 1123 4552 1157
rect 4618 1123 4646 1157
rect 4646 1123 4652 1157
rect 4718 1123 4724 1157
rect 4724 1123 4752 1157
rect 4818 1123 4852 1157
rect 4918 1123 4952 1157
rect 5018 1123 5052 1157
rect 5118 1123 5152 1157
rect 5218 1123 5252 1157
rect 5318 1123 5352 1157
rect 5418 1123 5446 1157
rect 5446 1123 5452 1157
rect 5518 1123 5524 1157
rect 5524 1123 5552 1157
rect 5618 1123 5652 1157
rect 5718 1123 5752 1157
rect 5818 1123 5852 1157
rect 5918 1123 5952 1157
rect 6018 1123 6052 1157
rect 6118 1123 6152 1157
rect 6218 1123 6252 1157
rect 6318 1123 6352 1157
rect 6418 1123 6452 1157
rect 6518 1123 6552 1157
rect 6618 1123 6652 1157
rect 6718 1123 6746 1157
rect 6746 1123 6752 1157
rect 6818 1123 6824 1157
rect 6824 1123 6852 1157
rect 6918 1123 6952 1157
rect 7018 1123 7052 1157
rect 7118 1123 7152 1157
rect 7218 1123 7252 1157
rect 7318 1123 7352 1157
rect 7418 1123 7452 1157
rect 7518 1123 7552 1157
rect 7618 1123 7652 1157
rect 7718 1123 7752 1157
rect 7818 1123 7852 1157
rect 7918 1123 7952 1157
rect 8018 1123 8052 1157
rect 8118 1123 8152 1157
rect 8218 1123 8252 1157
rect 8318 1123 8352 1157
rect 8418 1123 8452 1157
rect 8518 1123 8552 1157
rect 8618 1123 8652 1157
rect 8718 1123 8752 1157
rect 8818 1123 8852 1157
rect 8918 1123 8952 1157
rect 9018 1123 9052 1157
rect 9118 1123 9152 1157
rect 9218 1123 9252 1157
rect 9318 1123 9352 1157
rect 9418 1123 9452 1157
rect 9518 1123 9552 1157
rect 9618 1123 9646 1157
rect 9646 1123 9652 1157
rect 9718 1123 9724 1157
rect 9724 1123 9752 1157
rect 9818 1123 9852 1157
rect 9918 1123 9952 1157
rect 10018 1123 10052 1157
rect 10118 1123 10152 1157
rect 10218 1123 10252 1157
rect 10318 1123 10352 1157
rect 10418 1123 10452 1157
rect 10518 1123 10552 1157
rect 10618 1123 10652 1157
rect 10718 1123 10752 1157
rect 10818 1123 10852 1157
rect 10918 1123 10952 1157
rect 11018 1123 11046 1157
rect 11046 1123 11052 1157
rect 11118 1123 11124 1157
rect 11124 1123 11152 1157
rect 11218 1123 11246 1157
rect 11246 1123 11252 1157
rect 11318 1123 11324 1157
rect 11324 1123 11352 1157
rect 11418 1123 11446 1157
rect 11446 1123 11452 1157
rect 11518 1123 11524 1157
rect 11524 1123 11552 1157
rect 11618 1123 11652 1157
rect 11718 1123 11752 1157
rect 11818 1123 11852 1157
rect 11918 1123 11952 1157
rect 12018 1123 12046 1157
rect 12046 1123 12052 1157
rect 12118 1123 12124 1157
rect 12124 1123 12152 1157
rect 12218 1123 12252 1157
rect 12318 1123 12352 1157
rect 12418 1123 12452 1157
rect 12518 1123 12552 1157
rect 12618 1123 12646 1157
rect 12646 1123 12652 1157
rect 12718 1123 12724 1157
rect 12724 1123 12752 1157
rect 12818 1123 12846 1157
rect 12846 1123 12852 1157
rect 12916 1138 12924 1172
rect 12924 1138 12950 1172
rect 13120 1108 13146 1142
rect 13146 1108 13154 1142
rect 18 983 24 1017
rect 24 983 52 1017
rect 118 983 146 1017
rect 146 983 152 1017
rect 218 983 224 1017
rect 224 983 252 1017
rect 318 983 352 1017
rect 418 983 452 1017
rect 518 983 552 1017
rect 618 983 646 1017
rect 646 983 652 1017
rect 718 983 724 1017
rect 724 983 752 1017
rect 818 983 852 1017
rect 918 983 952 1017
rect 1018 983 1052 1017
rect 1118 983 1152 1017
rect 1218 983 1246 1017
rect 1246 983 1252 1017
rect 1318 983 1324 1017
rect 1324 983 1352 1017
rect 1418 983 1452 1017
rect 1518 983 1552 1017
rect 1618 983 1652 1017
rect 1718 983 1752 1017
rect 1818 983 1852 1017
rect 1918 983 1952 1017
rect 2018 983 2052 1017
rect 2118 983 2152 1017
rect 2218 983 2252 1017
rect 2318 983 2352 1017
rect 2418 983 2452 1017
rect 2518 983 2552 1017
rect 2618 983 2646 1017
rect 2646 983 2652 1017
rect 2718 983 2724 1017
rect 2724 983 2752 1017
rect 2818 983 2846 1017
rect 2846 983 2852 1017
rect 2918 983 2924 1017
rect 2924 983 2952 1017
rect 3018 983 3052 1017
rect 3118 983 3146 1017
rect 3146 983 3152 1017
rect 3218 983 3224 1017
rect 3224 983 3252 1017
rect 3318 983 3346 1017
rect 3346 983 3352 1017
rect 3418 983 3424 1017
rect 3424 983 3452 1017
rect 3518 983 3552 1017
rect 3618 983 3646 1017
rect 3646 983 3652 1017
rect 3718 983 3724 1017
rect 3724 983 3752 1017
rect 3818 983 3846 1017
rect 3846 983 3852 1017
rect 3918 983 3924 1017
rect 3924 983 3952 1017
rect 4018 983 4052 1017
rect 4118 983 4152 1017
rect 4218 983 4252 1017
rect 4318 983 4352 1017
rect 4418 983 4452 1017
rect 4518 983 4552 1017
rect 4618 983 4652 1017
rect 4718 983 4752 1017
rect 4818 983 4846 1017
rect 4846 983 4852 1017
rect 4918 983 4924 1017
rect 4924 983 4952 1017
rect 5018 983 5052 1017
rect 5118 983 5152 1017
rect 5218 983 5252 1017
rect 5318 983 5346 1017
rect 5346 983 5352 1017
rect 5418 983 5424 1017
rect 5424 983 5452 1017
rect 5518 983 5552 1017
rect 5618 983 5652 1017
rect 5718 983 5752 1017
rect 5818 983 5852 1017
rect 5918 983 5952 1017
rect 6018 983 6052 1017
rect 6118 983 6152 1017
rect 6218 983 6252 1017
rect 6318 983 6352 1017
rect 6418 983 6446 1017
rect 6446 983 6452 1017
rect 6518 983 6524 1017
rect 6524 983 6552 1017
rect 6618 983 6652 1017
rect 6718 983 6752 1017
rect 6818 983 6852 1017
rect 6918 983 6946 1017
rect 6946 983 6952 1017
rect 7018 983 7024 1017
rect 7024 983 7052 1017
rect 7118 983 7146 1017
rect 7146 983 7152 1017
rect 7218 983 7224 1017
rect 7224 983 7252 1017
rect 7318 983 7346 1017
rect 7346 983 7352 1017
rect 7418 983 7424 1017
rect 7424 983 7452 1017
rect 7518 983 7552 1017
rect 7618 983 7652 1017
rect 7718 983 7752 1017
rect 7818 983 7852 1017
rect 7918 983 7952 1017
rect 8018 983 8052 1017
rect 8118 983 8152 1017
rect 8218 983 8252 1017
rect 8318 983 8352 1017
rect 8418 983 8452 1017
rect 8518 983 8552 1017
rect 8618 983 8646 1017
rect 8646 983 8652 1017
rect 8718 983 8724 1017
rect 8724 983 8752 1017
rect 8818 983 8846 1017
rect 8846 983 8852 1017
rect 8918 983 8924 1017
rect 8924 983 8952 1017
rect 9018 983 9052 1017
rect 9118 983 9152 1017
rect 9218 983 9252 1017
rect 9318 983 9352 1017
rect 9418 983 9452 1017
rect 9518 983 9546 1017
rect 9546 983 9552 1017
rect 9618 983 9624 1017
rect 9624 983 9652 1017
rect 9718 983 9752 1017
rect 9818 983 9852 1017
rect 9918 983 9946 1017
rect 9946 983 9952 1017
rect 10018 983 10024 1017
rect 10024 983 10052 1017
rect 10118 983 10152 1017
rect 10218 983 10252 1017
rect 10318 983 10346 1017
rect 10346 983 10352 1017
rect 10418 983 10424 1017
rect 10424 983 10452 1017
rect 10518 983 10552 1017
rect 10618 983 10652 1017
rect 10718 983 10752 1017
rect 10818 983 10852 1017
rect 10918 983 10952 1017
rect 11018 983 11052 1017
rect 11118 983 11152 1017
rect 11218 983 11252 1017
rect 11318 983 11346 1017
rect 11346 983 11352 1017
rect 11418 983 11424 1017
rect 11424 983 11452 1017
rect 11518 983 11552 1017
rect 11618 983 11646 1017
rect 11646 983 11652 1017
rect 11718 983 11724 1017
rect 11724 983 11752 1017
rect 11818 983 11852 1017
rect 11918 983 11946 1017
rect 11946 983 11952 1017
rect 12018 983 12024 1017
rect 12024 983 12052 1017
rect 12118 983 12152 1017
rect 12218 983 12252 1017
rect 12318 983 12352 1017
rect 12418 983 12452 1017
rect 12518 983 12552 1017
rect 12618 983 12652 1017
rect 12718 983 12752 1017
rect 12818 983 12846 1017
rect 12846 983 12852 1017
rect 12916 998 12924 1032
rect 12924 998 12950 1032
rect 13120 968 13146 1002
rect 13146 968 13154 1002
rect 18 843 24 877
rect 24 843 52 877
rect 118 843 146 877
rect 146 843 152 877
rect 218 843 224 877
rect 224 843 252 877
rect 318 843 352 877
rect 418 843 452 877
rect 518 843 552 877
rect 618 843 652 877
rect 718 843 752 877
rect 818 843 852 877
rect 918 843 952 877
rect 1018 843 1052 877
rect 1118 843 1152 877
rect 1218 843 1252 877
rect 1318 843 1352 877
rect 1418 843 1452 877
rect 1518 843 1552 877
rect 1618 843 1652 877
rect 1718 843 1752 877
rect 1818 843 1852 877
rect 1918 843 1952 877
rect 2018 843 2052 877
rect 2118 843 2152 877
rect 2218 843 2252 877
rect 2318 843 2352 877
rect 2418 843 2452 877
rect 2518 843 2552 877
rect 2618 843 2652 877
rect 2718 843 2752 877
rect 2818 843 2852 877
rect 2918 843 2946 877
rect 2946 843 2952 877
rect 3018 843 3024 877
rect 3024 843 3052 877
rect 3118 843 3152 877
rect 3218 843 3252 877
rect 3318 843 3352 877
rect 3418 843 3452 877
rect 3518 843 3552 877
rect 3618 843 3652 877
rect 3718 843 3752 877
rect 3818 843 3846 877
rect 3846 843 3852 877
rect 3918 843 3924 877
rect 3924 843 3952 877
rect 4018 843 4052 877
rect 4118 843 4152 877
rect 4218 843 4252 877
rect 4318 843 4352 877
rect 4418 843 4452 877
rect 4518 843 4552 877
rect 4618 843 4652 877
rect 4718 843 4752 877
rect 4818 843 4852 877
rect 4918 843 4952 877
rect 5018 843 5052 877
rect 5118 843 5152 877
rect 5218 843 5252 877
rect 5318 843 5352 877
rect 5418 843 5452 877
rect 5518 843 5552 877
rect 5618 843 5652 877
rect 5718 843 5752 877
rect 5818 843 5852 877
rect 5918 843 5952 877
rect 6018 843 6052 877
rect 6118 843 6152 877
rect 6218 843 6252 877
rect 6318 843 6352 877
rect 6418 843 6452 877
rect 6518 843 6552 877
rect 6618 843 6646 877
rect 6646 843 6652 877
rect 6718 843 6724 877
rect 6724 843 6752 877
rect 6818 843 6852 877
rect 6918 843 6952 877
rect 7018 843 7052 877
rect 7118 843 7152 877
rect 7218 843 7252 877
rect 7318 843 7346 877
rect 7346 843 7352 877
rect 7418 843 7424 877
rect 7424 843 7452 877
rect 7518 843 7546 877
rect 7546 843 7552 877
rect 7618 843 7624 877
rect 7624 843 7652 877
rect 7718 843 7746 877
rect 7746 843 7752 877
rect 7818 843 7824 877
rect 7824 843 7852 877
rect 7918 843 7946 877
rect 7946 843 7952 877
rect 8018 843 8024 877
rect 8024 843 8052 877
rect 8118 843 8152 877
rect 8218 843 8252 877
rect 8318 843 8352 877
rect 8418 843 8452 877
rect 8518 843 8552 877
rect 8618 843 8646 877
rect 8646 843 8652 877
rect 8718 843 8724 877
rect 8724 843 8752 877
rect 8818 843 8846 877
rect 8846 843 8852 877
rect 8918 843 8924 877
rect 8924 843 8952 877
rect 9018 843 9052 877
rect 9118 843 9152 877
rect 9218 843 9252 877
rect 9318 843 9352 877
rect 9418 843 9452 877
rect 9518 843 9552 877
rect 9618 843 9652 877
rect 9718 843 9752 877
rect 9818 843 9852 877
rect 9918 843 9946 877
rect 9946 843 9952 877
rect 10018 843 10024 877
rect 10024 843 10052 877
rect 10118 843 10152 877
rect 10218 843 10252 877
rect 10318 843 10352 877
rect 10418 843 10452 877
rect 10518 843 10552 877
rect 10618 843 10652 877
rect 10718 843 10746 877
rect 10746 843 10752 877
rect 10818 843 10824 877
rect 10824 843 10852 877
rect 10918 843 10946 877
rect 10946 843 10952 877
rect 11018 843 11024 877
rect 11024 843 11052 877
rect 11118 843 11152 877
rect 11218 843 11252 877
rect 11318 843 11352 877
rect 11418 843 11452 877
rect 11518 843 11552 877
rect 11618 843 11652 877
rect 11718 843 11752 877
rect 11818 843 11852 877
rect 11918 843 11946 877
rect 11946 843 11952 877
rect 12018 843 12024 877
rect 12024 843 12052 877
rect 12118 843 12152 877
rect 12218 843 12252 877
rect 12318 843 12346 877
rect 12346 843 12352 877
rect 12418 843 12424 877
rect 12424 843 12452 877
rect 12518 843 12546 877
rect 12546 843 12552 877
rect 12618 843 12624 877
rect 12624 843 12652 877
rect 12718 843 12752 877
rect 12818 843 12852 877
rect 12916 858 12924 892
rect 12924 858 12950 892
rect 13120 828 13146 862
rect 13146 828 13154 862
rect 18 703 52 737
rect 118 703 152 737
rect 218 703 252 737
rect 318 703 352 737
rect 418 703 452 737
rect 518 703 546 737
rect 546 703 552 737
rect 618 703 624 737
rect 624 703 652 737
rect 718 703 746 737
rect 746 703 752 737
rect 818 703 824 737
rect 824 703 852 737
rect 918 703 952 737
rect 1018 703 1052 737
rect 1118 703 1152 737
rect 1218 703 1246 737
rect 1246 703 1252 737
rect 1318 703 1324 737
rect 1324 703 1352 737
rect 1418 703 1446 737
rect 1446 703 1452 737
rect 1518 703 1524 737
rect 1524 703 1552 737
rect 1618 703 1652 737
rect 1718 703 1752 737
rect 1818 703 1852 737
rect 1918 703 1952 737
rect 2018 703 2046 737
rect 2046 703 2052 737
rect 2118 703 2124 737
rect 2124 703 2152 737
rect 2218 703 2252 737
rect 2318 703 2352 737
rect 2418 703 2446 737
rect 2446 703 2452 737
rect 2518 703 2524 737
rect 2524 703 2552 737
rect 2618 703 2652 737
rect 2718 703 2752 737
rect 2818 703 2846 737
rect 2846 703 2852 737
rect 2918 703 2924 737
rect 2924 703 2952 737
rect 3018 703 3046 737
rect 3046 703 3052 737
rect 3118 703 3124 737
rect 3124 703 3152 737
rect 3218 703 3252 737
rect 3318 703 3346 737
rect 3346 703 3352 737
rect 3418 703 3424 737
rect 3424 703 3452 737
rect 3518 703 3552 737
rect 3618 703 3646 737
rect 3646 703 3652 737
rect 3718 703 3724 737
rect 3724 703 3752 737
rect 3818 703 3852 737
rect 3918 703 3952 737
rect 4018 703 4052 737
rect 4118 703 4152 737
rect 4218 703 4252 737
rect 4318 703 4352 737
rect 4418 703 4452 737
rect 4518 703 4552 737
rect 4618 703 4646 737
rect 4646 703 4652 737
rect 4718 703 4724 737
rect 4724 703 4752 737
rect 4818 703 4852 737
rect 4918 703 4952 737
rect 5018 703 5052 737
rect 5118 703 5146 737
rect 5146 703 5152 737
rect 5218 703 5224 737
rect 5224 703 5252 737
rect 5318 703 5352 737
rect 5418 703 5452 737
rect 5518 703 5552 737
rect 5618 703 5652 737
rect 5718 703 5746 737
rect 5746 703 5752 737
rect 5818 703 5824 737
rect 5824 703 5852 737
rect 5918 703 5952 737
rect 6018 703 6052 737
rect 6118 703 6152 737
rect 6218 703 6246 737
rect 6246 703 6252 737
rect 6318 703 6324 737
rect 6324 703 6352 737
rect 6418 703 6446 737
rect 6446 703 6452 737
rect 6518 703 6524 737
rect 6524 703 6552 737
rect 6618 703 6652 737
rect 6718 703 6752 737
rect 6818 703 6852 737
rect 6918 703 6952 737
rect 7018 703 7046 737
rect 7046 703 7052 737
rect 7118 703 7124 737
rect 7124 703 7152 737
rect 7218 703 7252 737
rect 7318 703 7352 737
rect 7418 703 7452 737
rect 7518 703 7552 737
rect 7618 703 7652 737
rect 7718 703 7752 737
rect 7818 703 7852 737
rect 7918 703 7952 737
rect 8018 703 8052 737
rect 8118 703 8152 737
rect 8218 703 8252 737
rect 8318 703 8352 737
rect 8418 703 8452 737
rect 8518 703 8552 737
rect 8618 703 8652 737
rect 8718 703 8752 737
rect 8818 703 8852 737
rect 8918 703 8952 737
rect 9018 703 9052 737
rect 9118 703 9146 737
rect 9146 703 9152 737
rect 9218 703 9224 737
rect 9224 703 9252 737
rect 9318 703 9346 737
rect 9346 703 9352 737
rect 9418 703 9424 737
rect 9424 703 9452 737
rect 9518 703 9552 737
rect 9618 703 9646 737
rect 9646 703 9652 737
rect 9718 703 9724 737
rect 9724 703 9752 737
rect 9818 703 9846 737
rect 9846 703 9852 737
rect 9918 703 9924 737
rect 9924 703 9952 737
rect 10018 703 10052 737
rect 10118 703 10146 737
rect 10146 703 10152 737
rect 10218 703 10224 737
rect 10224 703 10252 737
rect 10318 703 10352 737
rect 10418 703 10452 737
rect 10518 703 10552 737
rect 10618 703 10652 737
rect 10718 703 10752 737
rect 10818 703 10852 737
rect 10918 703 10946 737
rect 10946 703 10952 737
rect 11018 703 11024 737
rect 11024 703 11052 737
rect 11118 703 11152 737
rect 11218 703 11252 737
rect 11318 703 11352 737
rect 11418 703 11452 737
rect 11518 703 11552 737
rect 11618 703 11652 737
rect 11718 703 11746 737
rect 11746 703 11752 737
rect 11818 703 11824 737
rect 11824 703 11852 737
rect 11918 703 11952 737
rect 12018 703 12052 737
rect 12118 703 12146 737
rect 12146 703 12152 737
rect 12218 703 12224 737
rect 12224 703 12252 737
rect 12318 703 12352 737
rect 12418 703 12452 737
rect 12518 703 12552 737
rect 12618 703 12652 737
rect 12718 703 12752 737
rect 12818 703 12852 737
rect 12916 718 12924 752
rect 12924 718 12950 752
rect 13120 688 13146 722
rect 13146 688 13154 722
rect 18 563 52 597
rect 118 563 152 597
rect 218 563 252 597
rect 318 563 352 597
rect 418 563 452 597
rect 518 563 552 597
rect 618 563 652 597
rect 718 563 746 597
rect 746 563 752 597
rect 818 563 824 597
rect 824 563 852 597
rect 918 563 952 597
rect 1018 563 1052 597
rect 1118 563 1152 597
rect 1218 563 1246 597
rect 1246 563 1252 597
rect 1318 563 1324 597
rect 1324 563 1352 597
rect 1418 563 1452 597
rect 1518 563 1552 597
rect 1618 563 1652 597
rect 1718 563 1752 597
rect 1818 563 1852 597
rect 1918 563 1952 597
rect 2018 563 2052 597
rect 2118 563 2146 597
rect 2146 563 2152 597
rect 2218 563 2224 597
rect 2224 563 2252 597
rect 2318 563 2352 597
rect 2418 563 2452 597
rect 2518 563 2552 597
rect 2618 563 2652 597
rect 2718 563 2746 597
rect 2746 563 2752 597
rect 2818 563 2824 597
rect 2824 563 2852 597
rect 2918 563 2952 597
rect 3018 563 3052 597
rect 3118 563 3152 597
rect 3218 563 3252 597
rect 3318 563 3352 597
rect 3418 563 3452 597
rect 3518 563 3552 597
rect 3618 563 3652 597
rect 3718 563 3752 597
rect 3818 563 3852 597
rect 3918 563 3946 597
rect 3946 563 3952 597
rect 4018 563 4024 597
rect 4024 563 4052 597
rect 4118 563 4146 597
rect 4146 563 4152 597
rect 4218 563 4224 597
rect 4224 563 4252 597
rect 4318 563 4352 597
rect 4418 563 4452 597
rect 4518 563 4552 597
rect 4618 563 4652 597
rect 4718 563 4752 597
rect 4818 563 4846 597
rect 4846 563 4852 597
rect 4918 563 4924 597
rect 4924 563 4952 597
rect 5018 563 5046 597
rect 5046 563 5052 597
rect 5118 563 5124 597
rect 5124 563 5152 597
rect 5218 563 5246 597
rect 5246 563 5252 597
rect 5318 563 5324 597
rect 5324 563 5352 597
rect 5418 563 5452 597
rect 5518 563 5552 597
rect 5618 563 5652 597
rect 5718 563 5752 597
rect 5818 563 5852 597
rect 5918 563 5952 597
rect 6018 563 6052 597
rect 6118 563 6152 597
rect 6218 563 6252 597
rect 6318 563 6352 597
rect 6418 563 6452 597
rect 6518 563 6552 597
rect 6618 563 6652 597
rect 6718 563 6752 597
rect 6818 563 6852 597
rect 6918 563 6952 597
rect 7018 563 7052 597
rect 7118 563 7152 597
rect 7218 563 7252 597
rect 7318 563 7352 597
rect 7418 563 7452 597
rect 7518 563 7552 597
rect 7618 563 7652 597
rect 7718 563 7752 597
rect 7818 563 7852 597
rect 7918 563 7952 597
rect 8018 563 8052 597
rect 8118 563 8152 597
rect 8218 563 8252 597
rect 8318 563 8346 597
rect 8346 563 8352 597
rect 8418 563 8424 597
rect 8424 563 8452 597
rect 8518 563 8552 597
rect 8618 563 8652 597
rect 8718 563 8752 597
rect 8818 563 8852 597
rect 8918 563 8952 597
rect 9018 563 9052 597
rect 9118 563 9152 597
rect 9218 563 9252 597
rect 9318 563 9352 597
rect 9418 563 9452 597
rect 9518 563 9552 597
rect 9618 563 9652 597
rect 9718 563 9752 597
rect 9818 563 9852 597
rect 9918 563 9952 597
rect 10018 563 10052 597
rect 10118 563 10152 597
rect 10218 563 10246 597
rect 10246 563 10252 597
rect 10318 563 10324 597
rect 10324 563 10352 597
rect 10418 563 10446 597
rect 10446 563 10452 597
rect 10518 563 10524 597
rect 10524 563 10552 597
rect 10618 563 10652 597
rect 10718 563 10752 597
rect 10818 563 10852 597
rect 10918 563 10952 597
rect 11018 563 11052 597
rect 11118 563 11152 597
rect 11218 563 11246 597
rect 11246 563 11252 597
rect 11318 563 11324 597
rect 11324 563 11352 597
rect 11418 563 11452 597
rect 11518 563 11552 597
rect 11618 563 11652 597
rect 11718 563 11752 597
rect 11818 563 11852 597
rect 11918 563 11952 597
rect 12018 563 12052 597
rect 12118 563 12152 597
rect 12218 563 12252 597
rect 12318 563 12352 597
rect 12418 563 12452 597
rect 12518 563 12552 597
rect 12618 563 12652 597
rect 12718 563 12752 597
rect 12818 563 12846 597
rect 12846 563 12852 597
rect 12916 578 12924 612
rect 12924 578 12950 612
rect 13120 548 13146 582
rect 13146 548 13154 582
rect 18 423 52 457
rect 118 423 152 457
rect 218 423 252 457
rect 318 423 346 457
rect 346 423 352 457
rect 418 423 424 457
rect 424 423 452 457
rect 518 423 552 457
rect 618 423 652 457
rect 718 423 752 457
rect 818 423 852 457
rect 918 423 952 457
rect 1018 423 1052 457
rect 1118 423 1146 457
rect 1146 423 1152 457
rect 1218 423 1224 457
rect 1224 423 1252 457
rect 1318 423 1352 457
rect 1418 423 1452 457
rect 1518 423 1552 457
rect 1618 423 1652 457
rect 1718 423 1752 457
rect 1818 423 1846 457
rect 1846 423 1852 457
rect 1918 423 1924 457
rect 1924 423 1952 457
rect 2018 423 2052 457
rect 2118 423 2152 457
rect 2218 423 2252 457
rect 2318 423 2346 457
rect 2346 423 2352 457
rect 2418 423 2424 457
rect 2424 423 2452 457
rect 2518 423 2552 457
rect 2618 423 2646 457
rect 2646 423 2652 457
rect 2718 423 2724 457
rect 2724 423 2752 457
rect 2818 423 2852 457
rect 2918 423 2952 457
rect 3018 423 3052 457
rect 3118 423 3152 457
rect 3218 423 3252 457
rect 3318 423 3352 457
rect 3418 423 3452 457
rect 3518 423 3552 457
rect 3618 423 3652 457
rect 3718 423 3752 457
rect 3818 423 3852 457
rect 3918 423 3952 457
rect 4018 423 4052 457
rect 4118 423 4152 457
rect 4218 423 4252 457
rect 4318 423 4352 457
rect 4418 423 4446 457
rect 4446 423 4452 457
rect 4518 423 4524 457
rect 4524 423 4552 457
rect 4618 423 4652 457
rect 4718 423 4752 457
rect 4818 423 4852 457
rect 4918 423 4952 457
rect 5018 423 5052 457
rect 5118 423 5146 457
rect 5146 423 5152 457
rect 5218 423 5224 457
rect 5224 423 5252 457
rect 5318 423 5346 457
rect 5346 423 5352 457
rect 5418 423 5424 457
rect 5424 423 5452 457
rect 5518 423 5552 457
rect 5618 423 5652 457
rect 5718 423 5752 457
rect 5818 423 5852 457
rect 5918 423 5952 457
rect 6018 423 6052 457
rect 6118 423 6146 457
rect 6146 423 6152 457
rect 6218 423 6224 457
rect 6224 423 6252 457
rect 6318 423 6352 457
rect 6418 423 6446 457
rect 6446 423 6452 457
rect 6518 423 6524 457
rect 6524 423 6552 457
rect 6618 423 6652 457
rect 6718 423 6752 457
rect 6818 423 6852 457
rect 6918 423 6952 457
rect 7018 423 7052 457
rect 7118 423 7146 457
rect 7146 423 7152 457
rect 7218 423 7224 457
rect 7224 423 7252 457
rect 7318 423 7346 457
rect 7346 423 7352 457
rect 7418 423 7424 457
rect 7424 423 7452 457
rect 7518 423 7546 457
rect 7546 423 7552 457
rect 7618 423 7624 457
rect 7624 423 7652 457
rect 7718 423 7752 457
rect 7818 423 7852 457
rect 7918 423 7952 457
rect 8018 423 8052 457
rect 8118 423 8152 457
rect 8218 423 8252 457
rect 8318 423 8346 457
rect 8346 423 8352 457
rect 8418 423 8424 457
rect 8424 423 8452 457
rect 8518 423 8552 457
rect 8618 423 8652 457
rect 8718 423 8752 457
rect 8818 423 8852 457
rect 8918 423 8952 457
rect 9018 423 9052 457
rect 9118 423 9152 457
rect 9218 423 9252 457
rect 9318 423 9352 457
rect 9418 423 9452 457
rect 9518 423 9552 457
rect 9618 423 9652 457
rect 9718 423 9752 457
rect 9818 423 9852 457
rect 9918 423 9946 457
rect 9946 423 9952 457
rect 10018 423 10024 457
rect 10024 423 10052 457
rect 10118 423 10152 457
rect 10218 423 10246 457
rect 10246 423 10252 457
rect 10318 423 10324 457
rect 10324 423 10352 457
rect 10418 423 10452 457
rect 10518 423 10552 457
rect 10618 423 10652 457
rect 10718 423 10752 457
rect 10818 423 10846 457
rect 10846 423 10852 457
rect 10918 423 10924 457
rect 10924 423 10952 457
rect 11018 423 11052 457
rect 11118 423 11146 457
rect 11146 423 11152 457
rect 11218 423 11224 457
rect 11224 423 11252 457
rect 11318 423 11346 457
rect 11346 423 11352 457
rect 11418 423 11424 457
rect 11424 423 11452 457
rect 11518 423 11552 457
rect 11618 423 11652 457
rect 11718 423 11752 457
rect 11818 423 11852 457
rect 11918 423 11952 457
rect 12018 423 12052 457
rect 12118 423 12152 457
rect 12218 423 12252 457
rect 12318 423 12346 457
rect 12346 423 12352 457
rect 12418 423 12424 457
rect 12424 423 12452 457
rect 12518 423 12552 457
rect 12618 423 12652 457
rect 12718 423 12752 457
rect 12818 423 12846 457
rect 12846 423 12852 457
rect 12916 438 12924 472
rect 12924 438 12950 472
rect 13120 408 13146 442
rect 13146 408 13154 442
rect 18 283 52 317
rect 118 283 152 317
rect 218 283 252 317
rect 318 283 352 317
rect 418 283 452 317
rect 518 283 552 317
rect 618 283 652 317
rect 718 283 752 317
rect 818 283 852 317
rect 918 283 952 317
rect 1018 283 1052 317
rect 1118 283 1152 317
rect 1218 283 1252 317
rect 1318 283 1352 317
rect 1418 283 1452 317
rect 1518 283 1552 317
rect 1618 283 1652 317
rect 1718 283 1746 317
rect 1746 283 1752 317
rect 1818 283 1824 317
rect 1824 283 1852 317
rect 1918 283 1952 317
rect 2018 283 2052 317
rect 2118 283 2152 317
rect 2218 283 2252 317
rect 2318 283 2352 317
rect 2418 283 2452 317
rect 2518 283 2552 317
rect 2618 283 2652 317
rect 2718 283 2752 317
rect 2818 283 2846 317
rect 2846 283 2852 317
rect 2918 283 2924 317
rect 2924 283 2952 317
rect 3018 283 3046 317
rect 3046 283 3052 317
rect 3118 283 3124 317
rect 3124 283 3152 317
rect 3218 283 3252 317
rect 3318 283 3352 317
rect 3418 283 3452 317
rect 3518 283 3552 317
rect 3618 283 3652 317
rect 3718 283 3752 317
rect 3818 283 3852 317
rect 3918 283 3952 317
rect 4018 283 4052 317
rect 4118 283 4152 317
rect 4218 283 4252 317
rect 4318 283 4352 317
rect 4418 283 4452 317
rect 4518 283 4546 317
rect 4546 283 4552 317
rect 4618 283 4624 317
rect 4624 283 4652 317
rect 4718 283 4752 317
rect 4818 283 4846 317
rect 4846 283 4852 317
rect 4918 283 4924 317
rect 4924 283 4952 317
rect 5018 283 5046 317
rect 5046 283 5052 317
rect 5118 283 5124 317
rect 5124 283 5152 317
rect 5218 283 5252 317
rect 5318 283 5352 317
rect 5418 283 5452 317
rect 5518 283 5552 317
rect 5618 283 5652 317
rect 5718 283 5752 317
rect 5818 283 5846 317
rect 5846 283 5852 317
rect 5918 283 5924 317
rect 5924 283 5952 317
rect 6018 283 6046 317
rect 6046 283 6052 317
rect 6118 283 6124 317
rect 6124 283 6152 317
rect 6218 283 6246 317
rect 6246 283 6252 317
rect 6318 283 6324 317
rect 6324 283 6352 317
rect 6418 283 6446 317
rect 6446 283 6452 317
rect 6518 283 6524 317
rect 6524 283 6552 317
rect 6618 283 6646 317
rect 6646 283 6652 317
rect 6718 283 6724 317
rect 6724 283 6752 317
rect 6818 283 6846 317
rect 6846 283 6852 317
rect 6918 283 6924 317
rect 6924 283 6952 317
rect 7018 283 7052 317
rect 7118 283 7152 317
rect 7218 283 7252 317
rect 7318 283 7352 317
rect 7418 283 7452 317
rect 7518 283 7552 317
rect 7618 283 7652 317
rect 7718 283 7752 317
rect 7818 283 7846 317
rect 7846 283 7852 317
rect 7918 283 7924 317
rect 7924 283 7952 317
rect 8018 283 8046 317
rect 8046 283 8052 317
rect 8118 283 8124 317
rect 8124 283 8152 317
rect 8218 283 8252 317
rect 8318 283 8352 317
rect 8418 283 8452 317
rect 8518 283 8552 317
rect 8618 283 8652 317
rect 8718 283 8746 317
rect 8746 283 8752 317
rect 8818 283 8824 317
rect 8824 283 8852 317
rect 8918 283 8952 317
rect 9018 283 9046 317
rect 9046 283 9052 317
rect 9118 283 9124 317
rect 9124 283 9152 317
rect 9218 283 9246 317
rect 9246 283 9252 317
rect 9318 283 9324 317
rect 9324 283 9352 317
rect 9418 283 9452 317
rect 9518 283 9552 317
rect 9618 283 9652 317
rect 9718 283 9752 317
rect 9818 283 9852 317
rect 9918 283 9952 317
rect 10018 283 10052 317
rect 10118 283 10146 317
rect 10146 283 10152 317
rect 10218 283 10224 317
rect 10224 283 10252 317
rect 10318 283 10352 317
rect 10418 283 10452 317
rect 10518 283 10552 317
rect 10618 283 10652 317
rect 10718 283 10752 317
rect 10818 283 10852 317
rect 10918 283 10952 317
rect 11018 283 11052 317
rect 11118 283 11152 317
rect 11218 283 11252 317
rect 11318 283 11352 317
rect 11418 283 11446 317
rect 11446 283 11452 317
rect 11518 283 11524 317
rect 11524 283 11552 317
rect 11618 283 11652 317
rect 11718 283 11752 317
rect 11818 283 11852 317
rect 11918 283 11952 317
rect 12018 283 12052 317
rect 12118 283 12152 317
rect 12218 283 12246 317
rect 12246 283 12252 317
rect 12318 283 12324 317
rect 12324 283 12352 317
rect 12418 283 12452 317
rect 12518 283 12552 317
rect 12618 283 12652 317
rect 12718 283 12752 317
rect 12818 283 12852 317
rect 12916 298 12924 332
rect 12924 298 12950 332
rect 13120 268 13146 302
rect 13146 268 13154 302
rect 18 143 24 177
rect 24 143 52 177
rect 118 143 152 177
rect 218 143 252 177
rect 318 143 352 177
rect 418 143 452 177
rect 518 143 552 177
rect 618 143 652 177
rect 718 143 752 177
rect 818 143 852 177
rect 918 143 952 177
rect 1018 143 1052 177
rect 1118 143 1152 177
rect 1218 143 1252 177
rect 1318 143 1352 177
rect 1418 143 1452 177
rect 1518 143 1552 177
rect 1618 143 1646 177
rect 1646 143 1652 177
rect 1718 143 1724 177
rect 1724 143 1752 177
rect 1818 143 1846 177
rect 1846 143 1852 177
rect 1918 143 1924 177
rect 1924 143 1952 177
rect 2018 143 2052 177
rect 2118 143 2152 177
rect 2218 143 2252 177
rect 2318 143 2352 177
rect 2418 143 2452 177
rect 2518 143 2552 177
rect 2618 143 2652 177
rect 2718 143 2752 177
rect 2818 143 2852 177
rect 2918 143 2952 177
rect 3018 143 3052 177
rect 3118 143 3152 177
rect 3218 143 3252 177
rect 3318 143 3352 177
rect 3418 143 3452 177
rect 3518 143 3552 177
rect 3618 143 3652 177
rect 3718 143 3752 177
rect 3818 143 3852 177
rect 3918 143 3952 177
rect 4018 143 4052 177
rect 4118 143 4152 177
rect 4218 143 4252 177
rect 4318 143 4352 177
rect 4418 143 4452 177
rect 4518 143 4552 177
rect 4618 143 4652 177
rect 4718 143 4752 177
rect 4818 143 4852 177
rect 4918 143 4952 177
rect 5018 143 5052 177
rect 5118 143 5152 177
rect 5218 143 5252 177
rect 5318 143 5352 177
rect 5418 143 5452 177
rect 5518 143 5552 177
rect 5618 143 5652 177
rect 5718 143 5752 177
rect 5818 143 5852 177
rect 5918 143 5952 177
rect 6018 143 6052 177
rect 6118 143 6152 177
rect 6218 143 6252 177
rect 6318 143 6352 177
rect 6418 143 6452 177
rect 6518 143 6552 177
rect 6618 143 6652 177
rect 6718 143 6752 177
rect 6818 143 6852 177
rect 6918 143 6952 177
rect 7018 143 7046 177
rect 7046 143 7052 177
rect 7118 143 7124 177
rect 7124 143 7152 177
rect 7218 143 7252 177
rect 7318 143 7352 177
rect 7418 143 7452 177
rect 7518 143 7552 177
rect 7618 143 7652 177
rect 7718 143 7752 177
rect 7818 143 7852 177
rect 7918 143 7952 177
rect 8018 143 8052 177
rect 8118 143 8152 177
rect 8218 143 8252 177
rect 8318 143 8352 177
rect 8418 143 8452 177
rect 8518 143 8552 177
rect 8618 143 8652 177
rect 8718 143 8752 177
rect 8818 143 8852 177
rect 8918 143 8952 177
rect 9018 143 9052 177
rect 9118 143 9152 177
rect 9218 143 9252 177
rect 9318 143 9352 177
rect 9418 143 9452 177
rect 9518 143 9552 177
rect 9618 143 9652 177
rect 9718 143 9752 177
rect 9818 143 9852 177
rect 9918 143 9952 177
rect 10018 143 10052 177
rect 10118 143 10152 177
rect 10218 143 10252 177
rect 10318 143 10352 177
rect 10418 143 10452 177
rect 10518 143 10552 177
rect 10618 143 10652 177
rect 10718 143 10752 177
rect 10818 143 10852 177
rect 10918 143 10952 177
rect 11018 143 11052 177
rect 11118 143 11152 177
rect 11218 143 11252 177
rect 11318 143 11352 177
rect 11418 143 11446 177
rect 11446 143 11452 177
rect 11518 143 11524 177
rect 11524 143 11552 177
rect 11618 143 11652 177
rect 11718 143 11752 177
rect 11818 143 11852 177
rect 11918 143 11952 177
rect 12018 143 12052 177
rect 12118 143 12152 177
rect 12218 143 12252 177
rect 12318 143 12352 177
rect 12418 143 12452 177
rect 12518 143 12552 177
rect 12618 143 12652 177
rect 12718 143 12752 177
rect 12818 143 12852 177
rect 12916 158 12924 192
rect 12924 158 12950 192
rect 13120 128 13146 162
rect 13146 128 13154 162
rect 18 20 52 54
rect 218 36 252 70
rect 418 20 452 54
rect 618 36 652 70
rect 818 20 852 54
rect 1018 36 1052 70
rect 1218 20 1252 54
rect 1418 36 1452 70
rect 1618 20 1652 54
rect 1818 36 1852 70
rect 2018 20 2052 54
rect 2218 36 2252 70
rect 2418 20 2452 54
rect 2618 36 2652 70
rect 2818 20 2852 54
rect 3018 36 3052 70
rect 3218 20 3252 54
rect 3418 36 3452 70
rect 3618 20 3652 54
rect 3818 36 3852 70
rect 4018 20 4052 54
rect 4218 36 4252 70
rect 4418 20 4452 54
rect 4618 36 4652 70
rect 4818 20 4852 54
rect 5018 36 5052 70
rect 5218 20 5252 54
rect 5418 36 5452 70
rect 5618 20 5652 54
rect 5818 36 5852 70
rect 6018 20 6052 54
rect 6218 36 6252 70
rect 6418 20 6452 54
rect 6618 36 6652 70
rect 6818 20 6852 54
rect 7018 36 7052 70
rect 7218 20 7252 54
rect 7418 36 7452 70
rect 7618 20 7652 54
rect 7818 36 7852 70
rect 8018 20 8052 54
rect 8218 36 8252 70
rect 8418 20 8452 54
rect 8618 36 8652 70
rect 8818 20 8852 54
rect 9018 36 9052 70
rect 9218 20 9252 54
rect 9418 36 9452 70
rect 9618 20 9652 54
rect 9818 36 9852 70
rect 10018 20 10052 54
rect 10218 36 10252 70
rect 10418 20 10452 54
rect 10618 36 10652 70
rect 10818 20 10852 54
rect 11018 36 11052 70
rect 11218 20 11252 54
rect 11418 36 11452 70
rect 11618 20 11652 54
rect 11818 36 11852 70
rect 12018 20 12052 54
rect 12218 36 12252 70
rect 12418 20 12452 54
rect 12618 36 12652 70
rect 12916 17 12950 51
rect 13120 39 13154 73
rect 13278 34 13312 68
rect 13378 34 13412 68
rect 13478 34 13512 68
rect 13578 34 13612 68
rect -82 -94 -48 -60
rect 118 -94 152 -60
rect -82 -149 -48 -132
rect -82 -166 -48 -149
rect 18 -149 52 -133
rect 18 -167 52 -149
rect 318 -94 352 -60
rect 118 -149 152 -132
rect 118 -166 152 -149
rect 218 -149 252 -133
rect 218 -167 252 -149
rect 518 -94 552 -60
rect 318 -149 352 -132
rect 318 -166 352 -149
rect 418 -149 452 -133
rect 418 -167 452 -149
rect 718 -94 752 -60
rect 518 -149 552 -132
rect 518 -166 552 -149
rect 618 -149 652 -133
rect 618 -167 652 -149
rect 918 -94 952 -60
rect 718 -149 752 -132
rect 718 -166 752 -149
rect 818 -149 852 -133
rect 818 -167 852 -149
rect 1118 -94 1152 -60
rect 918 -149 952 -132
rect 918 -166 952 -149
rect 1018 -149 1052 -133
rect 1018 -167 1052 -149
rect 1318 -94 1352 -60
rect 1118 -149 1152 -132
rect 1118 -166 1152 -149
rect 1218 -149 1252 -133
rect 1218 -167 1252 -149
rect 1518 -94 1552 -60
rect 1318 -149 1352 -132
rect 1318 -166 1352 -149
rect 1418 -149 1452 -133
rect 1418 -167 1452 -149
rect 1718 -94 1752 -60
rect 1518 -149 1552 -132
rect 1518 -166 1552 -149
rect 1618 -149 1652 -133
rect 1618 -167 1652 -149
rect 1918 -94 1952 -60
rect 1718 -149 1752 -132
rect 1718 -166 1752 -149
rect 1818 -149 1852 -133
rect 1818 -167 1852 -149
rect 2118 -94 2152 -60
rect 1918 -149 1952 -132
rect 1918 -166 1952 -149
rect 2018 -149 2052 -133
rect 2018 -167 2052 -149
rect 2318 -94 2352 -60
rect 2118 -149 2152 -132
rect 2118 -166 2152 -149
rect 2218 -149 2252 -133
rect 2218 -167 2252 -149
rect 2518 -94 2552 -60
rect 2318 -149 2352 -132
rect 2318 -166 2352 -149
rect 2418 -149 2452 -133
rect 2418 -167 2452 -149
rect 2718 -94 2752 -60
rect 2518 -149 2552 -132
rect 2518 -166 2552 -149
rect 2618 -149 2652 -133
rect 2618 -167 2652 -149
rect 2918 -94 2952 -60
rect 2718 -149 2752 -132
rect 2718 -166 2752 -149
rect 2818 -149 2852 -133
rect 2818 -167 2852 -149
rect 3118 -94 3152 -60
rect 2918 -149 2952 -132
rect 2918 -166 2952 -149
rect 3018 -149 3052 -133
rect 3018 -167 3052 -149
rect 3318 -94 3352 -60
rect 3118 -149 3152 -132
rect 3118 -166 3152 -149
rect 3218 -149 3252 -133
rect 3218 -167 3252 -149
rect 3518 -94 3552 -60
rect 3318 -149 3352 -132
rect 3318 -166 3352 -149
rect 3418 -149 3452 -133
rect 3418 -167 3452 -149
rect 3718 -94 3752 -60
rect 3518 -149 3552 -132
rect 3518 -166 3552 -149
rect 3618 -149 3652 -133
rect 3618 -167 3652 -149
rect 3918 -94 3952 -60
rect 3718 -149 3752 -132
rect 3718 -166 3752 -149
rect 3818 -149 3852 -133
rect 3818 -167 3852 -149
rect 4118 -94 4152 -60
rect 3918 -149 3952 -132
rect 3918 -166 3952 -149
rect 4018 -149 4052 -133
rect 4018 -167 4052 -149
rect 4318 -94 4352 -60
rect 4118 -149 4152 -132
rect 4118 -166 4152 -149
rect 4218 -149 4252 -133
rect 4218 -167 4252 -149
rect 4518 -94 4552 -60
rect 4318 -149 4352 -132
rect 4318 -166 4352 -149
rect 4418 -149 4452 -133
rect 4418 -167 4452 -149
rect 4718 -94 4752 -60
rect 4518 -149 4552 -132
rect 4518 -166 4552 -149
rect 4618 -149 4652 -133
rect 4618 -167 4652 -149
rect 4918 -94 4952 -60
rect 4718 -149 4752 -132
rect 4718 -166 4752 -149
rect 4818 -149 4852 -133
rect 4818 -167 4852 -149
rect 5118 -94 5152 -60
rect 4918 -149 4952 -132
rect 4918 -166 4952 -149
rect 5018 -149 5052 -133
rect 5018 -167 5052 -149
rect 5318 -94 5352 -60
rect 5118 -149 5152 -132
rect 5118 -166 5152 -149
rect 5218 -149 5252 -133
rect 5218 -167 5252 -149
rect 5518 -94 5552 -60
rect 5318 -149 5352 -132
rect 5318 -166 5352 -149
rect 5418 -149 5452 -133
rect 5418 -167 5452 -149
rect 5718 -94 5752 -60
rect 5518 -149 5552 -132
rect 5518 -166 5552 -149
rect 5618 -149 5652 -133
rect 5618 -167 5652 -149
rect 5918 -94 5952 -60
rect 5718 -149 5752 -132
rect 5718 -166 5752 -149
rect 5818 -149 5852 -133
rect 5818 -167 5852 -149
rect 6118 -94 6152 -60
rect 5918 -149 5952 -132
rect 5918 -166 5952 -149
rect 6018 -149 6052 -133
rect 6018 -167 6052 -149
rect 6318 -94 6352 -60
rect 6118 -149 6152 -132
rect 6118 -166 6152 -149
rect 6218 -149 6252 -133
rect 6218 -167 6252 -149
rect 6518 -94 6552 -60
rect 6318 -149 6352 -132
rect 6318 -166 6352 -149
rect 6418 -149 6452 -133
rect 6418 -167 6452 -149
rect 6718 -94 6752 -60
rect 6518 -149 6552 -132
rect 6518 -166 6552 -149
rect 6618 -149 6652 -133
rect 6618 -167 6652 -149
rect 6918 -94 6952 -60
rect 6718 -149 6752 -132
rect 6718 -166 6752 -149
rect 6818 -149 6852 -133
rect 6818 -167 6852 -149
rect 7118 -94 7152 -60
rect 6918 -149 6952 -132
rect 6918 -166 6952 -149
rect 7018 -149 7052 -133
rect 7018 -167 7052 -149
rect 7318 -94 7352 -60
rect 7118 -149 7152 -132
rect 7118 -166 7152 -149
rect 7218 -149 7252 -133
rect 7218 -167 7252 -149
rect 7518 -94 7552 -60
rect 7318 -149 7352 -132
rect 7318 -166 7352 -149
rect 7418 -149 7452 -133
rect 7418 -167 7452 -149
rect 7718 -94 7752 -60
rect 7518 -149 7552 -132
rect 7518 -166 7552 -149
rect 7618 -149 7652 -133
rect 7618 -167 7652 -149
rect 7918 -94 7952 -60
rect 7718 -149 7752 -132
rect 7718 -166 7752 -149
rect 7818 -149 7852 -133
rect 7818 -167 7852 -149
rect 8118 -94 8152 -60
rect 7918 -149 7952 -132
rect 7918 -166 7952 -149
rect 8018 -149 8052 -133
rect 8018 -167 8052 -149
rect 8318 -94 8352 -60
rect 8118 -149 8152 -132
rect 8118 -166 8152 -149
rect 8218 -149 8252 -133
rect 8218 -167 8252 -149
rect 8518 -94 8552 -60
rect 8318 -149 8352 -132
rect 8318 -166 8352 -149
rect 8418 -149 8452 -133
rect 8418 -167 8452 -149
rect 8718 -94 8752 -60
rect 8518 -149 8552 -132
rect 8518 -166 8552 -149
rect 8618 -149 8652 -133
rect 8618 -167 8652 -149
rect 8918 -94 8952 -60
rect 8718 -149 8752 -132
rect 8718 -166 8752 -149
rect 8818 -149 8852 -133
rect 8818 -167 8852 -149
rect 9118 -94 9152 -60
rect 8918 -149 8952 -132
rect 8918 -166 8952 -149
rect 9018 -149 9052 -133
rect 9018 -167 9052 -149
rect 9318 -94 9352 -60
rect 9118 -149 9152 -132
rect 9118 -166 9152 -149
rect 9218 -149 9252 -133
rect 9218 -167 9252 -149
rect 9518 -94 9552 -60
rect 9318 -149 9352 -132
rect 9318 -166 9352 -149
rect 9418 -149 9452 -133
rect 9418 -167 9452 -149
rect 9718 -94 9752 -60
rect 9518 -149 9552 -132
rect 9518 -166 9552 -149
rect 9618 -149 9652 -133
rect 9618 -167 9652 -149
rect 9918 -94 9952 -60
rect 9718 -149 9752 -132
rect 9718 -166 9752 -149
rect 9818 -149 9852 -133
rect 9818 -167 9852 -149
rect 10118 -94 10152 -60
rect 9918 -149 9952 -132
rect 9918 -166 9952 -149
rect 10018 -149 10052 -133
rect 10018 -167 10052 -149
rect 10318 -94 10352 -60
rect 10118 -149 10152 -132
rect 10118 -166 10152 -149
rect 10218 -149 10252 -133
rect 10218 -167 10252 -149
rect 10518 -94 10552 -60
rect 10318 -149 10352 -132
rect 10318 -166 10352 -149
rect 10418 -149 10452 -133
rect 10418 -167 10452 -149
rect 10718 -94 10752 -60
rect 10518 -149 10552 -132
rect 10518 -166 10552 -149
rect 10618 -149 10652 -133
rect 10618 -167 10652 -149
rect 10918 -94 10952 -60
rect 10718 -149 10752 -132
rect 10718 -166 10752 -149
rect 10818 -149 10852 -133
rect 10818 -167 10852 -149
rect 11118 -94 11152 -60
rect 10918 -149 10952 -132
rect 10918 -166 10952 -149
rect 11018 -149 11052 -133
rect 11018 -167 11052 -149
rect 11318 -94 11352 -60
rect 11118 -149 11152 -132
rect 11118 -166 11152 -149
rect 11218 -149 11252 -133
rect 11218 -167 11252 -149
rect 11518 -94 11552 -60
rect 11318 -149 11352 -132
rect 11318 -166 11352 -149
rect 11418 -149 11452 -133
rect 11418 -167 11452 -149
rect 11718 -94 11752 -60
rect 11518 -149 11552 -132
rect 11518 -166 11552 -149
rect 11618 -149 11652 -133
rect 11618 -167 11652 -149
rect 11918 -94 11952 -60
rect 11718 -149 11752 -132
rect 11718 -166 11752 -149
rect 11818 -149 11852 -133
rect 11818 -167 11852 -149
rect 12118 -94 12152 -60
rect 11918 -149 11952 -132
rect 11918 -166 11952 -149
rect 12018 -149 12052 -133
rect 12018 -167 12052 -149
rect 12318 -94 12352 -60
rect 12118 -149 12152 -132
rect 12118 -166 12152 -149
rect 12218 -149 12252 -133
rect 12218 -167 12252 -149
rect 12518 -94 12552 -60
rect 12318 -149 12352 -132
rect 12318 -166 12352 -149
rect 12418 -149 12452 -133
rect 12418 -167 12452 -149
rect 12718 -94 12752 -60
rect 12518 -149 12552 -132
rect 12518 -166 12552 -149
rect 12618 -149 12652 -133
rect 12618 -167 12652 -149
rect 12718 -149 12752 -132
rect 12718 -166 12752 -149
rect 14558 -242 14562 -208
rect 14562 -242 14592 -208
rect 14630 -242 14664 -208
rect 14842 -242 14847 -208
rect 14847 -242 14876 -208
rect 14914 -242 14915 -208
rect 14915 -242 14948 -208
rect 14986 -242 15017 -208
rect 15017 -242 15020 -208
rect 15058 -242 15085 -208
rect 15085 -242 15092 -208
rect 15249 -242 15257 -208
rect 15257 -242 15283 -208
rect 15321 -242 15325 -208
rect 15325 -242 15355 -208
rect 15393 -242 15427 -208
rect 15465 -242 15495 -208
rect 15495 -242 15499 -208
rect 15677 -242 15678 -208
rect 15678 -242 15711 -208
rect 15749 -242 15780 -208
rect 15780 -242 15783 -208
rect -66 -282 -32 -248
rect 134 -282 168 -248
rect 334 -282 368 -248
rect 534 -282 568 -248
rect 734 -282 768 -248
rect 934 -282 968 -248
rect 1134 -282 1168 -248
rect 1334 -282 1368 -248
rect 1534 -282 1568 -248
rect 1734 -282 1768 -248
rect 1934 -282 1968 -248
rect 2134 -282 2168 -248
rect 2334 -282 2368 -248
rect 2534 -282 2568 -248
rect 2734 -282 2768 -248
rect 2934 -282 2968 -248
rect 3134 -282 3168 -248
rect 3334 -282 3368 -248
rect 3534 -282 3568 -248
rect 3734 -282 3768 -248
rect 3934 -282 3968 -248
rect 4134 -282 4168 -248
rect 4334 -282 4368 -248
rect 4534 -282 4568 -248
rect 4734 -282 4768 -248
rect 4934 -282 4968 -248
rect 5134 -282 5168 -248
rect 5334 -282 5368 -248
rect 5534 -282 5568 -248
rect 5734 -282 5768 -248
rect 5934 -282 5968 -248
rect 6134 -282 6168 -248
rect 6334 -282 6368 -248
rect 6534 -282 6568 -248
rect 6734 -282 6768 -248
rect 6934 -282 6968 -248
rect 7134 -282 7168 -248
rect 7334 -282 7368 -248
rect 7534 -282 7568 -248
rect 7734 -282 7768 -248
rect 7934 -282 7968 -248
rect 8134 -282 8168 -248
rect 8334 -282 8368 -248
rect 8534 -282 8568 -248
rect 8734 -282 8768 -248
rect 8934 -282 8968 -248
rect 9134 -282 9168 -248
rect 9334 -282 9368 -248
rect 9534 -282 9568 -248
rect 9734 -282 9768 -248
rect 9934 -282 9968 -248
rect 10134 -282 10168 -248
rect 10334 -282 10368 -248
rect 10534 -282 10568 -248
rect 10734 -282 10768 -248
rect 10934 -282 10968 -248
rect 11134 -282 11168 -248
rect 11334 -282 11368 -248
rect 11534 -282 11568 -248
rect 11734 -282 11768 -248
rect 11934 -282 11968 -248
rect 12134 -282 12168 -248
rect 12334 -282 12368 -248
rect 12534 -282 12568 -248
rect -82 -397 -48 -363
rect -82 -465 -48 -435
rect -82 -469 -48 -465
rect 18 -397 52 -363
rect 18 -465 52 -435
rect 18 -469 52 -465
rect 118 -397 152 -363
rect 118 -465 152 -435
rect 118 -469 152 -465
rect -118 -595 -84 -561
rect -46 -595 -12 -561
rect 44 -664 78 -630
rect 218 -397 252 -363
rect 218 -465 252 -435
rect 218 -469 252 -465
rect 318 -397 352 -363
rect 318 -465 352 -435
rect 318 -469 352 -465
rect 418 -397 452 -363
rect 418 -465 452 -435
rect 418 -469 452 -465
rect 518 -397 552 -363
rect 518 -465 552 -435
rect 518 -469 552 -465
rect 282 -595 316 -561
rect 354 -595 388 -561
rect 192 -664 226 -630
rect 444 -664 478 -630
rect 618 -397 652 -363
rect 618 -465 652 -435
rect 618 -469 652 -465
rect 718 -397 752 -363
rect 718 -465 752 -435
rect 718 -469 752 -465
rect 818 -397 852 -363
rect 818 -465 852 -435
rect 818 -469 852 -465
rect 918 -397 952 -363
rect 918 -465 952 -435
rect 918 -469 952 -465
rect 682 -595 716 -561
rect 754 -595 788 -561
rect 592 -664 626 -630
rect 844 -664 878 -630
rect 1018 -397 1052 -363
rect 1018 -465 1052 -435
rect 1018 -469 1052 -465
rect 1118 -397 1152 -363
rect 1118 -465 1152 -435
rect 1118 -469 1152 -465
rect 1218 -397 1252 -363
rect 1218 -465 1252 -435
rect 1218 -469 1252 -465
rect 1318 -397 1352 -363
rect 1318 -465 1352 -435
rect 1318 -469 1352 -465
rect 1082 -595 1116 -561
rect 1154 -595 1188 -561
rect 992 -664 1026 -630
rect 1244 -664 1278 -630
rect 1418 -397 1452 -363
rect 1418 -465 1452 -435
rect 1418 -469 1452 -465
rect 1518 -397 1552 -363
rect 1518 -465 1552 -435
rect 1518 -469 1552 -465
rect 1618 -397 1652 -363
rect 1618 -465 1652 -435
rect 1618 -469 1652 -465
rect 1718 -397 1752 -363
rect 1718 -465 1752 -435
rect 1718 -469 1752 -465
rect 1482 -595 1516 -561
rect 1554 -595 1588 -561
rect 1392 -664 1426 -630
rect 1644 -664 1678 -630
rect 1818 -397 1852 -363
rect 1818 -465 1852 -435
rect 1818 -469 1852 -465
rect 1918 -397 1952 -363
rect 1918 -465 1952 -435
rect 1918 -469 1952 -465
rect 2018 -397 2052 -363
rect 2018 -465 2052 -435
rect 2018 -469 2052 -465
rect 2118 -397 2152 -363
rect 2118 -465 2152 -435
rect 2118 -469 2152 -465
rect 1882 -595 1916 -561
rect 1954 -595 1988 -561
rect 1792 -664 1826 -630
rect 2044 -664 2078 -630
rect 2218 -397 2252 -363
rect 2218 -465 2252 -435
rect 2218 -469 2252 -465
rect 2318 -397 2352 -363
rect 2318 -465 2352 -435
rect 2318 -469 2352 -465
rect 2418 -397 2452 -363
rect 2418 -465 2452 -435
rect 2418 -469 2452 -465
rect 2518 -397 2552 -363
rect 2518 -465 2552 -435
rect 2518 -469 2552 -465
rect 2282 -595 2316 -561
rect 2354 -595 2388 -561
rect 2192 -664 2226 -630
rect 2444 -664 2478 -630
rect 2618 -397 2652 -363
rect 2618 -465 2652 -435
rect 2618 -469 2652 -465
rect 2718 -397 2752 -363
rect 2718 -465 2752 -435
rect 2718 -469 2752 -465
rect 2818 -397 2852 -363
rect 2818 -465 2852 -435
rect 2818 -469 2852 -465
rect 2918 -397 2952 -363
rect 2918 -465 2952 -435
rect 2918 -469 2952 -465
rect 2682 -595 2716 -561
rect 2754 -595 2788 -561
rect 2592 -664 2626 -630
rect 2844 -664 2878 -630
rect 3018 -397 3052 -363
rect 3018 -465 3052 -435
rect 3018 -469 3052 -465
rect 3118 -397 3152 -363
rect 3118 -465 3152 -435
rect 3118 -469 3152 -465
rect 3218 -397 3252 -363
rect 3218 -465 3252 -435
rect 3218 -469 3252 -465
rect 3318 -397 3352 -363
rect 3318 -465 3352 -435
rect 3318 -469 3352 -465
rect 3082 -595 3116 -561
rect 3154 -595 3188 -561
rect 2992 -664 3026 -630
rect 3244 -664 3278 -630
rect 3418 -397 3452 -363
rect 3418 -465 3452 -435
rect 3418 -469 3452 -465
rect 3518 -397 3552 -363
rect 3518 -465 3552 -435
rect 3518 -469 3552 -465
rect 3618 -397 3652 -363
rect 3618 -465 3652 -435
rect 3618 -469 3652 -465
rect 3718 -397 3752 -363
rect 3718 -465 3752 -435
rect 3718 -469 3752 -465
rect 3482 -595 3516 -561
rect 3554 -595 3588 -561
rect 3392 -664 3426 -630
rect 3644 -664 3678 -630
rect 3818 -397 3852 -363
rect 3818 -465 3852 -435
rect 3818 -469 3852 -465
rect 3918 -397 3952 -363
rect 3918 -465 3952 -435
rect 3918 -469 3952 -465
rect 4018 -397 4052 -363
rect 4018 -465 4052 -435
rect 4018 -469 4052 -465
rect 4118 -397 4152 -363
rect 4118 -465 4152 -435
rect 4118 -469 4152 -465
rect 3882 -595 3916 -561
rect 3954 -595 3988 -561
rect 3792 -664 3826 -630
rect 4044 -664 4078 -630
rect 4218 -397 4252 -363
rect 4218 -465 4252 -435
rect 4218 -469 4252 -465
rect 4318 -397 4352 -363
rect 4318 -465 4352 -435
rect 4318 -469 4352 -465
rect 4418 -397 4452 -363
rect 4418 -465 4452 -435
rect 4418 -469 4452 -465
rect 4518 -397 4552 -363
rect 4518 -465 4552 -435
rect 4518 -469 4552 -465
rect 4282 -595 4316 -561
rect 4354 -595 4388 -561
rect 4192 -664 4226 -630
rect 4444 -664 4478 -630
rect 4618 -397 4652 -363
rect 4618 -465 4652 -435
rect 4618 -469 4652 -465
rect 4718 -397 4752 -363
rect 4718 -465 4752 -435
rect 4718 -469 4752 -465
rect 4818 -397 4852 -363
rect 4818 -465 4852 -435
rect 4818 -469 4852 -465
rect 4918 -397 4952 -363
rect 4918 -465 4952 -435
rect 4918 -469 4952 -465
rect 4682 -595 4716 -561
rect 4754 -595 4788 -561
rect 4592 -664 4626 -630
rect 4844 -664 4878 -630
rect 5018 -397 5052 -363
rect 5018 -465 5052 -435
rect 5018 -469 5052 -465
rect 5118 -397 5152 -363
rect 5118 -465 5152 -435
rect 5118 -469 5152 -465
rect 5218 -397 5252 -363
rect 5218 -465 5252 -435
rect 5218 -469 5252 -465
rect 5318 -397 5352 -363
rect 5318 -465 5352 -435
rect 5318 -469 5352 -465
rect 5082 -595 5116 -561
rect 5154 -595 5188 -561
rect 4992 -664 5026 -630
rect 5244 -664 5278 -630
rect 5418 -397 5452 -363
rect 5418 -465 5452 -435
rect 5418 -469 5452 -465
rect 5518 -397 5552 -363
rect 5518 -465 5552 -435
rect 5518 -469 5552 -465
rect 5618 -397 5652 -363
rect 5618 -465 5652 -435
rect 5618 -469 5652 -465
rect 5718 -397 5752 -363
rect 5718 -465 5752 -435
rect 5718 -469 5752 -465
rect 5482 -595 5516 -561
rect 5554 -595 5588 -561
rect 5392 -664 5426 -630
rect 5644 -664 5678 -630
rect 5818 -397 5852 -363
rect 5818 -465 5852 -435
rect 5818 -469 5852 -465
rect 5918 -397 5952 -363
rect 5918 -465 5952 -435
rect 5918 -469 5952 -465
rect 6018 -397 6052 -363
rect 6018 -465 6052 -435
rect 6018 -469 6052 -465
rect 6118 -397 6152 -363
rect 6118 -465 6152 -435
rect 6118 -469 6152 -465
rect 5882 -595 5916 -561
rect 5954 -595 5988 -561
rect 5792 -664 5826 -630
rect 6044 -664 6078 -630
rect 6218 -397 6252 -363
rect 6218 -465 6252 -435
rect 6218 -469 6252 -465
rect 6318 -397 6352 -363
rect 6318 -465 6352 -435
rect 6318 -469 6352 -465
rect 6418 -397 6452 -363
rect 6418 -465 6452 -435
rect 6418 -469 6452 -465
rect 6518 -397 6552 -363
rect 6518 -465 6552 -435
rect 6518 -469 6552 -465
rect 6282 -595 6316 -561
rect 6354 -595 6388 -561
rect 6192 -664 6226 -630
rect 6444 -664 6478 -630
rect 6618 -397 6652 -363
rect 6618 -465 6652 -435
rect 6618 -469 6652 -465
rect 6718 -397 6752 -363
rect 6718 -465 6752 -435
rect 6718 -469 6752 -465
rect 6818 -397 6852 -363
rect 6818 -465 6852 -435
rect 6818 -469 6852 -465
rect 6918 -397 6952 -363
rect 6918 -465 6952 -435
rect 6918 -469 6952 -465
rect 6682 -595 6716 -561
rect 6754 -595 6788 -561
rect 6592 -664 6626 -630
rect 6844 -664 6878 -630
rect 7018 -397 7052 -363
rect 7018 -465 7052 -435
rect 7018 -469 7052 -465
rect 7118 -397 7152 -363
rect 7118 -465 7152 -435
rect 7118 -469 7152 -465
rect 7218 -397 7252 -363
rect 7218 -465 7252 -435
rect 7218 -469 7252 -465
rect 7318 -397 7352 -363
rect 7318 -465 7352 -435
rect 7318 -469 7352 -465
rect 7082 -595 7116 -561
rect 7154 -595 7188 -561
rect 6992 -664 7026 -630
rect 7244 -664 7278 -630
rect 7418 -397 7452 -363
rect 7418 -465 7452 -435
rect 7418 -469 7452 -465
rect 7518 -397 7552 -363
rect 7518 -465 7552 -435
rect 7518 -469 7552 -465
rect 7618 -397 7652 -363
rect 7618 -465 7652 -435
rect 7618 -469 7652 -465
rect 7718 -397 7752 -363
rect 7718 -465 7752 -435
rect 7718 -469 7752 -465
rect 7482 -595 7516 -561
rect 7554 -595 7588 -561
rect 7392 -664 7426 -630
rect 7644 -664 7678 -630
rect 7818 -397 7852 -363
rect 7818 -465 7852 -435
rect 7818 -469 7852 -465
rect 7918 -397 7952 -363
rect 7918 -465 7952 -435
rect 7918 -469 7952 -465
rect 8018 -397 8052 -363
rect 8018 -465 8052 -435
rect 8018 -469 8052 -465
rect 8118 -397 8152 -363
rect 8118 -465 8152 -435
rect 8118 -469 8152 -465
rect 7882 -595 7916 -561
rect 7954 -595 7988 -561
rect 7792 -664 7826 -630
rect 8044 -664 8078 -630
rect 8218 -397 8252 -363
rect 8218 -465 8252 -435
rect 8218 -469 8252 -465
rect 8318 -397 8352 -363
rect 8318 -465 8352 -435
rect 8318 -469 8352 -465
rect 8418 -397 8452 -363
rect 8418 -465 8452 -435
rect 8418 -469 8452 -465
rect 8518 -397 8552 -363
rect 8518 -465 8552 -435
rect 8518 -469 8552 -465
rect 8282 -595 8316 -561
rect 8354 -595 8388 -561
rect 8192 -664 8226 -630
rect 8444 -664 8478 -630
rect 8618 -397 8652 -363
rect 8618 -465 8652 -435
rect 8618 -469 8652 -465
rect 8718 -397 8752 -363
rect 8718 -465 8752 -435
rect 8718 -469 8752 -465
rect 8818 -397 8852 -363
rect 8818 -465 8852 -435
rect 8818 -469 8852 -465
rect 8918 -397 8952 -363
rect 8918 -465 8952 -435
rect 8918 -469 8952 -465
rect 8682 -595 8716 -561
rect 8754 -595 8788 -561
rect 8592 -664 8626 -630
rect 8844 -664 8878 -630
rect 9018 -397 9052 -363
rect 9018 -465 9052 -435
rect 9018 -469 9052 -465
rect 9118 -397 9152 -363
rect 9118 -465 9152 -435
rect 9118 -469 9152 -465
rect 9218 -397 9252 -363
rect 9218 -465 9252 -435
rect 9218 -469 9252 -465
rect 9318 -397 9352 -363
rect 9318 -465 9352 -435
rect 9318 -469 9352 -465
rect 9082 -595 9116 -561
rect 9154 -595 9188 -561
rect 8992 -664 9026 -630
rect 9244 -664 9278 -630
rect 9418 -397 9452 -363
rect 9418 -465 9452 -435
rect 9418 -469 9452 -465
rect 9518 -397 9552 -363
rect 9518 -465 9552 -435
rect 9518 -469 9552 -465
rect 9618 -397 9652 -363
rect 9618 -465 9652 -435
rect 9618 -469 9652 -465
rect 9718 -397 9752 -363
rect 9718 -465 9752 -435
rect 9718 -469 9752 -465
rect 9482 -595 9516 -561
rect 9554 -595 9588 -561
rect 9392 -664 9426 -630
rect 9644 -664 9678 -630
rect 9818 -397 9852 -363
rect 9818 -465 9852 -435
rect 9818 -469 9852 -465
rect 9918 -397 9952 -363
rect 9918 -465 9952 -435
rect 9918 -469 9952 -465
rect 10018 -397 10052 -363
rect 10018 -465 10052 -435
rect 10018 -469 10052 -465
rect 10118 -397 10152 -363
rect 10118 -465 10152 -435
rect 10118 -469 10152 -465
rect 9882 -595 9916 -561
rect 9954 -595 9988 -561
rect 9792 -664 9826 -630
rect 10044 -664 10078 -630
rect 10218 -397 10252 -363
rect 10218 -465 10252 -435
rect 10218 -469 10252 -465
rect 10318 -397 10352 -363
rect 10318 -465 10352 -435
rect 10318 -469 10352 -465
rect 10418 -397 10452 -363
rect 10418 -465 10452 -435
rect 10418 -469 10452 -465
rect 10518 -397 10552 -363
rect 10518 -465 10552 -435
rect 10518 -469 10552 -465
rect 10282 -595 10316 -561
rect 10354 -595 10388 -561
rect 10192 -664 10226 -630
rect 10444 -664 10478 -630
rect 10618 -397 10652 -363
rect 10618 -465 10652 -435
rect 10618 -469 10652 -465
rect 10718 -397 10752 -363
rect 10718 -465 10752 -435
rect 10718 -469 10752 -465
rect 10818 -397 10852 -363
rect 10818 -465 10852 -435
rect 10818 -469 10852 -465
rect 10918 -397 10952 -363
rect 10918 -465 10952 -435
rect 10918 -469 10952 -465
rect 10682 -595 10716 -561
rect 10754 -595 10788 -561
rect 10592 -664 10626 -630
rect 10844 -664 10878 -630
rect 11018 -397 11052 -363
rect 11018 -465 11052 -435
rect 11018 -469 11052 -465
rect 11118 -397 11152 -363
rect 11118 -465 11152 -435
rect 11118 -469 11152 -465
rect 11218 -397 11252 -363
rect 11218 -465 11252 -435
rect 11218 -469 11252 -465
rect 11318 -397 11352 -363
rect 11318 -465 11352 -435
rect 11318 -469 11352 -465
rect 11082 -595 11116 -561
rect 11154 -595 11188 -561
rect 10992 -664 11026 -630
rect 11244 -664 11278 -630
rect 11418 -397 11452 -363
rect 11418 -465 11452 -435
rect 11418 -469 11452 -465
rect 11518 -397 11552 -363
rect 11518 -465 11552 -435
rect 11518 -469 11552 -465
rect 11618 -397 11652 -363
rect 11618 -465 11652 -435
rect 11618 -469 11652 -465
rect 11718 -397 11752 -363
rect 11718 -465 11752 -435
rect 11718 -469 11752 -465
rect 11482 -595 11516 -561
rect 11554 -595 11588 -561
rect 11392 -664 11426 -630
rect 11644 -664 11678 -630
rect 11818 -397 11852 -363
rect 11818 -465 11852 -435
rect 11818 -469 11852 -465
rect 11918 -397 11952 -363
rect 11918 -465 11952 -435
rect 11918 -469 11952 -465
rect 12018 -397 12052 -363
rect 12018 -465 12052 -435
rect 12018 -469 12052 -465
rect 12118 -397 12152 -363
rect 12118 -465 12152 -435
rect 12118 -469 12152 -465
rect 11882 -595 11916 -561
rect 11954 -595 11988 -561
rect 11792 -664 11826 -630
rect 12044 -664 12078 -630
rect 12218 -397 12252 -363
rect 12218 -465 12252 -435
rect 12218 -469 12252 -465
rect 12318 -397 12352 -363
rect 12318 -465 12352 -435
rect 12318 -469 12352 -465
rect 12418 -397 12452 -363
rect 12418 -465 12452 -435
rect 12418 -469 12452 -465
rect 12518 -397 12552 -363
rect 12518 -465 12552 -435
rect 12518 -469 12552 -465
rect 12282 -595 12316 -561
rect 12354 -595 12388 -561
rect 12192 -664 12226 -630
rect 12444 -664 12478 -630
rect 12618 -397 12652 -363
rect 12618 -465 12652 -435
rect 12618 -469 12652 -465
rect 14560 -342 14562 -308
rect 14562 -342 14594 -308
rect 14632 -342 14664 -308
rect 14664 -342 14666 -308
rect 12718 -397 12752 -363
rect 14841 -342 14847 -308
rect 14847 -342 14875 -308
rect 14913 -342 14915 -308
rect 14915 -342 14947 -308
rect 14985 -342 15017 -308
rect 15017 -342 15019 -308
rect 15057 -342 15085 -308
rect 15085 -342 15091 -308
rect 15251 -342 15257 -308
rect 15257 -342 15285 -308
rect 15323 -342 15325 -308
rect 15325 -342 15357 -308
rect 15395 -342 15427 -308
rect 15427 -342 15429 -308
rect 15467 -342 15495 -308
rect 15495 -342 15501 -308
rect 15676 -342 15678 -308
rect 15678 -342 15710 -308
rect 15748 -342 15780 -308
rect 15780 -342 15782 -308
rect 12718 -465 12752 -435
rect 14558 -442 14562 -408
rect 14562 -442 14592 -408
rect 14630 -442 14664 -408
rect 14734 -442 14768 -408
rect 14842 -442 14847 -408
rect 14847 -442 14876 -408
rect 14914 -442 14915 -408
rect 14915 -442 14948 -408
rect 14986 -442 15017 -408
rect 15017 -442 15020 -408
rect 15058 -442 15085 -408
rect 15085 -442 15092 -408
rect 15249 -442 15257 -408
rect 15257 -442 15283 -408
rect 15321 -442 15325 -408
rect 15325 -442 15355 -408
rect 15393 -442 15427 -408
rect 15465 -442 15495 -408
rect 15495 -442 15499 -408
rect 15574 -442 15608 -408
rect 15677 -442 15678 -408
rect 15678 -442 15711 -408
rect 15749 -442 15780 -408
rect 15780 -442 15783 -408
rect 12718 -469 12752 -465
rect 14560 -542 14562 -508
rect 14562 -542 14594 -508
rect 14632 -542 14664 -508
rect 14664 -542 14666 -508
rect 14841 -542 14847 -508
rect 14847 -542 14875 -508
rect 14913 -542 14915 -508
rect 14915 -542 14947 -508
rect 14985 -542 15017 -508
rect 15017 -542 15019 -508
rect 15057 -542 15085 -508
rect 15085 -542 15091 -508
rect 15251 -542 15257 -508
rect 15257 -542 15285 -508
rect 15323 -542 15325 -508
rect 15325 -542 15357 -508
rect 15395 -542 15427 -508
rect 15427 -542 15429 -508
rect 15467 -542 15495 -508
rect 15495 -542 15501 -508
rect 12682 -595 12716 -561
rect 12754 -595 12788 -561
rect 15676 -542 15678 -508
rect 15678 -542 15710 -508
rect 15748 -542 15780 -508
rect 15780 -542 15782 -508
rect 12592 -664 12626 -630
rect 14558 -642 14562 -608
rect 14562 -642 14592 -608
rect 14630 -642 14664 -608
rect 14734 -642 14768 -608
rect 14842 -642 14847 -608
rect 14847 -642 14876 -608
rect 14914 -642 14915 -608
rect 14915 -642 14948 -608
rect 14986 -642 15017 -608
rect 15017 -642 15020 -608
rect 15058 -642 15085 -608
rect 15085 -642 15092 -608
rect 15249 -642 15257 -608
rect 15257 -642 15283 -608
rect 15321 -642 15325 -608
rect 15325 -642 15355 -608
rect 15393 -642 15427 -608
rect 15465 -642 15495 -608
rect 15495 -642 15499 -608
rect 15574 -642 15608 -608
rect 15677 -642 15678 -608
rect 15678 -642 15711 -608
rect 15749 -642 15780 -608
rect 15780 -642 15783 -608
rect 14560 -742 14562 -708
rect 14562 -742 14594 -708
rect 14632 -742 14664 -708
rect 14664 -742 14666 -708
rect 14841 -742 14847 -708
rect 14847 -742 14875 -708
rect 14913 -742 14915 -708
rect 14915 -742 14947 -708
rect 14985 -742 15017 -708
rect 15017 -742 15019 -708
rect 15057 -742 15085 -708
rect 15085 -742 15091 -708
rect 15251 -742 15257 -708
rect 15257 -742 15285 -708
rect 15323 -742 15325 -708
rect 15325 -742 15357 -708
rect 15395 -742 15427 -708
rect 15427 -742 15429 -708
rect 15467 -742 15495 -708
rect 15495 -742 15501 -708
rect 15676 -742 15678 -708
rect 15678 -742 15710 -708
rect 15748 -742 15780 -708
rect 15780 -742 15782 -708
rect -4 -858 30 -837
rect 68 -858 102 -837
rect -4 -871 -2 -858
rect -2 -871 30 -858
rect 68 -871 100 -858
rect 100 -871 102 -858
rect -82 -942 -48 -908
rect 168 -858 202 -837
rect 240 -858 274 -837
rect 168 -871 170 -858
rect 170 -871 202 -858
rect 240 -871 272 -858
rect 272 -871 274 -858
rect 396 -858 430 -837
rect 468 -858 502 -837
rect 396 -871 398 -858
rect 398 -871 430 -858
rect 468 -871 500 -858
rect 500 -871 502 -858
rect -82 -1042 -48 -1008
rect -82 -1142 -48 -1108
rect 568 -858 602 -837
rect 640 -858 674 -837
rect 568 -871 570 -858
rect 570 -871 602 -858
rect 640 -871 672 -858
rect 672 -871 674 -858
rect 796 -858 830 -837
rect 868 -858 902 -837
rect 796 -871 798 -858
rect 798 -871 830 -858
rect 868 -871 900 -858
rect 900 -871 902 -858
rect 718 -942 752 -908
rect 968 -858 1002 -837
rect 1040 -858 1074 -837
rect 968 -871 970 -858
rect 970 -871 1002 -858
rect 1040 -871 1072 -858
rect 1072 -871 1074 -858
rect 1196 -858 1230 -837
rect 1268 -858 1302 -837
rect 1196 -871 1198 -858
rect 1198 -871 1230 -858
rect 1268 -871 1300 -858
rect 1300 -871 1302 -858
rect 718 -1042 752 -1008
rect 718 -1142 752 -1108
rect -82 -1242 -48 -1208
rect -82 -1342 -48 -1308
rect 1368 -858 1402 -837
rect 1440 -858 1474 -837
rect 1368 -871 1370 -858
rect 1370 -871 1402 -858
rect 1440 -871 1472 -858
rect 1472 -871 1474 -858
rect 1596 -858 1630 -837
rect 1668 -858 1702 -837
rect 1596 -871 1598 -858
rect 1598 -871 1630 -858
rect 1668 -871 1700 -858
rect 1700 -871 1702 -858
rect 1518 -942 1552 -908
rect 1768 -858 1802 -837
rect 1840 -858 1874 -837
rect 1768 -871 1770 -858
rect 1770 -871 1802 -858
rect 1840 -871 1872 -858
rect 1872 -871 1874 -858
rect 1996 -858 2030 -837
rect 2068 -858 2102 -837
rect 1996 -871 1998 -858
rect 1998 -871 2030 -858
rect 2068 -871 2100 -858
rect 2100 -871 2102 -858
rect 1518 -1042 1552 -1008
rect 1518 -1142 1552 -1108
rect 718 -1242 752 -1208
rect 2168 -858 2202 -837
rect 2240 -858 2274 -837
rect 2168 -871 2170 -858
rect 2170 -871 2202 -858
rect 2240 -871 2272 -858
rect 2272 -871 2274 -858
rect 2396 -858 2430 -837
rect 2468 -858 2502 -837
rect 2396 -871 2398 -858
rect 2398 -871 2430 -858
rect 2468 -871 2500 -858
rect 2500 -871 2502 -858
rect 2318 -942 2352 -908
rect 2568 -858 2602 -837
rect 2640 -858 2674 -837
rect 2568 -871 2570 -858
rect 2570 -871 2602 -858
rect 2640 -871 2672 -858
rect 2672 -871 2674 -858
rect 2796 -858 2830 -837
rect 2868 -858 2902 -837
rect 2796 -871 2798 -858
rect 2798 -871 2830 -858
rect 2868 -871 2900 -858
rect 2900 -871 2902 -858
rect 2318 -1042 2352 -1008
rect 2318 -1142 2352 -1108
rect 1518 -1242 1552 -1208
rect 718 -1342 752 -1308
rect 1518 -1342 1552 -1308
rect -82 -1442 -48 -1408
rect 718 -1442 752 -1408
rect -82 -1542 -48 -1508
rect 718 -1542 752 -1508
rect 2968 -858 3002 -837
rect 3040 -858 3074 -837
rect 2968 -871 2970 -858
rect 2970 -871 3002 -858
rect 3040 -871 3072 -858
rect 3072 -871 3074 -858
rect 3196 -858 3230 -837
rect 3268 -858 3302 -837
rect 3196 -871 3198 -858
rect 3198 -871 3230 -858
rect 3268 -871 3300 -858
rect 3300 -871 3302 -858
rect 3118 -942 3152 -908
rect 3368 -858 3402 -837
rect 3440 -858 3474 -837
rect 3368 -871 3370 -858
rect 3370 -871 3402 -858
rect 3440 -871 3472 -858
rect 3472 -871 3474 -858
rect 3596 -858 3630 -837
rect 3668 -858 3702 -837
rect 3596 -871 3598 -858
rect 3598 -871 3630 -858
rect 3668 -871 3700 -858
rect 3700 -871 3702 -858
rect 3118 -1042 3152 -1008
rect 3118 -1142 3152 -1108
rect 2318 -1242 2352 -1208
rect 3768 -858 3802 -837
rect 3840 -858 3874 -837
rect 3768 -871 3770 -858
rect 3770 -871 3802 -858
rect 3840 -871 3872 -858
rect 3872 -871 3874 -858
rect 3996 -858 4030 -837
rect 4068 -858 4102 -837
rect 3996 -871 3998 -858
rect 3998 -871 4030 -858
rect 4068 -871 4100 -858
rect 4100 -871 4102 -858
rect 3918 -942 3952 -908
rect 4168 -858 4202 -837
rect 4240 -858 4274 -837
rect 4168 -871 4170 -858
rect 4170 -871 4202 -858
rect 4240 -871 4272 -858
rect 4272 -871 4274 -858
rect 4396 -858 4430 -837
rect 4468 -858 4502 -837
rect 4396 -871 4398 -858
rect 4398 -871 4430 -858
rect 4468 -871 4500 -858
rect 4500 -871 4502 -858
rect 3918 -1042 3952 -1008
rect 3918 -1142 3952 -1108
rect 3118 -1242 3152 -1208
rect 2318 -1342 2352 -1308
rect 3118 -1342 3152 -1308
rect 1518 -1442 1552 -1408
rect 2318 -1442 2352 -1408
rect 4568 -858 4602 -837
rect 4640 -858 4674 -837
rect 4568 -871 4570 -858
rect 4570 -871 4602 -858
rect 4640 -871 4672 -858
rect 4672 -871 4674 -858
rect 4796 -858 4830 -837
rect 4868 -858 4902 -837
rect 4796 -871 4798 -858
rect 4798 -871 4830 -858
rect 4868 -871 4900 -858
rect 4900 -871 4902 -858
rect 4718 -942 4752 -908
rect 4968 -858 5002 -837
rect 5040 -858 5074 -837
rect 4968 -871 4970 -858
rect 4970 -871 5002 -858
rect 5040 -871 5072 -858
rect 5072 -871 5074 -858
rect 5196 -858 5230 -837
rect 5268 -858 5302 -837
rect 5196 -871 5198 -858
rect 5198 -871 5230 -858
rect 5268 -871 5300 -858
rect 5300 -871 5302 -858
rect 4718 -1042 4752 -1008
rect 4718 -1142 4752 -1108
rect 3918 -1242 3952 -1208
rect 5368 -858 5402 -837
rect 5440 -858 5474 -837
rect 5368 -871 5370 -858
rect 5370 -871 5402 -858
rect 5440 -871 5472 -858
rect 5472 -871 5474 -858
rect 5596 -858 5630 -837
rect 5668 -858 5702 -837
rect 5596 -871 5598 -858
rect 5598 -871 5630 -858
rect 5668 -871 5700 -858
rect 5700 -871 5702 -858
rect 5518 -942 5552 -908
rect 5768 -858 5802 -837
rect 5840 -858 5874 -837
rect 5768 -871 5770 -858
rect 5770 -871 5802 -858
rect 5840 -871 5872 -858
rect 5872 -871 5874 -858
rect 5996 -858 6030 -837
rect 6068 -858 6102 -837
rect 5996 -871 5998 -858
rect 5998 -871 6030 -858
rect 6068 -871 6100 -858
rect 6100 -871 6102 -858
rect 5518 -1042 5552 -1008
rect 5518 -1142 5552 -1108
rect 4718 -1242 4752 -1208
rect 3918 -1342 3952 -1308
rect 4718 -1342 4752 -1308
rect 3118 -1442 3152 -1408
rect 3918 -1442 3952 -1408
rect 1518 -1542 1552 -1508
rect 2318 -1542 2352 -1508
rect 3118 -1542 3152 -1508
rect -82 -1642 -48 -1608
rect 718 -1642 752 -1608
rect 1518 -1642 1552 -1608
rect -82 -1742 -48 -1708
rect 718 -1742 752 -1708
rect 1518 -1742 1552 -1708
rect 2318 -1642 2352 -1608
rect 2318 -1742 2352 -1708
rect 3918 -1542 3952 -1508
rect 6168 -858 6202 -837
rect 6240 -858 6274 -837
rect 6168 -871 6170 -858
rect 6170 -871 6202 -858
rect 6240 -871 6272 -858
rect 6272 -871 6274 -858
rect 6396 -858 6430 -837
rect 6468 -858 6502 -837
rect 6396 -871 6398 -858
rect 6398 -871 6430 -858
rect 6468 -871 6500 -858
rect 6500 -871 6502 -858
rect 6318 -942 6352 -908
rect 6568 -858 6602 -837
rect 6640 -858 6674 -837
rect 6568 -871 6570 -858
rect 6570 -871 6602 -858
rect 6640 -871 6672 -858
rect 6672 -871 6674 -858
rect 6796 -858 6830 -837
rect 6868 -858 6902 -837
rect 6796 -871 6798 -858
rect 6798 -871 6830 -858
rect 6868 -871 6900 -858
rect 6900 -871 6902 -858
rect 6318 -1042 6352 -1008
rect 6318 -1142 6352 -1108
rect 5518 -1242 5552 -1208
rect 6968 -858 7002 -837
rect 7040 -858 7074 -837
rect 6968 -871 6970 -858
rect 6970 -871 7002 -858
rect 7040 -871 7072 -858
rect 7072 -871 7074 -858
rect 7196 -858 7230 -837
rect 7268 -858 7302 -837
rect 7196 -871 7198 -858
rect 7198 -871 7230 -858
rect 7268 -871 7300 -858
rect 7300 -871 7302 -858
rect 7118 -942 7152 -908
rect 7368 -858 7402 -837
rect 7440 -858 7474 -837
rect 7368 -871 7370 -858
rect 7370 -871 7402 -858
rect 7440 -871 7472 -858
rect 7472 -871 7474 -858
rect 7596 -858 7630 -837
rect 7668 -858 7702 -837
rect 7596 -871 7598 -858
rect 7598 -871 7630 -858
rect 7668 -871 7700 -858
rect 7700 -871 7702 -858
rect 7118 -1042 7152 -1008
rect 7118 -1142 7152 -1108
rect 6318 -1242 6352 -1208
rect 5518 -1342 5552 -1308
rect 6318 -1342 6352 -1308
rect 4718 -1442 4752 -1408
rect 5518 -1442 5552 -1408
rect 7768 -858 7802 -837
rect 7840 -858 7874 -837
rect 7768 -871 7770 -858
rect 7770 -871 7802 -858
rect 7840 -871 7872 -858
rect 7872 -871 7874 -858
rect 7996 -858 8030 -837
rect 8068 -858 8102 -837
rect 7996 -871 7998 -858
rect 7998 -871 8030 -858
rect 8068 -871 8100 -858
rect 8100 -871 8102 -858
rect 7918 -942 7952 -908
rect 8168 -858 8202 -837
rect 8240 -858 8274 -837
rect 8168 -871 8170 -858
rect 8170 -871 8202 -858
rect 8240 -871 8272 -858
rect 8272 -871 8274 -858
rect 8396 -858 8430 -837
rect 8468 -858 8502 -837
rect 8396 -871 8398 -858
rect 8398 -871 8430 -858
rect 8468 -871 8500 -858
rect 8500 -871 8502 -858
rect 7918 -1042 7952 -1008
rect 7918 -1142 7952 -1108
rect 7118 -1242 7152 -1208
rect 8568 -858 8602 -837
rect 8640 -858 8674 -837
rect 8568 -871 8570 -858
rect 8570 -871 8602 -858
rect 8640 -871 8672 -858
rect 8672 -871 8674 -858
rect 8796 -858 8830 -837
rect 8868 -858 8902 -837
rect 8796 -871 8798 -858
rect 8798 -871 8830 -858
rect 8868 -871 8900 -858
rect 8900 -871 8902 -858
rect 8718 -942 8752 -908
rect 8968 -858 9002 -837
rect 9040 -858 9074 -837
rect 8968 -871 8970 -858
rect 8970 -871 9002 -858
rect 9040 -871 9072 -858
rect 9072 -871 9074 -858
rect 9196 -858 9230 -837
rect 9268 -858 9302 -837
rect 9196 -871 9198 -858
rect 9198 -871 9230 -858
rect 9268 -871 9300 -858
rect 9300 -871 9302 -858
rect 8718 -1042 8752 -1008
rect 8718 -1142 8752 -1108
rect 7918 -1242 7952 -1208
rect 7118 -1342 7152 -1308
rect 7918 -1342 7952 -1308
rect 6318 -1442 6352 -1408
rect 7118 -1442 7152 -1408
rect 4718 -1542 4752 -1508
rect 5518 -1542 5552 -1508
rect 6318 -1542 6352 -1508
rect 3118 -1642 3152 -1608
rect 3918 -1642 3952 -1608
rect 4718 -1642 4752 -1608
rect 5518 -1642 5552 -1608
rect 7118 -1542 7152 -1508
rect 9368 -858 9402 -837
rect 9440 -858 9474 -837
rect 9368 -871 9370 -858
rect 9370 -871 9402 -858
rect 9440 -871 9472 -858
rect 9472 -871 9474 -858
rect 9596 -858 9630 -837
rect 9668 -858 9702 -837
rect 9596 -871 9598 -858
rect 9598 -871 9630 -858
rect 9668 -871 9700 -858
rect 9700 -871 9702 -858
rect 9518 -942 9552 -908
rect 9768 -858 9802 -837
rect 9840 -858 9874 -837
rect 9768 -871 9770 -858
rect 9770 -871 9802 -858
rect 9840 -871 9872 -858
rect 9872 -871 9874 -858
rect 9996 -858 10030 -837
rect 10068 -858 10102 -837
rect 9996 -871 9998 -858
rect 9998 -871 10030 -858
rect 10068 -871 10100 -858
rect 10100 -871 10102 -858
rect 9518 -1042 9552 -1008
rect 9518 -1142 9552 -1108
rect 8718 -1242 8752 -1208
rect 10168 -858 10202 -837
rect 10240 -858 10274 -837
rect 10168 -871 10170 -858
rect 10170 -871 10202 -858
rect 10240 -871 10272 -858
rect 10272 -871 10274 -858
rect 10396 -858 10430 -837
rect 10468 -858 10502 -837
rect 10396 -871 10398 -858
rect 10398 -871 10430 -858
rect 10468 -871 10500 -858
rect 10500 -871 10502 -858
rect 10318 -942 10352 -908
rect 10568 -858 10602 -837
rect 10640 -858 10674 -837
rect 10568 -871 10570 -858
rect 10570 -871 10602 -858
rect 10640 -871 10672 -858
rect 10672 -871 10674 -858
rect 10796 -858 10830 -837
rect 10868 -858 10902 -837
rect 10796 -871 10798 -858
rect 10798 -871 10830 -858
rect 10868 -871 10900 -858
rect 10900 -871 10902 -858
rect 10318 -1042 10352 -1008
rect 10318 -1142 10352 -1108
rect 9518 -1242 9552 -1208
rect 8718 -1342 8752 -1308
rect 9518 -1342 9552 -1308
rect 7918 -1442 7952 -1408
rect 8718 -1442 8752 -1408
rect 10968 -858 11002 -837
rect 11040 -858 11074 -837
rect 10968 -871 10970 -858
rect 10970 -871 11002 -858
rect 11040 -871 11072 -858
rect 11072 -871 11074 -858
rect 11196 -858 11230 -837
rect 11268 -858 11302 -837
rect 11196 -871 11198 -858
rect 11198 -871 11230 -858
rect 11268 -871 11300 -858
rect 11300 -871 11302 -858
rect 11118 -942 11152 -908
rect 11368 -858 11402 -837
rect 11440 -858 11474 -837
rect 11368 -871 11370 -858
rect 11370 -871 11402 -858
rect 11440 -871 11472 -858
rect 11472 -871 11474 -858
rect 11596 -858 11630 -837
rect 11668 -858 11702 -837
rect 11596 -871 11598 -858
rect 11598 -871 11630 -858
rect 11668 -871 11700 -858
rect 11700 -871 11702 -858
rect 11118 -1042 11152 -1008
rect 11118 -1142 11152 -1108
rect 10318 -1242 10352 -1208
rect 11768 -858 11802 -837
rect 11840 -858 11874 -837
rect 11768 -871 11770 -858
rect 11770 -871 11802 -858
rect 11840 -871 11872 -858
rect 11872 -871 11874 -858
rect 11996 -858 12030 -837
rect 12068 -858 12102 -837
rect 11996 -871 11998 -858
rect 11998 -871 12030 -858
rect 12068 -871 12100 -858
rect 12100 -871 12102 -858
rect 11918 -942 11952 -908
rect 12168 -858 12202 -837
rect 12240 -858 12274 -837
rect 12168 -871 12170 -858
rect 12170 -871 12202 -858
rect 12240 -871 12272 -858
rect 12272 -871 12274 -858
rect 12396 -858 12430 -837
rect 12468 -858 12502 -837
rect 12396 -871 12398 -858
rect 12398 -871 12430 -858
rect 12468 -871 12500 -858
rect 12500 -871 12502 -858
rect 11918 -1042 11952 -1008
rect 11918 -1142 11952 -1108
rect 11118 -1242 11152 -1208
rect 10318 -1342 10352 -1308
rect 11118 -1342 11152 -1308
rect 9518 -1442 9552 -1408
rect 10318 -1442 10352 -1408
rect 7918 -1542 7952 -1508
rect 8718 -1542 8752 -1508
rect 9518 -1542 9552 -1508
rect 6318 -1642 6352 -1608
rect 7118 -1642 7152 -1608
rect 7918 -1642 7952 -1608
rect 3118 -1742 3152 -1708
rect 3918 -1742 3952 -1708
rect 4718 -1742 4752 -1708
rect 5518 -1742 5552 -1708
rect 6318 -1742 6352 -1708
rect -82 -1842 -48 -1808
rect 718 -1842 752 -1808
rect 1518 -1842 1552 -1808
rect 2318 -1842 2352 -1808
rect 3118 -1842 3152 -1808
rect -82 -1942 -48 -1908
rect 718 -1942 752 -1908
rect 1518 -1942 1552 -1908
rect 2318 -1942 2352 -1908
rect 3118 -1942 3152 -1908
rect 3918 -1842 3952 -1808
rect 3918 -1942 3952 -1908
rect 4718 -1842 4752 -1808
rect 4718 -1942 4752 -1908
rect 5518 -1842 5552 -1808
rect 5518 -1942 5552 -1908
rect 7118 -1742 7152 -1708
rect 7918 -1742 7952 -1708
rect 8718 -1642 8752 -1608
rect 8718 -1742 8752 -1708
rect 10318 -1542 10352 -1508
rect 12568 -858 12602 -837
rect 12640 -858 12674 -837
rect 12568 -871 12570 -858
rect 12570 -871 12602 -858
rect 12640 -871 12672 -858
rect 12672 -871 12674 -858
rect 14558 -842 14562 -808
rect 14562 -842 14592 -808
rect 14630 -842 14664 -808
rect 14734 -842 14768 -808
rect 14842 -842 14847 -808
rect 14847 -842 14876 -808
rect 14914 -842 14915 -808
rect 14915 -842 14948 -808
rect 14986 -842 15017 -808
rect 15017 -842 15020 -808
rect 15058 -842 15085 -808
rect 15085 -842 15092 -808
rect 15249 -842 15257 -808
rect 15257 -842 15283 -808
rect 15321 -842 15325 -808
rect 15325 -842 15355 -808
rect 15393 -842 15427 -808
rect 15465 -842 15495 -808
rect 15495 -842 15499 -808
rect 15574 -842 15608 -808
rect 15677 -842 15678 -808
rect 15678 -842 15711 -808
rect 15749 -842 15780 -808
rect 15780 -842 15783 -808
rect 12718 -942 12752 -908
rect 14560 -942 14562 -908
rect 14562 -942 14594 -908
rect 14632 -942 14664 -908
rect 14664 -942 14666 -908
rect 14841 -942 14847 -908
rect 14847 -942 14875 -908
rect 14913 -942 14915 -908
rect 14915 -942 14947 -908
rect 14985 -942 15017 -908
rect 15017 -942 15019 -908
rect 15057 -942 15085 -908
rect 15085 -942 15091 -908
rect 15251 -942 15257 -908
rect 15257 -942 15285 -908
rect 15323 -942 15325 -908
rect 15325 -942 15357 -908
rect 15395 -942 15427 -908
rect 15427 -942 15429 -908
rect 15467 -942 15495 -908
rect 15495 -942 15501 -908
rect 15676 -942 15678 -908
rect 15678 -942 15710 -908
rect 15748 -942 15780 -908
rect 15780 -942 15782 -908
rect 12718 -1042 12752 -1008
rect 14558 -1042 14562 -1008
rect 14562 -1042 14592 -1008
rect 14630 -1042 14664 -1008
rect 14734 -1042 14768 -1008
rect 14842 -1042 14847 -1008
rect 14847 -1042 14876 -1008
rect 14914 -1042 14915 -1008
rect 14915 -1042 14948 -1008
rect 14986 -1042 15017 -1008
rect 15017 -1042 15020 -1008
rect 15058 -1042 15085 -1008
rect 15085 -1042 15092 -1008
rect 15249 -1042 15257 -1008
rect 15257 -1042 15283 -1008
rect 15321 -1042 15325 -1008
rect 15325 -1042 15355 -1008
rect 15393 -1042 15427 -1008
rect 15465 -1042 15495 -1008
rect 15495 -1042 15499 -1008
rect 15574 -1042 15608 -1008
rect 15677 -1042 15678 -1008
rect 15678 -1042 15711 -1008
rect 15749 -1042 15780 -1008
rect 15780 -1042 15783 -1008
rect 12718 -1142 12752 -1108
rect 14560 -1142 14562 -1108
rect 14562 -1142 14594 -1108
rect 14632 -1142 14664 -1108
rect 14664 -1142 14666 -1108
rect 11918 -1242 11952 -1208
rect 14841 -1142 14847 -1108
rect 14847 -1142 14875 -1108
rect 14913 -1142 14915 -1108
rect 14915 -1142 14947 -1108
rect 14985 -1142 15017 -1108
rect 15017 -1142 15019 -1108
rect 15057 -1142 15085 -1108
rect 15085 -1142 15091 -1108
rect 15251 -1142 15257 -1108
rect 15257 -1142 15285 -1108
rect 15323 -1142 15325 -1108
rect 15325 -1142 15357 -1108
rect 15395 -1142 15427 -1108
rect 15427 -1142 15429 -1108
rect 15467 -1142 15495 -1108
rect 15495 -1142 15501 -1108
rect 15676 -1142 15678 -1108
rect 15678 -1142 15710 -1108
rect 15748 -1142 15780 -1108
rect 15780 -1142 15782 -1108
rect 12718 -1242 12752 -1208
rect 14558 -1242 14562 -1208
rect 14562 -1242 14592 -1208
rect 14630 -1242 14664 -1208
rect 14734 -1242 14768 -1208
rect 14842 -1242 14847 -1208
rect 14847 -1242 14876 -1208
rect 14914 -1242 14915 -1208
rect 14915 -1242 14948 -1208
rect 14986 -1242 15017 -1208
rect 15017 -1242 15020 -1208
rect 15058 -1242 15085 -1208
rect 15085 -1242 15092 -1208
rect 15249 -1242 15257 -1208
rect 15257 -1242 15283 -1208
rect 15321 -1242 15325 -1208
rect 15325 -1242 15355 -1208
rect 15393 -1242 15427 -1208
rect 15465 -1242 15495 -1208
rect 15495 -1242 15499 -1208
rect 15574 -1242 15608 -1208
rect 15677 -1242 15678 -1208
rect 15678 -1242 15711 -1208
rect 15749 -1242 15780 -1208
rect 15780 -1242 15783 -1208
rect 11918 -1342 11952 -1308
rect 12718 -1342 12752 -1308
rect 14560 -1342 14562 -1308
rect 14562 -1342 14594 -1308
rect 14632 -1342 14664 -1308
rect 14664 -1342 14666 -1308
rect 11118 -1442 11152 -1408
rect 11918 -1442 11952 -1408
rect 14841 -1342 14847 -1308
rect 14847 -1342 14875 -1308
rect 14913 -1342 14915 -1308
rect 14915 -1342 14947 -1308
rect 14985 -1342 15017 -1308
rect 15017 -1342 15019 -1308
rect 15057 -1342 15085 -1308
rect 15085 -1342 15091 -1308
rect 15251 -1342 15257 -1308
rect 15257 -1342 15285 -1308
rect 15323 -1342 15325 -1308
rect 15325 -1342 15357 -1308
rect 15395 -1342 15427 -1308
rect 15427 -1342 15429 -1308
rect 15467 -1342 15495 -1308
rect 15495 -1342 15501 -1308
rect 15676 -1342 15678 -1308
rect 15678 -1342 15710 -1308
rect 15748 -1342 15780 -1308
rect 15780 -1342 15782 -1308
rect 12718 -1442 12752 -1408
rect 14558 -1442 14562 -1408
rect 14562 -1442 14592 -1408
rect 14630 -1442 14664 -1408
rect 14734 -1442 14768 -1408
rect 14842 -1442 14847 -1408
rect 14847 -1442 14876 -1408
rect 14914 -1442 14915 -1408
rect 14915 -1442 14948 -1408
rect 14986 -1442 15017 -1408
rect 15017 -1442 15020 -1408
rect 15058 -1442 15085 -1408
rect 15085 -1442 15092 -1408
rect 15249 -1442 15257 -1408
rect 15257 -1442 15283 -1408
rect 15321 -1442 15325 -1408
rect 15325 -1442 15355 -1408
rect 15393 -1442 15427 -1408
rect 15465 -1442 15495 -1408
rect 15495 -1442 15499 -1408
rect 15574 -1442 15608 -1408
rect 15677 -1442 15678 -1408
rect 15678 -1442 15711 -1408
rect 15749 -1442 15780 -1408
rect 15780 -1442 15783 -1408
rect 11118 -1542 11152 -1508
rect 11918 -1542 11952 -1508
rect 12718 -1542 12752 -1508
rect 14560 -1542 14562 -1508
rect 14562 -1542 14594 -1508
rect 14632 -1542 14664 -1508
rect 14664 -1542 14666 -1508
rect 9518 -1642 9552 -1608
rect 10318 -1642 10352 -1608
rect 11118 -1642 11152 -1608
rect 11918 -1642 11952 -1608
rect 14841 -1542 14847 -1508
rect 14847 -1542 14875 -1508
rect 14913 -1542 14915 -1508
rect 14915 -1542 14947 -1508
rect 14985 -1542 15017 -1508
rect 15017 -1542 15019 -1508
rect 15057 -1542 15085 -1508
rect 15085 -1542 15091 -1508
rect 15251 -1542 15257 -1508
rect 15257 -1542 15285 -1508
rect 15323 -1542 15325 -1508
rect 15325 -1542 15357 -1508
rect 15395 -1542 15427 -1508
rect 15427 -1542 15429 -1508
rect 15467 -1542 15495 -1508
rect 15495 -1542 15501 -1508
rect 15676 -1542 15678 -1508
rect 15678 -1542 15710 -1508
rect 15748 -1542 15780 -1508
rect 15780 -1542 15782 -1508
rect 12718 -1642 12752 -1608
rect 14558 -1642 14562 -1608
rect 14562 -1642 14592 -1608
rect 14630 -1642 14664 -1608
rect 14734 -1642 14768 -1608
rect 14842 -1642 14847 -1608
rect 14847 -1642 14876 -1608
rect 14914 -1642 14915 -1608
rect 14915 -1642 14948 -1608
rect 14986 -1642 15017 -1608
rect 15017 -1642 15020 -1608
rect 15058 -1642 15085 -1608
rect 15085 -1642 15092 -1608
rect 15249 -1642 15257 -1608
rect 15257 -1642 15283 -1608
rect 15321 -1642 15325 -1608
rect 15325 -1642 15355 -1608
rect 15393 -1642 15427 -1608
rect 15465 -1642 15495 -1608
rect 15495 -1642 15499 -1608
rect 15574 -1642 15608 -1608
rect 15677 -1642 15678 -1608
rect 15678 -1642 15711 -1608
rect 15749 -1642 15780 -1608
rect 15780 -1642 15783 -1608
rect 9518 -1742 9552 -1708
rect 10318 -1742 10352 -1708
rect 11118 -1742 11152 -1708
rect 11918 -1742 11952 -1708
rect 12718 -1742 12752 -1708
rect 14560 -1742 14562 -1708
rect 14562 -1742 14594 -1708
rect 14632 -1742 14664 -1708
rect 14664 -1742 14666 -1708
rect 6318 -1842 6352 -1808
rect 7118 -1842 7152 -1808
rect 7918 -1842 7952 -1808
rect 8718 -1842 8752 -1808
rect 9518 -1842 9552 -1808
rect 10318 -1842 10352 -1808
rect 11118 -1842 11152 -1808
rect 11918 -1842 11952 -1808
rect 14841 -1742 14847 -1708
rect 14847 -1742 14875 -1708
rect 14913 -1742 14915 -1708
rect 14915 -1742 14947 -1708
rect 14985 -1742 15017 -1708
rect 15017 -1742 15019 -1708
rect 15057 -1742 15085 -1708
rect 15085 -1742 15091 -1708
rect 15251 -1742 15257 -1708
rect 15257 -1742 15285 -1708
rect 15323 -1742 15325 -1708
rect 15325 -1742 15357 -1708
rect 15395 -1742 15427 -1708
rect 15427 -1742 15429 -1708
rect 15467 -1742 15495 -1708
rect 15495 -1742 15501 -1708
rect 15676 -1742 15678 -1708
rect 15678 -1742 15710 -1708
rect 15748 -1742 15780 -1708
rect 15780 -1742 15782 -1708
rect 12718 -1842 12752 -1808
rect 14558 -1842 14562 -1808
rect 14562 -1842 14592 -1808
rect 14630 -1842 14664 -1808
rect 14734 -1842 14768 -1808
rect 14842 -1842 14847 -1808
rect 14847 -1842 14876 -1808
rect 14914 -1842 14915 -1808
rect 14915 -1842 14948 -1808
rect 14986 -1842 15017 -1808
rect 15017 -1842 15020 -1808
rect 15058 -1842 15085 -1808
rect 15085 -1842 15092 -1808
rect 15249 -1842 15257 -1808
rect 15257 -1842 15283 -1808
rect 15321 -1842 15325 -1808
rect 15325 -1842 15355 -1808
rect 15393 -1842 15427 -1808
rect 15465 -1842 15495 -1808
rect 15495 -1842 15499 -1808
rect 15574 -1842 15608 -1808
rect 15677 -1842 15678 -1808
rect 15678 -1842 15711 -1808
rect 15749 -1842 15780 -1808
rect 15780 -1842 15783 -1808
rect 6318 -1942 6352 -1908
rect 7118 -1942 7152 -1908
rect 7918 -1942 7952 -1908
rect 8718 -1942 8752 -1908
rect 9518 -1942 9552 -1908
rect 10318 -1942 10352 -1908
rect 11118 -1942 11152 -1908
rect 11918 -1942 11952 -1908
rect 12718 -1942 12752 -1908
rect 14560 -1942 14562 -1908
rect 14562 -1942 14594 -1908
rect 14632 -1942 14664 -1908
rect 14664 -1942 14666 -1908
rect -82 -2042 -48 -2008
rect 718 -2042 752 -2008
rect 1518 -2042 1552 -2008
rect 2318 -2042 2352 -2008
rect 3118 -2042 3152 -2008
rect 3918 -2042 3952 -2008
rect 4718 -2042 4752 -2008
rect 5518 -2042 5552 -2008
rect 6318 -2042 6352 -2008
rect 7118 -2042 7152 -2008
rect 7918 -2042 7952 -2008
rect 8718 -2042 8752 -2008
rect 9518 -2042 9552 -2008
rect 10318 -2042 10352 -2008
rect 11118 -2042 11152 -2008
rect 11918 -2042 11952 -2008
rect 14841 -1942 14847 -1908
rect 14847 -1942 14875 -1908
rect 14913 -1942 14915 -1908
rect 14915 -1942 14947 -1908
rect 14985 -1942 15017 -1908
rect 15017 -1942 15019 -1908
rect 15057 -1942 15085 -1908
rect 15085 -1942 15091 -1908
rect 15251 -1942 15257 -1908
rect 15257 -1942 15285 -1908
rect 15323 -1942 15325 -1908
rect 15325 -1942 15357 -1908
rect 15395 -1942 15427 -1908
rect 15427 -1942 15429 -1908
rect 15467 -1942 15495 -1908
rect 15495 -1942 15501 -1908
rect 15676 -1942 15678 -1908
rect 15678 -1942 15710 -1908
rect 15748 -1942 15780 -1908
rect 15780 -1942 15782 -1908
rect 12718 -2042 12752 -2008
rect 14558 -2042 14562 -2008
rect 14562 -2042 14592 -2008
rect 14630 -2042 14664 -2008
rect 14734 -2042 14768 -2008
rect 14842 -2042 14847 -2008
rect 14847 -2042 14876 -2008
rect 14914 -2042 14915 -2008
rect 14915 -2042 14948 -2008
rect 14986 -2042 15017 -2008
rect 15017 -2042 15020 -2008
rect 15058 -2042 15085 -2008
rect 15085 -2042 15092 -2008
rect 15249 -2042 15257 -2008
rect 15257 -2042 15283 -2008
rect 15321 -2042 15325 -2008
rect 15325 -2042 15355 -2008
rect 15393 -2042 15427 -2008
rect 15465 -2042 15495 -2008
rect 15495 -2042 15499 -2008
rect 15574 -2042 15608 -2008
rect 15677 -2042 15678 -2008
rect 15678 -2042 15711 -2008
rect 15749 -2042 15780 -2008
rect 15780 -2042 15783 -2008
rect -4 -2169 30 -2135
rect 68 -2169 102 -2135
rect 168 -2169 202 -2135
rect 240 -2169 274 -2135
rect 396 -2169 430 -2135
rect 468 -2169 502 -2135
rect 568 -2169 602 -2135
rect 640 -2169 674 -2135
rect 796 -2169 830 -2135
rect 868 -2169 902 -2135
rect 968 -2169 1002 -2135
rect 1040 -2169 1074 -2135
rect 1196 -2169 1230 -2135
rect 1268 -2169 1302 -2135
rect 1368 -2169 1402 -2135
rect 1440 -2169 1474 -2135
rect 1596 -2169 1630 -2135
rect 1668 -2169 1702 -2135
rect 1768 -2169 1802 -2135
rect 1840 -2169 1874 -2135
rect 1996 -2169 2030 -2135
rect 2068 -2169 2102 -2135
rect 2168 -2169 2202 -2135
rect 2240 -2169 2274 -2135
rect 2396 -2169 2430 -2135
rect 2468 -2169 2502 -2135
rect 2568 -2169 2602 -2135
rect 2640 -2169 2674 -2135
rect 2796 -2169 2830 -2135
rect 2868 -2169 2902 -2135
rect 2968 -2169 3002 -2135
rect 3040 -2169 3074 -2135
rect 3196 -2169 3230 -2135
rect 3268 -2169 3302 -2135
rect 3368 -2169 3402 -2135
rect 3440 -2169 3474 -2135
rect 3596 -2169 3630 -2135
rect 3668 -2169 3702 -2135
rect 3768 -2169 3802 -2135
rect 3840 -2169 3874 -2135
rect 3996 -2169 4030 -2135
rect 4068 -2169 4102 -2135
rect 4168 -2169 4202 -2135
rect 4240 -2169 4274 -2135
rect 4396 -2169 4430 -2135
rect 4468 -2169 4502 -2135
rect 4568 -2169 4602 -2135
rect 4640 -2169 4674 -2135
rect 4796 -2169 4830 -2135
rect 4868 -2169 4902 -2135
rect 4968 -2169 5002 -2135
rect 5040 -2169 5074 -2135
rect 5196 -2169 5230 -2135
rect 5268 -2169 5302 -2135
rect 5368 -2169 5402 -2135
rect 5440 -2169 5474 -2135
rect 5596 -2169 5630 -2135
rect 5668 -2169 5702 -2135
rect 5768 -2169 5802 -2135
rect 5840 -2169 5874 -2135
rect 5996 -2169 6030 -2135
rect 6068 -2169 6102 -2135
rect 6168 -2169 6202 -2135
rect 6240 -2169 6274 -2135
rect 6396 -2169 6430 -2135
rect 6468 -2169 6502 -2135
rect 6568 -2169 6602 -2135
rect 6640 -2169 6674 -2135
rect 6796 -2169 6830 -2135
rect 6868 -2169 6902 -2135
rect 6968 -2169 7002 -2135
rect 7040 -2169 7074 -2135
rect 7196 -2169 7230 -2135
rect 7268 -2169 7302 -2135
rect 7368 -2169 7402 -2135
rect 7440 -2169 7474 -2135
rect 7596 -2169 7630 -2135
rect 7668 -2169 7702 -2135
rect 7768 -2169 7802 -2135
rect 7840 -2169 7874 -2135
rect 7996 -2169 8030 -2135
rect 8068 -2169 8102 -2135
rect 8168 -2169 8202 -2135
rect 8240 -2169 8274 -2135
rect 8396 -2169 8430 -2135
rect 8468 -2169 8502 -2135
rect 8568 -2169 8602 -2135
rect 8640 -2169 8674 -2135
rect 8796 -2169 8830 -2135
rect 8868 -2169 8902 -2135
rect 8968 -2169 9002 -2135
rect 9040 -2169 9074 -2135
rect 9196 -2169 9230 -2135
rect 9268 -2169 9302 -2135
rect 9368 -2169 9402 -2135
rect 9440 -2169 9474 -2135
rect 9596 -2169 9630 -2135
rect 9668 -2169 9702 -2135
rect 9768 -2169 9802 -2135
rect 9840 -2169 9874 -2135
rect 9996 -2169 10030 -2135
rect 10068 -2169 10102 -2135
rect 10168 -2169 10202 -2135
rect 10240 -2169 10274 -2135
rect 10396 -2169 10430 -2135
rect 10468 -2169 10502 -2135
rect 10568 -2169 10602 -2135
rect 10640 -2169 10674 -2135
rect 10796 -2169 10830 -2135
rect 10868 -2169 10902 -2135
rect 10968 -2169 11002 -2135
rect 11040 -2169 11074 -2135
rect 11196 -2169 11230 -2135
rect 11268 -2169 11302 -2135
rect 11368 -2169 11402 -2135
rect 11440 -2169 11474 -2135
rect 11596 -2169 11630 -2135
rect 11668 -2169 11702 -2135
rect 11768 -2169 11802 -2135
rect 11840 -2169 11874 -2135
rect 11996 -2169 12030 -2135
rect 12068 -2169 12102 -2135
rect 12168 -2169 12202 -2135
rect 12240 -2169 12274 -2135
rect 12396 -2169 12430 -2135
rect 12468 -2169 12502 -2135
rect 12568 -2169 12602 -2135
rect 12640 -2169 12674 -2135
<< metal1 >>
rect 108 5040 162 5070
rect 308 5040 362 5070
rect 508 5040 562 5070
rect 708 5040 762 5070
rect 908 5040 962 5070
rect 1108 5040 1162 5070
rect 1308 5040 1362 5070
rect 1508 5040 1562 5070
rect 1708 5040 1762 5070
rect 1908 5040 1962 5070
rect 2108 5040 2162 5070
rect 2308 5040 2362 5070
rect 2508 5040 2562 5070
rect 2708 5040 2762 5070
rect 2908 5040 2962 5070
rect 3108 5040 3162 5070
rect 3308 5040 3362 5070
rect 3508 5040 3562 5070
rect 3708 5040 3762 5070
rect 3908 5040 3962 5070
rect 4108 5040 4162 5070
rect 4308 5040 4362 5070
rect 4508 5040 4562 5070
rect 4708 5040 4762 5070
rect 4908 5040 4962 5070
rect 5108 5040 5162 5070
rect 5308 5040 5362 5070
rect 5508 5040 5562 5070
rect 5708 5040 5762 5070
rect 5908 5040 5962 5070
rect 6108 5040 6162 5070
rect 6308 5040 6362 5070
rect 6508 5040 6562 5070
rect 6708 5040 6762 5070
rect 6908 5040 6962 5070
rect 7108 5040 7162 5070
rect 7308 5040 7362 5070
rect 7508 5040 7562 5070
rect 7708 5040 7762 5070
rect 7908 5040 7962 5070
rect 8108 5040 8162 5070
rect 8308 5040 8362 5070
rect 8508 5040 8562 5070
rect 8708 5040 8762 5070
rect 8908 5040 8962 5070
rect 9108 5040 9162 5070
rect 9308 5040 9362 5070
rect 9508 5040 9562 5070
rect 9708 5040 9762 5070
rect 9908 5040 9962 5070
rect 10108 5040 10162 5070
rect 10308 5040 10362 5070
rect 10508 5040 10562 5070
rect 10708 5040 10762 5070
rect 10908 5040 10962 5070
rect 11108 5040 11162 5070
rect 11308 5040 11362 5070
rect 11508 5040 11562 5070
rect 11708 5040 11762 5070
rect 11908 5040 11962 5070
rect 12108 5040 12162 5070
rect 12308 5040 12362 5070
rect 12508 5040 12562 5070
rect 12708 5040 12762 5070
rect 35 5017 12835 5040
rect 35 4983 118 5017
rect 152 4983 318 5017
rect 352 4983 518 5017
rect 552 4983 718 5017
rect 752 4983 918 5017
rect 952 4983 1118 5017
rect 1152 4983 1318 5017
rect 1352 4983 1518 5017
rect 1552 4983 1718 5017
rect 1752 4983 1918 5017
rect 1952 4983 2118 5017
rect 2152 4983 2318 5017
rect 2352 4983 2518 5017
rect 2552 4983 2718 5017
rect 2752 4983 2918 5017
rect 2952 4983 3118 5017
rect 3152 4983 3318 5017
rect 3352 4983 3518 5017
rect 3552 4983 3718 5017
rect 3752 4983 3918 5017
rect 3952 4983 4118 5017
rect 4152 4983 4318 5017
rect 4352 4983 4518 5017
rect 4552 4983 4718 5017
rect 4752 4983 4918 5017
rect 4952 4983 5118 5017
rect 5152 4983 5318 5017
rect 5352 4983 5518 5017
rect 5552 4983 5718 5017
rect 5752 4983 5918 5017
rect 5952 4983 6118 5017
rect 6152 4983 6318 5017
rect 6352 4983 6518 5017
rect 6552 4983 6718 5017
rect 6752 4983 6918 5017
rect 6952 4983 7118 5017
rect 7152 4983 7318 5017
rect 7352 4983 7518 5017
rect 7552 4983 7718 5017
rect 7752 4983 7918 5017
rect 7952 4983 8118 5017
rect 8152 4983 8318 5017
rect 8352 4983 8518 5017
rect 8552 4983 8718 5017
rect 8752 4983 8918 5017
rect 8952 4983 9118 5017
rect 9152 4983 9318 5017
rect 9352 4983 9518 5017
rect 9552 4983 9718 5017
rect 9752 4983 9918 5017
rect 9952 4983 10118 5017
rect 10152 4983 10318 5017
rect 10352 4983 10518 5017
rect 10552 4983 10718 5017
rect 10752 4983 10918 5017
rect 10952 4983 11118 5017
rect 11152 4983 11318 5017
rect 11352 4983 11518 5017
rect 11552 4983 11718 5017
rect 11752 4983 11918 5017
rect 11952 4983 12118 5017
rect 12152 4983 12318 5017
rect 12352 4983 12518 5017
rect 12552 4983 12718 5017
rect 12752 4983 12835 5017
rect 35 4960 12835 4983
rect 2 4903 68 4904
rect 2 4851 9 4903
rect 61 4851 68 4903
rect 2 4850 68 4851
rect 8 4787 62 4799
rect 8 4761 18 4787
rect 52 4761 62 4787
rect 8 4709 9 4761
rect 61 4709 62 4761
rect 8 4702 62 4709
rect 108 4787 162 4960
rect 202 4919 268 4920
rect 202 4867 209 4919
rect 261 4867 268 4919
rect 202 4866 268 4867
rect 108 4753 118 4787
rect 152 4753 162 4787
rect 8 4647 62 4659
rect 8 4621 18 4647
rect 52 4621 62 4647
rect 8 4569 9 4621
rect 61 4569 62 4621
rect 8 4562 62 4569
rect 108 4647 162 4753
rect 208 4831 262 4838
rect 208 4779 209 4831
rect 261 4779 262 4831
rect 208 4753 218 4779
rect 252 4753 262 4779
rect 208 4741 262 4753
rect 308 4787 362 4960
rect 402 4903 468 4904
rect 402 4851 409 4903
rect 461 4851 468 4903
rect 402 4850 468 4851
rect 308 4753 318 4787
rect 352 4753 362 4787
rect 108 4613 118 4647
rect 152 4613 162 4647
rect 8 4507 62 4519
rect 8 4481 18 4507
rect 52 4481 62 4507
rect 8 4429 9 4481
rect 61 4429 62 4481
rect 8 4422 62 4429
rect 108 4507 162 4613
rect 208 4691 262 4698
rect 208 4639 209 4691
rect 261 4639 262 4691
rect 208 4613 218 4639
rect 252 4613 262 4639
rect 208 4601 262 4613
rect 308 4647 362 4753
rect 408 4787 462 4799
rect 408 4761 418 4787
rect 452 4761 462 4787
rect 408 4709 409 4761
rect 461 4709 462 4761
rect 408 4702 462 4709
rect 508 4787 562 4960
rect 602 4919 668 4920
rect 602 4867 609 4919
rect 661 4867 668 4919
rect 602 4866 668 4867
rect 508 4753 518 4787
rect 552 4753 562 4787
rect 308 4613 318 4647
rect 352 4613 362 4647
rect 108 4473 118 4507
rect 152 4473 162 4507
rect 8 4367 62 4379
rect 8 4341 18 4367
rect 52 4341 62 4367
rect 8 4289 9 4341
rect 61 4289 62 4341
rect 8 4282 62 4289
rect 108 4367 162 4473
rect 208 4551 262 4558
rect 208 4499 209 4551
rect 261 4499 262 4551
rect 208 4473 218 4499
rect 252 4473 262 4499
rect 208 4461 262 4473
rect 308 4507 362 4613
rect 408 4647 462 4659
rect 408 4621 418 4647
rect 452 4621 462 4647
rect 408 4569 409 4621
rect 461 4569 462 4621
rect 408 4562 462 4569
rect 508 4647 562 4753
rect 608 4831 662 4838
rect 608 4779 609 4831
rect 661 4779 662 4831
rect 608 4753 618 4779
rect 652 4753 662 4779
rect 608 4741 662 4753
rect 708 4787 762 4960
rect 802 4903 868 4904
rect 802 4851 809 4903
rect 861 4851 868 4903
rect 802 4850 868 4851
rect 708 4753 718 4787
rect 752 4753 762 4787
rect 508 4613 518 4647
rect 552 4613 562 4647
rect 308 4473 318 4507
rect 352 4473 362 4507
rect 108 4333 118 4367
rect 152 4333 162 4367
rect 8 4227 62 4239
rect 8 4201 18 4227
rect 52 4201 62 4227
rect 8 4149 9 4201
rect 61 4149 62 4201
rect 8 4142 62 4149
rect 108 4227 162 4333
rect 208 4411 262 4418
rect 208 4359 209 4411
rect 261 4359 262 4411
rect 208 4333 218 4359
rect 252 4333 262 4359
rect 208 4321 262 4333
rect 308 4367 362 4473
rect 408 4507 462 4519
rect 408 4481 418 4507
rect 452 4481 462 4507
rect 408 4429 409 4481
rect 461 4429 462 4481
rect 408 4422 462 4429
rect 508 4507 562 4613
rect 608 4691 662 4698
rect 608 4639 609 4691
rect 661 4639 662 4691
rect 608 4613 618 4639
rect 652 4613 662 4639
rect 608 4601 662 4613
rect 708 4647 762 4753
rect 808 4787 862 4799
rect 808 4761 818 4787
rect 852 4761 862 4787
rect 808 4709 809 4761
rect 861 4709 862 4761
rect 808 4702 862 4709
rect 908 4787 962 4960
rect 1002 4919 1068 4920
rect 1002 4867 1009 4919
rect 1061 4867 1068 4919
rect 1002 4866 1068 4867
rect 908 4753 918 4787
rect 952 4753 962 4787
rect 708 4613 718 4647
rect 752 4613 762 4647
rect 508 4473 518 4507
rect 552 4473 562 4507
rect 308 4333 318 4367
rect 352 4333 362 4367
rect 108 4193 118 4227
rect 152 4193 162 4227
rect 8 4087 62 4099
rect 8 4061 18 4087
rect 52 4061 62 4087
rect 8 4009 9 4061
rect 61 4009 62 4061
rect 8 4002 62 4009
rect 108 4087 162 4193
rect 208 4271 262 4278
rect 208 4219 209 4271
rect 261 4219 262 4271
rect 208 4193 218 4219
rect 252 4193 262 4219
rect 208 4181 262 4193
rect 308 4227 362 4333
rect 408 4367 462 4379
rect 408 4341 418 4367
rect 452 4341 462 4367
rect 408 4289 409 4341
rect 461 4289 462 4341
rect 408 4282 462 4289
rect 508 4367 562 4473
rect 608 4551 662 4558
rect 608 4499 609 4551
rect 661 4499 662 4551
rect 608 4473 618 4499
rect 652 4473 662 4499
rect 608 4461 662 4473
rect 708 4507 762 4613
rect 808 4647 862 4659
rect 808 4621 818 4647
rect 852 4621 862 4647
rect 808 4569 809 4621
rect 861 4569 862 4621
rect 808 4562 862 4569
rect 908 4647 962 4753
rect 1008 4831 1062 4838
rect 1008 4779 1009 4831
rect 1061 4779 1062 4831
rect 1008 4753 1018 4779
rect 1052 4753 1062 4779
rect 1008 4741 1062 4753
rect 1108 4787 1162 4960
rect 1202 4903 1268 4904
rect 1202 4851 1209 4903
rect 1261 4851 1268 4903
rect 1202 4850 1268 4851
rect 1108 4753 1118 4787
rect 1152 4753 1162 4787
rect 908 4613 918 4647
rect 952 4613 962 4647
rect 708 4473 718 4507
rect 752 4473 762 4507
rect 508 4333 518 4367
rect 552 4333 562 4367
rect 308 4193 318 4227
rect 352 4193 362 4227
rect 108 4053 118 4087
rect 152 4053 162 4087
rect 8 3947 62 3959
rect 8 3921 18 3947
rect 52 3921 62 3947
rect 8 3869 9 3921
rect 61 3869 62 3921
rect 8 3862 62 3869
rect 108 3947 162 4053
rect 208 4131 262 4138
rect 208 4079 209 4131
rect 261 4079 262 4131
rect 208 4053 218 4079
rect 252 4053 262 4079
rect 208 4041 262 4053
rect 308 4087 362 4193
rect 408 4227 462 4239
rect 408 4201 418 4227
rect 452 4201 462 4227
rect 408 4149 409 4201
rect 461 4149 462 4201
rect 408 4142 462 4149
rect 508 4227 562 4333
rect 608 4411 662 4418
rect 608 4359 609 4411
rect 661 4359 662 4411
rect 608 4333 618 4359
rect 652 4333 662 4359
rect 608 4321 662 4333
rect 708 4367 762 4473
rect 808 4507 862 4519
rect 808 4481 818 4507
rect 852 4481 862 4507
rect 808 4429 809 4481
rect 861 4429 862 4481
rect 808 4422 862 4429
rect 908 4507 962 4613
rect 1008 4691 1062 4698
rect 1008 4639 1009 4691
rect 1061 4639 1062 4691
rect 1008 4613 1018 4639
rect 1052 4613 1062 4639
rect 1008 4601 1062 4613
rect 1108 4647 1162 4753
rect 1208 4787 1262 4799
rect 1208 4761 1218 4787
rect 1252 4761 1262 4787
rect 1208 4709 1209 4761
rect 1261 4709 1262 4761
rect 1208 4702 1262 4709
rect 1308 4787 1362 4960
rect 1402 4919 1468 4920
rect 1402 4867 1409 4919
rect 1461 4867 1468 4919
rect 1402 4866 1468 4867
rect 1308 4753 1318 4787
rect 1352 4753 1362 4787
rect 1108 4613 1118 4647
rect 1152 4613 1162 4647
rect 908 4473 918 4507
rect 952 4473 962 4507
rect 708 4333 718 4367
rect 752 4333 762 4367
rect 508 4193 518 4227
rect 552 4193 562 4227
rect 308 4053 318 4087
rect 352 4053 362 4087
rect 108 3913 118 3947
rect 152 3913 162 3947
rect 8 3807 62 3819
rect 8 3781 18 3807
rect 52 3781 62 3807
rect 8 3729 9 3781
rect 61 3729 62 3781
rect 8 3722 62 3729
rect 108 3807 162 3913
rect 208 3991 262 3998
rect 208 3939 209 3991
rect 261 3939 262 3991
rect 208 3913 218 3939
rect 252 3913 262 3939
rect 208 3901 262 3913
rect 308 3947 362 4053
rect 408 4087 462 4099
rect 408 4061 418 4087
rect 452 4061 462 4087
rect 408 4009 409 4061
rect 461 4009 462 4061
rect 408 4002 462 4009
rect 508 4087 562 4193
rect 608 4271 662 4278
rect 608 4219 609 4271
rect 661 4219 662 4271
rect 608 4193 618 4219
rect 652 4193 662 4219
rect 608 4181 662 4193
rect 708 4227 762 4333
rect 808 4367 862 4379
rect 808 4341 818 4367
rect 852 4341 862 4367
rect 808 4289 809 4341
rect 861 4289 862 4341
rect 808 4282 862 4289
rect 908 4367 962 4473
rect 1008 4551 1062 4558
rect 1008 4499 1009 4551
rect 1061 4499 1062 4551
rect 1008 4473 1018 4499
rect 1052 4473 1062 4499
rect 1008 4461 1062 4473
rect 1108 4507 1162 4613
rect 1208 4647 1262 4659
rect 1208 4621 1218 4647
rect 1252 4621 1262 4647
rect 1208 4569 1209 4621
rect 1261 4569 1262 4621
rect 1208 4562 1262 4569
rect 1308 4647 1362 4753
rect 1408 4831 1462 4838
rect 1408 4779 1409 4831
rect 1461 4779 1462 4831
rect 1408 4753 1418 4779
rect 1452 4753 1462 4779
rect 1408 4741 1462 4753
rect 1508 4787 1562 4960
rect 1602 4903 1668 4904
rect 1602 4851 1609 4903
rect 1661 4851 1668 4903
rect 1602 4850 1668 4851
rect 1508 4753 1518 4787
rect 1552 4753 1562 4787
rect 1308 4613 1318 4647
rect 1352 4613 1362 4647
rect 1108 4473 1118 4507
rect 1152 4473 1162 4507
rect 908 4333 918 4367
rect 952 4333 962 4367
rect 708 4193 718 4227
rect 752 4193 762 4227
rect 508 4053 518 4087
rect 552 4053 562 4087
rect 308 3913 318 3947
rect 352 3913 362 3947
rect 108 3773 118 3807
rect 152 3773 162 3807
rect 2 3693 68 3694
rect 2 3641 9 3693
rect 61 3641 68 3693
rect 2 3640 68 3641
rect 8 3577 62 3589
rect 8 3551 18 3577
rect 52 3551 62 3577
rect 8 3499 9 3551
rect 61 3499 62 3551
rect 8 3492 62 3499
rect 108 3577 162 3773
rect 208 3851 262 3858
rect 208 3799 209 3851
rect 261 3799 262 3851
rect 208 3773 218 3799
rect 252 3773 262 3799
rect 208 3761 262 3773
rect 308 3807 362 3913
rect 408 3947 462 3959
rect 408 3921 418 3947
rect 452 3921 462 3947
rect 408 3869 409 3921
rect 461 3869 462 3921
rect 408 3862 462 3869
rect 508 3947 562 4053
rect 608 4131 662 4138
rect 608 4079 609 4131
rect 661 4079 662 4131
rect 608 4053 618 4079
rect 652 4053 662 4079
rect 608 4041 662 4053
rect 708 4087 762 4193
rect 808 4227 862 4239
rect 808 4201 818 4227
rect 852 4201 862 4227
rect 808 4149 809 4201
rect 861 4149 862 4201
rect 808 4142 862 4149
rect 908 4227 962 4333
rect 1008 4411 1062 4418
rect 1008 4359 1009 4411
rect 1061 4359 1062 4411
rect 1008 4333 1018 4359
rect 1052 4333 1062 4359
rect 1008 4321 1062 4333
rect 1108 4367 1162 4473
rect 1208 4507 1262 4519
rect 1208 4481 1218 4507
rect 1252 4481 1262 4507
rect 1208 4429 1209 4481
rect 1261 4429 1262 4481
rect 1208 4422 1262 4429
rect 1308 4507 1362 4613
rect 1408 4691 1462 4698
rect 1408 4639 1409 4691
rect 1461 4639 1462 4691
rect 1408 4613 1418 4639
rect 1452 4613 1462 4639
rect 1408 4601 1462 4613
rect 1508 4647 1562 4753
rect 1608 4787 1662 4799
rect 1608 4761 1618 4787
rect 1652 4761 1662 4787
rect 1608 4709 1609 4761
rect 1661 4709 1662 4761
rect 1608 4702 1662 4709
rect 1708 4787 1762 4960
rect 1802 4919 1868 4920
rect 1802 4867 1809 4919
rect 1861 4867 1868 4919
rect 1802 4866 1868 4867
rect 1708 4753 1718 4787
rect 1752 4753 1762 4787
rect 1508 4613 1518 4647
rect 1552 4613 1562 4647
rect 1308 4473 1318 4507
rect 1352 4473 1362 4507
rect 1108 4333 1118 4367
rect 1152 4333 1162 4367
rect 908 4193 918 4227
rect 952 4193 962 4227
rect 708 4053 718 4087
rect 752 4053 762 4087
rect 508 3913 518 3947
rect 552 3913 562 3947
rect 308 3773 318 3807
rect 352 3773 362 3807
rect 202 3709 268 3710
rect 202 3657 209 3709
rect 261 3657 268 3709
rect 202 3656 268 3657
rect 108 3543 118 3577
rect 152 3543 162 3577
rect 8 3437 62 3449
rect 8 3411 18 3437
rect 52 3411 62 3437
rect 8 3359 9 3411
rect 61 3359 62 3411
rect 8 3352 62 3359
rect 108 3437 162 3543
rect 208 3621 262 3628
rect 208 3569 209 3621
rect 261 3569 262 3621
rect 208 3543 218 3569
rect 252 3543 262 3569
rect 208 3531 262 3543
rect 308 3577 362 3773
rect 408 3807 462 3819
rect 408 3781 418 3807
rect 452 3781 462 3807
rect 408 3729 409 3781
rect 461 3729 462 3781
rect 408 3722 462 3729
rect 508 3807 562 3913
rect 608 3991 662 3998
rect 608 3939 609 3991
rect 661 3939 662 3991
rect 608 3913 618 3939
rect 652 3913 662 3939
rect 608 3901 662 3913
rect 708 3947 762 4053
rect 808 4087 862 4099
rect 808 4061 818 4087
rect 852 4061 862 4087
rect 808 4009 809 4061
rect 861 4009 862 4061
rect 808 4002 862 4009
rect 908 4087 962 4193
rect 1008 4271 1062 4278
rect 1008 4219 1009 4271
rect 1061 4219 1062 4271
rect 1008 4193 1018 4219
rect 1052 4193 1062 4219
rect 1008 4181 1062 4193
rect 1108 4227 1162 4333
rect 1208 4367 1262 4379
rect 1208 4341 1218 4367
rect 1252 4341 1262 4367
rect 1208 4289 1209 4341
rect 1261 4289 1262 4341
rect 1208 4282 1262 4289
rect 1308 4367 1362 4473
rect 1408 4551 1462 4558
rect 1408 4499 1409 4551
rect 1461 4499 1462 4551
rect 1408 4473 1418 4499
rect 1452 4473 1462 4499
rect 1408 4461 1462 4473
rect 1508 4507 1562 4613
rect 1608 4647 1662 4659
rect 1608 4621 1618 4647
rect 1652 4621 1662 4647
rect 1608 4569 1609 4621
rect 1661 4569 1662 4621
rect 1608 4562 1662 4569
rect 1708 4647 1762 4753
rect 1808 4831 1862 4838
rect 1808 4779 1809 4831
rect 1861 4779 1862 4831
rect 1808 4753 1818 4779
rect 1852 4753 1862 4779
rect 1808 4741 1862 4753
rect 1908 4787 1962 4960
rect 2002 4903 2068 4904
rect 2002 4851 2009 4903
rect 2061 4851 2068 4903
rect 2002 4850 2068 4851
rect 1908 4753 1918 4787
rect 1952 4753 1962 4787
rect 1708 4613 1718 4647
rect 1752 4613 1762 4647
rect 1508 4473 1518 4507
rect 1552 4473 1562 4507
rect 1308 4333 1318 4367
rect 1352 4333 1362 4367
rect 1108 4193 1118 4227
rect 1152 4193 1162 4227
rect 908 4053 918 4087
rect 952 4053 962 4087
rect 708 3913 718 3947
rect 752 3913 762 3947
rect 508 3773 518 3807
rect 552 3773 562 3807
rect 402 3693 468 3694
rect 402 3641 409 3693
rect 461 3641 468 3693
rect 402 3640 468 3641
rect 308 3543 318 3577
rect 352 3543 362 3577
rect 108 3403 118 3437
rect 152 3403 162 3437
rect 8 3297 62 3309
rect 8 3271 18 3297
rect 52 3271 62 3297
rect 8 3219 9 3271
rect 61 3219 62 3271
rect 8 3212 62 3219
rect 108 3297 162 3403
rect 208 3481 262 3488
rect 208 3429 209 3481
rect 261 3429 262 3481
rect 208 3403 218 3429
rect 252 3403 262 3429
rect 208 3391 262 3403
rect 308 3437 362 3543
rect 408 3577 462 3589
rect 408 3551 418 3577
rect 452 3551 462 3577
rect 408 3499 409 3551
rect 461 3499 462 3551
rect 408 3492 462 3499
rect 508 3577 562 3773
rect 608 3851 662 3858
rect 608 3799 609 3851
rect 661 3799 662 3851
rect 608 3773 618 3799
rect 652 3773 662 3799
rect 608 3761 662 3773
rect 708 3807 762 3913
rect 808 3947 862 3959
rect 808 3921 818 3947
rect 852 3921 862 3947
rect 808 3869 809 3921
rect 861 3869 862 3921
rect 808 3862 862 3869
rect 908 3947 962 4053
rect 1008 4131 1062 4138
rect 1008 4079 1009 4131
rect 1061 4079 1062 4131
rect 1008 4053 1018 4079
rect 1052 4053 1062 4079
rect 1008 4041 1062 4053
rect 1108 4087 1162 4193
rect 1208 4227 1262 4239
rect 1208 4201 1218 4227
rect 1252 4201 1262 4227
rect 1208 4149 1209 4201
rect 1261 4149 1262 4201
rect 1208 4142 1262 4149
rect 1308 4227 1362 4333
rect 1408 4411 1462 4418
rect 1408 4359 1409 4411
rect 1461 4359 1462 4411
rect 1408 4333 1418 4359
rect 1452 4333 1462 4359
rect 1408 4321 1462 4333
rect 1508 4367 1562 4473
rect 1608 4507 1662 4519
rect 1608 4481 1618 4507
rect 1652 4481 1662 4507
rect 1608 4429 1609 4481
rect 1661 4429 1662 4481
rect 1608 4422 1662 4429
rect 1708 4507 1762 4613
rect 1808 4691 1862 4698
rect 1808 4639 1809 4691
rect 1861 4639 1862 4691
rect 1808 4613 1818 4639
rect 1852 4613 1862 4639
rect 1808 4601 1862 4613
rect 1908 4647 1962 4753
rect 2008 4787 2062 4799
rect 2008 4761 2018 4787
rect 2052 4761 2062 4787
rect 2008 4709 2009 4761
rect 2061 4709 2062 4761
rect 2008 4702 2062 4709
rect 2108 4787 2162 4960
rect 2202 4919 2268 4920
rect 2202 4867 2209 4919
rect 2261 4867 2268 4919
rect 2202 4866 2268 4867
rect 2108 4753 2118 4787
rect 2152 4753 2162 4787
rect 1908 4613 1918 4647
rect 1952 4613 1962 4647
rect 1708 4473 1718 4507
rect 1752 4473 1762 4507
rect 1508 4333 1518 4367
rect 1552 4333 1562 4367
rect 1308 4193 1318 4227
rect 1352 4193 1362 4227
rect 1108 4053 1118 4087
rect 1152 4053 1162 4087
rect 908 3913 918 3947
rect 952 3913 962 3947
rect 708 3773 718 3807
rect 752 3773 762 3807
rect 602 3709 668 3710
rect 602 3657 609 3709
rect 661 3657 668 3709
rect 602 3656 668 3657
rect 508 3543 518 3577
rect 552 3543 562 3577
rect 308 3403 318 3437
rect 352 3403 362 3437
rect 108 3263 118 3297
rect 152 3263 162 3297
rect 8 3157 62 3169
rect 8 3131 18 3157
rect 52 3131 62 3157
rect 8 3079 9 3131
rect 61 3079 62 3131
rect 8 3072 62 3079
rect 108 3157 162 3263
rect 208 3341 262 3348
rect 208 3289 209 3341
rect 261 3289 262 3341
rect 208 3263 218 3289
rect 252 3263 262 3289
rect 208 3251 262 3263
rect 308 3297 362 3403
rect 408 3437 462 3449
rect 408 3411 418 3437
rect 452 3411 462 3437
rect 408 3359 409 3411
rect 461 3359 462 3411
rect 408 3352 462 3359
rect 508 3437 562 3543
rect 608 3621 662 3628
rect 608 3569 609 3621
rect 661 3569 662 3621
rect 608 3543 618 3569
rect 652 3543 662 3569
rect 608 3531 662 3543
rect 708 3577 762 3773
rect 808 3807 862 3819
rect 808 3781 818 3807
rect 852 3781 862 3807
rect 808 3729 809 3781
rect 861 3729 862 3781
rect 808 3722 862 3729
rect 908 3807 962 3913
rect 1008 3991 1062 3998
rect 1008 3939 1009 3991
rect 1061 3939 1062 3991
rect 1008 3913 1018 3939
rect 1052 3913 1062 3939
rect 1008 3901 1062 3913
rect 1108 3947 1162 4053
rect 1208 4087 1262 4099
rect 1208 4061 1218 4087
rect 1252 4061 1262 4087
rect 1208 4009 1209 4061
rect 1261 4009 1262 4061
rect 1208 4002 1262 4009
rect 1308 4087 1362 4193
rect 1408 4271 1462 4278
rect 1408 4219 1409 4271
rect 1461 4219 1462 4271
rect 1408 4193 1418 4219
rect 1452 4193 1462 4219
rect 1408 4181 1462 4193
rect 1508 4227 1562 4333
rect 1608 4367 1662 4379
rect 1608 4341 1618 4367
rect 1652 4341 1662 4367
rect 1608 4289 1609 4341
rect 1661 4289 1662 4341
rect 1608 4282 1662 4289
rect 1708 4367 1762 4473
rect 1808 4551 1862 4558
rect 1808 4499 1809 4551
rect 1861 4499 1862 4551
rect 1808 4473 1818 4499
rect 1852 4473 1862 4499
rect 1808 4461 1862 4473
rect 1908 4507 1962 4613
rect 2008 4647 2062 4659
rect 2008 4621 2018 4647
rect 2052 4621 2062 4647
rect 2008 4569 2009 4621
rect 2061 4569 2062 4621
rect 2008 4562 2062 4569
rect 2108 4647 2162 4753
rect 2208 4831 2262 4838
rect 2208 4779 2209 4831
rect 2261 4779 2262 4831
rect 2208 4753 2218 4779
rect 2252 4753 2262 4779
rect 2208 4741 2262 4753
rect 2308 4787 2362 4960
rect 2402 4903 2468 4904
rect 2402 4851 2409 4903
rect 2461 4851 2468 4903
rect 2402 4850 2468 4851
rect 2308 4753 2318 4787
rect 2352 4753 2362 4787
rect 2108 4613 2118 4647
rect 2152 4613 2162 4647
rect 1908 4473 1918 4507
rect 1952 4473 1962 4507
rect 1708 4333 1718 4367
rect 1752 4333 1762 4367
rect 1508 4193 1518 4227
rect 1552 4193 1562 4227
rect 1308 4053 1318 4087
rect 1352 4053 1362 4087
rect 1108 3913 1118 3947
rect 1152 3913 1162 3947
rect 908 3773 918 3807
rect 952 3773 962 3807
rect 802 3693 868 3694
rect 802 3641 809 3693
rect 861 3641 868 3693
rect 802 3640 868 3641
rect 708 3543 718 3577
rect 752 3543 762 3577
rect 508 3403 518 3437
rect 552 3403 562 3437
rect 308 3263 318 3297
rect 352 3263 362 3297
rect 108 3123 118 3157
rect 152 3123 162 3157
rect 8 3017 62 3029
rect 8 2991 18 3017
rect 52 2991 62 3017
rect 8 2939 9 2991
rect 61 2939 62 2991
rect 8 2932 62 2939
rect 108 3017 162 3123
rect 208 3201 262 3208
rect 208 3149 209 3201
rect 261 3149 262 3201
rect 208 3123 218 3149
rect 252 3123 262 3149
rect 208 3111 262 3123
rect 308 3157 362 3263
rect 408 3297 462 3309
rect 408 3271 418 3297
rect 452 3271 462 3297
rect 408 3219 409 3271
rect 461 3219 462 3271
rect 408 3212 462 3219
rect 508 3297 562 3403
rect 608 3481 662 3488
rect 608 3429 609 3481
rect 661 3429 662 3481
rect 608 3403 618 3429
rect 652 3403 662 3429
rect 608 3391 662 3403
rect 708 3437 762 3543
rect 808 3577 862 3589
rect 808 3551 818 3577
rect 852 3551 862 3577
rect 808 3499 809 3551
rect 861 3499 862 3551
rect 808 3492 862 3499
rect 908 3577 962 3773
rect 1008 3851 1062 3858
rect 1008 3799 1009 3851
rect 1061 3799 1062 3851
rect 1008 3773 1018 3799
rect 1052 3773 1062 3799
rect 1008 3761 1062 3773
rect 1108 3807 1162 3913
rect 1208 3947 1262 3959
rect 1208 3921 1218 3947
rect 1252 3921 1262 3947
rect 1208 3869 1209 3921
rect 1261 3869 1262 3921
rect 1208 3862 1262 3869
rect 1308 3947 1362 4053
rect 1408 4131 1462 4138
rect 1408 4079 1409 4131
rect 1461 4079 1462 4131
rect 1408 4053 1418 4079
rect 1452 4053 1462 4079
rect 1408 4041 1462 4053
rect 1508 4087 1562 4193
rect 1608 4227 1662 4239
rect 1608 4201 1618 4227
rect 1652 4201 1662 4227
rect 1608 4149 1609 4201
rect 1661 4149 1662 4201
rect 1608 4142 1662 4149
rect 1708 4227 1762 4333
rect 1808 4411 1862 4418
rect 1808 4359 1809 4411
rect 1861 4359 1862 4411
rect 1808 4333 1818 4359
rect 1852 4333 1862 4359
rect 1808 4321 1862 4333
rect 1908 4367 1962 4473
rect 2008 4507 2062 4519
rect 2008 4481 2018 4507
rect 2052 4481 2062 4507
rect 2008 4429 2009 4481
rect 2061 4429 2062 4481
rect 2008 4422 2062 4429
rect 2108 4507 2162 4613
rect 2208 4691 2262 4698
rect 2208 4639 2209 4691
rect 2261 4639 2262 4691
rect 2208 4613 2218 4639
rect 2252 4613 2262 4639
rect 2208 4601 2262 4613
rect 2308 4647 2362 4753
rect 2408 4787 2462 4799
rect 2408 4761 2418 4787
rect 2452 4761 2462 4787
rect 2408 4709 2409 4761
rect 2461 4709 2462 4761
rect 2408 4702 2462 4709
rect 2508 4787 2562 4960
rect 2602 4919 2668 4920
rect 2602 4867 2609 4919
rect 2661 4867 2668 4919
rect 2602 4866 2668 4867
rect 2508 4753 2518 4787
rect 2552 4753 2562 4787
rect 2308 4613 2318 4647
rect 2352 4613 2362 4647
rect 2108 4473 2118 4507
rect 2152 4473 2162 4507
rect 1908 4333 1918 4367
rect 1952 4333 1962 4367
rect 1708 4193 1718 4227
rect 1752 4193 1762 4227
rect 1508 4053 1518 4087
rect 1552 4053 1562 4087
rect 1308 3913 1318 3947
rect 1352 3913 1362 3947
rect 1108 3773 1118 3807
rect 1152 3773 1162 3807
rect 1002 3709 1068 3710
rect 1002 3657 1009 3709
rect 1061 3657 1068 3709
rect 1002 3656 1068 3657
rect 908 3543 918 3577
rect 952 3543 962 3577
rect 708 3403 718 3437
rect 752 3403 762 3437
rect 508 3263 518 3297
rect 552 3263 562 3297
rect 308 3123 318 3157
rect 352 3123 362 3157
rect 108 2983 118 3017
rect 152 2983 162 3017
rect 8 2877 62 2889
rect 8 2851 18 2877
rect 52 2851 62 2877
rect 8 2799 9 2851
rect 61 2799 62 2851
rect 8 2792 62 2799
rect 108 2877 162 2983
rect 208 3061 262 3068
rect 208 3009 209 3061
rect 261 3009 262 3061
rect 208 2983 218 3009
rect 252 2983 262 3009
rect 208 2971 262 2983
rect 308 3017 362 3123
rect 408 3157 462 3169
rect 408 3131 418 3157
rect 452 3131 462 3157
rect 408 3079 409 3131
rect 461 3079 462 3131
rect 408 3072 462 3079
rect 508 3157 562 3263
rect 608 3341 662 3348
rect 608 3289 609 3341
rect 661 3289 662 3341
rect 608 3263 618 3289
rect 652 3263 662 3289
rect 608 3251 662 3263
rect 708 3297 762 3403
rect 808 3437 862 3449
rect 808 3411 818 3437
rect 852 3411 862 3437
rect 808 3359 809 3411
rect 861 3359 862 3411
rect 808 3352 862 3359
rect 908 3437 962 3543
rect 1008 3621 1062 3628
rect 1008 3569 1009 3621
rect 1061 3569 1062 3621
rect 1008 3543 1018 3569
rect 1052 3543 1062 3569
rect 1008 3531 1062 3543
rect 1108 3577 1162 3773
rect 1208 3807 1262 3819
rect 1208 3781 1218 3807
rect 1252 3781 1262 3807
rect 1208 3729 1209 3781
rect 1261 3729 1262 3781
rect 1208 3722 1262 3729
rect 1308 3807 1362 3913
rect 1408 3991 1462 3998
rect 1408 3939 1409 3991
rect 1461 3939 1462 3991
rect 1408 3913 1418 3939
rect 1452 3913 1462 3939
rect 1408 3901 1462 3913
rect 1508 3947 1562 4053
rect 1608 4087 1662 4099
rect 1608 4061 1618 4087
rect 1652 4061 1662 4087
rect 1608 4009 1609 4061
rect 1661 4009 1662 4061
rect 1608 4002 1662 4009
rect 1708 4087 1762 4193
rect 1808 4271 1862 4278
rect 1808 4219 1809 4271
rect 1861 4219 1862 4271
rect 1808 4193 1818 4219
rect 1852 4193 1862 4219
rect 1808 4181 1862 4193
rect 1908 4227 1962 4333
rect 2008 4367 2062 4379
rect 2008 4341 2018 4367
rect 2052 4341 2062 4367
rect 2008 4289 2009 4341
rect 2061 4289 2062 4341
rect 2008 4282 2062 4289
rect 2108 4367 2162 4473
rect 2208 4551 2262 4558
rect 2208 4499 2209 4551
rect 2261 4499 2262 4551
rect 2208 4473 2218 4499
rect 2252 4473 2262 4499
rect 2208 4461 2262 4473
rect 2308 4507 2362 4613
rect 2408 4647 2462 4659
rect 2408 4621 2418 4647
rect 2452 4621 2462 4647
rect 2408 4569 2409 4621
rect 2461 4569 2462 4621
rect 2408 4562 2462 4569
rect 2508 4647 2562 4753
rect 2608 4831 2662 4838
rect 2608 4779 2609 4831
rect 2661 4779 2662 4831
rect 2608 4753 2618 4779
rect 2652 4753 2662 4779
rect 2608 4741 2662 4753
rect 2708 4787 2762 4960
rect 2802 4903 2868 4904
rect 2802 4851 2809 4903
rect 2861 4851 2868 4903
rect 2802 4850 2868 4851
rect 2708 4753 2718 4787
rect 2752 4753 2762 4787
rect 2508 4613 2518 4647
rect 2552 4613 2562 4647
rect 2308 4473 2318 4507
rect 2352 4473 2362 4507
rect 2108 4333 2118 4367
rect 2152 4333 2162 4367
rect 1908 4193 1918 4227
rect 1952 4193 1962 4227
rect 1708 4053 1718 4087
rect 1752 4053 1762 4087
rect 1508 3913 1518 3947
rect 1552 3913 1562 3947
rect 1308 3773 1318 3807
rect 1352 3773 1362 3807
rect 1202 3693 1268 3694
rect 1202 3641 1209 3693
rect 1261 3641 1268 3693
rect 1202 3640 1268 3641
rect 1108 3543 1118 3577
rect 1152 3543 1162 3577
rect 908 3403 918 3437
rect 952 3403 962 3437
rect 708 3263 718 3297
rect 752 3263 762 3297
rect 508 3123 518 3157
rect 552 3123 562 3157
rect 308 2983 318 3017
rect 352 2983 362 3017
rect 108 2843 118 2877
rect 152 2843 162 2877
rect 8 2737 62 2749
rect 8 2711 18 2737
rect 52 2711 62 2737
rect 8 2659 9 2711
rect 61 2659 62 2711
rect 8 2652 62 2659
rect 108 2737 162 2843
rect 208 2921 262 2928
rect 208 2869 209 2921
rect 261 2869 262 2921
rect 208 2843 218 2869
rect 252 2843 262 2869
rect 208 2831 262 2843
rect 308 2877 362 2983
rect 408 3017 462 3029
rect 408 2991 418 3017
rect 452 2991 462 3017
rect 408 2939 409 2991
rect 461 2939 462 2991
rect 408 2932 462 2939
rect 508 3017 562 3123
rect 608 3201 662 3208
rect 608 3149 609 3201
rect 661 3149 662 3201
rect 608 3123 618 3149
rect 652 3123 662 3149
rect 608 3111 662 3123
rect 708 3157 762 3263
rect 808 3297 862 3309
rect 808 3271 818 3297
rect 852 3271 862 3297
rect 808 3219 809 3271
rect 861 3219 862 3271
rect 808 3212 862 3219
rect 908 3297 962 3403
rect 1008 3481 1062 3488
rect 1008 3429 1009 3481
rect 1061 3429 1062 3481
rect 1008 3403 1018 3429
rect 1052 3403 1062 3429
rect 1008 3391 1062 3403
rect 1108 3437 1162 3543
rect 1208 3577 1262 3589
rect 1208 3551 1218 3577
rect 1252 3551 1262 3577
rect 1208 3499 1209 3551
rect 1261 3499 1262 3551
rect 1208 3492 1262 3499
rect 1308 3577 1362 3773
rect 1408 3851 1462 3858
rect 1408 3799 1409 3851
rect 1461 3799 1462 3851
rect 1408 3773 1418 3799
rect 1452 3773 1462 3799
rect 1408 3761 1462 3773
rect 1508 3807 1562 3913
rect 1608 3947 1662 3959
rect 1608 3921 1618 3947
rect 1652 3921 1662 3947
rect 1608 3869 1609 3921
rect 1661 3869 1662 3921
rect 1608 3862 1662 3869
rect 1708 3947 1762 4053
rect 1808 4131 1862 4138
rect 1808 4079 1809 4131
rect 1861 4079 1862 4131
rect 1808 4053 1818 4079
rect 1852 4053 1862 4079
rect 1808 4041 1862 4053
rect 1908 4087 1962 4193
rect 2008 4227 2062 4239
rect 2008 4201 2018 4227
rect 2052 4201 2062 4227
rect 2008 4149 2009 4201
rect 2061 4149 2062 4201
rect 2008 4142 2062 4149
rect 2108 4227 2162 4333
rect 2208 4411 2262 4418
rect 2208 4359 2209 4411
rect 2261 4359 2262 4411
rect 2208 4333 2218 4359
rect 2252 4333 2262 4359
rect 2208 4321 2262 4333
rect 2308 4367 2362 4473
rect 2408 4507 2462 4519
rect 2408 4481 2418 4507
rect 2452 4481 2462 4507
rect 2408 4429 2409 4481
rect 2461 4429 2462 4481
rect 2408 4422 2462 4429
rect 2508 4507 2562 4613
rect 2608 4691 2662 4698
rect 2608 4639 2609 4691
rect 2661 4639 2662 4691
rect 2608 4613 2618 4639
rect 2652 4613 2662 4639
rect 2608 4601 2662 4613
rect 2708 4647 2762 4753
rect 2808 4787 2862 4799
rect 2808 4761 2818 4787
rect 2852 4761 2862 4787
rect 2808 4709 2809 4761
rect 2861 4709 2862 4761
rect 2808 4702 2862 4709
rect 2908 4787 2962 4960
rect 3002 4919 3068 4920
rect 3002 4867 3009 4919
rect 3061 4867 3068 4919
rect 3002 4866 3068 4867
rect 2908 4753 2918 4787
rect 2952 4753 2962 4787
rect 2708 4613 2718 4647
rect 2752 4613 2762 4647
rect 2508 4473 2518 4507
rect 2552 4473 2562 4507
rect 2308 4333 2318 4367
rect 2352 4333 2362 4367
rect 2108 4193 2118 4227
rect 2152 4193 2162 4227
rect 1908 4053 1918 4087
rect 1952 4053 1962 4087
rect 1708 3913 1718 3947
rect 1752 3913 1762 3947
rect 1508 3773 1518 3807
rect 1552 3773 1562 3807
rect 1402 3709 1468 3710
rect 1402 3657 1409 3709
rect 1461 3657 1468 3709
rect 1402 3656 1468 3657
rect 1308 3543 1318 3577
rect 1352 3543 1362 3577
rect 1108 3403 1118 3437
rect 1152 3403 1162 3437
rect 908 3263 918 3297
rect 952 3263 962 3297
rect 708 3123 718 3157
rect 752 3123 762 3157
rect 508 2983 518 3017
rect 552 2983 562 3017
rect 308 2843 318 2877
rect 352 2843 362 2877
rect 108 2703 118 2737
rect 152 2703 162 2737
rect 8 2597 62 2609
rect 8 2571 18 2597
rect 52 2571 62 2597
rect 8 2519 9 2571
rect 61 2519 62 2571
rect 8 2512 62 2519
rect 108 2597 162 2703
rect 208 2781 262 2788
rect 208 2729 209 2781
rect 261 2729 262 2781
rect 208 2703 218 2729
rect 252 2703 262 2729
rect 208 2691 262 2703
rect 308 2737 362 2843
rect 408 2877 462 2889
rect 408 2851 418 2877
rect 452 2851 462 2877
rect 408 2799 409 2851
rect 461 2799 462 2851
rect 408 2792 462 2799
rect 508 2877 562 2983
rect 608 3061 662 3068
rect 608 3009 609 3061
rect 661 3009 662 3061
rect 608 2983 618 3009
rect 652 2983 662 3009
rect 608 2971 662 2983
rect 708 3017 762 3123
rect 808 3157 862 3169
rect 808 3131 818 3157
rect 852 3131 862 3157
rect 808 3079 809 3131
rect 861 3079 862 3131
rect 808 3072 862 3079
rect 908 3157 962 3263
rect 1008 3341 1062 3348
rect 1008 3289 1009 3341
rect 1061 3289 1062 3341
rect 1008 3263 1018 3289
rect 1052 3263 1062 3289
rect 1008 3251 1062 3263
rect 1108 3297 1162 3403
rect 1208 3437 1262 3449
rect 1208 3411 1218 3437
rect 1252 3411 1262 3437
rect 1208 3359 1209 3411
rect 1261 3359 1262 3411
rect 1208 3352 1262 3359
rect 1308 3437 1362 3543
rect 1408 3621 1462 3628
rect 1408 3569 1409 3621
rect 1461 3569 1462 3621
rect 1408 3543 1418 3569
rect 1452 3543 1462 3569
rect 1408 3531 1462 3543
rect 1508 3577 1562 3773
rect 1608 3807 1662 3819
rect 1608 3781 1618 3807
rect 1652 3781 1662 3807
rect 1608 3729 1609 3781
rect 1661 3729 1662 3781
rect 1608 3722 1662 3729
rect 1708 3807 1762 3913
rect 1808 3991 1862 3998
rect 1808 3939 1809 3991
rect 1861 3939 1862 3991
rect 1808 3913 1818 3939
rect 1852 3913 1862 3939
rect 1808 3901 1862 3913
rect 1908 3947 1962 4053
rect 2008 4087 2062 4099
rect 2008 4061 2018 4087
rect 2052 4061 2062 4087
rect 2008 4009 2009 4061
rect 2061 4009 2062 4061
rect 2008 4002 2062 4009
rect 2108 4087 2162 4193
rect 2208 4271 2262 4278
rect 2208 4219 2209 4271
rect 2261 4219 2262 4271
rect 2208 4193 2218 4219
rect 2252 4193 2262 4219
rect 2208 4181 2262 4193
rect 2308 4227 2362 4333
rect 2408 4367 2462 4379
rect 2408 4341 2418 4367
rect 2452 4341 2462 4367
rect 2408 4289 2409 4341
rect 2461 4289 2462 4341
rect 2408 4282 2462 4289
rect 2508 4367 2562 4473
rect 2608 4551 2662 4558
rect 2608 4499 2609 4551
rect 2661 4499 2662 4551
rect 2608 4473 2618 4499
rect 2652 4473 2662 4499
rect 2608 4461 2662 4473
rect 2708 4507 2762 4613
rect 2808 4647 2862 4659
rect 2808 4621 2818 4647
rect 2852 4621 2862 4647
rect 2808 4569 2809 4621
rect 2861 4569 2862 4621
rect 2808 4562 2862 4569
rect 2908 4647 2962 4753
rect 3008 4831 3062 4838
rect 3008 4779 3009 4831
rect 3061 4779 3062 4831
rect 3008 4753 3018 4779
rect 3052 4753 3062 4779
rect 3008 4741 3062 4753
rect 3108 4787 3162 4960
rect 3202 4903 3268 4904
rect 3202 4851 3209 4903
rect 3261 4851 3268 4903
rect 3202 4850 3268 4851
rect 3108 4753 3118 4787
rect 3152 4753 3162 4787
rect 2908 4613 2918 4647
rect 2952 4613 2962 4647
rect 2708 4473 2718 4507
rect 2752 4473 2762 4507
rect 2508 4333 2518 4367
rect 2552 4333 2562 4367
rect 2308 4193 2318 4227
rect 2352 4193 2362 4227
rect 2108 4053 2118 4087
rect 2152 4053 2162 4087
rect 1908 3913 1918 3947
rect 1952 3913 1962 3947
rect 1708 3773 1718 3807
rect 1752 3773 1762 3807
rect 1602 3693 1668 3694
rect 1602 3641 1609 3693
rect 1661 3641 1668 3693
rect 1602 3640 1668 3641
rect 1508 3543 1518 3577
rect 1552 3543 1562 3577
rect 1308 3403 1318 3437
rect 1352 3403 1362 3437
rect 1108 3263 1118 3297
rect 1152 3263 1162 3297
rect 908 3123 918 3157
rect 952 3123 962 3157
rect 708 2983 718 3017
rect 752 2983 762 3017
rect 508 2843 518 2877
rect 552 2843 562 2877
rect 308 2703 318 2737
rect 352 2703 362 2737
rect 108 2563 118 2597
rect 152 2563 162 2597
rect 2 2483 68 2484
rect 2 2431 9 2483
rect 61 2431 68 2483
rect 2 2430 68 2431
rect 8 2367 62 2379
rect 8 2341 18 2367
rect 52 2341 62 2367
rect 8 2289 9 2341
rect 61 2289 62 2341
rect 8 2282 62 2289
rect 108 2367 162 2563
rect 208 2641 262 2648
rect 208 2589 209 2641
rect 261 2589 262 2641
rect 208 2563 218 2589
rect 252 2563 262 2589
rect 208 2551 262 2563
rect 308 2597 362 2703
rect 408 2737 462 2749
rect 408 2711 418 2737
rect 452 2711 462 2737
rect 408 2659 409 2711
rect 461 2659 462 2711
rect 408 2652 462 2659
rect 508 2737 562 2843
rect 608 2921 662 2928
rect 608 2869 609 2921
rect 661 2869 662 2921
rect 608 2843 618 2869
rect 652 2843 662 2869
rect 608 2831 662 2843
rect 708 2877 762 2983
rect 808 3017 862 3029
rect 808 2991 818 3017
rect 852 2991 862 3017
rect 808 2939 809 2991
rect 861 2939 862 2991
rect 808 2932 862 2939
rect 908 3017 962 3123
rect 1008 3201 1062 3208
rect 1008 3149 1009 3201
rect 1061 3149 1062 3201
rect 1008 3123 1018 3149
rect 1052 3123 1062 3149
rect 1008 3111 1062 3123
rect 1108 3157 1162 3263
rect 1208 3297 1262 3309
rect 1208 3271 1218 3297
rect 1252 3271 1262 3297
rect 1208 3219 1209 3271
rect 1261 3219 1262 3271
rect 1208 3212 1262 3219
rect 1308 3297 1362 3403
rect 1408 3481 1462 3488
rect 1408 3429 1409 3481
rect 1461 3429 1462 3481
rect 1408 3403 1418 3429
rect 1452 3403 1462 3429
rect 1408 3391 1462 3403
rect 1508 3437 1562 3543
rect 1608 3577 1662 3589
rect 1608 3551 1618 3577
rect 1652 3551 1662 3577
rect 1608 3499 1609 3551
rect 1661 3499 1662 3551
rect 1608 3492 1662 3499
rect 1708 3577 1762 3773
rect 1808 3851 1862 3858
rect 1808 3799 1809 3851
rect 1861 3799 1862 3851
rect 1808 3773 1818 3799
rect 1852 3773 1862 3799
rect 1808 3761 1862 3773
rect 1908 3807 1962 3913
rect 2008 3947 2062 3959
rect 2008 3921 2018 3947
rect 2052 3921 2062 3947
rect 2008 3869 2009 3921
rect 2061 3869 2062 3921
rect 2008 3862 2062 3869
rect 2108 3947 2162 4053
rect 2208 4131 2262 4138
rect 2208 4079 2209 4131
rect 2261 4079 2262 4131
rect 2208 4053 2218 4079
rect 2252 4053 2262 4079
rect 2208 4041 2262 4053
rect 2308 4087 2362 4193
rect 2408 4227 2462 4239
rect 2408 4201 2418 4227
rect 2452 4201 2462 4227
rect 2408 4149 2409 4201
rect 2461 4149 2462 4201
rect 2408 4142 2462 4149
rect 2508 4227 2562 4333
rect 2608 4411 2662 4418
rect 2608 4359 2609 4411
rect 2661 4359 2662 4411
rect 2608 4333 2618 4359
rect 2652 4333 2662 4359
rect 2608 4321 2662 4333
rect 2708 4367 2762 4473
rect 2808 4507 2862 4519
rect 2808 4481 2818 4507
rect 2852 4481 2862 4507
rect 2808 4429 2809 4481
rect 2861 4429 2862 4481
rect 2808 4422 2862 4429
rect 2908 4507 2962 4613
rect 3008 4691 3062 4698
rect 3008 4639 3009 4691
rect 3061 4639 3062 4691
rect 3008 4613 3018 4639
rect 3052 4613 3062 4639
rect 3008 4601 3062 4613
rect 3108 4647 3162 4753
rect 3208 4787 3262 4799
rect 3208 4761 3218 4787
rect 3252 4761 3262 4787
rect 3208 4709 3209 4761
rect 3261 4709 3262 4761
rect 3208 4702 3262 4709
rect 3308 4787 3362 4960
rect 3402 4919 3468 4920
rect 3402 4867 3409 4919
rect 3461 4867 3468 4919
rect 3402 4866 3468 4867
rect 3308 4753 3318 4787
rect 3352 4753 3362 4787
rect 3108 4613 3118 4647
rect 3152 4613 3162 4647
rect 2908 4473 2918 4507
rect 2952 4473 2962 4507
rect 2708 4333 2718 4367
rect 2752 4333 2762 4367
rect 2508 4193 2518 4227
rect 2552 4193 2562 4227
rect 2308 4053 2318 4087
rect 2352 4053 2362 4087
rect 2108 3913 2118 3947
rect 2152 3913 2162 3947
rect 1908 3773 1918 3807
rect 1952 3773 1962 3807
rect 1802 3709 1868 3710
rect 1802 3657 1809 3709
rect 1861 3657 1868 3709
rect 1802 3656 1868 3657
rect 1708 3543 1718 3577
rect 1752 3543 1762 3577
rect 1508 3403 1518 3437
rect 1552 3403 1562 3437
rect 1308 3263 1318 3297
rect 1352 3263 1362 3297
rect 1108 3123 1118 3157
rect 1152 3123 1162 3157
rect 908 2983 918 3017
rect 952 2983 962 3017
rect 708 2843 718 2877
rect 752 2843 762 2877
rect 508 2703 518 2737
rect 552 2703 562 2737
rect 308 2563 318 2597
rect 352 2563 362 2597
rect 202 2499 268 2500
rect 202 2447 209 2499
rect 261 2447 268 2499
rect 202 2446 268 2447
rect 108 2333 118 2367
rect 152 2333 162 2367
rect 8 2227 62 2239
rect 8 2201 18 2227
rect 52 2201 62 2227
rect 8 2149 9 2201
rect 61 2149 62 2201
rect 8 2142 62 2149
rect 108 2227 162 2333
rect 208 2411 262 2418
rect 208 2359 209 2411
rect 261 2359 262 2411
rect 208 2333 218 2359
rect 252 2333 262 2359
rect 208 2321 262 2333
rect 308 2367 362 2563
rect 408 2597 462 2609
rect 408 2571 418 2597
rect 452 2571 462 2597
rect 408 2519 409 2571
rect 461 2519 462 2571
rect 408 2512 462 2519
rect 508 2597 562 2703
rect 608 2781 662 2788
rect 608 2729 609 2781
rect 661 2729 662 2781
rect 608 2703 618 2729
rect 652 2703 662 2729
rect 608 2691 662 2703
rect 708 2737 762 2843
rect 808 2877 862 2889
rect 808 2851 818 2877
rect 852 2851 862 2877
rect 808 2799 809 2851
rect 861 2799 862 2851
rect 808 2792 862 2799
rect 908 2877 962 2983
rect 1008 3061 1062 3068
rect 1008 3009 1009 3061
rect 1061 3009 1062 3061
rect 1008 2983 1018 3009
rect 1052 2983 1062 3009
rect 1008 2971 1062 2983
rect 1108 3017 1162 3123
rect 1208 3157 1262 3169
rect 1208 3131 1218 3157
rect 1252 3131 1262 3157
rect 1208 3079 1209 3131
rect 1261 3079 1262 3131
rect 1208 3072 1262 3079
rect 1308 3157 1362 3263
rect 1408 3341 1462 3348
rect 1408 3289 1409 3341
rect 1461 3289 1462 3341
rect 1408 3263 1418 3289
rect 1452 3263 1462 3289
rect 1408 3251 1462 3263
rect 1508 3297 1562 3403
rect 1608 3437 1662 3449
rect 1608 3411 1618 3437
rect 1652 3411 1662 3437
rect 1608 3359 1609 3411
rect 1661 3359 1662 3411
rect 1608 3352 1662 3359
rect 1708 3437 1762 3543
rect 1808 3621 1862 3628
rect 1808 3569 1809 3621
rect 1861 3569 1862 3621
rect 1808 3543 1818 3569
rect 1852 3543 1862 3569
rect 1808 3531 1862 3543
rect 1908 3577 1962 3773
rect 2008 3807 2062 3819
rect 2008 3781 2018 3807
rect 2052 3781 2062 3807
rect 2008 3729 2009 3781
rect 2061 3729 2062 3781
rect 2008 3722 2062 3729
rect 2108 3807 2162 3913
rect 2208 3991 2262 3998
rect 2208 3939 2209 3991
rect 2261 3939 2262 3991
rect 2208 3913 2218 3939
rect 2252 3913 2262 3939
rect 2208 3901 2262 3913
rect 2308 3947 2362 4053
rect 2408 4087 2462 4099
rect 2408 4061 2418 4087
rect 2452 4061 2462 4087
rect 2408 4009 2409 4061
rect 2461 4009 2462 4061
rect 2408 4002 2462 4009
rect 2508 4087 2562 4193
rect 2608 4271 2662 4278
rect 2608 4219 2609 4271
rect 2661 4219 2662 4271
rect 2608 4193 2618 4219
rect 2652 4193 2662 4219
rect 2608 4181 2662 4193
rect 2708 4227 2762 4333
rect 2808 4367 2862 4379
rect 2808 4341 2818 4367
rect 2852 4341 2862 4367
rect 2808 4289 2809 4341
rect 2861 4289 2862 4341
rect 2808 4282 2862 4289
rect 2908 4367 2962 4473
rect 3008 4551 3062 4558
rect 3008 4499 3009 4551
rect 3061 4499 3062 4551
rect 3008 4473 3018 4499
rect 3052 4473 3062 4499
rect 3008 4461 3062 4473
rect 3108 4507 3162 4613
rect 3208 4647 3262 4659
rect 3208 4621 3218 4647
rect 3252 4621 3262 4647
rect 3208 4569 3209 4621
rect 3261 4569 3262 4621
rect 3208 4562 3262 4569
rect 3308 4647 3362 4753
rect 3408 4831 3462 4838
rect 3408 4779 3409 4831
rect 3461 4779 3462 4831
rect 3408 4753 3418 4779
rect 3452 4753 3462 4779
rect 3408 4741 3462 4753
rect 3508 4787 3562 4960
rect 3602 4903 3668 4904
rect 3602 4851 3609 4903
rect 3661 4851 3668 4903
rect 3602 4850 3668 4851
rect 3508 4753 3518 4787
rect 3552 4753 3562 4787
rect 3308 4613 3318 4647
rect 3352 4613 3362 4647
rect 3108 4473 3118 4507
rect 3152 4473 3162 4507
rect 2908 4333 2918 4367
rect 2952 4333 2962 4367
rect 2708 4193 2718 4227
rect 2752 4193 2762 4227
rect 2508 4053 2518 4087
rect 2552 4053 2562 4087
rect 2308 3913 2318 3947
rect 2352 3913 2362 3947
rect 2108 3773 2118 3807
rect 2152 3773 2162 3807
rect 2002 3693 2068 3694
rect 2002 3641 2009 3693
rect 2061 3641 2068 3693
rect 2002 3640 2068 3641
rect 1908 3543 1918 3577
rect 1952 3543 1962 3577
rect 1708 3403 1718 3437
rect 1752 3403 1762 3437
rect 1508 3263 1518 3297
rect 1552 3263 1562 3297
rect 1308 3123 1318 3157
rect 1352 3123 1362 3157
rect 1108 2983 1118 3017
rect 1152 2983 1162 3017
rect 908 2843 918 2877
rect 952 2843 962 2877
rect 708 2703 718 2737
rect 752 2703 762 2737
rect 508 2563 518 2597
rect 552 2563 562 2597
rect 402 2483 468 2484
rect 402 2431 409 2483
rect 461 2431 468 2483
rect 402 2430 468 2431
rect 308 2333 318 2367
rect 352 2333 362 2367
rect 108 2193 118 2227
rect 152 2193 162 2227
rect 8 2087 62 2099
rect 8 2061 18 2087
rect 52 2061 62 2087
rect 8 2009 9 2061
rect 61 2009 62 2061
rect 8 2002 62 2009
rect 108 2087 162 2193
rect 208 2271 262 2278
rect 208 2219 209 2271
rect 261 2219 262 2271
rect 208 2193 218 2219
rect 252 2193 262 2219
rect 208 2181 262 2193
rect 308 2227 362 2333
rect 408 2367 462 2379
rect 408 2341 418 2367
rect 452 2341 462 2367
rect 408 2289 409 2341
rect 461 2289 462 2341
rect 408 2282 462 2289
rect 508 2367 562 2563
rect 608 2641 662 2648
rect 608 2589 609 2641
rect 661 2589 662 2641
rect 608 2563 618 2589
rect 652 2563 662 2589
rect 608 2551 662 2563
rect 708 2597 762 2703
rect 808 2737 862 2749
rect 808 2711 818 2737
rect 852 2711 862 2737
rect 808 2659 809 2711
rect 861 2659 862 2711
rect 808 2652 862 2659
rect 908 2737 962 2843
rect 1008 2921 1062 2928
rect 1008 2869 1009 2921
rect 1061 2869 1062 2921
rect 1008 2843 1018 2869
rect 1052 2843 1062 2869
rect 1008 2831 1062 2843
rect 1108 2877 1162 2983
rect 1208 3017 1262 3029
rect 1208 2991 1218 3017
rect 1252 2991 1262 3017
rect 1208 2939 1209 2991
rect 1261 2939 1262 2991
rect 1208 2932 1262 2939
rect 1308 3017 1362 3123
rect 1408 3201 1462 3208
rect 1408 3149 1409 3201
rect 1461 3149 1462 3201
rect 1408 3123 1418 3149
rect 1452 3123 1462 3149
rect 1408 3111 1462 3123
rect 1508 3157 1562 3263
rect 1608 3297 1662 3309
rect 1608 3271 1618 3297
rect 1652 3271 1662 3297
rect 1608 3219 1609 3271
rect 1661 3219 1662 3271
rect 1608 3212 1662 3219
rect 1708 3297 1762 3403
rect 1808 3481 1862 3488
rect 1808 3429 1809 3481
rect 1861 3429 1862 3481
rect 1808 3403 1818 3429
rect 1852 3403 1862 3429
rect 1808 3391 1862 3403
rect 1908 3437 1962 3543
rect 2008 3577 2062 3589
rect 2008 3551 2018 3577
rect 2052 3551 2062 3577
rect 2008 3499 2009 3551
rect 2061 3499 2062 3551
rect 2008 3492 2062 3499
rect 2108 3577 2162 3773
rect 2208 3851 2262 3858
rect 2208 3799 2209 3851
rect 2261 3799 2262 3851
rect 2208 3773 2218 3799
rect 2252 3773 2262 3799
rect 2208 3761 2262 3773
rect 2308 3807 2362 3913
rect 2408 3947 2462 3959
rect 2408 3921 2418 3947
rect 2452 3921 2462 3947
rect 2408 3869 2409 3921
rect 2461 3869 2462 3921
rect 2408 3862 2462 3869
rect 2508 3947 2562 4053
rect 2608 4131 2662 4138
rect 2608 4079 2609 4131
rect 2661 4079 2662 4131
rect 2608 4053 2618 4079
rect 2652 4053 2662 4079
rect 2608 4041 2662 4053
rect 2708 4087 2762 4193
rect 2808 4227 2862 4239
rect 2808 4201 2818 4227
rect 2852 4201 2862 4227
rect 2808 4149 2809 4201
rect 2861 4149 2862 4201
rect 2808 4142 2862 4149
rect 2908 4227 2962 4333
rect 3008 4411 3062 4418
rect 3008 4359 3009 4411
rect 3061 4359 3062 4411
rect 3008 4333 3018 4359
rect 3052 4333 3062 4359
rect 3008 4321 3062 4333
rect 3108 4367 3162 4473
rect 3208 4507 3262 4519
rect 3208 4481 3218 4507
rect 3252 4481 3262 4507
rect 3208 4429 3209 4481
rect 3261 4429 3262 4481
rect 3208 4422 3262 4429
rect 3308 4507 3362 4613
rect 3408 4691 3462 4698
rect 3408 4639 3409 4691
rect 3461 4639 3462 4691
rect 3408 4613 3418 4639
rect 3452 4613 3462 4639
rect 3408 4601 3462 4613
rect 3508 4647 3562 4753
rect 3608 4787 3662 4799
rect 3608 4761 3618 4787
rect 3652 4761 3662 4787
rect 3608 4709 3609 4761
rect 3661 4709 3662 4761
rect 3608 4702 3662 4709
rect 3708 4787 3762 4960
rect 3802 4919 3868 4920
rect 3802 4867 3809 4919
rect 3861 4867 3868 4919
rect 3802 4866 3868 4867
rect 3708 4753 3718 4787
rect 3752 4753 3762 4787
rect 3508 4613 3518 4647
rect 3552 4613 3562 4647
rect 3308 4473 3318 4507
rect 3352 4473 3362 4507
rect 3108 4333 3118 4367
rect 3152 4333 3162 4367
rect 2908 4193 2918 4227
rect 2952 4193 2962 4227
rect 2708 4053 2718 4087
rect 2752 4053 2762 4087
rect 2508 3913 2518 3947
rect 2552 3913 2562 3947
rect 2308 3773 2318 3807
rect 2352 3773 2362 3807
rect 2202 3709 2268 3710
rect 2202 3657 2209 3709
rect 2261 3657 2268 3709
rect 2202 3656 2268 3657
rect 2108 3543 2118 3577
rect 2152 3543 2162 3577
rect 1908 3403 1918 3437
rect 1952 3403 1962 3437
rect 1708 3263 1718 3297
rect 1752 3263 1762 3297
rect 1508 3123 1518 3157
rect 1552 3123 1562 3157
rect 1308 2983 1318 3017
rect 1352 2983 1362 3017
rect 1108 2843 1118 2877
rect 1152 2843 1162 2877
rect 908 2703 918 2737
rect 952 2703 962 2737
rect 708 2563 718 2597
rect 752 2563 762 2597
rect 602 2499 668 2500
rect 602 2447 609 2499
rect 661 2447 668 2499
rect 602 2446 668 2447
rect 508 2333 518 2367
rect 552 2333 562 2367
rect 308 2193 318 2227
rect 352 2193 362 2227
rect 108 2053 118 2087
rect 152 2053 162 2087
rect 8 1947 62 1959
rect 8 1921 18 1947
rect 52 1921 62 1947
rect 8 1869 9 1921
rect 61 1869 62 1921
rect 8 1862 62 1869
rect 108 1947 162 2053
rect 208 2131 262 2138
rect 208 2079 209 2131
rect 261 2079 262 2131
rect 208 2053 218 2079
rect 252 2053 262 2079
rect 208 2041 262 2053
rect 308 2087 362 2193
rect 408 2227 462 2239
rect 408 2201 418 2227
rect 452 2201 462 2227
rect 408 2149 409 2201
rect 461 2149 462 2201
rect 408 2142 462 2149
rect 508 2227 562 2333
rect 608 2411 662 2418
rect 608 2359 609 2411
rect 661 2359 662 2411
rect 608 2333 618 2359
rect 652 2333 662 2359
rect 608 2321 662 2333
rect 708 2367 762 2563
rect 808 2597 862 2609
rect 808 2571 818 2597
rect 852 2571 862 2597
rect 808 2519 809 2571
rect 861 2519 862 2571
rect 808 2512 862 2519
rect 908 2597 962 2703
rect 1008 2781 1062 2788
rect 1008 2729 1009 2781
rect 1061 2729 1062 2781
rect 1008 2703 1018 2729
rect 1052 2703 1062 2729
rect 1008 2691 1062 2703
rect 1108 2737 1162 2843
rect 1208 2877 1262 2889
rect 1208 2851 1218 2877
rect 1252 2851 1262 2877
rect 1208 2799 1209 2851
rect 1261 2799 1262 2851
rect 1208 2792 1262 2799
rect 1308 2877 1362 2983
rect 1408 3061 1462 3068
rect 1408 3009 1409 3061
rect 1461 3009 1462 3061
rect 1408 2983 1418 3009
rect 1452 2983 1462 3009
rect 1408 2971 1462 2983
rect 1508 3017 1562 3123
rect 1608 3157 1662 3169
rect 1608 3131 1618 3157
rect 1652 3131 1662 3157
rect 1608 3079 1609 3131
rect 1661 3079 1662 3131
rect 1608 3072 1662 3079
rect 1708 3157 1762 3263
rect 1808 3341 1862 3348
rect 1808 3289 1809 3341
rect 1861 3289 1862 3341
rect 1808 3263 1818 3289
rect 1852 3263 1862 3289
rect 1808 3251 1862 3263
rect 1908 3297 1962 3403
rect 2008 3437 2062 3449
rect 2008 3411 2018 3437
rect 2052 3411 2062 3437
rect 2008 3359 2009 3411
rect 2061 3359 2062 3411
rect 2008 3352 2062 3359
rect 2108 3437 2162 3543
rect 2208 3621 2262 3628
rect 2208 3569 2209 3621
rect 2261 3569 2262 3621
rect 2208 3543 2218 3569
rect 2252 3543 2262 3569
rect 2208 3531 2262 3543
rect 2308 3577 2362 3773
rect 2408 3807 2462 3819
rect 2408 3781 2418 3807
rect 2452 3781 2462 3807
rect 2408 3729 2409 3781
rect 2461 3729 2462 3781
rect 2408 3722 2462 3729
rect 2508 3807 2562 3913
rect 2608 3991 2662 3998
rect 2608 3939 2609 3991
rect 2661 3939 2662 3991
rect 2608 3913 2618 3939
rect 2652 3913 2662 3939
rect 2608 3901 2662 3913
rect 2708 3947 2762 4053
rect 2808 4087 2862 4099
rect 2808 4061 2818 4087
rect 2852 4061 2862 4087
rect 2808 4009 2809 4061
rect 2861 4009 2862 4061
rect 2808 4002 2862 4009
rect 2908 4087 2962 4193
rect 3008 4271 3062 4278
rect 3008 4219 3009 4271
rect 3061 4219 3062 4271
rect 3008 4193 3018 4219
rect 3052 4193 3062 4219
rect 3008 4181 3062 4193
rect 3108 4227 3162 4333
rect 3208 4367 3262 4379
rect 3208 4341 3218 4367
rect 3252 4341 3262 4367
rect 3208 4289 3209 4341
rect 3261 4289 3262 4341
rect 3208 4282 3262 4289
rect 3308 4367 3362 4473
rect 3408 4551 3462 4558
rect 3408 4499 3409 4551
rect 3461 4499 3462 4551
rect 3408 4473 3418 4499
rect 3452 4473 3462 4499
rect 3408 4461 3462 4473
rect 3508 4507 3562 4613
rect 3608 4647 3662 4659
rect 3608 4621 3618 4647
rect 3652 4621 3662 4647
rect 3608 4569 3609 4621
rect 3661 4569 3662 4621
rect 3608 4562 3662 4569
rect 3708 4647 3762 4753
rect 3808 4831 3862 4838
rect 3808 4779 3809 4831
rect 3861 4779 3862 4831
rect 3808 4753 3818 4779
rect 3852 4753 3862 4779
rect 3808 4741 3862 4753
rect 3908 4787 3962 4960
rect 4002 4903 4068 4904
rect 4002 4851 4009 4903
rect 4061 4851 4068 4903
rect 4002 4850 4068 4851
rect 3908 4753 3918 4787
rect 3952 4753 3962 4787
rect 3708 4613 3718 4647
rect 3752 4613 3762 4647
rect 3508 4473 3518 4507
rect 3552 4473 3562 4507
rect 3308 4333 3318 4367
rect 3352 4333 3362 4367
rect 3108 4193 3118 4227
rect 3152 4193 3162 4227
rect 2908 4053 2918 4087
rect 2952 4053 2962 4087
rect 2708 3913 2718 3947
rect 2752 3913 2762 3947
rect 2508 3773 2518 3807
rect 2552 3773 2562 3807
rect 2402 3693 2468 3694
rect 2402 3641 2409 3693
rect 2461 3641 2468 3693
rect 2402 3640 2468 3641
rect 2308 3543 2318 3577
rect 2352 3543 2362 3577
rect 2108 3403 2118 3437
rect 2152 3403 2162 3437
rect 1908 3263 1918 3297
rect 1952 3263 1962 3297
rect 1708 3123 1718 3157
rect 1752 3123 1762 3157
rect 1508 2983 1518 3017
rect 1552 2983 1562 3017
rect 1308 2843 1318 2877
rect 1352 2843 1362 2877
rect 1108 2703 1118 2737
rect 1152 2703 1162 2737
rect 908 2563 918 2597
rect 952 2563 962 2597
rect 802 2483 868 2484
rect 802 2431 809 2483
rect 861 2431 868 2483
rect 802 2430 868 2431
rect 708 2333 718 2367
rect 752 2333 762 2367
rect 508 2193 518 2227
rect 552 2193 562 2227
rect 308 2053 318 2087
rect 352 2053 362 2087
rect 108 1913 118 1947
rect 152 1913 162 1947
rect 8 1807 62 1819
rect 8 1781 18 1807
rect 52 1781 62 1807
rect 8 1729 9 1781
rect 61 1729 62 1781
rect 8 1722 62 1729
rect 108 1807 162 1913
rect 208 1991 262 1998
rect 208 1939 209 1991
rect 261 1939 262 1991
rect 208 1913 218 1939
rect 252 1913 262 1939
rect 208 1901 262 1913
rect 308 1947 362 2053
rect 408 2087 462 2099
rect 408 2061 418 2087
rect 452 2061 462 2087
rect 408 2009 409 2061
rect 461 2009 462 2061
rect 408 2002 462 2009
rect 508 2087 562 2193
rect 608 2271 662 2278
rect 608 2219 609 2271
rect 661 2219 662 2271
rect 608 2193 618 2219
rect 652 2193 662 2219
rect 608 2181 662 2193
rect 708 2227 762 2333
rect 808 2367 862 2379
rect 808 2341 818 2367
rect 852 2341 862 2367
rect 808 2289 809 2341
rect 861 2289 862 2341
rect 808 2282 862 2289
rect 908 2367 962 2563
rect 1008 2641 1062 2648
rect 1008 2589 1009 2641
rect 1061 2589 1062 2641
rect 1008 2563 1018 2589
rect 1052 2563 1062 2589
rect 1008 2551 1062 2563
rect 1108 2597 1162 2703
rect 1208 2737 1262 2749
rect 1208 2711 1218 2737
rect 1252 2711 1262 2737
rect 1208 2659 1209 2711
rect 1261 2659 1262 2711
rect 1208 2652 1262 2659
rect 1308 2737 1362 2843
rect 1408 2921 1462 2928
rect 1408 2869 1409 2921
rect 1461 2869 1462 2921
rect 1408 2843 1418 2869
rect 1452 2843 1462 2869
rect 1408 2831 1462 2843
rect 1508 2877 1562 2983
rect 1608 3017 1662 3029
rect 1608 2991 1618 3017
rect 1652 2991 1662 3017
rect 1608 2939 1609 2991
rect 1661 2939 1662 2991
rect 1608 2932 1662 2939
rect 1708 3017 1762 3123
rect 1808 3201 1862 3208
rect 1808 3149 1809 3201
rect 1861 3149 1862 3201
rect 1808 3123 1818 3149
rect 1852 3123 1862 3149
rect 1808 3111 1862 3123
rect 1908 3157 1962 3263
rect 2008 3297 2062 3309
rect 2008 3271 2018 3297
rect 2052 3271 2062 3297
rect 2008 3219 2009 3271
rect 2061 3219 2062 3271
rect 2008 3212 2062 3219
rect 2108 3297 2162 3403
rect 2208 3481 2262 3488
rect 2208 3429 2209 3481
rect 2261 3429 2262 3481
rect 2208 3403 2218 3429
rect 2252 3403 2262 3429
rect 2208 3391 2262 3403
rect 2308 3437 2362 3543
rect 2408 3577 2462 3589
rect 2408 3551 2418 3577
rect 2452 3551 2462 3577
rect 2408 3499 2409 3551
rect 2461 3499 2462 3551
rect 2408 3492 2462 3499
rect 2508 3577 2562 3773
rect 2608 3851 2662 3858
rect 2608 3799 2609 3851
rect 2661 3799 2662 3851
rect 2608 3773 2618 3799
rect 2652 3773 2662 3799
rect 2608 3761 2662 3773
rect 2708 3807 2762 3913
rect 2808 3947 2862 3959
rect 2808 3921 2818 3947
rect 2852 3921 2862 3947
rect 2808 3869 2809 3921
rect 2861 3869 2862 3921
rect 2808 3862 2862 3869
rect 2908 3947 2962 4053
rect 3008 4131 3062 4138
rect 3008 4079 3009 4131
rect 3061 4079 3062 4131
rect 3008 4053 3018 4079
rect 3052 4053 3062 4079
rect 3008 4041 3062 4053
rect 3108 4087 3162 4193
rect 3208 4227 3262 4239
rect 3208 4201 3218 4227
rect 3252 4201 3262 4227
rect 3208 4149 3209 4201
rect 3261 4149 3262 4201
rect 3208 4142 3262 4149
rect 3308 4227 3362 4333
rect 3408 4411 3462 4418
rect 3408 4359 3409 4411
rect 3461 4359 3462 4411
rect 3408 4333 3418 4359
rect 3452 4333 3462 4359
rect 3408 4321 3462 4333
rect 3508 4367 3562 4473
rect 3608 4507 3662 4519
rect 3608 4481 3618 4507
rect 3652 4481 3662 4507
rect 3608 4429 3609 4481
rect 3661 4429 3662 4481
rect 3608 4422 3662 4429
rect 3708 4507 3762 4613
rect 3808 4691 3862 4698
rect 3808 4639 3809 4691
rect 3861 4639 3862 4691
rect 3808 4613 3818 4639
rect 3852 4613 3862 4639
rect 3808 4601 3862 4613
rect 3908 4647 3962 4753
rect 4008 4787 4062 4799
rect 4008 4761 4018 4787
rect 4052 4761 4062 4787
rect 4008 4709 4009 4761
rect 4061 4709 4062 4761
rect 4008 4702 4062 4709
rect 4108 4787 4162 4960
rect 4202 4919 4268 4920
rect 4202 4867 4209 4919
rect 4261 4867 4268 4919
rect 4202 4866 4268 4867
rect 4108 4753 4118 4787
rect 4152 4753 4162 4787
rect 3908 4613 3918 4647
rect 3952 4613 3962 4647
rect 3708 4473 3718 4507
rect 3752 4473 3762 4507
rect 3508 4333 3518 4367
rect 3552 4333 3562 4367
rect 3308 4193 3318 4227
rect 3352 4193 3362 4227
rect 3108 4053 3118 4087
rect 3152 4053 3162 4087
rect 2908 3913 2918 3947
rect 2952 3913 2962 3947
rect 2708 3773 2718 3807
rect 2752 3773 2762 3807
rect 2602 3709 2668 3710
rect 2602 3657 2609 3709
rect 2661 3657 2668 3709
rect 2602 3656 2668 3657
rect 2508 3543 2518 3577
rect 2552 3543 2562 3577
rect 2308 3403 2318 3437
rect 2352 3403 2362 3437
rect 2108 3263 2118 3297
rect 2152 3263 2162 3297
rect 1908 3123 1918 3157
rect 1952 3123 1962 3157
rect 1708 2983 1718 3017
rect 1752 2983 1762 3017
rect 1508 2843 1518 2877
rect 1552 2843 1562 2877
rect 1308 2703 1318 2737
rect 1352 2703 1362 2737
rect 1108 2563 1118 2597
rect 1152 2563 1162 2597
rect 1002 2499 1068 2500
rect 1002 2447 1009 2499
rect 1061 2447 1068 2499
rect 1002 2446 1068 2447
rect 908 2333 918 2367
rect 952 2333 962 2367
rect 708 2193 718 2227
rect 752 2193 762 2227
rect 508 2053 518 2087
rect 552 2053 562 2087
rect 308 1913 318 1947
rect 352 1913 362 1947
rect 108 1773 118 1807
rect 152 1773 162 1807
rect 8 1667 62 1679
rect 8 1641 18 1667
rect 52 1641 62 1667
rect 8 1589 9 1641
rect 61 1589 62 1641
rect 8 1582 62 1589
rect 108 1667 162 1773
rect 208 1851 262 1858
rect 208 1799 209 1851
rect 261 1799 262 1851
rect 208 1773 218 1799
rect 252 1773 262 1799
rect 208 1761 262 1773
rect 308 1807 362 1913
rect 408 1947 462 1959
rect 408 1921 418 1947
rect 452 1921 462 1947
rect 408 1869 409 1921
rect 461 1869 462 1921
rect 408 1862 462 1869
rect 508 1947 562 2053
rect 608 2131 662 2138
rect 608 2079 609 2131
rect 661 2079 662 2131
rect 608 2053 618 2079
rect 652 2053 662 2079
rect 608 2041 662 2053
rect 708 2087 762 2193
rect 808 2227 862 2239
rect 808 2201 818 2227
rect 852 2201 862 2227
rect 808 2149 809 2201
rect 861 2149 862 2201
rect 808 2142 862 2149
rect 908 2227 962 2333
rect 1008 2411 1062 2418
rect 1008 2359 1009 2411
rect 1061 2359 1062 2411
rect 1008 2333 1018 2359
rect 1052 2333 1062 2359
rect 1008 2321 1062 2333
rect 1108 2367 1162 2563
rect 1208 2597 1262 2609
rect 1208 2571 1218 2597
rect 1252 2571 1262 2597
rect 1208 2519 1209 2571
rect 1261 2519 1262 2571
rect 1208 2512 1262 2519
rect 1308 2597 1362 2703
rect 1408 2781 1462 2788
rect 1408 2729 1409 2781
rect 1461 2729 1462 2781
rect 1408 2703 1418 2729
rect 1452 2703 1462 2729
rect 1408 2691 1462 2703
rect 1508 2737 1562 2843
rect 1608 2877 1662 2889
rect 1608 2851 1618 2877
rect 1652 2851 1662 2877
rect 1608 2799 1609 2851
rect 1661 2799 1662 2851
rect 1608 2792 1662 2799
rect 1708 2877 1762 2983
rect 1808 3061 1862 3068
rect 1808 3009 1809 3061
rect 1861 3009 1862 3061
rect 1808 2983 1818 3009
rect 1852 2983 1862 3009
rect 1808 2971 1862 2983
rect 1908 3017 1962 3123
rect 2008 3157 2062 3169
rect 2008 3131 2018 3157
rect 2052 3131 2062 3157
rect 2008 3079 2009 3131
rect 2061 3079 2062 3131
rect 2008 3072 2062 3079
rect 2108 3157 2162 3263
rect 2208 3341 2262 3348
rect 2208 3289 2209 3341
rect 2261 3289 2262 3341
rect 2208 3263 2218 3289
rect 2252 3263 2262 3289
rect 2208 3251 2262 3263
rect 2308 3297 2362 3403
rect 2408 3437 2462 3449
rect 2408 3411 2418 3437
rect 2452 3411 2462 3437
rect 2408 3359 2409 3411
rect 2461 3359 2462 3411
rect 2408 3352 2462 3359
rect 2508 3437 2562 3543
rect 2608 3621 2662 3628
rect 2608 3569 2609 3621
rect 2661 3569 2662 3621
rect 2608 3543 2618 3569
rect 2652 3543 2662 3569
rect 2608 3531 2662 3543
rect 2708 3577 2762 3773
rect 2808 3807 2862 3819
rect 2808 3781 2818 3807
rect 2852 3781 2862 3807
rect 2808 3729 2809 3781
rect 2861 3729 2862 3781
rect 2808 3722 2862 3729
rect 2908 3807 2962 3913
rect 3008 3991 3062 3998
rect 3008 3939 3009 3991
rect 3061 3939 3062 3991
rect 3008 3913 3018 3939
rect 3052 3913 3062 3939
rect 3008 3901 3062 3913
rect 3108 3947 3162 4053
rect 3208 4087 3262 4099
rect 3208 4061 3218 4087
rect 3252 4061 3262 4087
rect 3208 4009 3209 4061
rect 3261 4009 3262 4061
rect 3208 4002 3262 4009
rect 3308 4087 3362 4193
rect 3408 4271 3462 4278
rect 3408 4219 3409 4271
rect 3461 4219 3462 4271
rect 3408 4193 3418 4219
rect 3452 4193 3462 4219
rect 3408 4181 3462 4193
rect 3508 4227 3562 4333
rect 3608 4367 3662 4379
rect 3608 4341 3618 4367
rect 3652 4341 3662 4367
rect 3608 4289 3609 4341
rect 3661 4289 3662 4341
rect 3608 4282 3662 4289
rect 3708 4367 3762 4473
rect 3808 4551 3862 4558
rect 3808 4499 3809 4551
rect 3861 4499 3862 4551
rect 3808 4473 3818 4499
rect 3852 4473 3862 4499
rect 3808 4461 3862 4473
rect 3908 4507 3962 4613
rect 4008 4647 4062 4659
rect 4008 4621 4018 4647
rect 4052 4621 4062 4647
rect 4008 4569 4009 4621
rect 4061 4569 4062 4621
rect 4008 4562 4062 4569
rect 4108 4647 4162 4753
rect 4208 4831 4262 4838
rect 4208 4779 4209 4831
rect 4261 4779 4262 4831
rect 4208 4753 4218 4779
rect 4252 4753 4262 4779
rect 4208 4741 4262 4753
rect 4308 4787 4362 4960
rect 4402 4903 4468 4904
rect 4402 4851 4409 4903
rect 4461 4851 4468 4903
rect 4402 4850 4468 4851
rect 4308 4753 4318 4787
rect 4352 4753 4362 4787
rect 4108 4613 4118 4647
rect 4152 4613 4162 4647
rect 3908 4473 3918 4507
rect 3952 4473 3962 4507
rect 3708 4333 3718 4367
rect 3752 4333 3762 4367
rect 3508 4193 3518 4227
rect 3552 4193 3562 4227
rect 3308 4053 3318 4087
rect 3352 4053 3362 4087
rect 3108 3913 3118 3947
rect 3152 3913 3162 3947
rect 2908 3773 2918 3807
rect 2952 3773 2962 3807
rect 2802 3693 2868 3694
rect 2802 3641 2809 3693
rect 2861 3641 2868 3693
rect 2802 3640 2868 3641
rect 2708 3543 2718 3577
rect 2752 3543 2762 3577
rect 2508 3403 2518 3437
rect 2552 3403 2562 3437
rect 2308 3263 2318 3297
rect 2352 3263 2362 3297
rect 2108 3123 2118 3157
rect 2152 3123 2162 3157
rect 1908 2983 1918 3017
rect 1952 2983 1962 3017
rect 1708 2843 1718 2877
rect 1752 2843 1762 2877
rect 1508 2703 1518 2737
rect 1552 2703 1562 2737
rect 1308 2563 1318 2597
rect 1352 2563 1362 2597
rect 1202 2483 1268 2484
rect 1202 2431 1209 2483
rect 1261 2431 1268 2483
rect 1202 2430 1268 2431
rect 1108 2333 1118 2367
rect 1152 2333 1162 2367
rect 908 2193 918 2227
rect 952 2193 962 2227
rect 708 2053 718 2087
rect 752 2053 762 2087
rect 508 1913 518 1947
rect 552 1913 562 1947
rect 308 1773 318 1807
rect 352 1773 362 1807
rect 108 1633 118 1667
rect 152 1633 162 1667
rect 8 1527 62 1539
rect 8 1501 18 1527
rect 52 1501 62 1527
rect 8 1449 9 1501
rect 61 1449 62 1501
rect 8 1442 62 1449
rect 108 1527 162 1633
rect 208 1711 262 1718
rect 208 1659 209 1711
rect 261 1659 262 1711
rect 208 1633 218 1659
rect 252 1633 262 1659
rect 208 1621 262 1633
rect 308 1667 362 1773
rect 408 1807 462 1819
rect 408 1781 418 1807
rect 452 1781 462 1807
rect 408 1729 409 1781
rect 461 1729 462 1781
rect 408 1722 462 1729
rect 508 1807 562 1913
rect 608 1991 662 1998
rect 608 1939 609 1991
rect 661 1939 662 1991
rect 608 1913 618 1939
rect 652 1913 662 1939
rect 608 1901 662 1913
rect 708 1947 762 2053
rect 808 2087 862 2099
rect 808 2061 818 2087
rect 852 2061 862 2087
rect 808 2009 809 2061
rect 861 2009 862 2061
rect 808 2002 862 2009
rect 908 2087 962 2193
rect 1008 2271 1062 2278
rect 1008 2219 1009 2271
rect 1061 2219 1062 2271
rect 1008 2193 1018 2219
rect 1052 2193 1062 2219
rect 1008 2181 1062 2193
rect 1108 2227 1162 2333
rect 1208 2367 1262 2379
rect 1208 2341 1218 2367
rect 1252 2341 1262 2367
rect 1208 2289 1209 2341
rect 1261 2289 1262 2341
rect 1208 2282 1262 2289
rect 1308 2367 1362 2563
rect 1408 2641 1462 2648
rect 1408 2589 1409 2641
rect 1461 2589 1462 2641
rect 1408 2563 1418 2589
rect 1452 2563 1462 2589
rect 1408 2551 1462 2563
rect 1508 2597 1562 2703
rect 1608 2737 1662 2749
rect 1608 2711 1618 2737
rect 1652 2711 1662 2737
rect 1608 2659 1609 2711
rect 1661 2659 1662 2711
rect 1608 2652 1662 2659
rect 1708 2737 1762 2843
rect 1808 2921 1862 2928
rect 1808 2869 1809 2921
rect 1861 2869 1862 2921
rect 1808 2843 1818 2869
rect 1852 2843 1862 2869
rect 1808 2831 1862 2843
rect 1908 2877 1962 2983
rect 2008 3017 2062 3029
rect 2008 2991 2018 3017
rect 2052 2991 2062 3017
rect 2008 2939 2009 2991
rect 2061 2939 2062 2991
rect 2008 2932 2062 2939
rect 2108 3017 2162 3123
rect 2208 3201 2262 3208
rect 2208 3149 2209 3201
rect 2261 3149 2262 3201
rect 2208 3123 2218 3149
rect 2252 3123 2262 3149
rect 2208 3111 2262 3123
rect 2308 3157 2362 3263
rect 2408 3297 2462 3309
rect 2408 3271 2418 3297
rect 2452 3271 2462 3297
rect 2408 3219 2409 3271
rect 2461 3219 2462 3271
rect 2408 3212 2462 3219
rect 2508 3297 2562 3403
rect 2608 3481 2662 3488
rect 2608 3429 2609 3481
rect 2661 3429 2662 3481
rect 2608 3403 2618 3429
rect 2652 3403 2662 3429
rect 2608 3391 2662 3403
rect 2708 3437 2762 3543
rect 2808 3577 2862 3589
rect 2808 3551 2818 3577
rect 2852 3551 2862 3577
rect 2808 3499 2809 3551
rect 2861 3499 2862 3551
rect 2808 3492 2862 3499
rect 2908 3577 2962 3773
rect 3008 3851 3062 3858
rect 3008 3799 3009 3851
rect 3061 3799 3062 3851
rect 3008 3773 3018 3799
rect 3052 3773 3062 3799
rect 3008 3761 3062 3773
rect 3108 3807 3162 3913
rect 3208 3947 3262 3959
rect 3208 3921 3218 3947
rect 3252 3921 3262 3947
rect 3208 3869 3209 3921
rect 3261 3869 3262 3921
rect 3208 3862 3262 3869
rect 3308 3947 3362 4053
rect 3408 4131 3462 4138
rect 3408 4079 3409 4131
rect 3461 4079 3462 4131
rect 3408 4053 3418 4079
rect 3452 4053 3462 4079
rect 3408 4041 3462 4053
rect 3508 4087 3562 4193
rect 3608 4227 3662 4239
rect 3608 4201 3618 4227
rect 3652 4201 3662 4227
rect 3608 4149 3609 4201
rect 3661 4149 3662 4201
rect 3608 4142 3662 4149
rect 3708 4227 3762 4333
rect 3808 4411 3862 4418
rect 3808 4359 3809 4411
rect 3861 4359 3862 4411
rect 3808 4333 3818 4359
rect 3852 4333 3862 4359
rect 3808 4321 3862 4333
rect 3908 4367 3962 4473
rect 4008 4507 4062 4519
rect 4008 4481 4018 4507
rect 4052 4481 4062 4507
rect 4008 4429 4009 4481
rect 4061 4429 4062 4481
rect 4008 4422 4062 4429
rect 4108 4507 4162 4613
rect 4208 4691 4262 4698
rect 4208 4639 4209 4691
rect 4261 4639 4262 4691
rect 4208 4613 4218 4639
rect 4252 4613 4262 4639
rect 4208 4601 4262 4613
rect 4308 4647 4362 4753
rect 4408 4787 4462 4799
rect 4408 4761 4418 4787
rect 4452 4761 4462 4787
rect 4408 4709 4409 4761
rect 4461 4709 4462 4761
rect 4408 4702 4462 4709
rect 4508 4787 4562 4960
rect 4602 4919 4668 4920
rect 4602 4867 4609 4919
rect 4661 4867 4668 4919
rect 4602 4866 4668 4867
rect 4508 4753 4518 4787
rect 4552 4753 4562 4787
rect 4308 4613 4318 4647
rect 4352 4613 4362 4647
rect 4108 4473 4118 4507
rect 4152 4473 4162 4507
rect 3908 4333 3918 4367
rect 3952 4333 3962 4367
rect 3708 4193 3718 4227
rect 3752 4193 3762 4227
rect 3508 4053 3518 4087
rect 3552 4053 3562 4087
rect 3308 3913 3318 3947
rect 3352 3913 3362 3947
rect 3108 3773 3118 3807
rect 3152 3773 3162 3807
rect 3002 3709 3068 3710
rect 3002 3657 3009 3709
rect 3061 3657 3068 3709
rect 3002 3656 3068 3657
rect 2908 3543 2918 3577
rect 2952 3543 2962 3577
rect 2708 3403 2718 3437
rect 2752 3403 2762 3437
rect 2508 3263 2518 3297
rect 2552 3263 2562 3297
rect 2308 3123 2318 3157
rect 2352 3123 2362 3157
rect 2108 2983 2118 3017
rect 2152 2983 2162 3017
rect 1908 2843 1918 2877
rect 1952 2843 1962 2877
rect 1708 2703 1718 2737
rect 1752 2703 1762 2737
rect 1508 2563 1518 2597
rect 1552 2563 1562 2597
rect 1402 2499 1468 2500
rect 1402 2447 1409 2499
rect 1461 2447 1468 2499
rect 1402 2446 1468 2447
rect 1308 2333 1318 2367
rect 1352 2333 1362 2367
rect 1108 2193 1118 2227
rect 1152 2193 1162 2227
rect 908 2053 918 2087
rect 952 2053 962 2087
rect 708 1913 718 1947
rect 752 1913 762 1947
rect 508 1773 518 1807
rect 552 1773 562 1807
rect 308 1633 318 1667
rect 352 1633 362 1667
rect 108 1493 118 1527
rect 152 1493 162 1527
rect 8 1387 62 1399
rect 8 1361 18 1387
rect 52 1361 62 1387
rect 8 1309 9 1361
rect 61 1309 62 1361
rect 8 1302 62 1309
rect 108 1387 162 1493
rect 208 1571 262 1578
rect 208 1519 209 1571
rect 261 1519 262 1571
rect 208 1493 218 1519
rect 252 1493 262 1519
rect 208 1481 262 1493
rect 308 1527 362 1633
rect 408 1667 462 1679
rect 408 1641 418 1667
rect 452 1641 462 1667
rect 408 1589 409 1641
rect 461 1589 462 1641
rect 408 1582 462 1589
rect 508 1667 562 1773
rect 608 1851 662 1858
rect 608 1799 609 1851
rect 661 1799 662 1851
rect 608 1773 618 1799
rect 652 1773 662 1799
rect 608 1761 662 1773
rect 708 1807 762 1913
rect 808 1947 862 1959
rect 808 1921 818 1947
rect 852 1921 862 1947
rect 808 1869 809 1921
rect 861 1869 862 1921
rect 808 1862 862 1869
rect 908 1947 962 2053
rect 1008 2131 1062 2138
rect 1008 2079 1009 2131
rect 1061 2079 1062 2131
rect 1008 2053 1018 2079
rect 1052 2053 1062 2079
rect 1008 2041 1062 2053
rect 1108 2087 1162 2193
rect 1208 2227 1262 2239
rect 1208 2201 1218 2227
rect 1252 2201 1262 2227
rect 1208 2149 1209 2201
rect 1261 2149 1262 2201
rect 1208 2142 1262 2149
rect 1308 2227 1362 2333
rect 1408 2411 1462 2418
rect 1408 2359 1409 2411
rect 1461 2359 1462 2411
rect 1408 2333 1418 2359
rect 1452 2333 1462 2359
rect 1408 2321 1462 2333
rect 1508 2367 1562 2563
rect 1608 2597 1662 2609
rect 1608 2571 1618 2597
rect 1652 2571 1662 2597
rect 1608 2519 1609 2571
rect 1661 2519 1662 2571
rect 1608 2512 1662 2519
rect 1708 2597 1762 2703
rect 1808 2781 1862 2788
rect 1808 2729 1809 2781
rect 1861 2729 1862 2781
rect 1808 2703 1818 2729
rect 1852 2703 1862 2729
rect 1808 2691 1862 2703
rect 1908 2737 1962 2843
rect 2008 2877 2062 2889
rect 2008 2851 2018 2877
rect 2052 2851 2062 2877
rect 2008 2799 2009 2851
rect 2061 2799 2062 2851
rect 2008 2792 2062 2799
rect 2108 2877 2162 2983
rect 2208 3061 2262 3068
rect 2208 3009 2209 3061
rect 2261 3009 2262 3061
rect 2208 2983 2218 3009
rect 2252 2983 2262 3009
rect 2208 2971 2262 2983
rect 2308 3017 2362 3123
rect 2408 3157 2462 3169
rect 2408 3131 2418 3157
rect 2452 3131 2462 3157
rect 2408 3079 2409 3131
rect 2461 3079 2462 3131
rect 2408 3072 2462 3079
rect 2508 3157 2562 3263
rect 2608 3341 2662 3348
rect 2608 3289 2609 3341
rect 2661 3289 2662 3341
rect 2608 3263 2618 3289
rect 2652 3263 2662 3289
rect 2608 3251 2662 3263
rect 2708 3297 2762 3403
rect 2808 3437 2862 3449
rect 2808 3411 2818 3437
rect 2852 3411 2862 3437
rect 2808 3359 2809 3411
rect 2861 3359 2862 3411
rect 2808 3352 2862 3359
rect 2908 3437 2962 3543
rect 3008 3621 3062 3628
rect 3008 3569 3009 3621
rect 3061 3569 3062 3621
rect 3008 3543 3018 3569
rect 3052 3543 3062 3569
rect 3008 3531 3062 3543
rect 3108 3577 3162 3773
rect 3208 3807 3262 3819
rect 3208 3781 3218 3807
rect 3252 3781 3262 3807
rect 3208 3729 3209 3781
rect 3261 3729 3262 3781
rect 3208 3722 3262 3729
rect 3308 3807 3362 3913
rect 3408 3991 3462 3998
rect 3408 3939 3409 3991
rect 3461 3939 3462 3991
rect 3408 3913 3418 3939
rect 3452 3913 3462 3939
rect 3408 3901 3462 3913
rect 3508 3947 3562 4053
rect 3608 4087 3662 4099
rect 3608 4061 3618 4087
rect 3652 4061 3662 4087
rect 3608 4009 3609 4061
rect 3661 4009 3662 4061
rect 3608 4002 3662 4009
rect 3708 4087 3762 4193
rect 3808 4271 3862 4278
rect 3808 4219 3809 4271
rect 3861 4219 3862 4271
rect 3808 4193 3818 4219
rect 3852 4193 3862 4219
rect 3808 4181 3862 4193
rect 3908 4227 3962 4333
rect 4008 4367 4062 4379
rect 4008 4341 4018 4367
rect 4052 4341 4062 4367
rect 4008 4289 4009 4341
rect 4061 4289 4062 4341
rect 4008 4282 4062 4289
rect 4108 4367 4162 4473
rect 4208 4551 4262 4558
rect 4208 4499 4209 4551
rect 4261 4499 4262 4551
rect 4208 4473 4218 4499
rect 4252 4473 4262 4499
rect 4208 4461 4262 4473
rect 4308 4507 4362 4613
rect 4408 4647 4462 4659
rect 4408 4621 4418 4647
rect 4452 4621 4462 4647
rect 4408 4569 4409 4621
rect 4461 4569 4462 4621
rect 4408 4562 4462 4569
rect 4508 4647 4562 4753
rect 4608 4831 4662 4838
rect 4608 4779 4609 4831
rect 4661 4779 4662 4831
rect 4608 4753 4618 4779
rect 4652 4753 4662 4779
rect 4608 4741 4662 4753
rect 4708 4787 4762 4960
rect 4802 4903 4868 4904
rect 4802 4851 4809 4903
rect 4861 4851 4868 4903
rect 4802 4850 4868 4851
rect 4708 4753 4718 4787
rect 4752 4753 4762 4787
rect 4508 4613 4518 4647
rect 4552 4613 4562 4647
rect 4308 4473 4318 4507
rect 4352 4473 4362 4507
rect 4108 4333 4118 4367
rect 4152 4333 4162 4367
rect 3908 4193 3918 4227
rect 3952 4193 3962 4227
rect 3708 4053 3718 4087
rect 3752 4053 3762 4087
rect 3508 3913 3518 3947
rect 3552 3913 3562 3947
rect 3308 3773 3318 3807
rect 3352 3773 3362 3807
rect 3202 3693 3268 3694
rect 3202 3641 3209 3693
rect 3261 3641 3268 3693
rect 3202 3640 3268 3641
rect 3108 3543 3118 3577
rect 3152 3543 3162 3577
rect 2908 3403 2918 3437
rect 2952 3403 2962 3437
rect 2708 3263 2718 3297
rect 2752 3263 2762 3297
rect 2508 3123 2518 3157
rect 2552 3123 2562 3157
rect 2308 2983 2318 3017
rect 2352 2983 2362 3017
rect 2108 2843 2118 2877
rect 2152 2843 2162 2877
rect 1908 2703 1918 2737
rect 1952 2703 1962 2737
rect 1708 2563 1718 2597
rect 1752 2563 1762 2597
rect 1602 2483 1668 2484
rect 1602 2431 1609 2483
rect 1661 2431 1668 2483
rect 1602 2430 1668 2431
rect 1508 2333 1518 2367
rect 1552 2333 1562 2367
rect 1308 2193 1318 2227
rect 1352 2193 1362 2227
rect 1108 2053 1118 2087
rect 1152 2053 1162 2087
rect 908 1913 918 1947
rect 952 1913 962 1947
rect 708 1773 718 1807
rect 752 1773 762 1807
rect 508 1633 518 1667
rect 552 1633 562 1667
rect 308 1493 318 1527
rect 352 1493 362 1527
rect 108 1353 118 1387
rect 152 1353 162 1387
rect 2 1273 68 1274
rect 2 1221 9 1273
rect 61 1221 68 1273
rect 2 1220 68 1221
rect 8 1157 62 1169
rect 8 1131 18 1157
rect 52 1131 62 1157
rect 8 1079 9 1131
rect 61 1079 62 1131
rect 8 1072 62 1079
rect 108 1157 162 1353
rect 208 1431 262 1438
rect 208 1379 209 1431
rect 261 1379 262 1431
rect 208 1353 218 1379
rect 252 1353 262 1379
rect 208 1341 262 1353
rect 308 1387 362 1493
rect 408 1527 462 1539
rect 408 1501 418 1527
rect 452 1501 462 1527
rect 408 1449 409 1501
rect 461 1449 462 1501
rect 408 1442 462 1449
rect 508 1527 562 1633
rect 608 1711 662 1718
rect 608 1659 609 1711
rect 661 1659 662 1711
rect 608 1633 618 1659
rect 652 1633 662 1659
rect 608 1621 662 1633
rect 708 1667 762 1773
rect 808 1807 862 1819
rect 808 1781 818 1807
rect 852 1781 862 1807
rect 808 1729 809 1781
rect 861 1729 862 1781
rect 808 1722 862 1729
rect 908 1807 962 1913
rect 1008 1991 1062 1998
rect 1008 1939 1009 1991
rect 1061 1939 1062 1991
rect 1008 1913 1018 1939
rect 1052 1913 1062 1939
rect 1008 1901 1062 1913
rect 1108 1947 1162 2053
rect 1208 2087 1262 2099
rect 1208 2061 1218 2087
rect 1252 2061 1262 2087
rect 1208 2009 1209 2061
rect 1261 2009 1262 2061
rect 1208 2002 1262 2009
rect 1308 2087 1362 2193
rect 1408 2271 1462 2278
rect 1408 2219 1409 2271
rect 1461 2219 1462 2271
rect 1408 2193 1418 2219
rect 1452 2193 1462 2219
rect 1408 2181 1462 2193
rect 1508 2227 1562 2333
rect 1608 2367 1662 2379
rect 1608 2341 1618 2367
rect 1652 2341 1662 2367
rect 1608 2289 1609 2341
rect 1661 2289 1662 2341
rect 1608 2282 1662 2289
rect 1708 2367 1762 2563
rect 1808 2641 1862 2648
rect 1808 2589 1809 2641
rect 1861 2589 1862 2641
rect 1808 2563 1818 2589
rect 1852 2563 1862 2589
rect 1808 2551 1862 2563
rect 1908 2597 1962 2703
rect 2008 2737 2062 2749
rect 2008 2711 2018 2737
rect 2052 2711 2062 2737
rect 2008 2659 2009 2711
rect 2061 2659 2062 2711
rect 2008 2652 2062 2659
rect 2108 2737 2162 2843
rect 2208 2921 2262 2928
rect 2208 2869 2209 2921
rect 2261 2869 2262 2921
rect 2208 2843 2218 2869
rect 2252 2843 2262 2869
rect 2208 2831 2262 2843
rect 2308 2877 2362 2983
rect 2408 3017 2462 3029
rect 2408 2991 2418 3017
rect 2452 2991 2462 3017
rect 2408 2939 2409 2991
rect 2461 2939 2462 2991
rect 2408 2932 2462 2939
rect 2508 3017 2562 3123
rect 2608 3201 2662 3208
rect 2608 3149 2609 3201
rect 2661 3149 2662 3201
rect 2608 3123 2618 3149
rect 2652 3123 2662 3149
rect 2608 3111 2662 3123
rect 2708 3157 2762 3263
rect 2808 3297 2862 3309
rect 2808 3271 2818 3297
rect 2852 3271 2862 3297
rect 2808 3219 2809 3271
rect 2861 3219 2862 3271
rect 2808 3212 2862 3219
rect 2908 3297 2962 3403
rect 3008 3481 3062 3488
rect 3008 3429 3009 3481
rect 3061 3429 3062 3481
rect 3008 3403 3018 3429
rect 3052 3403 3062 3429
rect 3008 3391 3062 3403
rect 3108 3437 3162 3543
rect 3208 3577 3262 3589
rect 3208 3551 3218 3577
rect 3252 3551 3262 3577
rect 3208 3499 3209 3551
rect 3261 3499 3262 3551
rect 3208 3492 3262 3499
rect 3308 3577 3362 3773
rect 3408 3851 3462 3858
rect 3408 3799 3409 3851
rect 3461 3799 3462 3851
rect 3408 3773 3418 3799
rect 3452 3773 3462 3799
rect 3408 3761 3462 3773
rect 3508 3807 3562 3913
rect 3608 3947 3662 3959
rect 3608 3921 3618 3947
rect 3652 3921 3662 3947
rect 3608 3869 3609 3921
rect 3661 3869 3662 3921
rect 3608 3862 3662 3869
rect 3708 3947 3762 4053
rect 3808 4131 3862 4138
rect 3808 4079 3809 4131
rect 3861 4079 3862 4131
rect 3808 4053 3818 4079
rect 3852 4053 3862 4079
rect 3808 4041 3862 4053
rect 3908 4087 3962 4193
rect 4008 4227 4062 4239
rect 4008 4201 4018 4227
rect 4052 4201 4062 4227
rect 4008 4149 4009 4201
rect 4061 4149 4062 4201
rect 4008 4142 4062 4149
rect 4108 4227 4162 4333
rect 4208 4411 4262 4418
rect 4208 4359 4209 4411
rect 4261 4359 4262 4411
rect 4208 4333 4218 4359
rect 4252 4333 4262 4359
rect 4208 4321 4262 4333
rect 4308 4367 4362 4473
rect 4408 4507 4462 4519
rect 4408 4481 4418 4507
rect 4452 4481 4462 4507
rect 4408 4429 4409 4481
rect 4461 4429 4462 4481
rect 4408 4422 4462 4429
rect 4508 4507 4562 4613
rect 4608 4691 4662 4698
rect 4608 4639 4609 4691
rect 4661 4639 4662 4691
rect 4608 4613 4618 4639
rect 4652 4613 4662 4639
rect 4608 4601 4662 4613
rect 4708 4647 4762 4753
rect 4808 4787 4862 4799
rect 4808 4761 4818 4787
rect 4852 4761 4862 4787
rect 4808 4709 4809 4761
rect 4861 4709 4862 4761
rect 4808 4702 4862 4709
rect 4908 4787 4962 4960
rect 5002 4919 5068 4920
rect 5002 4867 5009 4919
rect 5061 4867 5068 4919
rect 5002 4866 5068 4867
rect 4908 4753 4918 4787
rect 4952 4753 4962 4787
rect 4708 4613 4718 4647
rect 4752 4613 4762 4647
rect 4508 4473 4518 4507
rect 4552 4473 4562 4507
rect 4308 4333 4318 4367
rect 4352 4333 4362 4367
rect 4108 4193 4118 4227
rect 4152 4193 4162 4227
rect 3908 4053 3918 4087
rect 3952 4053 3962 4087
rect 3708 3913 3718 3947
rect 3752 3913 3762 3947
rect 3508 3773 3518 3807
rect 3552 3773 3562 3807
rect 3402 3709 3468 3710
rect 3402 3657 3409 3709
rect 3461 3657 3468 3709
rect 3402 3656 3468 3657
rect 3308 3543 3318 3577
rect 3352 3543 3362 3577
rect 3108 3403 3118 3437
rect 3152 3403 3162 3437
rect 2908 3263 2918 3297
rect 2952 3263 2962 3297
rect 2708 3123 2718 3157
rect 2752 3123 2762 3157
rect 2508 2983 2518 3017
rect 2552 2983 2562 3017
rect 2308 2843 2318 2877
rect 2352 2843 2362 2877
rect 2108 2703 2118 2737
rect 2152 2703 2162 2737
rect 1908 2563 1918 2597
rect 1952 2563 1962 2597
rect 1802 2499 1868 2500
rect 1802 2447 1809 2499
rect 1861 2447 1868 2499
rect 1802 2446 1868 2447
rect 1708 2333 1718 2367
rect 1752 2333 1762 2367
rect 1508 2193 1518 2227
rect 1552 2193 1562 2227
rect 1308 2053 1318 2087
rect 1352 2053 1362 2087
rect 1108 1913 1118 1947
rect 1152 1913 1162 1947
rect 908 1773 918 1807
rect 952 1773 962 1807
rect 708 1633 718 1667
rect 752 1633 762 1667
rect 508 1493 518 1527
rect 552 1493 562 1527
rect 308 1353 318 1387
rect 352 1353 362 1387
rect 202 1289 268 1290
rect 202 1237 209 1289
rect 261 1237 268 1289
rect 202 1236 268 1237
rect 108 1123 118 1157
rect 152 1123 162 1157
rect 8 1017 62 1029
rect 8 991 18 1017
rect 52 991 62 1017
rect 8 939 9 991
rect 61 939 62 991
rect 8 932 62 939
rect 108 1017 162 1123
rect 208 1201 262 1208
rect 208 1149 209 1201
rect 261 1149 262 1201
rect 208 1123 218 1149
rect 252 1123 262 1149
rect 208 1111 262 1123
rect 308 1157 362 1353
rect 408 1387 462 1399
rect 408 1361 418 1387
rect 452 1361 462 1387
rect 408 1309 409 1361
rect 461 1309 462 1361
rect 408 1302 462 1309
rect 508 1387 562 1493
rect 608 1571 662 1578
rect 608 1519 609 1571
rect 661 1519 662 1571
rect 608 1493 618 1519
rect 652 1493 662 1519
rect 608 1481 662 1493
rect 708 1527 762 1633
rect 808 1667 862 1679
rect 808 1641 818 1667
rect 852 1641 862 1667
rect 808 1589 809 1641
rect 861 1589 862 1641
rect 808 1582 862 1589
rect 908 1667 962 1773
rect 1008 1851 1062 1858
rect 1008 1799 1009 1851
rect 1061 1799 1062 1851
rect 1008 1773 1018 1799
rect 1052 1773 1062 1799
rect 1008 1761 1062 1773
rect 1108 1807 1162 1913
rect 1208 1947 1262 1959
rect 1208 1921 1218 1947
rect 1252 1921 1262 1947
rect 1208 1869 1209 1921
rect 1261 1869 1262 1921
rect 1208 1862 1262 1869
rect 1308 1947 1362 2053
rect 1408 2131 1462 2138
rect 1408 2079 1409 2131
rect 1461 2079 1462 2131
rect 1408 2053 1418 2079
rect 1452 2053 1462 2079
rect 1408 2041 1462 2053
rect 1508 2087 1562 2193
rect 1608 2227 1662 2239
rect 1608 2201 1618 2227
rect 1652 2201 1662 2227
rect 1608 2149 1609 2201
rect 1661 2149 1662 2201
rect 1608 2142 1662 2149
rect 1708 2227 1762 2333
rect 1808 2411 1862 2418
rect 1808 2359 1809 2411
rect 1861 2359 1862 2411
rect 1808 2333 1818 2359
rect 1852 2333 1862 2359
rect 1808 2321 1862 2333
rect 1908 2367 1962 2563
rect 2008 2597 2062 2609
rect 2008 2571 2018 2597
rect 2052 2571 2062 2597
rect 2008 2519 2009 2571
rect 2061 2519 2062 2571
rect 2008 2512 2062 2519
rect 2108 2597 2162 2703
rect 2208 2781 2262 2788
rect 2208 2729 2209 2781
rect 2261 2729 2262 2781
rect 2208 2703 2218 2729
rect 2252 2703 2262 2729
rect 2208 2691 2262 2703
rect 2308 2737 2362 2843
rect 2408 2877 2462 2889
rect 2408 2851 2418 2877
rect 2452 2851 2462 2877
rect 2408 2799 2409 2851
rect 2461 2799 2462 2851
rect 2408 2792 2462 2799
rect 2508 2877 2562 2983
rect 2608 3061 2662 3068
rect 2608 3009 2609 3061
rect 2661 3009 2662 3061
rect 2608 2983 2618 3009
rect 2652 2983 2662 3009
rect 2608 2971 2662 2983
rect 2708 3017 2762 3123
rect 2808 3157 2862 3169
rect 2808 3131 2818 3157
rect 2852 3131 2862 3157
rect 2808 3079 2809 3131
rect 2861 3079 2862 3131
rect 2808 3072 2862 3079
rect 2908 3157 2962 3263
rect 3008 3341 3062 3348
rect 3008 3289 3009 3341
rect 3061 3289 3062 3341
rect 3008 3263 3018 3289
rect 3052 3263 3062 3289
rect 3008 3251 3062 3263
rect 3108 3297 3162 3403
rect 3208 3437 3262 3449
rect 3208 3411 3218 3437
rect 3252 3411 3262 3437
rect 3208 3359 3209 3411
rect 3261 3359 3262 3411
rect 3208 3352 3262 3359
rect 3308 3437 3362 3543
rect 3408 3621 3462 3628
rect 3408 3569 3409 3621
rect 3461 3569 3462 3621
rect 3408 3543 3418 3569
rect 3452 3543 3462 3569
rect 3408 3531 3462 3543
rect 3508 3577 3562 3773
rect 3608 3807 3662 3819
rect 3608 3781 3618 3807
rect 3652 3781 3662 3807
rect 3608 3729 3609 3781
rect 3661 3729 3662 3781
rect 3608 3722 3662 3729
rect 3708 3807 3762 3913
rect 3808 3991 3862 3998
rect 3808 3939 3809 3991
rect 3861 3939 3862 3991
rect 3808 3913 3818 3939
rect 3852 3913 3862 3939
rect 3808 3901 3862 3913
rect 3908 3947 3962 4053
rect 4008 4087 4062 4099
rect 4008 4061 4018 4087
rect 4052 4061 4062 4087
rect 4008 4009 4009 4061
rect 4061 4009 4062 4061
rect 4008 4002 4062 4009
rect 4108 4087 4162 4193
rect 4208 4271 4262 4278
rect 4208 4219 4209 4271
rect 4261 4219 4262 4271
rect 4208 4193 4218 4219
rect 4252 4193 4262 4219
rect 4208 4181 4262 4193
rect 4308 4227 4362 4333
rect 4408 4367 4462 4379
rect 4408 4341 4418 4367
rect 4452 4341 4462 4367
rect 4408 4289 4409 4341
rect 4461 4289 4462 4341
rect 4408 4282 4462 4289
rect 4508 4367 4562 4473
rect 4608 4551 4662 4558
rect 4608 4499 4609 4551
rect 4661 4499 4662 4551
rect 4608 4473 4618 4499
rect 4652 4473 4662 4499
rect 4608 4461 4662 4473
rect 4708 4507 4762 4613
rect 4808 4647 4862 4659
rect 4808 4621 4818 4647
rect 4852 4621 4862 4647
rect 4808 4569 4809 4621
rect 4861 4569 4862 4621
rect 4808 4562 4862 4569
rect 4908 4647 4962 4753
rect 5008 4831 5062 4838
rect 5008 4779 5009 4831
rect 5061 4779 5062 4831
rect 5008 4753 5018 4779
rect 5052 4753 5062 4779
rect 5008 4741 5062 4753
rect 5108 4787 5162 4960
rect 5202 4903 5268 4904
rect 5202 4851 5209 4903
rect 5261 4851 5268 4903
rect 5202 4850 5268 4851
rect 5108 4753 5118 4787
rect 5152 4753 5162 4787
rect 4908 4613 4918 4647
rect 4952 4613 4962 4647
rect 4708 4473 4718 4507
rect 4752 4473 4762 4507
rect 4508 4333 4518 4367
rect 4552 4333 4562 4367
rect 4308 4193 4318 4227
rect 4352 4193 4362 4227
rect 4108 4053 4118 4087
rect 4152 4053 4162 4087
rect 3908 3913 3918 3947
rect 3952 3913 3962 3947
rect 3708 3773 3718 3807
rect 3752 3773 3762 3807
rect 3602 3693 3668 3694
rect 3602 3641 3609 3693
rect 3661 3641 3668 3693
rect 3602 3640 3668 3641
rect 3508 3543 3518 3577
rect 3552 3543 3562 3577
rect 3308 3403 3318 3437
rect 3352 3403 3362 3437
rect 3108 3263 3118 3297
rect 3152 3263 3162 3297
rect 2908 3123 2918 3157
rect 2952 3123 2962 3157
rect 2708 2983 2718 3017
rect 2752 2983 2762 3017
rect 2508 2843 2518 2877
rect 2552 2843 2562 2877
rect 2308 2703 2318 2737
rect 2352 2703 2362 2737
rect 2108 2563 2118 2597
rect 2152 2563 2162 2597
rect 2002 2483 2068 2484
rect 2002 2431 2009 2483
rect 2061 2431 2068 2483
rect 2002 2430 2068 2431
rect 1908 2333 1918 2367
rect 1952 2333 1962 2367
rect 1708 2193 1718 2227
rect 1752 2193 1762 2227
rect 1508 2053 1518 2087
rect 1552 2053 1562 2087
rect 1308 1913 1318 1947
rect 1352 1913 1362 1947
rect 1108 1773 1118 1807
rect 1152 1773 1162 1807
rect 908 1633 918 1667
rect 952 1633 962 1667
rect 708 1493 718 1527
rect 752 1493 762 1527
rect 508 1353 518 1387
rect 552 1353 562 1387
rect 402 1273 468 1274
rect 402 1221 409 1273
rect 461 1221 468 1273
rect 402 1220 468 1221
rect 308 1123 318 1157
rect 352 1123 362 1157
rect 108 983 118 1017
rect 152 983 162 1017
rect 8 877 62 889
rect 8 851 18 877
rect 52 851 62 877
rect 8 799 9 851
rect 61 799 62 851
rect 8 792 62 799
rect 108 877 162 983
rect 208 1061 262 1068
rect 208 1009 209 1061
rect 261 1009 262 1061
rect 208 983 218 1009
rect 252 983 262 1009
rect 208 971 262 983
rect 308 1017 362 1123
rect 408 1157 462 1169
rect 408 1131 418 1157
rect 452 1131 462 1157
rect 408 1079 409 1131
rect 461 1079 462 1131
rect 408 1072 462 1079
rect 508 1157 562 1353
rect 608 1431 662 1438
rect 608 1379 609 1431
rect 661 1379 662 1431
rect 608 1353 618 1379
rect 652 1353 662 1379
rect 608 1341 662 1353
rect 708 1387 762 1493
rect 808 1527 862 1539
rect 808 1501 818 1527
rect 852 1501 862 1527
rect 808 1449 809 1501
rect 861 1449 862 1501
rect 808 1442 862 1449
rect 908 1527 962 1633
rect 1008 1711 1062 1718
rect 1008 1659 1009 1711
rect 1061 1659 1062 1711
rect 1008 1633 1018 1659
rect 1052 1633 1062 1659
rect 1008 1621 1062 1633
rect 1108 1667 1162 1773
rect 1208 1807 1262 1819
rect 1208 1781 1218 1807
rect 1252 1781 1262 1807
rect 1208 1729 1209 1781
rect 1261 1729 1262 1781
rect 1208 1722 1262 1729
rect 1308 1807 1362 1913
rect 1408 1991 1462 1998
rect 1408 1939 1409 1991
rect 1461 1939 1462 1991
rect 1408 1913 1418 1939
rect 1452 1913 1462 1939
rect 1408 1901 1462 1913
rect 1508 1947 1562 2053
rect 1608 2087 1662 2099
rect 1608 2061 1618 2087
rect 1652 2061 1662 2087
rect 1608 2009 1609 2061
rect 1661 2009 1662 2061
rect 1608 2002 1662 2009
rect 1708 2087 1762 2193
rect 1808 2271 1862 2278
rect 1808 2219 1809 2271
rect 1861 2219 1862 2271
rect 1808 2193 1818 2219
rect 1852 2193 1862 2219
rect 1808 2181 1862 2193
rect 1908 2227 1962 2333
rect 2008 2367 2062 2379
rect 2008 2341 2018 2367
rect 2052 2341 2062 2367
rect 2008 2289 2009 2341
rect 2061 2289 2062 2341
rect 2008 2282 2062 2289
rect 2108 2367 2162 2563
rect 2208 2641 2262 2648
rect 2208 2589 2209 2641
rect 2261 2589 2262 2641
rect 2208 2563 2218 2589
rect 2252 2563 2262 2589
rect 2208 2551 2262 2563
rect 2308 2597 2362 2703
rect 2408 2737 2462 2749
rect 2408 2711 2418 2737
rect 2452 2711 2462 2737
rect 2408 2659 2409 2711
rect 2461 2659 2462 2711
rect 2408 2652 2462 2659
rect 2508 2737 2562 2843
rect 2608 2921 2662 2928
rect 2608 2869 2609 2921
rect 2661 2869 2662 2921
rect 2608 2843 2618 2869
rect 2652 2843 2662 2869
rect 2608 2831 2662 2843
rect 2708 2877 2762 2983
rect 2808 3017 2862 3029
rect 2808 2991 2818 3017
rect 2852 2991 2862 3017
rect 2808 2939 2809 2991
rect 2861 2939 2862 2991
rect 2808 2932 2862 2939
rect 2908 3017 2962 3123
rect 3008 3201 3062 3208
rect 3008 3149 3009 3201
rect 3061 3149 3062 3201
rect 3008 3123 3018 3149
rect 3052 3123 3062 3149
rect 3008 3111 3062 3123
rect 3108 3157 3162 3263
rect 3208 3297 3262 3309
rect 3208 3271 3218 3297
rect 3252 3271 3262 3297
rect 3208 3219 3209 3271
rect 3261 3219 3262 3271
rect 3208 3212 3262 3219
rect 3308 3297 3362 3403
rect 3408 3481 3462 3488
rect 3408 3429 3409 3481
rect 3461 3429 3462 3481
rect 3408 3403 3418 3429
rect 3452 3403 3462 3429
rect 3408 3391 3462 3403
rect 3508 3437 3562 3543
rect 3608 3577 3662 3589
rect 3608 3551 3618 3577
rect 3652 3551 3662 3577
rect 3608 3499 3609 3551
rect 3661 3499 3662 3551
rect 3608 3492 3662 3499
rect 3708 3577 3762 3773
rect 3808 3851 3862 3858
rect 3808 3799 3809 3851
rect 3861 3799 3862 3851
rect 3808 3773 3818 3799
rect 3852 3773 3862 3799
rect 3808 3761 3862 3773
rect 3908 3807 3962 3913
rect 4008 3947 4062 3959
rect 4008 3921 4018 3947
rect 4052 3921 4062 3947
rect 4008 3869 4009 3921
rect 4061 3869 4062 3921
rect 4008 3862 4062 3869
rect 4108 3947 4162 4053
rect 4208 4131 4262 4138
rect 4208 4079 4209 4131
rect 4261 4079 4262 4131
rect 4208 4053 4218 4079
rect 4252 4053 4262 4079
rect 4208 4041 4262 4053
rect 4308 4087 4362 4193
rect 4408 4227 4462 4239
rect 4408 4201 4418 4227
rect 4452 4201 4462 4227
rect 4408 4149 4409 4201
rect 4461 4149 4462 4201
rect 4408 4142 4462 4149
rect 4508 4227 4562 4333
rect 4608 4411 4662 4418
rect 4608 4359 4609 4411
rect 4661 4359 4662 4411
rect 4608 4333 4618 4359
rect 4652 4333 4662 4359
rect 4608 4321 4662 4333
rect 4708 4367 4762 4473
rect 4808 4507 4862 4519
rect 4808 4481 4818 4507
rect 4852 4481 4862 4507
rect 4808 4429 4809 4481
rect 4861 4429 4862 4481
rect 4808 4422 4862 4429
rect 4908 4507 4962 4613
rect 5008 4691 5062 4698
rect 5008 4639 5009 4691
rect 5061 4639 5062 4691
rect 5008 4613 5018 4639
rect 5052 4613 5062 4639
rect 5008 4601 5062 4613
rect 5108 4647 5162 4753
rect 5208 4787 5262 4799
rect 5208 4761 5218 4787
rect 5252 4761 5262 4787
rect 5208 4709 5209 4761
rect 5261 4709 5262 4761
rect 5208 4702 5262 4709
rect 5308 4787 5362 4960
rect 5402 4919 5468 4920
rect 5402 4867 5409 4919
rect 5461 4867 5468 4919
rect 5402 4866 5468 4867
rect 5308 4753 5318 4787
rect 5352 4753 5362 4787
rect 5108 4613 5118 4647
rect 5152 4613 5162 4647
rect 4908 4473 4918 4507
rect 4952 4473 4962 4507
rect 4708 4333 4718 4367
rect 4752 4333 4762 4367
rect 4508 4193 4518 4227
rect 4552 4193 4562 4227
rect 4308 4053 4318 4087
rect 4352 4053 4362 4087
rect 4108 3913 4118 3947
rect 4152 3913 4162 3947
rect 3908 3773 3918 3807
rect 3952 3773 3962 3807
rect 3802 3709 3868 3710
rect 3802 3657 3809 3709
rect 3861 3657 3868 3709
rect 3802 3656 3868 3657
rect 3708 3543 3718 3577
rect 3752 3543 3762 3577
rect 3508 3403 3518 3437
rect 3552 3403 3562 3437
rect 3308 3263 3318 3297
rect 3352 3263 3362 3297
rect 3108 3123 3118 3157
rect 3152 3123 3162 3157
rect 2908 2983 2918 3017
rect 2952 2983 2962 3017
rect 2708 2843 2718 2877
rect 2752 2843 2762 2877
rect 2508 2703 2518 2737
rect 2552 2703 2562 2737
rect 2308 2563 2318 2597
rect 2352 2563 2362 2597
rect 2202 2499 2268 2500
rect 2202 2447 2209 2499
rect 2261 2447 2268 2499
rect 2202 2446 2268 2447
rect 2108 2333 2118 2367
rect 2152 2333 2162 2367
rect 1908 2193 1918 2227
rect 1952 2193 1962 2227
rect 1708 2053 1718 2087
rect 1752 2053 1762 2087
rect 1508 1913 1518 1947
rect 1552 1913 1562 1947
rect 1308 1773 1318 1807
rect 1352 1773 1362 1807
rect 1108 1633 1118 1667
rect 1152 1633 1162 1667
rect 908 1493 918 1527
rect 952 1493 962 1527
rect 708 1353 718 1387
rect 752 1353 762 1387
rect 602 1289 668 1290
rect 602 1237 609 1289
rect 661 1237 668 1289
rect 602 1236 668 1237
rect 508 1123 518 1157
rect 552 1123 562 1157
rect 308 983 318 1017
rect 352 983 362 1017
rect 108 843 118 877
rect 152 843 162 877
rect 8 737 62 749
rect 8 711 18 737
rect 52 711 62 737
rect 8 659 9 711
rect 61 659 62 711
rect 8 652 62 659
rect 108 737 162 843
rect 208 921 262 928
rect 208 869 209 921
rect 261 869 262 921
rect 208 843 218 869
rect 252 843 262 869
rect 208 831 262 843
rect 308 877 362 983
rect 408 1017 462 1029
rect 408 991 418 1017
rect 452 991 462 1017
rect 408 939 409 991
rect 461 939 462 991
rect 408 932 462 939
rect 508 1017 562 1123
rect 608 1201 662 1208
rect 608 1149 609 1201
rect 661 1149 662 1201
rect 608 1123 618 1149
rect 652 1123 662 1149
rect 608 1111 662 1123
rect 708 1157 762 1353
rect 808 1387 862 1399
rect 808 1361 818 1387
rect 852 1361 862 1387
rect 808 1309 809 1361
rect 861 1309 862 1361
rect 808 1302 862 1309
rect 908 1387 962 1493
rect 1008 1571 1062 1578
rect 1008 1519 1009 1571
rect 1061 1519 1062 1571
rect 1008 1493 1018 1519
rect 1052 1493 1062 1519
rect 1008 1481 1062 1493
rect 1108 1527 1162 1633
rect 1208 1667 1262 1679
rect 1208 1641 1218 1667
rect 1252 1641 1262 1667
rect 1208 1589 1209 1641
rect 1261 1589 1262 1641
rect 1208 1582 1262 1589
rect 1308 1667 1362 1773
rect 1408 1851 1462 1858
rect 1408 1799 1409 1851
rect 1461 1799 1462 1851
rect 1408 1773 1418 1799
rect 1452 1773 1462 1799
rect 1408 1761 1462 1773
rect 1508 1807 1562 1913
rect 1608 1947 1662 1959
rect 1608 1921 1618 1947
rect 1652 1921 1662 1947
rect 1608 1869 1609 1921
rect 1661 1869 1662 1921
rect 1608 1862 1662 1869
rect 1708 1947 1762 2053
rect 1808 2131 1862 2138
rect 1808 2079 1809 2131
rect 1861 2079 1862 2131
rect 1808 2053 1818 2079
rect 1852 2053 1862 2079
rect 1808 2041 1862 2053
rect 1908 2087 1962 2193
rect 2008 2227 2062 2239
rect 2008 2201 2018 2227
rect 2052 2201 2062 2227
rect 2008 2149 2009 2201
rect 2061 2149 2062 2201
rect 2008 2142 2062 2149
rect 2108 2227 2162 2333
rect 2208 2411 2262 2418
rect 2208 2359 2209 2411
rect 2261 2359 2262 2411
rect 2208 2333 2218 2359
rect 2252 2333 2262 2359
rect 2208 2321 2262 2333
rect 2308 2367 2362 2563
rect 2408 2597 2462 2609
rect 2408 2571 2418 2597
rect 2452 2571 2462 2597
rect 2408 2519 2409 2571
rect 2461 2519 2462 2571
rect 2408 2512 2462 2519
rect 2508 2597 2562 2703
rect 2608 2781 2662 2788
rect 2608 2729 2609 2781
rect 2661 2729 2662 2781
rect 2608 2703 2618 2729
rect 2652 2703 2662 2729
rect 2608 2691 2662 2703
rect 2708 2737 2762 2843
rect 2808 2877 2862 2889
rect 2808 2851 2818 2877
rect 2852 2851 2862 2877
rect 2808 2799 2809 2851
rect 2861 2799 2862 2851
rect 2808 2792 2862 2799
rect 2908 2877 2962 2983
rect 3008 3061 3062 3068
rect 3008 3009 3009 3061
rect 3061 3009 3062 3061
rect 3008 2983 3018 3009
rect 3052 2983 3062 3009
rect 3008 2971 3062 2983
rect 3108 3017 3162 3123
rect 3208 3157 3262 3169
rect 3208 3131 3218 3157
rect 3252 3131 3262 3157
rect 3208 3079 3209 3131
rect 3261 3079 3262 3131
rect 3208 3072 3262 3079
rect 3308 3157 3362 3263
rect 3408 3341 3462 3348
rect 3408 3289 3409 3341
rect 3461 3289 3462 3341
rect 3408 3263 3418 3289
rect 3452 3263 3462 3289
rect 3408 3251 3462 3263
rect 3508 3297 3562 3403
rect 3608 3437 3662 3449
rect 3608 3411 3618 3437
rect 3652 3411 3662 3437
rect 3608 3359 3609 3411
rect 3661 3359 3662 3411
rect 3608 3352 3662 3359
rect 3708 3437 3762 3543
rect 3808 3621 3862 3628
rect 3808 3569 3809 3621
rect 3861 3569 3862 3621
rect 3808 3543 3818 3569
rect 3852 3543 3862 3569
rect 3808 3531 3862 3543
rect 3908 3577 3962 3773
rect 4008 3807 4062 3819
rect 4008 3781 4018 3807
rect 4052 3781 4062 3807
rect 4008 3729 4009 3781
rect 4061 3729 4062 3781
rect 4008 3722 4062 3729
rect 4108 3807 4162 3913
rect 4208 3991 4262 3998
rect 4208 3939 4209 3991
rect 4261 3939 4262 3991
rect 4208 3913 4218 3939
rect 4252 3913 4262 3939
rect 4208 3901 4262 3913
rect 4308 3947 4362 4053
rect 4408 4087 4462 4099
rect 4408 4061 4418 4087
rect 4452 4061 4462 4087
rect 4408 4009 4409 4061
rect 4461 4009 4462 4061
rect 4408 4002 4462 4009
rect 4508 4087 4562 4193
rect 4608 4271 4662 4278
rect 4608 4219 4609 4271
rect 4661 4219 4662 4271
rect 4608 4193 4618 4219
rect 4652 4193 4662 4219
rect 4608 4181 4662 4193
rect 4708 4227 4762 4333
rect 4808 4367 4862 4379
rect 4808 4341 4818 4367
rect 4852 4341 4862 4367
rect 4808 4289 4809 4341
rect 4861 4289 4862 4341
rect 4808 4282 4862 4289
rect 4908 4367 4962 4473
rect 5008 4551 5062 4558
rect 5008 4499 5009 4551
rect 5061 4499 5062 4551
rect 5008 4473 5018 4499
rect 5052 4473 5062 4499
rect 5008 4461 5062 4473
rect 5108 4507 5162 4613
rect 5208 4647 5262 4659
rect 5208 4621 5218 4647
rect 5252 4621 5262 4647
rect 5208 4569 5209 4621
rect 5261 4569 5262 4621
rect 5208 4562 5262 4569
rect 5308 4647 5362 4753
rect 5408 4831 5462 4838
rect 5408 4779 5409 4831
rect 5461 4779 5462 4831
rect 5408 4753 5418 4779
rect 5452 4753 5462 4779
rect 5408 4741 5462 4753
rect 5508 4787 5562 4960
rect 5602 4903 5668 4904
rect 5602 4851 5609 4903
rect 5661 4851 5668 4903
rect 5602 4850 5668 4851
rect 5508 4753 5518 4787
rect 5552 4753 5562 4787
rect 5308 4613 5318 4647
rect 5352 4613 5362 4647
rect 5108 4473 5118 4507
rect 5152 4473 5162 4507
rect 4908 4333 4918 4367
rect 4952 4333 4962 4367
rect 4708 4193 4718 4227
rect 4752 4193 4762 4227
rect 4508 4053 4518 4087
rect 4552 4053 4562 4087
rect 4308 3913 4318 3947
rect 4352 3913 4362 3947
rect 4108 3773 4118 3807
rect 4152 3773 4162 3807
rect 4002 3693 4068 3694
rect 4002 3641 4009 3693
rect 4061 3641 4068 3693
rect 4002 3640 4068 3641
rect 3908 3543 3918 3577
rect 3952 3543 3962 3577
rect 3708 3403 3718 3437
rect 3752 3403 3762 3437
rect 3508 3263 3518 3297
rect 3552 3263 3562 3297
rect 3308 3123 3318 3157
rect 3352 3123 3362 3157
rect 3108 2983 3118 3017
rect 3152 2983 3162 3017
rect 2908 2843 2918 2877
rect 2952 2843 2962 2877
rect 2708 2703 2718 2737
rect 2752 2703 2762 2737
rect 2508 2563 2518 2597
rect 2552 2563 2562 2597
rect 2402 2483 2468 2484
rect 2402 2431 2409 2483
rect 2461 2431 2468 2483
rect 2402 2430 2468 2431
rect 2308 2333 2318 2367
rect 2352 2333 2362 2367
rect 2108 2193 2118 2227
rect 2152 2193 2162 2227
rect 1908 2053 1918 2087
rect 1952 2053 1962 2087
rect 1708 1913 1718 1947
rect 1752 1913 1762 1947
rect 1508 1773 1518 1807
rect 1552 1773 1562 1807
rect 1308 1633 1318 1667
rect 1352 1633 1362 1667
rect 1108 1493 1118 1527
rect 1152 1493 1162 1527
rect 908 1353 918 1387
rect 952 1353 962 1387
rect 802 1273 868 1274
rect 802 1221 809 1273
rect 861 1221 868 1273
rect 802 1220 868 1221
rect 708 1123 718 1157
rect 752 1123 762 1157
rect 508 983 518 1017
rect 552 983 562 1017
rect 308 843 318 877
rect 352 843 362 877
rect 108 703 118 737
rect 152 703 162 737
rect 8 597 62 609
rect 8 571 18 597
rect 52 571 62 597
rect 8 519 9 571
rect 61 519 62 571
rect 8 512 62 519
rect 108 597 162 703
rect 208 781 262 788
rect 208 729 209 781
rect 261 729 262 781
rect 208 703 218 729
rect 252 703 262 729
rect 208 691 262 703
rect 308 737 362 843
rect 408 877 462 889
rect 408 851 418 877
rect 452 851 462 877
rect 408 799 409 851
rect 461 799 462 851
rect 408 792 462 799
rect 508 877 562 983
rect 608 1061 662 1068
rect 608 1009 609 1061
rect 661 1009 662 1061
rect 608 983 618 1009
rect 652 983 662 1009
rect 608 971 662 983
rect 708 1017 762 1123
rect 808 1157 862 1169
rect 808 1131 818 1157
rect 852 1131 862 1157
rect 808 1079 809 1131
rect 861 1079 862 1131
rect 808 1072 862 1079
rect 908 1157 962 1353
rect 1008 1431 1062 1438
rect 1008 1379 1009 1431
rect 1061 1379 1062 1431
rect 1008 1353 1018 1379
rect 1052 1353 1062 1379
rect 1008 1341 1062 1353
rect 1108 1387 1162 1493
rect 1208 1527 1262 1539
rect 1208 1501 1218 1527
rect 1252 1501 1262 1527
rect 1208 1449 1209 1501
rect 1261 1449 1262 1501
rect 1208 1442 1262 1449
rect 1308 1527 1362 1633
rect 1408 1711 1462 1718
rect 1408 1659 1409 1711
rect 1461 1659 1462 1711
rect 1408 1633 1418 1659
rect 1452 1633 1462 1659
rect 1408 1621 1462 1633
rect 1508 1667 1562 1773
rect 1608 1807 1662 1819
rect 1608 1781 1618 1807
rect 1652 1781 1662 1807
rect 1608 1729 1609 1781
rect 1661 1729 1662 1781
rect 1608 1722 1662 1729
rect 1708 1807 1762 1913
rect 1808 1991 1862 1998
rect 1808 1939 1809 1991
rect 1861 1939 1862 1991
rect 1808 1913 1818 1939
rect 1852 1913 1862 1939
rect 1808 1901 1862 1913
rect 1908 1947 1962 2053
rect 2008 2087 2062 2099
rect 2008 2061 2018 2087
rect 2052 2061 2062 2087
rect 2008 2009 2009 2061
rect 2061 2009 2062 2061
rect 2008 2002 2062 2009
rect 2108 2087 2162 2193
rect 2208 2271 2262 2278
rect 2208 2219 2209 2271
rect 2261 2219 2262 2271
rect 2208 2193 2218 2219
rect 2252 2193 2262 2219
rect 2208 2181 2262 2193
rect 2308 2227 2362 2333
rect 2408 2367 2462 2379
rect 2408 2341 2418 2367
rect 2452 2341 2462 2367
rect 2408 2289 2409 2341
rect 2461 2289 2462 2341
rect 2408 2282 2462 2289
rect 2508 2367 2562 2563
rect 2608 2641 2662 2648
rect 2608 2589 2609 2641
rect 2661 2589 2662 2641
rect 2608 2563 2618 2589
rect 2652 2563 2662 2589
rect 2608 2551 2662 2563
rect 2708 2597 2762 2703
rect 2808 2737 2862 2749
rect 2808 2711 2818 2737
rect 2852 2711 2862 2737
rect 2808 2659 2809 2711
rect 2861 2659 2862 2711
rect 2808 2652 2862 2659
rect 2908 2737 2962 2843
rect 3008 2921 3062 2928
rect 3008 2869 3009 2921
rect 3061 2869 3062 2921
rect 3008 2843 3018 2869
rect 3052 2843 3062 2869
rect 3008 2831 3062 2843
rect 3108 2877 3162 2983
rect 3208 3017 3262 3029
rect 3208 2991 3218 3017
rect 3252 2991 3262 3017
rect 3208 2939 3209 2991
rect 3261 2939 3262 2991
rect 3208 2932 3262 2939
rect 3308 3017 3362 3123
rect 3408 3201 3462 3208
rect 3408 3149 3409 3201
rect 3461 3149 3462 3201
rect 3408 3123 3418 3149
rect 3452 3123 3462 3149
rect 3408 3111 3462 3123
rect 3508 3157 3562 3263
rect 3608 3297 3662 3309
rect 3608 3271 3618 3297
rect 3652 3271 3662 3297
rect 3608 3219 3609 3271
rect 3661 3219 3662 3271
rect 3608 3212 3662 3219
rect 3708 3297 3762 3403
rect 3808 3481 3862 3488
rect 3808 3429 3809 3481
rect 3861 3429 3862 3481
rect 3808 3403 3818 3429
rect 3852 3403 3862 3429
rect 3808 3391 3862 3403
rect 3908 3437 3962 3543
rect 4008 3577 4062 3589
rect 4008 3551 4018 3577
rect 4052 3551 4062 3577
rect 4008 3499 4009 3551
rect 4061 3499 4062 3551
rect 4008 3492 4062 3499
rect 4108 3577 4162 3773
rect 4208 3851 4262 3858
rect 4208 3799 4209 3851
rect 4261 3799 4262 3851
rect 4208 3773 4218 3799
rect 4252 3773 4262 3799
rect 4208 3761 4262 3773
rect 4308 3807 4362 3913
rect 4408 3947 4462 3959
rect 4408 3921 4418 3947
rect 4452 3921 4462 3947
rect 4408 3869 4409 3921
rect 4461 3869 4462 3921
rect 4408 3862 4462 3869
rect 4508 3947 4562 4053
rect 4608 4131 4662 4138
rect 4608 4079 4609 4131
rect 4661 4079 4662 4131
rect 4608 4053 4618 4079
rect 4652 4053 4662 4079
rect 4608 4041 4662 4053
rect 4708 4087 4762 4193
rect 4808 4227 4862 4239
rect 4808 4201 4818 4227
rect 4852 4201 4862 4227
rect 4808 4149 4809 4201
rect 4861 4149 4862 4201
rect 4808 4142 4862 4149
rect 4908 4227 4962 4333
rect 5008 4411 5062 4418
rect 5008 4359 5009 4411
rect 5061 4359 5062 4411
rect 5008 4333 5018 4359
rect 5052 4333 5062 4359
rect 5008 4321 5062 4333
rect 5108 4367 5162 4473
rect 5208 4507 5262 4519
rect 5208 4481 5218 4507
rect 5252 4481 5262 4507
rect 5208 4429 5209 4481
rect 5261 4429 5262 4481
rect 5208 4422 5262 4429
rect 5308 4507 5362 4613
rect 5408 4691 5462 4698
rect 5408 4639 5409 4691
rect 5461 4639 5462 4691
rect 5408 4613 5418 4639
rect 5452 4613 5462 4639
rect 5408 4601 5462 4613
rect 5508 4647 5562 4753
rect 5608 4787 5662 4799
rect 5608 4761 5618 4787
rect 5652 4761 5662 4787
rect 5608 4709 5609 4761
rect 5661 4709 5662 4761
rect 5608 4702 5662 4709
rect 5708 4787 5762 4960
rect 5802 4919 5868 4920
rect 5802 4867 5809 4919
rect 5861 4867 5868 4919
rect 5802 4866 5868 4867
rect 5708 4753 5718 4787
rect 5752 4753 5762 4787
rect 5508 4613 5518 4647
rect 5552 4613 5562 4647
rect 5308 4473 5318 4507
rect 5352 4473 5362 4507
rect 5108 4333 5118 4367
rect 5152 4333 5162 4367
rect 4908 4193 4918 4227
rect 4952 4193 4962 4227
rect 4708 4053 4718 4087
rect 4752 4053 4762 4087
rect 4508 3913 4518 3947
rect 4552 3913 4562 3947
rect 4308 3773 4318 3807
rect 4352 3773 4362 3807
rect 4202 3709 4268 3710
rect 4202 3657 4209 3709
rect 4261 3657 4268 3709
rect 4202 3656 4268 3657
rect 4108 3543 4118 3577
rect 4152 3543 4162 3577
rect 3908 3403 3918 3437
rect 3952 3403 3962 3437
rect 3708 3263 3718 3297
rect 3752 3263 3762 3297
rect 3508 3123 3518 3157
rect 3552 3123 3562 3157
rect 3308 2983 3318 3017
rect 3352 2983 3362 3017
rect 3108 2843 3118 2877
rect 3152 2843 3162 2877
rect 2908 2703 2918 2737
rect 2952 2703 2962 2737
rect 2708 2563 2718 2597
rect 2752 2563 2762 2597
rect 2602 2499 2668 2500
rect 2602 2447 2609 2499
rect 2661 2447 2668 2499
rect 2602 2446 2668 2447
rect 2508 2333 2518 2367
rect 2552 2333 2562 2367
rect 2308 2193 2318 2227
rect 2352 2193 2362 2227
rect 2108 2053 2118 2087
rect 2152 2053 2162 2087
rect 1908 1913 1918 1947
rect 1952 1913 1962 1947
rect 1708 1773 1718 1807
rect 1752 1773 1762 1807
rect 1508 1633 1518 1667
rect 1552 1633 1562 1667
rect 1308 1493 1318 1527
rect 1352 1493 1362 1527
rect 1108 1353 1118 1387
rect 1152 1353 1162 1387
rect 1002 1289 1068 1290
rect 1002 1237 1009 1289
rect 1061 1237 1068 1289
rect 1002 1236 1068 1237
rect 908 1123 918 1157
rect 952 1123 962 1157
rect 708 983 718 1017
rect 752 983 762 1017
rect 508 843 518 877
rect 552 843 562 877
rect 308 703 318 737
rect 352 703 362 737
rect 108 563 118 597
rect 152 563 162 597
rect 8 457 62 469
rect 8 431 18 457
rect 52 431 62 457
rect 8 379 9 431
rect 61 379 62 431
rect 8 372 62 379
rect 108 457 162 563
rect 208 641 262 648
rect 208 589 209 641
rect 261 589 262 641
rect 208 563 218 589
rect 252 563 262 589
rect 208 551 262 563
rect 308 597 362 703
rect 408 737 462 749
rect 408 711 418 737
rect 452 711 462 737
rect 408 659 409 711
rect 461 659 462 711
rect 408 652 462 659
rect 508 737 562 843
rect 608 921 662 928
rect 608 869 609 921
rect 661 869 662 921
rect 608 843 618 869
rect 652 843 662 869
rect 608 831 662 843
rect 708 877 762 983
rect 808 1017 862 1029
rect 808 991 818 1017
rect 852 991 862 1017
rect 808 939 809 991
rect 861 939 862 991
rect 808 932 862 939
rect 908 1017 962 1123
rect 1008 1201 1062 1208
rect 1008 1149 1009 1201
rect 1061 1149 1062 1201
rect 1008 1123 1018 1149
rect 1052 1123 1062 1149
rect 1008 1111 1062 1123
rect 1108 1157 1162 1353
rect 1208 1387 1262 1399
rect 1208 1361 1218 1387
rect 1252 1361 1262 1387
rect 1208 1309 1209 1361
rect 1261 1309 1262 1361
rect 1208 1302 1262 1309
rect 1308 1387 1362 1493
rect 1408 1571 1462 1578
rect 1408 1519 1409 1571
rect 1461 1519 1462 1571
rect 1408 1493 1418 1519
rect 1452 1493 1462 1519
rect 1408 1481 1462 1493
rect 1508 1527 1562 1633
rect 1608 1667 1662 1679
rect 1608 1641 1618 1667
rect 1652 1641 1662 1667
rect 1608 1589 1609 1641
rect 1661 1589 1662 1641
rect 1608 1582 1662 1589
rect 1708 1667 1762 1773
rect 1808 1851 1862 1858
rect 1808 1799 1809 1851
rect 1861 1799 1862 1851
rect 1808 1773 1818 1799
rect 1852 1773 1862 1799
rect 1808 1761 1862 1773
rect 1908 1807 1962 1913
rect 2008 1947 2062 1959
rect 2008 1921 2018 1947
rect 2052 1921 2062 1947
rect 2008 1869 2009 1921
rect 2061 1869 2062 1921
rect 2008 1862 2062 1869
rect 2108 1947 2162 2053
rect 2208 2131 2262 2138
rect 2208 2079 2209 2131
rect 2261 2079 2262 2131
rect 2208 2053 2218 2079
rect 2252 2053 2262 2079
rect 2208 2041 2262 2053
rect 2308 2087 2362 2193
rect 2408 2227 2462 2239
rect 2408 2201 2418 2227
rect 2452 2201 2462 2227
rect 2408 2149 2409 2201
rect 2461 2149 2462 2201
rect 2408 2142 2462 2149
rect 2508 2227 2562 2333
rect 2608 2411 2662 2418
rect 2608 2359 2609 2411
rect 2661 2359 2662 2411
rect 2608 2333 2618 2359
rect 2652 2333 2662 2359
rect 2608 2321 2662 2333
rect 2708 2367 2762 2563
rect 2808 2597 2862 2609
rect 2808 2571 2818 2597
rect 2852 2571 2862 2597
rect 2808 2519 2809 2571
rect 2861 2519 2862 2571
rect 2808 2512 2862 2519
rect 2908 2597 2962 2703
rect 3008 2781 3062 2788
rect 3008 2729 3009 2781
rect 3061 2729 3062 2781
rect 3008 2703 3018 2729
rect 3052 2703 3062 2729
rect 3008 2691 3062 2703
rect 3108 2737 3162 2843
rect 3208 2877 3262 2889
rect 3208 2851 3218 2877
rect 3252 2851 3262 2877
rect 3208 2799 3209 2851
rect 3261 2799 3262 2851
rect 3208 2792 3262 2799
rect 3308 2877 3362 2983
rect 3408 3061 3462 3068
rect 3408 3009 3409 3061
rect 3461 3009 3462 3061
rect 3408 2983 3418 3009
rect 3452 2983 3462 3009
rect 3408 2971 3462 2983
rect 3508 3017 3562 3123
rect 3608 3157 3662 3169
rect 3608 3131 3618 3157
rect 3652 3131 3662 3157
rect 3608 3079 3609 3131
rect 3661 3079 3662 3131
rect 3608 3072 3662 3079
rect 3708 3157 3762 3263
rect 3808 3341 3862 3348
rect 3808 3289 3809 3341
rect 3861 3289 3862 3341
rect 3808 3263 3818 3289
rect 3852 3263 3862 3289
rect 3808 3251 3862 3263
rect 3908 3297 3962 3403
rect 4008 3437 4062 3449
rect 4008 3411 4018 3437
rect 4052 3411 4062 3437
rect 4008 3359 4009 3411
rect 4061 3359 4062 3411
rect 4008 3352 4062 3359
rect 4108 3437 4162 3543
rect 4208 3621 4262 3628
rect 4208 3569 4209 3621
rect 4261 3569 4262 3621
rect 4208 3543 4218 3569
rect 4252 3543 4262 3569
rect 4208 3531 4262 3543
rect 4308 3577 4362 3773
rect 4408 3807 4462 3819
rect 4408 3781 4418 3807
rect 4452 3781 4462 3807
rect 4408 3729 4409 3781
rect 4461 3729 4462 3781
rect 4408 3722 4462 3729
rect 4508 3807 4562 3913
rect 4608 3991 4662 3998
rect 4608 3939 4609 3991
rect 4661 3939 4662 3991
rect 4608 3913 4618 3939
rect 4652 3913 4662 3939
rect 4608 3901 4662 3913
rect 4708 3947 4762 4053
rect 4808 4087 4862 4099
rect 4808 4061 4818 4087
rect 4852 4061 4862 4087
rect 4808 4009 4809 4061
rect 4861 4009 4862 4061
rect 4808 4002 4862 4009
rect 4908 4087 4962 4193
rect 5008 4271 5062 4278
rect 5008 4219 5009 4271
rect 5061 4219 5062 4271
rect 5008 4193 5018 4219
rect 5052 4193 5062 4219
rect 5008 4181 5062 4193
rect 5108 4227 5162 4333
rect 5208 4367 5262 4379
rect 5208 4341 5218 4367
rect 5252 4341 5262 4367
rect 5208 4289 5209 4341
rect 5261 4289 5262 4341
rect 5208 4282 5262 4289
rect 5308 4367 5362 4473
rect 5408 4551 5462 4558
rect 5408 4499 5409 4551
rect 5461 4499 5462 4551
rect 5408 4473 5418 4499
rect 5452 4473 5462 4499
rect 5408 4461 5462 4473
rect 5508 4507 5562 4613
rect 5608 4647 5662 4659
rect 5608 4621 5618 4647
rect 5652 4621 5662 4647
rect 5608 4569 5609 4621
rect 5661 4569 5662 4621
rect 5608 4562 5662 4569
rect 5708 4647 5762 4753
rect 5808 4831 5862 4838
rect 5808 4779 5809 4831
rect 5861 4779 5862 4831
rect 5808 4753 5818 4779
rect 5852 4753 5862 4779
rect 5808 4741 5862 4753
rect 5908 4787 5962 4960
rect 6002 4903 6068 4904
rect 6002 4851 6009 4903
rect 6061 4851 6068 4903
rect 6002 4850 6068 4851
rect 5908 4753 5918 4787
rect 5952 4753 5962 4787
rect 5708 4613 5718 4647
rect 5752 4613 5762 4647
rect 5508 4473 5518 4507
rect 5552 4473 5562 4507
rect 5308 4333 5318 4367
rect 5352 4333 5362 4367
rect 5108 4193 5118 4227
rect 5152 4193 5162 4227
rect 4908 4053 4918 4087
rect 4952 4053 4962 4087
rect 4708 3913 4718 3947
rect 4752 3913 4762 3947
rect 4508 3773 4518 3807
rect 4552 3773 4562 3807
rect 4402 3693 4468 3694
rect 4402 3641 4409 3693
rect 4461 3641 4468 3693
rect 4402 3640 4468 3641
rect 4308 3543 4318 3577
rect 4352 3543 4362 3577
rect 4108 3403 4118 3437
rect 4152 3403 4162 3437
rect 3908 3263 3918 3297
rect 3952 3263 3962 3297
rect 3708 3123 3718 3157
rect 3752 3123 3762 3157
rect 3508 2983 3518 3017
rect 3552 2983 3562 3017
rect 3308 2843 3318 2877
rect 3352 2843 3362 2877
rect 3108 2703 3118 2737
rect 3152 2703 3162 2737
rect 2908 2563 2918 2597
rect 2952 2563 2962 2597
rect 2802 2483 2868 2484
rect 2802 2431 2809 2483
rect 2861 2431 2868 2483
rect 2802 2430 2868 2431
rect 2708 2333 2718 2367
rect 2752 2333 2762 2367
rect 2508 2193 2518 2227
rect 2552 2193 2562 2227
rect 2308 2053 2318 2087
rect 2352 2053 2362 2087
rect 2108 1913 2118 1947
rect 2152 1913 2162 1947
rect 1908 1773 1918 1807
rect 1952 1773 1962 1807
rect 1708 1633 1718 1667
rect 1752 1633 1762 1667
rect 1508 1493 1518 1527
rect 1552 1493 1562 1527
rect 1308 1353 1318 1387
rect 1352 1353 1362 1387
rect 1202 1273 1268 1274
rect 1202 1221 1209 1273
rect 1261 1221 1268 1273
rect 1202 1220 1268 1221
rect 1108 1123 1118 1157
rect 1152 1123 1162 1157
rect 908 983 918 1017
rect 952 983 962 1017
rect 708 843 718 877
rect 752 843 762 877
rect 508 703 518 737
rect 552 703 562 737
rect 308 563 318 597
rect 352 563 362 597
rect 108 423 118 457
rect 152 423 162 457
rect 8 317 62 329
rect 8 291 18 317
rect 52 291 62 317
rect 8 239 9 291
rect 61 239 62 291
rect 8 232 62 239
rect 108 317 162 423
rect 208 501 262 508
rect 208 449 209 501
rect 261 449 262 501
rect 208 423 218 449
rect 252 423 262 449
rect 208 411 262 423
rect 308 457 362 563
rect 408 597 462 609
rect 408 571 418 597
rect 452 571 462 597
rect 408 519 409 571
rect 461 519 462 571
rect 408 512 462 519
rect 508 597 562 703
rect 608 781 662 788
rect 608 729 609 781
rect 661 729 662 781
rect 608 703 618 729
rect 652 703 662 729
rect 608 691 662 703
rect 708 737 762 843
rect 808 877 862 889
rect 808 851 818 877
rect 852 851 862 877
rect 808 799 809 851
rect 861 799 862 851
rect 808 792 862 799
rect 908 877 962 983
rect 1008 1061 1062 1068
rect 1008 1009 1009 1061
rect 1061 1009 1062 1061
rect 1008 983 1018 1009
rect 1052 983 1062 1009
rect 1008 971 1062 983
rect 1108 1017 1162 1123
rect 1208 1157 1262 1169
rect 1208 1131 1218 1157
rect 1252 1131 1262 1157
rect 1208 1079 1209 1131
rect 1261 1079 1262 1131
rect 1208 1072 1262 1079
rect 1308 1157 1362 1353
rect 1408 1431 1462 1438
rect 1408 1379 1409 1431
rect 1461 1379 1462 1431
rect 1408 1353 1418 1379
rect 1452 1353 1462 1379
rect 1408 1341 1462 1353
rect 1508 1387 1562 1493
rect 1608 1527 1662 1539
rect 1608 1501 1618 1527
rect 1652 1501 1662 1527
rect 1608 1449 1609 1501
rect 1661 1449 1662 1501
rect 1608 1442 1662 1449
rect 1708 1527 1762 1633
rect 1808 1711 1862 1718
rect 1808 1659 1809 1711
rect 1861 1659 1862 1711
rect 1808 1633 1818 1659
rect 1852 1633 1862 1659
rect 1808 1621 1862 1633
rect 1908 1667 1962 1773
rect 2008 1807 2062 1819
rect 2008 1781 2018 1807
rect 2052 1781 2062 1807
rect 2008 1729 2009 1781
rect 2061 1729 2062 1781
rect 2008 1722 2062 1729
rect 2108 1807 2162 1913
rect 2208 1991 2262 1998
rect 2208 1939 2209 1991
rect 2261 1939 2262 1991
rect 2208 1913 2218 1939
rect 2252 1913 2262 1939
rect 2208 1901 2262 1913
rect 2308 1947 2362 2053
rect 2408 2087 2462 2099
rect 2408 2061 2418 2087
rect 2452 2061 2462 2087
rect 2408 2009 2409 2061
rect 2461 2009 2462 2061
rect 2408 2002 2462 2009
rect 2508 2087 2562 2193
rect 2608 2271 2662 2278
rect 2608 2219 2609 2271
rect 2661 2219 2662 2271
rect 2608 2193 2618 2219
rect 2652 2193 2662 2219
rect 2608 2181 2662 2193
rect 2708 2227 2762 2333
rect 2808 2367 2862 2379
rect 2808 2341 2818 2367
rect 2852 2341 2862 2367
rect 2808 2289 2809 2341
rect 2861 2289 2862 2341
rect 2808 2282 2862 2289
rect 2908 2367 2962 2563
rect 3008 2641 3062 2648
rect 3008 2589 3009 2641
rect 3061 2589 3062 2641
rect 3008 2563 3018 2589
rect 3052 2563 3062 2589
rect 3008 2551 3062 2563
rect 3108 2597 3162 2703
rect 3208 2737 3262 2749
rect 3208 2711 3218 2737
rect 3252 2711 3262 2737
rect 3208 2659 3209 2711
rect 3261 2659 3262 2711
rect 3208 2652 3262 2659
rect 3308 2737 3362 2843
rect 3408 2921 3462 2928
rect 3408 2869 3409 2921
rect 3461 2869 3462 2921
rect 3408 2843 3418 2869
rect 3452 2843 3462 2869
rect 3408 2831 3462 2843
rect 3508 2877 3562 2983
rect 3608 3017 3662 3029
rect 3608 2991 3618 3017
rect 3652 2991 3662 3017
rect 3608 2939 3609 2991
rect 3661 2939 3662 2991
rect 3608 2932 3662 2939
rect 3708 3017 3762 3123
rect 3808 3201 3862 3208
rect 3808 3149 3809 3201
rect 3861 3149 3862 3201
rect 3808 3123 3818 3149
rect 3852 3123 3862 3149
rect 3808 3111 3862 3123
rect 3908 3157 3962 3263
rect 4008 3297 4062 3309
rect 4008 3271 4018 3297
rect 4052 3271 4062 3297
rect 4008 3219 4009 3271
rect 4061 3219 4062 3271
rect 4008 3212 4062 3219
rect 4108 3297 4162 3403
rect 4208 3481 4262 3488
rect 4208 3429 4209 3481
rect 4261 3429 4262 3481
rect 4208 3403 4218 3429
rect 4252 3403 4262 3429
rect 4208 3391 4262 3403
rect 4308 3437 4362 3543
rect 4408 3577 4462 3589
rect 4408 3551 4418 3577
rect 4452 3551 4462 3577
rect 4408 3499 4409 3551
rect 4461 3499 4462 3551
rect 4408 3492 4462 3499
rect 4508 3577 4562 3773
rect 4608 3851 4662 3858
rect 4608 3799 4609 3851
rect 4661 3799 4662 3851
rect 4608 3773 4618 3799
rect 4652 3773 4662 3799
rect 4608 3761 4662 3773
rect 4708 3807 4762 3913
rect 4808 3947 4862 3959
rect 4808 3921 4818 3947
rect 4852 3921 4862 3947
rect 4808 3869 4809 3921
rect 4861 3869 4862 3921
rect 4808 3862 4862 3869
rect 4908 3947 4962 4053
rect 5008 4131 5062 4138
rect 5008 4079 5009 4131
rect 5061 4079 5062 4131
rect 5008 4053 5018 4079
rect 5052 4053 5062 4079
rect 5008 4041 5062 4053
rect 5108 4087 5162 4193
rect 5208 4227 5262 4239
rect 5208 4201 5218 4227
rect 5252 4201 5262 4227
rect 5208 4149 5209 4201
rect 5261 4149 5262 4201
rect 5208 4142 5262 4149
rect 5308 4227 5362 4333
rect 5408 4411 5462 4418
rect 5408 4359 5409 4411
rect 5461 4359 5462 4411
rect 5408 4333 5418 4359
rect 5452 4333 5462 4359
rect 5408 4321 5462 4333
rect 5508 4367 5562 4473
rect 5608 4507 5662 4519
rect 5608 4481 5618 4507
rect 5652 4481 5662 4507
rect 5608 4429 5609 4481
rect 5661 4429 5662 4481
rect 5608 4422 5662 4429
rect 5708 4507 5762 4613
rect 5808 4691 5862 4698
rect 5808 4639 5809 4691
rect 5861 4639 5862 4691
rect 5808 4613 5818 4639
rect 5852 4613 5862 4639
rect 5808 4601 5862 4613
rect 5908 4647 5962 4753
rect 6008 4787 6062 4799
rect 6008 4761 6018 4787
rect 6052 4761 6062 4787
rect 6008 4709 6009 4761
rect 6061 4709 6062 4761
rect 6008 4702 6062 4709
rect 6108 4787 6162 4960
rect 6202 4919 6268 4920
rect 6202 4867 6209 4919
rect 6261 4867 6268 4919
rect 6202 4866 6268 4867
rect 6108 4753 6118 4787
rect 6152 4753 6162 4787
rect 5908 4613 5918 4647
rect 5952 4613 5962 4647
rect 5708 4473 5718 4507
rect 5752 4473 5762 4507
rect 5508 4333 5518 4367
rect 5552 4333 5562 4367
rect 5308 4193 5318 4227
rect 5352 4193 5362 4227
rect 5108 4053 5118 4087
rect 5152 4053 5162 4087
rect 4908 3913 4918 3947
rect 4952 3913 4962 3947
rect 4708 3773 4718 3807
rect 4752 3773 4762 3807
rect 4602 3709 4668 3710
rect 4602 3657 4609 3709
rect 4661 3657 4668 3709
rect 4602 3656 4668 3657
rect 4508 3543 4518 3577
rect 4552 3543 4562 3577
rect 4308 3403 4318 3437
rect 4352 3403 4362 3437
rect 4108 3263 4118 3297
rect 4152 3263 4162 3297
rect 3908 3123 3918 3157
rect 3952 3123 3962 3157
rect 3708 2983 3718 3017
rect 3752 2983 3762 3017
rect 3508 2843 3518 2877
rect 3552 2843 3562 2877
rect 3308 2703 3318 2737
rect 3352 2703 3362 2737
rect 3108 2563 3118 2597
rect 3152 2563 3162 2597
rect 3002 2499 3068 2500
rect 3002 2447 3009 2499
rect 3061 2447 3068 2499
rect 3002 2446 3068 2447
rect 2908 2333 2918 2367
rect 2952 2333 2962 2367
rect 2708 2193 2718 2227
rect 2752 2193 2762 2227
rect 2508 2053 2518 2087
rect 2552 2053 2562 2087
rect 2308 1913 2318 1947
rect 2352 1913 2362 1947
rect 2108 1773 2118 1807
rect 2152 1773 2162 1807
rect 1908 1633 1918 1667
rect 1952 1633 1962 1667
rect 1708 1493 1718 1527
rect 1752 1493 1762 1527
rect 1508 1353 1518 1387
rect 1552 1353 1562 1387
rect 1402 1289 1468 1290
rect 1402 1237 1409 1289
rect 1461 1237 1468 1289
rect 1402 1236 1468 1237
rect 1308 1123 1318 1157
rect 1352 1123 1362 1157
rect 1108 983 1118 1017
rect 1152 983 1162 1017
rect 908 843 918 877
rect 952 843 962 877
rect 708 703 718 737
rect 752 703 762 737
rect 508 563 518 597
rect 552 563 562 597
rect 308 423 318 457
rect 352 423 362 457
rect 108 283 118 317
rect 152 283 162 317
rect 8 177 62 189
rect 8 151 18 177
rect 52 151 62 177
rect 8 99 9 151
rect 61 99 62 151
rect 8 92 62 99
rect 108 177 162 283
rect 208 361 262 368
rect 208 309 209 361
rect 261 309 262 361
rect 208 283 218 309
rect 252 283 262 309
rect 208 271 262 283
rect 308 317 362 423
rect 408 457 462 469
rect 408 431 418 457
rect 452 431 462 457
rect 408 379 409 431
rect 461 379 462 431
rect 408 372 462 379
rect 508 457 562 563
rect 608 641 662 648
rect 608 589 609 641
rect 661 589 662 641
rect 608 563 618 589
rect 652 563 662 589
rect 608 551 662 563
rect 708 597 762 703
rect 808 737 862 749
rect 808 711 818 737
rect 852 711 862 737
rect 808 659 809 711
rect 861 659 862 711
rect 808 652 862 659
rect 908 737 962 843
rect 1008 921 1062 928
rect 1008 869 1009 921
rect 1061 869 1062 921
rect 1008 843 1018 869
rect 1052 843 1062 869
rect 1008 831 1062 843
rect 1108 877 1162 983
rect 1208 1017 1262 1029
rect 1208 991 1218 1017
rect 1252 991 1262 1017
rect 1208 939 1209 991
rect 1261 939 1262 991
rect 1208 932 1262 939
rect 1308 1017 1362 1123
rect 1408 1201 1462 1208
rect 1408 1149 1409 1201
rect 1461 1149 1462 1201
rect 1408 1123 1418 1149
rect 1452 1123 1462 1149
rect 1408 1111 1462 1123
rect 1508 1157 1562 1353
rect 1608 1387 1662 1399
rect 1608 1361 1618 1387
rect 1652 1361 1662 1387
rect 1608 1309 1609 1361
rect 1661 1309 1662 1361
rect 1608 1302 1662 1309
rect 1708 1387 1762 1493
rect 1808 1571 1862 1578
rect 1808 1519 1809 1571
rect 1861 1519 1862 1571
rect 1808 1493 1818 1519
rect 1852 1493 1862 1519
rect 1808 1481 1862 1493
rect 1908 1527 1962 1633
rect 2008 1667 2062 1679
rect 2008 1641 2018 1667
rect 2052 1641 2062 1667
rect 2008 1589 2009 1641
rect 2061 1589 2062 1641
rect 2008 1582 2062 1589
rect 2108 1667 2162 1773
rect 2208 1851 2262 1858
rect 2208 1799 2209 1851
rect 2261 1799 2262 1851
rect 2208 1773 2218 1799
rect 2252 1773 2262 1799
rect 2208 1761 2262 1773
rect 2308 1807 2362 1913
rect 2408 1947 2462 1959
rect 2408 1921 2418 1947
rect 2452 1921 2462 1947
rect 2408 1869 2409 1921
rect 2461 1869 2462 1921
rect 2408 1862 2462 1869
rect 2508 1947 2562 2053
rect 2608 2131 2662 2138
rect 2608 2079 2609 2131
rect 2661 2079 2662 2131
rect 2608 2053 2618 2079
rect 2652 2053 2662 2079
rect 2608 2041 2662 2053
rect 2708 2087 2762 2193
rect 2808 2227 2862 2239
rect 2808 2201 2818 2227
rect 2852 2201 2862 2227
rect 2808 2149 2809 2201
rect 2861 2149 2862 2201
rect 2808 2142 2862 2149
rect 2908 2227 2962 2333
rect 3008 2411 3062 2418
rect 3008 2359 3009 2411
rect 3061 2359 3062 2411
rect 3008 2333 3018 2359
rect 3052 2333 3062 2359
rect 3008 2321 3062 2333
rect 3108 2367 3162 2563
rect 3208 2597 3262 2609
rect 3208 2571 3218 2597
rect 3252 2571 3262 2597
rect 3208 2519 3209 2571
rect 3261 2519 3262 2571
rect 3208 2512 3262 2519
rect 3308 2597 3362 2703
rect 3408 2781 3462 2788
rect 3408 2729 3409 2781
rect 3461 2729 3462 2781
rect 3408 2703 3418 2729
rect 3452 2703 3462 2729
rect 3408 2691 3462 2703
rect 3508 2737 3562 2843
rect 3608 2877 3662 2889
rect 3608 2851 3618 2877
rect 3652 2851 3662 2877
rect 3608 2799 3609 2851
rect 3661 2799 3662 2851
rect 3608 2792 3662 2799
rect 3708 2877 3762 2983
rect 3808 3061 3862 3068
rect 3808 3009 3809 3061
rect 3861 3009 3862 3061
rect 3808 2983 3818 3009
rect 3852 2983 3862 3009
rect 3808 2971 3862 2983
rect 3908 3017 3962 3123
rect 4008 3157 4062 3169
rect 4008 3131 4018 3157
rect 4052 3131 4062 3157
rect 4008 3079 4009 3131
rect 4061 3079 4062 3131
rect 4008 3072 4062 3079
rect 4108 3157 4162 3263
rect 4208 3341 4262 3348
rect 4208 3289 4209 3341
rect 4261 3289 4262 3341
rect 4208 3263 4218 3289
rect 4252 3263 4262 3289
rect 4208 3251 4262 3263
rect 4308 3297 4362 3403
rect 4408 3437 4462 3449
rect 4408 3411 4418 3437
rect 4452 3411 4462 3437
rect 4408 3359 4409 3411
rect 4461 3359 4462 3411
rect 4408 3352 4462 3359
rect 4508 3437 4562 3543
rect 4608 3621 4662 3628
rect 4608 3569 4609 3621
rect 4661 3569 4662 3621
rect 4608 3543 4618 3569
rect 4652 3543 4662 3569
rect 4608 3531 4662 3543
rect 4708 3577 4762 3773
rect 4808 3807 4862 3819
rect 4808 3781 4818 3807
rect 4852 3781 4862 3807
rect 4808 3729 4809 3781
rect 4861 3729 4862 3781
rect 4808 3722 4862 3729
rect 4908 3807 4962 3913
rect 5008 3991 5062 3998
rect 5008 3939 5009 3991
rect 5061 3939 5062 3991
rect 5008 3913 5018 3939
rect 5052 3913 5062 3939
rect 5008 3901 5062 3913
rect 5108 3947 5162 4053
rect 5208 4087 5262 4099
rect 5208 4061 5218 4087
rect 5252 4061 5262 4087
rect 5208 4009 5209 4061
rect 5261 4009 5262 4061
rect 5208 4002 5262 4009
rect 5308 4087 5362 4193
rect 5408 4271 5462 4278
rect 5408 4219 5409 4271
rect 5461 4219 5462 4271
rect 5408 4193 5418 4219
rect 5452 4193 5462 4219
rect 5408 4181 5462 4193
rect 5508 4227 5562 4333
rect 5608 4367 5662 4379
rect 5608 4341 5618 4367
rect 5652 4341 5662 4367
rect 5608 4289 5609 4341
rect 5661 4289 5662 4341
rect 5608 4282 5662 4289
rect 5708 4367 5762 4473
rect 5808 4551 5862 4558
rect 5808 4499 5809 4551
rect 5861 4499 5862 4551
rect 5808 4473 5818 4499
rect 5852 4473 5862 4499
rect 5808 4461 5862 4473
rect 5908 4507 5962 4613
rect 6008 4647 6062 4659
rect 6008 4621 6018 4647
rect 6052 4621 6062 4647
rect 6008 4569 6009 4621
rect 6061 4569 6062 4621
rect 6008 4562 6062 4569
rect 6108 4647 6162 4753
rect 6208 4831 6262 4838
rect 6208 4779 6209 4831
rect 6261 4779 6262 4831
rect 6208 4753 6218 4779
rect 6252 4753 6262 4779
rect 6208 4741 6262 4753
rect 6308 4787 6362 4960
rect 6402 4903 6468 4904
rect 6402 4851 6409 4903
rect 6461 4851 6468 4903
rect 6402 4850 6468 4851
rect 6308 4753 6318 4787
rect 6352 4753 6362 4787
rect 6108 4613 6118 4647
rect 6152 4613 6162 4647
rect 5908 4473 5918 4507
rect 5952 4473 5962 4507
rect 5708 4333 5718 4367
rect 5752 4333 5762 4367
rect 5508 4193 5518 4227
rect 5552 4193 5562 4227
rect 5308 4053 5318 4087
rect 5352 4053 5362 4087
rect 5108 3913 5118 3947
rect 5152 3913 5162 3947
rect 4908 3773 4918 3807
rect 4952 3773 4962 3807
rect 4802 3693 4868 3694
rect 4802 3641 4809 3693
rect 4861 3641 4868 3693
rect 4802 3640 4868 3641
rect 4708 3543 4718 3577
rect 4752 3543 4762 3577
rect 4508 3403 4518 3437
rect 4552 3403 4562 3437
rect 4308 3263 4318 3297
rect 4352 3263 4362 3297
rect 4108 3123 4118 3157
rect 4152 3123 4162 3157
rect 3908 2983 3918 3017
rect 3952 2983 3962 3017
rect 3708 2843 3718 2877
rect 3752 2843 3762 2877
rect 3508 2703 3518 2737
rect 3552 2703 3562 2737
rect 3308 2563 3318 2597
rect 3352 2563 3362 2597
rect 3202 2483 3268 2484
rect 3202 2431 3209 2483
rect 3261 2431 3268 2483
rect 3202 2430 3268 2431
rect 3108 2333 3118 2367
rect 3152 2333 3162 2367
rect 2908 2193 2918 2227
rect 2952 2193 2962 2227
rect 2708 2053 2718 2087
rect 2752 2053 2762 2087
rect 2508 1913 2518 1947
rect 2552 1913 2562 1947
rect 2308 1773 2318 1807
rect 2352 1773 2362 1807
rect 2108 1633 2118 1667
rect 2152 1633 2162 1667
rect 1908 1493 1918 1527
rect 1952 1493 1962 1527
rect 1708 1353 1718 1387
rect 1752 1353 1762 1387
rect 1602 1273 1668 1274
rect 1602 1221 1609 1273
rect 1661 1221 1668 1273
rect 1602 1220 1668 1221
rect 1508 1123 1518 1157
rect 1552 1123 1562 1157
rect 1308 983 1318 1017
rect 1352 983 1362 1017
rect 1108 843 1118 877
rect 1152 843 1162 877
rect 908 703 918 737
rect 952 703 962 737
rect 708 563 718 597
rect 752 563 762 597
rect 508 423 518 457
rect 552 423 562 457
rect 308 283 318 317
rect 352 283 362 317
rect 108 143 118 177
rect 152 143 162 177
rect 2 63 68 64
rect 2 11 9 63
rect 61 11 68 63
rect 2 10 68 11
rect -92 -15 -38 0
rect -92 -67 -91 -15
rect -39 -67 -38 -15
rect -92 -79 -82 -67
rect -48 -79 -38 -67
rect -92 -131 -91 -79
rect -39 -131 -38 -79
rect 8 -22 62 10
rect 8 -74 9 -22
rect 61 -74 62 -22
rect 8 -81 62 -74
rect 108 -15 162 143
rect 208 221 262 228
rect 208 169 209 221
rect 261 169 262 221
rect 208 143 218 169
rect 252 143 262 169
rect 208 131 262 143
rect 308 177 362 283
rect 408 317 462 329
rect 408 291 418 317
rect 452 291 462 317
rect 408 239 409 291
rect 461 239 462 291
rect 408 232 462 239
rect 508 317 562 423
rect 608 501 662 508
rect 608 449 609 501
rect 661 449 662 501
rect 608 423 618 449
rect 652 423 662 449
rect 608 411 662 423
rect 708 457 762 563
rect 808 597 862 609
rect 808 571 818 597
rect 852 571 862 597
rect 808 519 809 571
rect 861 519 862 571
rect 808 512 862 519
rect 908 597 962 703
rect 1008 781 1062 788
rect 1008 729 1009 781
rect 1061 729 1062 781
rect 1008 703 1018 729
rect 1052 703 1062 729
rect 1008 691 1062 703
rect 1108 737 1162 843
rect 1208 877 1262 889
rect 1208 851 1218 877
rect 1252 851 1262 877
rect 1208 799 1209 851
rect 1261 799 1262 851
rect 1208 792 1262 799
rect 1308 877 1362 983
rect 1408 1061 1462 1068
rect 1408 1009 1409 1061
rect 1461 1009 1462 1061
rect 1408 983 1418 1009
rect 1452 983 1462 1009
rect 1408 971 1462 983
rect 1508 1017 1562 1123
rect 1608 1157 1662 1169
rect 1608 1131 1618 1157
rect 1652 1131 1662 1157
rect 1608 1079 1609 1131
rect 1661 1079 1662 1131
rect 1608 1072 1662 1079
rect 1708 1157 1762 1353
rect 1808 1431 1862 1438
rect 1808 1379 1809 1431
rect 1861 1379 1862 1431
rect 1808 1353 1818 1379
rect 1852 1353 1862 1379
rect 1808 1341 1862 1353
rect 1908 1387 1962 1493
rect 2008 1527 2062 1539
rect 2008 1501 2018 1527
rect 2052 1501 2062 1527
rect 2008 1449 2009 1501
rect 2061 1449 2062 1501
rect 2008 1442 2062 1449
rect 2108 1527 2162 1633
rect 2208 1711 2262 1718
rect 2208 1659 2209 1711
rect 2261 1659 2262 1711
rect 2208 1633 2218 1659
rect 2252 1633 2262 1659
rect 2208 1621 2262 1633
rect 2308 1667 2362 1773
rect 2408 1807 2462 1819
rect 2408 1781 2418 1807
rect 2452 1781 2462 1807
rect 2408 1729 2409 1781
rect 2461 1729 2462 1781
rect 2408 1722 2462 1729
rect 2508 1807 2562 1913
rect 2608 1991 2662 1998
rect 2608 1939 2609 1991
rect 2661 1939 2662 1991
rect 2608 1913 2618 1939
rect 2652 1913 2662 1939
rect 2608 1901 2662 1913
rect 2708 1947 2762 2053
rect 2808 2087 2862 2099
rect 2808 2061 2818 2087
rect 2852 2061 2862 2087
rect 2808 2009 2809 2061
rect 2861 2009 2862 2061
rect 2808 2002 2862 2009
rect 2908 2087 2962 2193
rect 3008 2271 3062 2278
rect 3008 2219 3009 2271
rect 3061 2219 3062 2271
rect 3008 2193 3018 2219
rect 3052 2193 3062 2219
rect 3008 2181 3062 2193
rect 3108 2227 3162 2333
rect 3208 2367 3262 2379
rect 3208 2341 3218 2367
rect 3252 2341 3262 2367
rect 3208 2289 3209 2341
rect 3261 2289 3262 2341
rect 3208 2282 3262 2289
rect 3308 2367 3362 2563
rect 3408 2641 3462 2648
rect 3408 2589 3409 2641
rect 3461 2589 3462 2641
rect 3408 2563 3418 2589
rect 3452 2563 3462 2589
rect 3408 2551 3462 2563
rect 3508 2597 3562 2703
rect 3608 2737 3662 2749
rect 3608 2711 3618 2737
rect 3652 2711 3662 2737
rect 3608 2659 3609 2711
rect 3661 2659 3662 2711
rect 3608 2652 3662 2659
rect 3708 2737 3762 2843
rect 3808 2921 3862 2928
rect 3808 2869 3809 2921
rect 3861 2869 3862 2921
rect 3808 2843 3818 2869
rect 3852 2843 3862 2869
rect 3808 2831 3862 2843
rect 3908 2877 3962 2983
rect 4008 3017 4062 3029
rect 4008 2991 4018 3017
rect 4052 2991 4062 3017
rect 4008 2939 4009 2991
rect 4061 2939 4062 2991
rect 4008 2932 4062 2939
rect 4108 3017 4162 3123
rect 4208 3201 4262 3208
rect 4208 3149 4209 3201
rect 4261 3149 4262 3201
rect 4208 3123 4218 3149
rect 4252 3123 4262 3149
rect 4208 3111 4262 3123
rect 4308 3157 4362 3263
rect 4408 3297 4462 3309
rect 4408 3271 4418 3297
rect 4452 3271 4462 3297
rect 4408 3219 4409 3271
rect 4461 3219 4462 3271
rect 4408 3212 4462 3219
rect 4508 3297 4562 3403
rect 4608 3481 4662 3488
rect 4608 3429 4609 3481
rect 4661 3429 4662 3481
rect 4608 3403 4618 3429
rect 4652 3403 4662 3429
rect 4608 3391 4662 3403
rect 4708 3437 4762 3543
rect 4808 3577 4862 3589
rect 4808 3551 4818 3577
rect 4852 3551 4862 3577
rect 4808 3499 4809 3551
rect 4861 3499 4862 3551
rect 4808 3492 4862 3499
rect 4908 3577 4962 3773
rect 5008 3851 5062 3858
rect 5008 3799 5009 3851
rect 5061 3799 5062 3851
rect 5008 3773 5018 3799
rect 5052 3773 5062 3799
rect 5008 3761 5062 3773
rect 5108 3807 5162 3913
rect 5208 3947 5262 3959
rect 5208 3921 5218 3947
rect 5252 3921 5262 3947
rect 5208 3869 5209 3921
rect 5261 3869 5262 3921
rect 5208 3862 5262 3869
rect 5308 3947 5362 4053
rect 5408 4131 5462 4138
rect 5408 4079 5409 4131
rect 5461 4079 5462 4131
rect 5408 4053 5418 4079
rect 5452 4053 5462 4079
rect 5408 4041 5462 4053
rect 5508 4087 5562 4193
rect 5608 4227 5662 4239
rect 5608 4201 5618 4227
rect 5652 4201 5662 4227
rect 5608 4149 5609 4201
rect 5661 4149 5662 4201
rect 5608 4142 5662 4149
rect 5708 4227 5762 4333
rect 5808 4411 5862 4418
rect 5808 4359 5809 4411
rect 5861 4359 5862 4411
rect 5808 4333 5818 4359
rect 5852 4333 5862 4359
rect 5808 4321 5862 4333
rect 5908 4367 5962 4473
rect 6008 4507 6062 4519
rect 6008 4481 6018 4507
rect 6052 4481 6062 4507
rect 6008 4429 6009 4481
rect 6061 4429 6062 4481
rect 6008 4422 6062 4429
rect 6108 4507 6162 4613
rect 6208 4691 6262 4698
rect 6208 4639 6209 4691
rect 6261 4639 6262 4691
rect 6208 4613 6218 4639
rect 6252 4613 6262 4639
rect 6208 4601 6262 4613
rect 6308 4647 6362 4753
rect 6408 4787 6462 4799
rect 6408 4761 6418 4787
rect 6452 4761 6462 4787
rect 6408 4709 6409 4761
rect 6461 4709 6462 4761
rect 6408 4702 6462 4709
rect 6508 4787 6562 4960
rect 6602 4919 6668 4920
rect 6602 4867 6609 4919
rect 6661 4867 6668 4919
rect 6602 4866 6668 4867
rect 6508 4753 6518 4787
rect 6552 4753 6562 4787
rect 6308 4613 6318 4647
rect 6352 4613 6362 4647
rect 6108 4473 6118 4507
rect 6152 4473 6162 4507
rect 5908 4333 5918 4367
rect 5952 4333 5962 4367
rect 5708 4193 5718 4227
rect 5752 4193 5762 4227
rect 5508 4053 5518 4087
rect 5552 4053 5562 4087
rect 5308 3913 5318 3947
rect 5352 3913 5362 3947
rect 5108 3773 5118 3807
rect 5152 3773 5162 3807
rect 5002 3709 5068 3710
rect 5002 3657 5009 3709
rect 5061 3657 5068 3709
rect 5002 3656 5068 3657
rect 4908 3543 4918 3577
rect 4952 3543 4962 3577
rect 4708 3403 4718 3437
rect 4752 3403 4762 3437
rect 4508 3263 4518 3297
rect 4552 3263 4562 3297
rect 4308 3123 4318 3157
rect 4352 3123 4362 3157
rect 4108 2983 4118 3017
rect 4152 2983 4162 3017
rect 3908 2843 3918 2877
rect 3952 2843 3962 2877
rect 3708 2703 3718 2737
rect 3752 2703 3762 2737
rect 3508 2563 3518 2597
rect 3552 2563 3562 2597
rect 3402 2499 3468 2500
rect 3402 2447 3409 2499
rect 3461 2447 3468 2499
rect 3402 2446 3468 2447
rect 3308 2333 3318 2367
rect 3352 2333 3362 2367
rect 3108 2193 3118 2227
rect 3152 2193 3162 2227
rect 2908 2053 2918 2087
rect 2952 2053 2962 2087
rect 2708 1913 2718 1947
rect 2752 1913 2762 1947
rect 2508 1773 2518 1807
rect 2552 1773 2562 1807
rect 2308 1633 2318 1667
rect 2352 1633 2362 1667
rect 2108 1493 2118 1527
rect 2152 1493 2162 1527
rect 1908 1353 1918 1387
rect 1952 1353 1962 1387
rect 1802 1289 1868 1290
rect 1802 1237 1809 1289
rect 1861 1237 1868 1289
rect 1802 1236 1868 1237
rect 1708 1123 1718 1157
rect 1752 1123 1762 1157
rect 1508 983 1518 1017
rect 1552 983 1562 1017
rect 1308 843 1318 877
rect 1352 843 1362 877
rect 1108 703 1118 737
rect 1152 703 1162 737
rect 908 563 918 597
rect 952 563 962 597
rect 708 423 718 457
rect 752 423 762 457
rect 508 283 518 317
rect 552 283 562 317
rect 308 143 318 177
rect 352 143 362 177
rect 202 79 268 80
rect 202 27 209 79
rect 261 27 268 79
rect 202 26 268 27
rect 108 -67 109 -15
rect 161 -67 162 -15
rect 108 -79 118 -67
rect 152 -79 162 -67
rect -92 -132 -38 -131
rect -92 -143 -82 -132
rect -48 -143 -38 -132
rect -92 -195 -91 -143
rect -39 -195 -38 -143
rect -92 -210 -38 -195
rect 12 -133 58 -81
rect 12 -167 18 -133
rect 52 -167 58 -133
rect -82 -291 -75 -239
rect -23 -291 -16 -239
rect -91 -326 -39 -320
rect -91 -390 -82 -378
rect -48 -390 -39 -378
rect -91 -454 -82 -442
rect -48 -454 -39 -442
rect -91 -555 -39 -506
rect 12 -363 58 -167
rect 108 -131 109 -79
rect 161 -131 162 -79
rect 208 -22 262 26
rect 208 -74 209 -22
rect 261 -74 262 -22
rect 208 -81 262 -74
rect 308 -15 362 143
rect 408 177 462 189
rect 408 151 418 177
rect 452 151 462 177
rect 408 99 409 151
rect 461 99 462 151
rect 408 92 462 99
rect 508 177 562 283
rect 608 361 662 368
rect 608 309 609 361
rect 661 309 662 361
rect 608 283 618 309
rect 652 283 662 309
rect 608 271 662 283
rect 708 317 762 423
rect 808 457 862 469
rect 808 431 818 457
rect 852 431 862 457
rect 808 379 809 431
rect 861 379 862 431
rect 808 372 862 379
rect 908 457 962 563
rect 1008 641 1062 648
rect 1008 589 1009 641
rect 1061 589 1062 641
rect 1008 563 1018 589
rect 1052 563 1062 589
rect 1008 551 1062 563
rect 1108 597 1162 703
rect 1208 737 1262 749
rect 1208 711 1218 737
rect 1252 711 1262 737
rect 1208 659 1209 711
rect 1261 659 1262 711
rect 1208 652 1262 659
rect 1308 737 1362 843
rect 1408 921 1462 928
rect 1408 869 1409 921
rect 1461 869 1462 921
rect 1408 843 1418 869
rect 1452 843 1462 869
rect 1408 831 1462 843
rect 1508 877 1562 983
rect 1608 1017 1662 1029
rect 1608 991 1618 1017
rect 1652 991 1662 1017
rect 1608 939 1609 991
rect 1661 939 1662 991
rect 1608 932 1662 939
rect 1708 1017 1762 1123
rect 1808 1201 1862 1208
rect 1808 1149 1809 1201
rect 1861 1149 1862 1201
rect 1808 1123 1818 1149
rect 1852 1123 1862 1149
rect 1808 1111 1862 1123
rect 1908 1157 1962 1353
rect 2008 1387 2062 1399
rect 2008 1361 2018 1387
rect 2052 1361 2062 1387
rect 2008 1309 2009 1361
rect 2061 1309 2062 1361
rect 2008 1302 2062 1309
rect 2108 1387 2162 1493
rect 2208 1571 2262 1578
rect 2208 1519 2209 1571
rect 2261 1519 2262 1571
rect 2208 1493 2218 1519
rect 2252 1493 2262 1519
rect 2208 1481 2262 1493
rect 2308 1527 2362 1633
rect 2408 1667 2462 1679
rect 2408 1641 2418 1667
rect 2452 1641 2462 1667
rect 2408 1589 2409 1641
rect 2461 1589 2462 1641
rect 2408 1582 2462 1589
rect 2508 1667 2562 1773
rect 2608 1851 2662 1858
rect 2608 1799 2609 1851
rect 2661 1799 2662 1851
rect 2608 1773 2618 1799
rect 2652 1773 2662 1799
rect 2608 1761 2662 1773
rect 2708 1807 2762 1913
rect 2808 1947 2862 1959
rect 2808 1921 2818 1947
rect 2852 1921 2862 1947
rect 2808 1869 2809 1921
rect 2861 1869 2862 1921
rect 2808 1862 2862 1869
rect 2908 1947 2962 2053
rect 3008 2131 3062 2138
rect 3008 2079 3009 2131
rect 3061 2079 3062 2131
rect 3008 2053 3018 2079
rect 3052 2053 3062 2079
rect 3008 2041 3062 2053
rect 3108 2087 3162 2193
rect 3208 2227 3262 2239
rect 3208 2201 3218 2227
rect 3252 2201 3262 2227
rect 3208 2149 3209 2201
rect 3261 2149 3262 2201
rect 3208 2142 3262 2149
rect 3308 2227 3362 2333
rect 3408 2411 3462 2418
rect 3408 2359 3409 2411
rect 3461 2359 3462 2411
rect 3408 2333 3418 2359
rect 3452 2333 3462 2359
rect 3408 2321 3462 2333
rect 3508 2367 3562 2563
rect 3608 2597 3662 2609
rect 3608 2571 3618 2597
rect 3652 2571 3662 2597
rect 3608 2519 3609 2571
rect 3661 2519 3662 2571
rect 3608 2512 3662 2519
rect 3708 2597 3762 2703
rect 3808 2781 3862 2788
rect 3808 2729 3809 2781
rect 3861 2729 3862 2781
rect 3808 2703 3818 2729
rect 3852 2703 3862 2729
rect 3808 2691 3862 2703
rect 3908 2737 3962 2843
rect 4008 2877 4062 2889
rect 4008 2851 4018 2877
rect 4052 2851 4062 2877
rect 4008 2799 4009 2851
rect 4061 2799 4062 2851
rect 4008 2792 4062 2799
rect 4108 2877 4162 2983
rect 4208 3061 4262 3068
rect 4208 3009 4209 3061
rect 4261 3009 4262 3061
rect 4208 2983 4218 3009
rect 4252 2983 4262 3009
rect 4208 2971 4262 2983
rect 4308 3017 4362 3123
rect 4408 3157 4462 3169
rect 4408 3131 4418 3157
rect 4452 3131 4462 3157
rect 4408 3079 4409 3131
rect 4461 3079 4462 3131
rect 4408 3072 4462 3079
rect 4508 3157 4562 3263
rect 4608 3341 4662 3348
rect 4608 3289 4609 3341
rect 4661 3289 4662 3341
rect 4608 3263 4618 3289
rect 4652 3263 4662 3289
rect 4608 3251 4662 3263
rect 4708 3297 4762 3403
rect 4808 3437 4862 3449
rect 4808 3411 4818 3437
rect 4852 3411 4862 3437
rect 4808 3359 4809 3411
rect 4861 3359 4862 3411
rect 4808 3352 4862 3359
rect 4908 3437 4962 3543
rect 5008 3621 5062 3628
rect 5008 3569 5009 3621
rect 5061 3569 5062 3621
rect 5008 3543 5018 3569
rect 5052 3543 5062 3569
rect 5008 3531 5062 3543
rect 5108 3577 5162 3773
rect 5208 3807 5262 3819
rect 5208 3781 5218 3807
rect 5252 3781 5262 3807
rect 5208 3729 5209 3781
rect 5261 3729 5262 3781
rect 5208 3722 5262 3729
rect 5308 3807 5362 3913
rect 5408 3991 5462 3998
rect 5408 3939 5409 3991
rect 5461 3939 5462 3991
rect 5408 3913 5418 3939
rect 5452 3913 5462 3939
rect 5408 3901 5462 3913
rect 5508 3947 5562 4053
rect 5608 4087 5662 4099
rect 5608 4061 5618 4087
rect 5652 4061 5662 4087
rect 5608 4009 5609 4061
rect 5661 4009 5662 4061
rect 5608 4002 5662 4009
rect 5708 4087 5762 4193
rect 5808 4271 5862 4278
rect 5808 4219 5809 4271
rect 5861 4219 5862 4271
rect 5808 4193 5818 4219
rect 5852 4193 5862 4219
rect 5808 4181 5862 4193
rect 5908 4227 5962 4333
rect 6008 4367 6062 4379
rect 6008 4341 6018 4367
rect 6052 4341 6062 4367
rect 6008 4289 6009 4341
rect 6061 4289 6062 4341
rect 6008 4282 6062 4289
rect 6108 4367 6162 4473
rect 6208 4551 6262 4558
rect 6208 4499 6209 4551
rect 6261 4499 6262 4551
rect 6208 4473 6218 4499
rect 6252 4473 6262 4499
rect 6208 4461 6262 4473
rect 6308 4507 6362 4613
rect 6408 4647 6462 4659
rect 6408 4621 6418 4647
rect 6452 4621 6462 4647
rect 6408 4569 6409 4621
rect 6461 4569 6462 4621
rect 6408 4562 6462 4569
rect 6508 4647 6562 4753
rect 6608 4831 6662 4838
rect 6608 4779 6609 4831
rect 6661 4779 6662 4831
rect 6608 4753 6618 4779
rect 6652 4753 6662 4779
rect 6608 4741 6662 4753
rect 6708 4787 6762 4960
rect 6802 4903 6868 4904
rect 6802 4851 6809 4903
rect 6861 4851 6868 4903
rect 6802 4850 6868 4851
rect 6708 4753 6718 4787
rect 6752 4753 6762 4787
rect 6508 4613 6518 4647
rect 6552 4613 6562 4647
rect 6308 4473 6318 4507
rect 6352 4473 6362 4507
rect 6108 4333 6118 4367
rect 6152 4333 6162 4367
rect 5908 4193 5918 4227
rect 5952 4193 5962 4227
rect 5708 4053 5718 4087
rect 5752 4053 5762 4087
rect 5508 3913 5518 3947
rect 5552 3913 5562 3947
rect 5308 3773 5318 3807
rect 5352 3773 5362 3807
rect 5202 3693 5268 3694
rect 5202 3641 5209 3693
rect 5261 3641 5268 3693
rect 5202 3640 5268 3641
rect 5108 3543 5118 3577
rect 5152 3543 5162 3577
rect 4908 3403 4918 3437
rect 4952 3403 4962 3437
rect 4708 3263 4718 3297
rect 4752 3263 4762 3297
rect 4508 3123 4518 3157
rect 4552 3123 4562 3157
rect 4308 2983 4318 3017
rect 4352 2983 4362 3017
rect 4108 2843 4118 2877
rect 4152 2843 4162 2877
rect 3908 2703 3918 2737
rect 3952 2703 3962 2737
rect 3708 2563 3718 2597
rect 3752 2563 3762 2597
rect 3602 2483 3668 2484
rect 3602 2431 3609 2483
rect 3661 2431 3668 2483
rect 3602 2430 3668 2431
rect 3508 2333 3518 2367
rect 3552 2333 3562 2367
rect 3308 2193 3318 2227
rect 3352 2193 3362 2227
rect 3108 2053 3118 2087
rect 3152 2053 3162 2087
rect 2908 1913 2918 1947
rect 2952 1913 2962 1947
rect 2708 1773 2718 1807
rect 2752 1773 2762 1807
rect 2508 1633 2518 1667
rect 2552 1633 2562 1667
rect 2308 1493 2318 1527
rect 2352 1493 2362 1527
rect 2108 1353 2118 1387
rect 2152 1353 2162 1387
rect 2002 1273 2068 1274
rect 2002 1221 2009 1273
rect 2061 1221 2068 1273
rect 2002 1220 2068 1221
rect 1908 1123 1918 1157
rect 1952 1123 1962 1157
rect 1708 983 1718 1017
rect 1752 983 1762 1017
rect 1508 843 1518 877
rect 1552 843 1562 877
rect 1308 703 1318 737
rect 1352 703 1362 737
rect 1108 563 1118 597
rect 1152 563 1162 597
rect 908 423 918 457
rect 952 423 962 457
rect 708 283 718 317
rect 752 283 762 317
rect 508 143 518 177
rect 552 143 562 177
rect 402 63 468 64
rect 402 11 409 63
rect 461 11 468 63
rect 402 10 468 11
rect 308 -67 309 -15
rect 361 -67 362 -15
rect 308 -79 318 -67
rect 352 -79 362 -67
rect 108 -132 162 -131
rect 108 -143 118 -132
rect 152 -143 162 -132
rect 108 -195 109 -143
rect 161 -195 162 -143
rect 108 -210 162 -195
rect 212 -133 258 -81
rect 212 -167 218 -133
rect 252 -167 258 -133
rect 118 -291 125 -239
rect 177 -291 184 -239
rect 12 -397 18 -363
rect 52 -397 58 -363
rect 12 -435 58 -397
rect 12 -469 18 -435
rect 52 -469 58 -435
rect 12 -512 58 -469
rect 109 -326 161 -320
rect 109 -390 118 -378
rect 152 -390 161 -378
rect 109 -454 118 -442
rect 152 -454 161 -442
rect 109 -512 161 -506
rect 212 -363 258 -167
rect 308 -131 309 -79
rect 361 -131 362 -79
rect 408 -22 462 10
rect 408 -74 409 -22
rect 461 -74 462 -22
rect 408 -81 462 -74
rect 508 -15 562 143
rect 608 221 662 228
rect 608 169 609 221
rect 661 169 662 221
rect 608 143 618 169
rect 652 143 662 169
rect 608 131 662 143
rect 708 177 762 283
rect 808 317 862 329
rect 808 291 818 317
rect 852 291 862 317
rect 808 239 809 291
rect 861 239 862 291
rect 808 232 862 239
rect 908 317 962 423
rect 1008 501 1062 508
rect 1008 449 1009 501
rect 1061 449 1062 501
rect 1008 423 1018 449
rect 1052 423 1062 449
rect 1008 411 1062 423
rect 1108 457 1162 563
rect 1208 597 1262 609
rect 1208 571 1218 597
rect 1252 571 1262 597
rect 1208 519 1209 571
rect 1261 519 1262 571
rect 1208 512 1262 519
rect 1308 597 1362 703
rect 1408 781 1462 788
rect 1408 729 1409 781
rect 1461 729 1462 781
rect 1408 703 1418 729
rect 1452 703 1462 729
rect 1408 691 1462 703
rect 1508 737 1562 843
rect 1608 877 1662 889
rect 1608 851 1618 877
rect 1652 851 1662 877
rect 1608 799 1609 851
rect 1661 799 1662 851
rect 1608 792 1662 799
rect 1708 877 1762 983
rect 1808 1061 1862 1068
rect 1808 1009 1809 1061
rect 1861 1009 1862 1061
rect 1808 983 1818 1009
rect 1852 983 1862 1009
rect 1808 971 1862 983
rect 1908 1017 1962 1123
rect 2008 1157 2062 1169
rect 2008 1131 2018 1157
rect 2052 1131 2062 1157
rect 2008 1079 2009 1131
rect 2061 1079 2062 1131
rect 2008 1072 2062 1079
rect 2108 1157 2162 1353
rect 2208 1431 2262 1438
rect 2208 1379 2209 1431
rect 2261 1379 2262 1431
rect 2208 1353 2218 1379
rect 2252 1353 2262 1379
rect 2208 1341 2262 1353
rect 2308 1387 2362 1493
rect 2408 1527 2462 1539
rect 2408 1501 2418 1527
rect 2452 1501 2462 1527
rect 2408 1449 2409 1501
rect 2461 1449 2462 1501
rect 2408 1442 2462 1449
rect 2508 1527 2562 1633
rect 2608 1711 2662 1718
rect 2608 1659 2609 1711
rect 2661 1659 2662 1711
rect 2608 1633 2618 1659
rect 2652 1633 2662 1659
rect 2608 1621 2662 1633
rect 2708 1667 2762 1773
rect 2808 1807 2862 1819
rect 2808 1781 2818 1807
rect 2852 1781 2862 1807
rect 2808 1729 2809 1781
rect 2861 1729 2862 1781
rect 2808 1722 2862 1729
rect 2908 1807 2962 1913
rect 3008 1991 3062 1998
rect 3008 1939 3009 1991
rect 3061 1939 3062 1991
rect 3008 1913 3018 1939
rect 3052 1913 3062 1939
rect 3008 1901 3062 1913
rect 3108 1947 3162 2053
rect 3208 2087 3262 2099
rect 3208 2061 3218 2087
rect 3252 2061 3262 2087
rect 3208 2009 3209 2061
rect 3261 2009 3262 2061
rect 3208 2002 3262 2009
rect 3308 2087 3362 2193
rect 3408 2271 3462 2278
rect 3408 2219 3409 2271
rect 3461 2219 3462 2271
rect 3408 2193 3418 2219
rect 3452 2193 3462 2219
rect 3408 2181 3462 2193
rect 3508 2227 3562 2333
rect 3608 2367 3662 2379
rect 3608 2341 3618 2367
rect 3652 2341 3662 2367
rect 3608 2289 3609 2341
rect 3661 2289 3662 2341
rect 3608 2282 3662 2289
rect 3708 2367 3762 2563
rect 3808 2641 3862 2648
rect 3808 2589 3809 2641
rect 3861 2589 3862 2641
rect 3808 2563 3818 2589
rect 3852 2563 3862 2589
rect 3808 2551 3862 2563
rect 3908 2597 3962 2703
rect 4008 2737 4062 2749
rect 4008 2711 4018 2737
rect 4052 2711 4062 2737
rect 4008 2659 4009 2711
rect 4061 2659 4062 2711
rect 4008 2652 4062 2659
rect 4108 2737 4162 2843
rect 4208 2921 4262 2928
rect 4208 2869 4209 2921
rect 4261 2869 4262 2921
rect 4208 2843 4218 2869
rect 4252 2843 4262 2869
rect 4208 2831 4262 2843
rect 4308 2877 4362 2983
rect 4408 3017 4462 3029
rect 4408 2991 4418 3017
rect 4452 2991 4462 3017
rect 4408 2939 4409 2991
rect 4461 2939 4462 2991
rect 4408 2932 4462 2939
rect 4508 3017 4562 3123
rect 4608 3201 4662 3208
rect 4608 3149 4609 3201
rect 4661 3149 4662 3201
rect 4608 3123 4618 3149
rect 4652 3123 4662 3149
rect 4608 3111 4662 3123
rect 4708 3157 4762 3263
rect 4808 3297 4862 3309
rect 4808 3271 4818 3297
rect 4852 3271 4862 3297
rect 4808 3219 4809 3271
rect 4861 3219 4862 3271
rect 4808 3212 4862 3219
rect 4908 3297 4962 3403
rect 5008 3481 5062 3488
rect 5008 3429 5009 3481
rect 5061 3429 5062 3481
rect 5008 3403 5018 3429
rect 5052 3403 5062 3429
rect 5008 3391 5062 3403
rect 5108 3437 5162 3543
rect 5208 3577 5262 3589
rect 5208 3551 5218 3577
rect 5252 3551 5262 3577
rect 5208 3499 5209 3551
rect 5261 3499 5262 3551
rect 5208 3492 5262 3499
rect 5308 3577 5362 3773
rect 5408 3851 5462 3858
rect 5408 3799 5409 3851
rect 5461 3799 5462 3851
rect 5408 3773 5418 3799
rect 5452 3773 5462 3799
rect 5408 3761 5462 3773
rect 5508 3807 5562 3913
rect 5608 3947 5662 3959
rect 5608 3921 5618 3947
rect 5652 3921 5662 3947
rect 5608 3869 5609 3921
rect 5661 3869 5662 3921
rect 5608 3862 5662 3869
rect 5708 3947 5762 4053
rect 5808 4131 5862 4138
rect 5808 4079 5809 4131
rect 5861 4079 5862 4131
rect 5808 4053 5818 4079
rect 5852 4053 5862 4079
rect 5808 4041 5862 4053
rect 5908 4087 5962 4193
rect 6008 4227 6062 4239
rect 6008 4201 6018 4227
rect 6052 4201 6062 4227
rect 6008 4149 6009 4201
rect 6061 4149 6062 4201
rect 6008 4142 6062 4149
rect 6108 4227 6162 4333
rect 6208 4411 6262 4418
rect 6208 4359 6209 4411
rect 6261 4359 6262 4411
rect 6208 4333 6218 4359
rect 6252 4333 6262 4359
rect 6208 4321 6262 4333
rect 6308 4367 6362 4473
rect 6408 4507 6462 4519
rect 6408 4481 6418 4507
rect 6452 4481 6462 4507
rect 6408 4429 6409 4481
rect 6461 4429 6462 4481
rect 6408 4422 6462 4429
rect 6508 4507 6562 4613
rect 6608 4691 6662 4698
rect 6608 4639 6609 4691
rect 6661 4639 6662 4691
rect 6608 4613 6618 4639
rect 6652 4613 6662 4639
rect 6608 4601 6662 4613
rect 6708 4647 6762 4753
rect 6808 4787 6862 4799
rect 6808 4761 6818 4787
rect 6852 4761 6862 4787
rect 6808 4709 6809 4761
rect 6861 4709 6862 4761
rect 6808 4702 6862 4709
rect 6908 4787 6962 4960
rect 7002 4919 7068 4920
rect 7002 4867 7009 4919
rect 7061 4867 7068 4919
rect 7002 4866 7068 4867
rect 6908 4753 6918 4787
rect 6952 4753 6962 4787
rect 6708 4613 6718 4647
rect 6752 4613 6762 4647
rect 6508 4473 6518 4507
rect 6552 4473 6562 4507
rect 6308 4333 6318 4367
rect 6352 4333 6362 4367
rect 6108 4193 6118 4227
rect 6152 4193 6162 4227
rect 5908 4053 5918 4087
rect 5952 4053 5962 4087
rect 5708 3913 5718 3947
rect 5752 3913 5762 3947
rect 5508 3773 5518 3807
rect 5552 3773 5562 3807
rect 5402 3709 5468 3710
rect 5402 3657 5409 3709
rect 5461 3657 5468 3709
rect 5402 3656 5468 3657
rect 5308 3543 5318 3577
rect 5352 3543 5362 3577
rect 5108 3403 5118 3437
rect 5152 3403 5162 3437
rect 4908 3263 4918 3297
rect 4952 3263 4962 3297
rect 4708 3123 4718 3157
rect 4752 3123 4762 3157
rect 4508 2983 4518 3017
rect 4552 2983 4562 3017
rect 4308 2843 4318 2877
rect 4352 2843 4362 2877
rect 4108 2703 4118 2737
rect 4152 2703 4162 2737
rect 3908 2563 3918 2597
rect 3952 2563 3962 2597
rect 3802 2499 3868 2500
rect 3802 2447 3809 2499
rect 3861 2447 3868 2499
rect 3802 2446 3868 2447
rect 3708 2333 3718 2367
rect 3752 2333 3762 2367
rect 3508 2193 3518 2227
rect 3552 2193 3562 2227
rect 3308 2053 3318 2087
rect 3352 2053 3362 2087
rect 3108 1913 3118 1947
rect 3152 1913 3162 1947
rect 2908 1773 2918 1807
rect 2952 1773 2962 1807
rect 2708 1633 2718 1667
rect 2752 1633 2762 1667
rect 2508 1493 2518 1527
rect 2552 1493 2562 1527
rect 2308 1353 2318 1387
rect 2352 1353 2362 1387
rect 2202 1289 2268 1290
rect 2202 1237 2209 1289
rect 2261 1237 2268 1289
rect 2202 1236 2268 1237
rect 2108 1123 2118 1157
rect 2152 1123 2162 1157
rect 1908 983 1918 1017
rect 1952 983 1962 1017
rect 1708 843 1718 877
rect 1752 843 1762 877
rect 1508 703 1518 737
rect 1552 703 1562 737
rect 1308 563 1318 597
rect 1352 563 1362 597
rect 1108 423 1118 457
rect 1152 423 1162 457
rect 908 283 918 317
rect 952 283 962 317
rect 708 143 718 177
rect 752 143 762 177
rect 602 79 668 80
rect 602 27 609 79
rect 661 27 668 79
rect 602 26 668 27
rect 508 -67 509 -15
rect 561 -67 562 -15
rect 508 -79 518 -67
rect 552 -79 562 -67
rect 308 -132 362 -131
rect 308 -143 318 -132
rect 352 -143 362 -132
rect 308 -195 309 -143
rect 361 -195 362 -143
rect 308 -210 362 -195
rect 412 -133 458 -81
rect 412 -167 418 -133
rect 452 -167 458 -133
rect 318 -291 325 -239
rect 377 -291 384 -239
rect 212 -397 218 -363
rect 252 -397 258 -363
rect 212 -435 258 -397
rect 212 -469 218 -435
rect 252 -469 258 -435
rect 212 -512 258 -469
rect 309 -326 361 -320
rect 309 -390 318 -378
rect 352 -390 361 -378
rect 309 -454 318 -442
rect 352 -454 361 -442
rect 309 -555 361 -506
rect 412 -363 458 -167
rect 508 -131 509 -79
rect 561 -131 562 -79
rect 608 -22 662 26
rect 608 -74 609 -22
rect 661 -74 662 -22
rect 608 -81 662 -74
rect 708 -15 762 143
rect 808 177 862 189
rect 808 151 818 177
rect 852 151 862 177
rect 808 99 809 151
rect 861 99 862 151
rect 808 92 862 99
rect 908 177 962 283
rect 1008 361 1062 368
rect 1008 309 1009 361
rect 1061 309 1062 361
rect 1008 283 1018 309
rect 1052 283 1062 309
rect 1008 271 1062 283
rect 1108 317 1162 423
rect 1208 457 1262 469
rect 1208 431 1218 457
rect 1252 431 1262 457
rect 1208 379 1209 431
rect 1261 379 1262 431
rect 1208 372 1262 379
rect 1308 457 1362 563
rect 1408 641 1462 648
rect 1408 589 1409 641
rect 1461 589 1462 641
rect 1408 563 1418 589
rect 1452 563 1462 589
rect 1408 551 1462 563
rect 1508 597 1562 703
rect 1608 737 1662 749
rect 1608 711 1618 737
rect 1652 711 1662 737
rect 1608 659 1609 711
rect 1661 659 1662 711
rect 1608 652 1662 659
rect 1708 737 1762 843
rect 1808 921 1862 928
rect 1808 869 1809 921
rect 1861 869 1862 921
rect 1808 843 1818 869
rect 1852 843 1862 869
rect 1808 831 1862 843
rect 1908 877 1962 983
rect 2008 1017 2062 1029
rect 2008 991 2018 1017
rect 2052 991 2062 1017
rect 2008 939 2009 991
rect 2061 939 2062 991
rect 2008 932 2062 939
rect 2108 1017 2162 1123
rect 2208 1201 2262 1208
rect 2208 1149 2209 1201
rect 2261 1149 2262 1201
rect 2208 1123 2218 1149
rect 2252 1123 2262 1149
rect 2208 1111 2262 1123
rect 2308 1157 2362 1353
rect 2408 1387 2462 1399
rect 2408 1361 2418 1387
rect 2452 1361 2462 1387
rect 2408 1309 2409 1361
rect 2461 1309 2462 1361
rect 2408 1302 2462 1309
rect 2508 1387 2562 1493
rect 2608 1571 2662 1578
rect 2608 1519 2609 1571
rect 2661 1519 2662 1571
rect 2608 1493 2618 1519
rect 2652 1493 2662 1519
rect 2608 1481 2662 1493
rect 2708 1527 2762 1633
rect 2808 1667 2862 1679
rect 2808 1641 2818 1667
rect 2852 1641 2862 1667
rect 2808 1589 2809 1641
rect 2861 1589 2862 1641
rect 2808 1582 2862 1589
rect 2908 1667 2962 1773
rect 3008 1851 3062 1858
rect 3008 1799 3009 1851
rect 3061 1799 3062 1851
rect 3008 1773 3018 1799
rect 3052 1773 3062 1799
rect 3008 1761 3062 1773
rect 3108 1807 3162 1913
rect 3208 1947 3262 1959
rect 3208 1921 3218 1947
rect 3252 1921 3262 1947
rect 3208 1869 3209 1921
rect 3261 1869 3262 1921
rect 3208 1862 3262 1869
rect 3308 1947 3362 2053
rect 3408 2131 3462 2138
rect 3408 2079 3409 2131
rect 3461 2079 3462 2131
rect 3408 2053 3418 2079
rect 3452 2053 3462 2079
rect 3408 2041 3462 2053
rect 3508 2087 3562 2193
rect 3608 2227 3662 2239
rect 3608 2201 3618 2227
rect 3652 2201 3662 2227
rect 3608 2149 3609 2201
rect 3661 2149 3662 2201
rect 3608 2142 3662 2149
rect 3708 2227 3762 2333
rect 3808 2411 3862 2418
rect 3808 2359 3809 2411
rect 3861 2359 3862 2411
rect 3808 2333 3818 2359
rect 3852 2333 3862 2359
rect 3808 2321 3862 2333
rect 3908 2367 3962 2563
rect 4008 2597 4062 2609
rect 4008 2571 4018 2597
rect 4052 2571 4062 2597
rect 4008 2519 4009 2571
rect 4061 2519 4062 2571
rect 4008 2512 4062 2519
rect 4108 2597 4162 2703
rect 4208 2781 4262 2788
rect 4208 2729 4209 2781
rect 4261 2729 4262 2781
rect 4208 2703 4218 2729
rect 4252 2703 4262 2729
rect 4208 2691 4262 2703
rect 4308 2737 4362 2843
rect 4408 2877 4462 2889
rect 4408 2851 4418 2877
rect 4452 2851 4462 2877
rect 4408 2799 4409 2851
rect 4461 2799 4462 2851
rect 4408 2792 4462 2799
rect 4508 2877 4562 2983
rect 4608 3061 4662 3068
rect 4608 3009 4609 3061
rect 4661 3009 4662 3061
rect 4608 2983 4618 3009
rect 4652 2983 4662 3009
rect 4608 2971 4662 2983
rect 4708 3017 4762 3123
rect 4808 3157 4862 3169
rect 4808 3131 4818 3157
rect 4852 3131 4862 3157
rect 4808 3079 4809 3131
rect 4861 3079 4862 3131
rect 4808 3072 4862 3079
rect 4908 3157 4962 3263
rect 5008 3341 5062 3348
rect 5008 3289 5009 3341
rect 5061 3289 5062 3341
rect 5008 3263 5018 3289
rect 5052 3263 5062 3289
rect 5008 3251 5062 3263
rect 5108 3297 5162 3403
rect 5208 3437 5262 3449
rect 5208 3411 5218 3437
rect 5252 3411 5262 3437
rect 5208 3359 5209 3411
rect 5261 3359 5262 3411
rect 5208 3352 5262 3359
rect 5308 3437 5362 3543
rect 5408 3621 5462 3628
rect 5408 3569 5409 3621
rect 5461 3569 5462 3621
rect 5408 3543 5418 3569
rect 5452 3543 5462 3569
rect 5408 3531 5462 3543
rect 5508 3577 5562 3773
rect 5608 3807 5662 3819
rect 5608 3781 5618 3807
rect 5652 3781 5662 3807
rect 5608 3729 5609 3781
rect 5661 3729 5662 3781
rect 5608 3722 5662 3729
rect 5708 3807 5762 3913
rect 5808 3991 5862 3998
rect 5808 3939 5809 3991
rect 5861 3939 5862 3991
rect 5808 3913 5818 3939
rect 5852 3913 5862 3939
rect 5808 3901 5862 3913
rect 5908 3947 5962 4053
rect 6008 4087 6062 4099
rect 6008 4061 6018 4087
rect 6052 4061 6062 4087
rect 6008 4009 6009 4061
rect 6061 4009 6062 4061
rect 6008 4002 6062 4009
rect 6108 4087 6162 4193
rect 6208 4271 6262 4278
rect 6208 4219 6209 4271
rect 6261 4219 6262 4271
rect 6208 4193 6218 4219
rect 6252 4193 6262 4219
rect 6208 4181 6262 4193
rect 6308 4227 6362 4333
rect 6408 4367 6462 4379
rect 6408 4341 6418 4367
rect 6452 4341 6462 4367
rect 6408 4289 6409 4341
rect 6461 4289 6462 4341
rect 6408 4282 6462 4289
rect 6508 4367 6562 4473
rect 6608 4551 6662 4558
rect 6608 4499 6609 4551
rect 6661 4499 6662 4551
rect 6608 4473 6618 4499
rect 6652 4473 6662 4499
rect 6608 4461 6662 4473
rect 6708 4507 6762 4613
rect 6808 4647 6862 4659
rect 6808 4621 6818 4647
rect 6852 4621 6862 4647
rect 6808 4569 6809 4621
rect 6861 4569 6862 4621
rect 6808 4562 6862 4569
rect 6908 4647 6962 4753
rect 7008 4831 7062 4838
rect 7008 4779 7009 4831
rect 7061 4779 7062 4831
rect 7008 4753 7018 4779
rect 7052 4753 7062 4779
rect 7008 4741 7062 4753
rect 7108 4787 7162 4960
rect 7202 4903 7268 4904
rect 7202 4851 7209 4903
rect 7261 4851 7268 4903
rect 7202 4850 7268 4851
rect 7108 4753 7118 4787
rect 7152 4753 7162 4787
rect 6908 4613 6918 4647
rect 6952 4613 6962 4647
rect 6708 4473 6718 4507
rect 6752 4473 6762 4507
rect 6508 4333 6518 4367
rect 6552 4333 6562 4367
rect 6308 4193 6318 4227
rect 6352 4193 6362 4227
rect 6108 4053 6118 4087
rect 6152 4053 6162 4087
rect 5908 3913 5918 3947
rect 5952 3913 5962 3947
rect 5708 3773 5718 3807
rect 5752 3773 5762 3807
rect 5602 3693 5668 3694
rect 5602 3641 5609 3693
rect 5661 3641 5668 3693
rect 5602 3640 5668 3641
rect 5508 3543 5518 3577
rect 5552 3543 5562 3577
rect 5308 3403 5318 3437
rect 5352 3403 5362 3437
rect 5108 3263 5118 3297
rect 5152 3263 5162 3297
rect 4908 3123 4918 3157
rect 4952 3123 4962 3157
rect 4708 2983 4718 3017
rect 4752 2983 4762 3017
rect 4508 2843 4518 2877
rect 4552 2843 4562 2877
rect 4308 2703 4318 2737
rect 4352 2703 4362 2737
rect 4108 2563 4118 2597
rect 4152 2563 4162 2597
rect 4002 2483 4068 2484
rect 4002 2431 4009 2483
rect 4061 2431 4068 2483
rect 4002 2430 4068 2431
rect 3908 2333 3918 2367
rect 3952 2333 3962 2367
rect 3708 2193 3718 2227
rect 3752 2193 3762 2227
rect 3508 2053 3518 2087
rect 3552 2053 3562 2087
rect 3308 1913 3318 1947
rect 3352 1913 3362 1947
rect 3108 1773 3118 1807
rect 3152 1773 3162 1807
rect 2908 1633 2918 1667
rect 2952 1633 2962 1667
rect 2708 1493 2718 1527
rect 2752 1493 2762 1527
rect 2508 1353 2518 1387
rect 2552 1353 2562 1387
rect 2402 1273 2468 1274
rect 2402 1221 2409 1273
rect 2461 1221 2468 1273
rect 2402 1220 2468 1221
rect 2308 1123 2318 1157
rect 2352 1123 2362 1157
rect 2108 983 2118 1017
rect 2152 983 2162 1017
rect 1908 843 1918 877
rect 1952 843 1962 877
rect 1708 703 1718 737
rect 1752 703 1762 737
rect 1508 563 1518 597
rect 1552 563 1562 597
rect 1308 423 1318 457
rect 1352 423 1362 457
rect 1108 283 1118 317
rect 1152 283 1162 317
rect 908 143 918 177
rect 952 143 962 177
rect 802 63 868 64
rect 802 11 809 63
rect 861 11 868 63
rect 802 10 868 11
rect 708 -67 709 -15
rect 761 -67 762 -15
rect 708 -79 718 -67
rect 752 -79 762 -67
rect 508 -132 562 -131
rect 508 -143 518 -132
rect 552 -143 562 -132
rect 508 -195 509 -143
rect 561 -195 562 -143
rect 508 -210 562 -195
rect 612 -133 658 -81
rect 612 -167 618 -133
rect 652 -167 658 -133
rect 518 -291 525 -239
rect 577 -291 584 -239
rect 412 -397 418 -363
rect 452 -397 458 -363
rect 412 -435 458 -397
rect 412 -469 418 -435
rect 452 -469 458 -435
rect 412 -512 458 -469
rect 509 -326 561 -320
rect 509 -390 518 -378
rect 552 -390 561 -378
rect 509 -454 518 -442
rect 552 -454 561 -442
rect 509 -512 561 -506
rect 612 -363 658 -167
rect 708 -131 709 -79
rect 761 -131 762 -79
rect 808 -22 862 10
rect 808 -74 809 -22
rect 861 -74 862 -22
rect 808 -81 862 -74
rect 908 -15 962 143
rect 1008 221 1062 228
rect 1008 169 1009 221
rect 1061 169 1062 221
rect 1008 143 1018 169
rect 1052 143 1062 169
rect 1008 131 1062 143
rect 1108 177 1162 283
rect 1208 317 1262 329
rect 1208 291 1218 317
rect 1252 291 1262 317
rect 1208 239 1209 291
rect 1261 239 1262 291
rect 1208 232 1262 239
rect 1308 317 1362 423
rect 1408 501 1462 508
rect 1408 449 1409 501
rect 1461 449 1462 501
rect 1408 423 1418 449
rect 1452 423 1462 449
rect 1408 411 1462 423
rect 1508 457 1562 563
rect 1608 597 1662 609
rect 1608 571 1618 597
rect 1652 571 1662 597
rect 1608 519 1609 571
rect 1661 519 1662 571
rect 1608 512 1662 519
rect 1708 597 1762 703
rect 1808 781 1862 788
rect 1808 729 1809 781
rect 1861 729 1862 781
rect 1808 703 1818 729
rect 1852 703 1862 729
rect 1808 691 1862 703
rect 1908 737 1962 843
rect 2008 877 2062 889
rect 2008 851 2018 877
rect 2052 851 2062 877
rect 2008 799 2009 851
rect 2061 799 2062 851
rect 2008 792 2062 799
rect 2108 877 2162 983
rect 2208 1061 2262 1068
rect 2208 1009 2209 1061
rect 2261 1009 2262 1061
rect 2208 983 2218 1009
rect 2252 983 2262 1009
rect 2208 971 2262 983
rect 2308 1017 2362 1123
rect 2408 1157 2462 1169
rect 2408 1131 2418 1157
rect 2452 1131 2462 1157
rect 2408 1079 2409 1131
rect 2461 1079 2462 1131
rect 2408 1072 2462 1079
rect 2508 1157 2562 1353
rect 2608 1431 2662 1438
rect 2608 1379 2609 1431
rect 2661 1379 2662 1431
rect 2608 1353 2618 1379
rect 2652 1353 2662 1379
rect 2608 1341 2662 1353
rect 2708 1387 2762 1493
rect 2808 1527 2862 1539
rect 2808 1501 2818 1527
rect 2852 1501 2862 1527
rect 2808 1449 2809 1501
rect 2861 1449 2862 1501
rect 2808 1442 2862 1449
rect 2908 1527 2962 1633
rect 3008 1711 3062 1718
rect 3008 1659 3009 1711
rect 3061 1659 3062 1711
rect 3008 1633 3018 1659
rect 3052 1633 3062 1659
rect 3008 1621 3062 1633
rect 3108 1667 3162 1773
rect 3208 1807 3262 1819
rect 3208 1781 3218 1807
rect 3252 1781 3262 1807
rect 3208 1729 3209 1781
rect 3261 1729 3262 1781
rect 3208 1722 3262 1729
rect 3308 1807 3362 1913
rect 3408 1991 3462 1998
rect 3408 1939 3409 1991
rect 3461 1939 3462 1991
rect 3408 1913 3418 1939
rect 3452 1913 3462 1939
rect 3408 1901 3462 1913
rect 3508 1947 3562 2053
rect 3608 2087 3662 2099
rect 3608 2061 3618 2087
rect 3652 2061 3662 2087
rect 3608 2009 3609 2061
rect 3661 2009 3662 2061
rect 3608 2002 3662 2009
rect 3708 2087 3762 2193
rect 3808 2271 3862 2278
rect 3808 2219 3809 2271
rect 3861 2219 3862 2271
rect 3808 2193 3818 2219
rect 3852 2193 3862 2219
rect 3808 2181 3862 2193
rect 3908 2227 3962 2333
rect 4008 2367 4062 2379
rect 4008 2341 4018 2367
rect 4052 2341 4062 2367
rect 4008 2289 4009 2341
rect 4061 2289 4062 2341
rect 4008 2282 4062 2289
rect 4108 2367 4162 2563
rect 4208 2641 4262 2648
rect 4208 2589 4209 2641
rect 4261 2589 4262 2641
rect 4208 2563 4218 2589
rect 4252 2563 4262 2589
rect 4208 2551 4262 2563
rect 4308 2597 4362 2703
rect 4408 2737 4462 2749
rect 4408 2711 4418 2737
rect 4452 2711 4462 2737
rect 4408 2659 4409 2711
rect 4461 2659 4462 2711
rect 4408 2652 4462 2659
rect 4508 2737 4562 2843
rect 4608 2921 4662 2928
rect 4608 2869 4609 2921
rect 4661 2869 4662 2921
rect 4608 2843 4618 2869
rect 4652 2843 4662 2869
rect 4608 2831 4662 2843
rect 4708 2877 4762 2983
rect 4808 3017 4862 3029
rect 4808 2991 4818 3017
rect 4852 2991 4862 3017
rect 4808 2939 4809 2991
rect 4861 2939 4862 2991
rect 4808 2932 4862 2939
rect 4908 3017 4962 3123
rect 5008 3201 5062 3208
rect 5008 3149 5009 3201
rect 5061 3149 5062 3201
rect 5008 3123 5018 3149
rect 5052 3123 5062 3149
rect 5008 3111 5062 3123
rect 5108 3157 5162 3263
rect 5208 3297 5262 3309
rect 5208 3271 5218 3297
rect 5252 3271 5262 3297
rect 5208 3219 5209 3271
rect 5261 3219 5262 3271
rect 5208 3212 5262 3219
rect 5308 3297 5362 3403
rect 5408 3481 5462 3488
rect 5408 3429 5409 3481
rect 5461 3429 5462 3481
rect 5408 3403 5418 3429
rect 5452 3403 5462 3429
rect 5408 3391 5462 3403
rect 5508 3437 5562 3543
rect 5608 3577 5662 3589
rect 5608 3551 5618 3577
rect 5652 3551 5662 3577
rect 5608 3499 5609 3551
rect 5661 3499 5662 3551
rect 5608 3492 5662 3499
rect 5708 3577 5762 3773
rect 5808 3851 5862 3858
rect 5808 3799 5809 3851
rect 5861 3799 5862 3851
rect 5808 3773 5818 3799
rect 5852 3773 5862 3799
rect 5808 3761 5862 3773
rect 5908 3807 5962 3913
rect 6008 3947 6062 3959
rect 6008 3921 6018 3947
rect 6052 3921 6062 3947
rect 6008 3869 6009 3921
rect 6061 3869 6062 3921
rect 6008 3862 6062 3869
rect 6108 3947 6162 4053
rect 6208 4131 6262 4138
rect 6208 4079 6209 4131
rect 6261 4079 6262 4131
rect 6208 4053 6218 4079
rect 6252 4053 6262 4079
rect 6208 4041 6262 4053
rect 6308 4087 6362 4193
rect 6408 4227 6462 4239
rect 6408 4201 6418 4227
rect 6452 4201 6462 4227
rect 6408 4149 6409 4201
rect 6461 4149 6462 4201
rect 6408 4142 6462 4149
rect 6508 4227 6562 4333
rect 6608 4411 6662 4418
rect 6608 4359 6609 4411
rect 6661 4359 6662 4411
rect 6608 4333 6618 4359
rect 6652 4333 6662 4359
rect 6608 4321 6662 4333
rect 6708 4367 6762 4473
rect 6808 4507 6862 4519
rect 6808 4481 6818 4507
rect 6852 4481 6862 4507
rect 6808 4429 6809 4481
rect 6861 4429 6862 4481
rect 6808 4422 6862 4429
rect 6908 4507 6962 4613
rect 7008 4691 7062 4698
rect 7008 4639 7009 4691
rect 7061 4639 7062 4691
rect 7008 4613 7018 4639
rect 7052 4613 7062 4639
rect 7008 4601 7062 4613
rect 7108 4647 7162 4753
rect 7208 4787 7262 4799
rect 7208 4761 7218 4787
rect 7252 4761 7262 4787
rect 7208 4709 7209 4761
rect 7261 4709 7262 4761
rect 7208 4702 7262 4709
rect 7308 4787 7362 4960
rect 7402 4919 7468 4920
rect 7402 4867 7409 4919
rect 7461 4867 7468 4919
rect 7402 4866 7468 4867
rect 7308 4753 7318 4787
rect 7352 4753 7362 4787
rect 7108 4613 7118 4647
rect 7152 4613 7162 4647
rect 6908 4473 6918 4507
rect 6952 4473 6962 4507
rect 6708 4333 6718 4367
rect 6752 4333 6762 4367
rect 6508 4193 6518 4227
rect 6552 4193 6562 4227
rect 6308 4053 6318 4087
rect 6352 4053 6362 4087
rect 6108 3913 6118 3947
rect 6152 3913 6162 3947
rect 5908 3773 5918 3807
rect 5952 3773 5962 3807
rect 5802 3709 5868 3710
rect 5802 3657 5809 3709
rect 5861 3657 5868 3709
rect 5802 3656 5868 3657
rect 5708 3543 5718 3577
rect 5752 3543 5762 3577
rect 5508 3403 5518 3437
rect 5552 3403 5562 3437
rect 5308 3263 5318 3297
rect 5352 3263 5362 3297
rect 5108 3123 5118 3157
rect 5152 3123 5162 3157
rect 4908 2983 4918 3017
rect 4952 2983 4962 3017
rect 4708 2843 4718 2877
rect 4752 2843 4762 2877
rect 4508 2703 4518 2737
rect 4552 2703 4562 2737
rect 4308 2563 4318 2597
rect 4352 2563 4362 2597
rect 4202 2499 4268 2500
rect 4202 2447 4209 2499
rect 4261 2447 4268 2499
rect 4202 2446 4268 2447
rect 4108 2333 4118 2367
rect 4152 2333 4162 2367
rect 3908 2193 3918 2227
rect 3952 2193 3962 2227
rect 3708 2053 3718 2087
rect 3752 2053 3762 2087
rect 3508 1913 3518 1947
rect 3552 1913 3562 1947
rect 3308 1773 3318 1807
rect 3352 1773 3362 1807
rect 3108 1633 3118 1667
rect 3152 1633 3162 1667
rect 2908 1493 2918 1527
rect 2952 1493 2962 1527
rect 2708 1353 2718 1387
rect 2752 1353 2762 1387
rect 2602 1289 2668 1290
rect 2602 1237 2609 1289
rect 2661 1237 2668 1289
rect 2602 1236 2668 1237
rect 2508 1123 2518 1157
rect 2552 1123 2562 1157
rect 2308 983 2318 1017
rect 2352 983 2362 1017
rect 2108 843 2118 877
rect 2152 843 2162 877
rect 1908 703 1918 737
rect 1952 703 1962 737
rect 1708 563 1718 597
rect 1752 563 1762 597
rect 1508 423 1518 457
rect 1552 423 1562 457
rect 1308 283 1318 317
rect 1352 283 1362 317
rect 1108 143 1118 177
rect 1152 143 1162 177
rect 1002 79 1068 80
rect 1002 27 1009 79
rect 1061 27 1068 79
rect 1002 26 1068 27
rect 908 -67 909 -15
rect 961 -67 962 -15
rect 908 -79 918 -67
rect 952 -79 962 -67
rect 708 -132 762 -131
rect 708 -143 718 -132
rect 752 -143 762 -132
rect 708 -195 709 -143
rect 761 -195 762 -143
rect 708 -210 762 -195
rect 812 -133 858 -81
rect 812 -167 818 -133
rect 852 -167 858 -133
rect 718 -291 725 -239
rect 777 -291 784 -239
rect 612 -397 618 -363
rect 652 -397 658 -363
rect 612 -435 658 -397
rect 612 -469 618 -435
rect 652 -469 658 -435
rect 612 -512 658 -469
rect 709 -326 761 -320
rect 709 -390 718 -378
rect 752 -390 761 -378
rect 709 -454 718 -442
rect 752 -454 761 -442
rect 709 -555 761 -506
rect 812 -363 858 -167
rect 908 -131 909 -79
rect 961 -131 962 -79
rect 1008 -22 1062 26
rect 1008 -74 1009 -22
rect 1061 -74 1062 -22
rect 1008 -81 1062 -74
rect 1108 -15 1162 143
rect 1208 177 1262 189
rect 1208 151 1218 177
rect 1252 151 1262 177
rect 1208 99 1209 151
rect 1261 99 1262 151
rect 1208 92 1262 99
rect 1308 177 1362 283
rect 1408 361 1462 368
rect 1408 309 1409 361
rect 1461 309 1462 361
rect 1408 283 1418 309
rect 1452 283 1462 309
rect 1408 271 1462 283
rect 1508 317 1562 423
rect 1608 457 1662 469
rect 1608 431 1618 457
rect 1652 431 1662 457
rect 1608 379 1609 431
rect 1661 379 1662 431
rect 1608 372 1662 379
rect 1708 457 1762 563
rect 1808 641 1862 648
rect 1808 589 1809 641
rect 1861 589 1862 641
rect 1808 563 1818 589
rect 1852 563 1862 589
rect 1808 551 1862 563
rect 1908 597 1962 703
rect 2008 737 2062 749
rect 2008 711 2018 737
rect 2052 711 2062 737
rect 2008 659 2009 711
rect 2061 659 2062 711
rect 2008 652 2062 659
rect 2108 737 2162 843
rect 2208 921 2262 928
rect 2208 869 2209 921
rect 2261 869 2262 921
rect 2208 843 2218 869
rect 2252 843 2262 869
rect 2208 831 2262 843
rect 2308 877 2362 983
rect 2408 1017 2462 1029
rect 2408 991 2418 1017
rect 2452 991 2462 1017
rect 2408 939 2409 991
rect 2461 939 2462 991
rect 2408 932 2462 939
rect 2508 1017 2562 1123
rect 2608 1201 2662 1208
rect 2608 1149 2609 1201
rect 2661 1149 2662 1201
rect 2608 1123 2618 1149
rect 2652 1123 2662 1149
rect 2608 1111 2662 1123
rect 2708 1157 2762 1353
rect 2808 1387 2862 1399
rect 2808 1361 2818 1387
rect 2852 1361 2862 1387
rect 2808 1309 2809 1361
rect 2861 1309 2862 1361
rect 2808 1302 2862 1309
rect 2908 1387 2962 1493
rect 3008 1571 3062 1578
rect 3008 1519 3009 1571
rect 3061 1519 3062 1571
rect 3008 1493 3018 1519
rect 3052 1493 3062 1519
rect 3008 1481 3062 1493
rect 3108 1527 3162 1633
rect 3208 1667 3262 1679
rect 3208 1641 3218 1667
rect 3252 1641 3262 1667
rect 3208 1589 3209 1641
rect 3261 1589 3262 1641
rect 3208 1582 3262 1589
rect 3308 1667 3362 1773
rect 3408 1851 3462 1858
rect 3408 1799 3409 1851
rect 3461 1799 3462 1851
rect 3408 1773 3418 1799
rect 3452 1773 3462 1799
rect 3408 1761 3462 1773
rect 3508 1807 3562 1913
rect 3608 1947 3662 1959
rect 3608 1921 3618 1947
rect 3652 1921 3662 1947
rect 3608 1869 3609 1921
rect 3661 1869 3662 1921
rect 3608 1862 3662 1869
rect 3708 1947 3762 2053
rect 3808 2131 3862 2138
rect 3808 2079 3809 2131
rect 3861 2079 3862 2131
rect 3808 2053 3818 2079
rect 3852 2053 3862 2079
rect 3808 2041 3862 2053
rect 3908 2087 3962 2193
rect 4008 2227 4062 2239
rect 4008 2201 4018 2227
rect 4052 2201 4062 2227
rect 4008 2149 4009 2201
rect 4061 2149 4062 2201
rect 4008 2142 4062 2149
rect 4108 2227 4162 2333
rect 4208 2411 4262 2418
rect 4208 2359 4209 2411
rect 4261 2359 4262 2411
rect 4208 2333 4218 2359
rect 4252 2333 4262 2359
rect 4208 2321 4262 2333
rect 4308 2367 4362 2563
rect 4408 2597 4462 2609
rect 4408 2571 4418 2597
rect 4452 2571 4462 2597
rect 4408 2519 4409 2571
rect 4461 2519 4462 2571
rect 4408 2512 4462 2519
rect 4508 2597 4562 2703
rect 4608 2781 4662 2788
rect 4608 2729 4609 2781
rect 4661 2729 4662 2781
rect 4608 2703 4618 2729
rect 4652 2703 4662 2729
rect 4608 2691 4662 2703
rect 4708 2737 4762 2843
rect 4808 2877 4862 2889
rect 4808 2851 4818 2877
rect 4852 2851 4862 2877
rect 4808 2799 4809 2851
rect 4861 2799 4862 2851
rect 4808 2792 4862 2799
rect 4908 2877 4962 2983
rect 5008 3061 5062 3068
rect 5008 3009 5009 3061
rect 5061 3009 5062 3061
rect 5008 2983 5018 3009
rect 5052 2983 5062 3009
rect 5008 2971 5062 2983
rect 5108 3017 5162 3123
rect 5208 3157 5262 3169
rect 5208 3131 5218 3157
rect 5252 3131 5262 3157
rect 5208 3079 5209 3131
rect 5261 3079 5262 3131
rect 5208 3072 5262 3079
rect 5308 3157 5362 3263
rect 5408 3341 5462 3348
rect 5408 3289 5409 3341
rect 5461 3289 5462 3341
rect 5408 3263 5418 3289
rect 5452 3263 5462 3289
rect 5408 3251 5462 3263
rect 5508 3297 5562 3403
rect 5608 3437 5662 3449
rect 5608 3411 5618 3437
rect 5652 3411 5662 3437
rect 5608 3359 5609 3411
rect 5661 3359 5662 3411
rect 5608 3352 5662 3359
rect 5708 3437 5762 3543
rect 5808 3621 5862 3628
rect 5808 3569 5809 3621
rect 5861 3569 5862 3621
rect 5808 3543 5818 3569
rect 5852 3543 5862 3569
rect 5808 3531 5862 3543
rect 5908 3577 5962 3773
rect 6008 3807 6062 3819
rect 6008 3781 6018 3807
rect 6052 3781 6062 3807
rect 6008 3729 6009 3781
rect 6061 3729 6062 3781
rect 6008 3722 6062 3729
rect 6108 3807 6162 3913
rect 6208 3991 6262 3998
rect 6208 3939 6209 3991
rect 6261 3939 6262 3991
rect 6208 3913 6218 3939
rect 6252 3913 6262 3939
rect 6208 3901 6262 3913
rect 6308 3947 6362 4053
rect 6408 4087 6462 4099
rect 6408 4061 6418 4087
rect 6452 4061 6462 4087
rect 6408 4009 6409 4061
rect 6461 4009 6462 4061
rect 6408 4002 6462 4009
rect 6508 4087 6562 4193
rect 6608 4271 6662 4278
rect 6608 4219 6609 4271
rect 6661 4219 6662 4271
rect 6608 4193 6618 4219
rect 6652 4193 6662 4219
rect 6608 4181 6662 4193
rect 6708 4227 6762 4333
rect 6808 4367 6862 4379
rect 6808 4341 6818 4367
rect 6852 4341 6862 4367
rect 6808 4289 6809 4341
rect 6861 4289 6862 4341
rect 6808 4282 6862 4289
rect 6908 4367 6962 4473
rect 7008 4551 7062 4558
rect 7008 4499 7009 4551
rect 7061 4499 7062 4551
rect 7008 4473 7018 4499
rect 7052 4473 7062 4499
rect 7008 4461 7062 4473
rect 7108 4507 7162 4613
rect 7208 4647 7262 4659
rect 7208 4621 7218 4647
rect 7252 4621 7262 4647
rect 7208 4569 7209 4621
rect 7261 4569 7262 4621
rect 7208 4562 7262 4569
rect 7308 4647 7362 4753
rect 7408 4831 7462 4838
rect 7408 4779 7409 4831
rect 7461 4779 7462 4831
rect 7408 4753 7418 4779
rect 7452 4753 7462 4779
rect 7408 4741 7462 4753
rect 7508 4787 7562 4960
rect 7602 4903 7668 4904
rect 7602 4851 7609 4903
rect 7661 4851 7668 4903
rect 7602 4850 7668 4851
rect 7508 4753 7518 4787
rect 7552 4753 7562 4787
rect 7308 4613 7318 4647
rect 7352 4613 7362 4647
rect 7108 4473 7118 4507
rect 7152 4473 7162 4507
rect 6908 4333 6918 4367
rect 6952 4333 6962 4367
rect 6708 4193 6718 4227
rect 6752 4193 6762 4227
rect 6508 4053 6518 4087
rect 6552 4053 6562 4087
rect 6308 3913 6318 3947
rect 6352 3913 6362 3947
rect 6108 3773 6118 3807
rect 6152 3773 6162 3807
rect 6002 3693 6068 3694
rect 6002 3641 6009 3693
rect 6061 3641 6068 3693
rect 6002 3640 6068 3641
rect 5908 3543 5918 3577
rect 5952 3543 5962 3577
rect 5708 3403 5718 3437
rect 5752 3403 5762 3437
rect 5508 3263 5518 3297
rect 5552 3263 5562 3297
rect 5308 3123 5318 3157
rect 5352 3123 5362 3157
rect 5108 2983 5118 3017
rect 5152 2983 5162 3017
rect 4908 2843 4918 2877
rect 4952 2843 4962 2877
rect 4708 2703 4718 2737
rect 4752 2703 4762 2737
rect 4508 2563 4518 2597
rect 4552 2563 4562 2597
rect 4402 2483 4468 2484
rect 4402 2431 4409 2483
rect 4461 2431 4468 2483
rect 4402 2430 4468 2431
rect 4308 2333 4318 2367
rect 4352 2333 4362 2367
rect 4108 2193 4118 2227
rect 4152 2193 4162 2227
rect 3908 2053 3918 2087
rect 3952 2053 3962 2087
rect 3708 1913 3718 1947
rect 3752 1913 3762 1947
rect 3508 1773 3518 1807
rect 3552 1773 3562 1807
rect 3308 1633 3318 1667
rect 3352 1633 3362 1667
rect 3108 1493 3118 1527
rect 3152 1493 3162 1527
rect 2908 1353 2918 1387
rect 2952 1353 2962 1387
rect 2802 1273 2868 1274
rect 2802 1221 2809 1273
rect 2861 1221 2868 1273
rect 2802 1220 2868 1221
rect 2708 1123 2718 1157
rect 2752 1123 2762 1157
rect 2508 983 2518 1017
rect 2552 983 2562 1017
rect 2308 843 2318 877
rect 2352 843 2362 877
rect 2108 703 2118 737
rect 2152 703 2162 737
rect 1908 563 1918 597
rect 1952 563 1962 597
rect 1708 423 1718 457
rect 1752 423 1762 457
rect 1508 283 1518 317
rect 1552 283 1562 317
rect 1308 143 1318 177
rect 1352 143 1362 177
rect 1202 63 1268 64
rect 1202 11 1209 63
rect 1261 11 1268 63
rect 1202 10 1268 11
rect 1108 -67 1109 -15
rect 1161 -67 1162 -15
rect 1108 -79 1118 -67
rect 1152 -79 1162 -67
rect 908 -132 962 -131
rect 908 -143 918 -132
rect 952 -143 962 -132
rect 908 -195 909 -143
rect 961 -195 962 -143
rect 908 -210 962 -195
rect 1012 -133 1058 -81
rect 1012 -167 1018 -133
rect 1052 -167 1058 -133
rect 918 -291 925 -239
rect 977 -291 984 -239
rect 812 -397 818 -363
rect 852 -397 858 -363
rect 812 -435 858 -397
rect 812 -469 818 -435
rect 852 -469 858 -435
rect 812 -512 858 -469
rect 909 -326 961 -320
rect 909 -390 918 -378
rect 952 -390 961 -378
rect 909 -454 918 -442
rect 952 -454 961 -442
rect 909 -512 961 -506
rect 1012 -363 1058 -167
rect 1108 -131 1109 -79
rect 1161 -131 1162 -79
rect 1208 -22 1262 10
rect 1208 -74 1209 -22
rect 1261 -74 1262 -22
rect 1208 -81 1262 -74
rect 1308 -15 1362 143
rect 1408 221 1462 228
rect 1408 169 1409 221
rect 1461 169 1462 221
rect 1408 143 1418 169
rect 1452 143 1462 169
rect 1408 131 1462 143
rect 1508 177 1562 283
rect 1608 317 1662 329
rect 1608 291 1618 317
rect 1652 291 1662 317
rect 1608 239 1609 291
rect 1661 239 1662 291
rect 1608 232 1662 239
rect 1708 317 1762 423
rect 1808 501 1862 508
rect 1808 449 1809 501
rect 1861 449 1862 501
rect 1808 423 1818 449
rect 1852 423 1862 449
rect 1808 411 1862 423
rect 1908 457 1962 563
rect 2008 597 2062 609
rect 2008 571 2018 597
rect 2052 571 2062 597
rect 2008 519 2009 571
rect 2061 519 2062 571
rect 2008 512 2062 519
rect 2108 597 2162 703
rect 2208 781 2262 788
rect 2208 729 2209 781
rect 2261 729 2262 781
rect 2208 703 2218 729
rect 2252 703 2262 729
rect 2208 691 2262 703
rect 2308 737 2362 843
rect 2408 877 2462 889
rect 2408 851 2418 877
rect 2452 851 2462 877
rect 2408 799 2409 851
rect 2461 799 2462 851
rect 2408 792 2462 799
rect 2508 877 2562 983
rect 2608 1061 2662 1068
rect 2608 1009 2609 1061
rect 2661 1009 2662 1061
rect 2608 983 2618 1009
rect 2652 983 2662 1009
rect 2608 971 2662 983
rect 2708 1017 2762 1123
rect 2808 1157 2862 1169
rect 2808 1131 2818 1157
rect 2852 1131 2862 1157
rect 2808 1079 2809 1131
rect 2861 1079 2862 1131
rect 2808 1072 2862 1079
rect 2908 1157 2962 1353
rect 3008 1431 3062 1438
rect 3008 1379 3009 1431
rect 3061 1379 3062 1431
rect 3008 1353 3018 1379
rect 3052 1353 3062 1379
rect 3008 1341 3062 1353
rect 3108 1387 3162 1493
rect 3208 1527 3262 1539
rect 3208 1501 3218 1527
rect 3252 1501 3262 1527
rect 3208 1449 3209 1501
rect 3261 1449 3262 1501
rect 3208 1442 3262 1449
rect 3308 1527 3362 1633
rect 3408 1711 3462 1718
rect 3408 1659 3409 1711
rect 3461 1659 3462 1711
rect 3408 1633 3418 1659
rect 3452 1633 3462 1659
rect 3408 1621 3462 1633
rect 3508 1667 3562 1773
rect 3608 1807 3662 1819
rect 3608 1781 3618 1807
rect 3652 1781 3662 1807
rect 3608 1729 3609 1781
rect 3661 1729 3662 1781
rect 3608 1722 3662 1729
rect 3708 1807 3762 1913
rect 3808 1991 3862 1998
rect 3808 1939 3809 1991
rect 3861 1939 3862 1991
rect 3808 1913 3818 1939
rect 3852 1913 3862 1939
rect 3808 1901 3862 1913
rect 3908 1947 3962 2053
rect 4008 2087 4062 2099
rect 4008 2061 4018 2087
rect 4052 2061 4062 2087
rect 4008 2009 4009 2061
rect 4061 2009 4062 2061
rect 4008 2002 4062 2009
rect 4108 2087 4162 2193
rect 4208 2271 4262 2278
rect 4208 2219 4209 2271
rect 4261 2219 4262 2271
rect 4208 2193 4218 2219
rect 4252 2193 4262 2219
rect 4208 2181 4262 2193
rect 4308 2227 4362 2333
rect 4408 2367 4462 2379
rect 4408 2341 4418 2367
rect 4452 2341 4462 2367
rect 4408 2289 4409 2341
rect 4461 2289 4462 2341
rect 4408 2282 4462 2289
rect 4508 2367 4562 2563
rect 4608 2641 4662 2648
rect 4608 2589 4609 2641
rect 4661 2589 4662 2641
rect 4608 2563 4618 2589
rect 4652 2563 4662 2589
rect 4608 2551 4662 2563
rect 4708 2597 4762 2703
rect 4808 2737 4862 2749
rect 4808 2711 4818 2737
rect 4852 2711 4862 2737
rect 4808 2659 4809 2711
rect 4861 2659 4862 2711
rect 4808 2652 4862 2659
rect 4908 2737 4962 2843
rect 5008 2921 5062 2928
rect 5008 2869 5009 2921
rect 5061 2869 5062 2921
rect 5008 2843 5018 2869
rect 5052 2843 5062 2869
rect 5008 2831 5062 2843
rect 5108 2877 5162 2983
rect 5208 3017 5262 3029
rect 5208 2991 5218 3017
rect 5252 2991 5262 3017
rect 5208 2939 5209 2991
rect 5261 2939 5262 2991
rect 5208 2932 5262 2939
rect 5308 3017 5362 3123
rect 5408 3201 5462 3208
rect 5408 3149 5409 3201
rect 5461 3149 5462 3201
rect 5408 3123 5418 3149
rect 5452 3123 5462 3149
rect 5408 3111 5462 3123
rect 5508 3157 5562 3263
rect 5608 3297 5662 3309
rect 5608 3271 5618 3297
rect 5652 3271 5662 3297
rect 5608 3219 5609 3271
rect 5661 3219 5662 3271
rect 5608 3212 5662 3219
rect 5708 3297 5762 3403
rect 5808 3481 5862 3488
rect 5808 3429 5809 3481
rect 5861 3429 5862 3481
rect 5808 3403 5818 3429
rect 5852 3403 5862 3429
rect 5808 3391 5862 3403
rect 5908 3437 5962 3543
rect 6008 3577 6062 3589
rect 6008 3551 6018 3577
rect 6052 3551 6062 3577
rect 6008 3499 6009 3551
rect 6061 3499 6062 3551
rect 6008 3492 6062 3499
rect 6108 3577 6162 3773
rect 6208 3851 6262 3858
rect 6208 3799 6209 3851
rect 6261 3799 6262 3851
rect 6208 3773 6218 3799
rect 6252 3773 6262 3799
rect 6208 3761 6262 3773
rect 6308 3807 6362 3913
rect 6408 3947 6462 3959
rect 6408 3921 6418 3947
rect 6452 3921 6462 3947
rect 6408 3869 6409 3921
rect 6461 3869 6462 3921
rect 6408 3862 6462 3869
rect 6508 3947 6562 4053
rect 6608 4131 6662 4138
rect 6608 4079 6609 4131
rect 6661 4079 6662 4131
rect 6608 4053 6618 4079
rect 6652 4053 6662 4079
rect 6608 4041 6662 4053
rect 6708 4087 6762 4193
rect 6808 4227 6862 4239
rect 6808 4201 6818 4227
rect 6852 4201 6862 4227
rect 6808 4149 6809 4201
rect 6861 4149 6862 4201
rect 6808 4142 6862 4149
rect 6908 4227 6962 4333
rect 7008 4411 7062 4418
rect 7008 4359 7009 4411
rect 7061 4359 7062 4411
rect 7008 4333 7018 4359
rect 7052 4333 7062 4359
rect 7008 4321 7062 4333
rect 7108 4367 7162 4473
rect 7208 4507 7262 4519
rect 7208 4481 7218 4507
rect 7252 4481 7262 4507
rect 7208 4429 7209 4481
rect 7261 4429 7262 4481
rect 7208 4422 7262 4429
rect 7308 4507 7362 4613
rect 7408 4691 7462 4698
rect 7408 4639 7409 4691
rect 7461 4639 7462 4691
rect 7408 4613 7418 4639
rect 7452 4613 7462 4639
rect 7408 4601 7462 4613
rect 7508 4647 7562 4753
rect 7608 4787 7662 4799
rect 7608 4761 7618 4787
rect 7652 4761 7662 4787
rect 7608 4709 7609 4761
rect 7661 4709 7662 4761
rect 7608 4702 7662 4709
rect 7708 4787 7762 4960
rect 7802 4919 7868 4920
rect 7802 4867 7809 4919
rect 7861 4867 7868 4919
rect 7802 4866 7868 4867
rect 7708 4753 7718 4787
rect 7752 4753 7762 4787
rect 7508 4613 7518 4647
rect 7552 4613 7562 4647
rect 7308 4473 7318 4507
rect 7352 4473 7362 4507
rect 7108 4333 7118 4367
rect 7152 4333 7162 4367
rect 6908 4193 6918 4227
rect 6952 4193 6962 4227
rect 6708 4053 6718 4087
rect 6752 4053 6762 4087
rect 6508 3913 6518 3947
rect 6552 3913 6562 3947
rect 6308 3773 6318 3807
rect 6352 3773 6362 3807
rect 6202 3709 6268 3710
rect 6202 3657 6209 3709
rect 6261 3657 6268 3709
rect 6202 3656 6268 3657
rect 6108 3543 6118 3577
rect 6152 3543 6162 3577
rect 5908 3403 5918 3437
rect 5952 3403 5962 3437
rect 5708 3263 5718 3297
rect 5752 3263 5762 3297
rect 5508 3123 5518 3157
rect 5552 3123 5562 3157
rect 5308 2983 5318 3017
rect 5352 2983 5362 3017
rect 5108 2843 5118 2877
rect 5152 2843 5162 2877
rect 4908 2703 4918 2737
rect 4952 2703 4962 2737
rect 4708 2563 4718 2597
rect 4752 2563 4762 2597
rect 4602 2499 4668 2500
rect 4602 2447 4609 2499
rect 4661 2447 4668 2499
rect 4602 2446 4668 2447
rect 4508 2333 4518 2367
rect 4552 2333 4562 2367
rect 4308 2193 4318 2227
rect 4352 2193 4362 2227
rect 4108 2053 4118 2087
rect 4152 2053 4162 2087
rect 3908 1913 3918 1947
rect 3952 1913 3962 1947
rect 3708 1773 3718 1807
rect 3752 1773 3762 1807
rect 3508 1633 3518 1667
rect 3552 1633 3562 1667
rect 3308 1493 3318 1527
rect 3352 1493 3362 1527
rect 3108 1353 3118 1387
rect 3152 1353 3162 1387
rect 3002 1289 3068 1290
rect 3002 1237 3009 1289
rect 3061 1237 3068 1289
rect 3002 1236 3068 1237
rect 2908 1123 2918 1157
rect 2952 1123 2962 1157
rect 2708 983 2718 1017
rect 2752 983 2762 1017
rect 2508 843 2518 877
rect 2552 843 2562 877
rect 2308 703 2318 737
rect 2352 703 2362 737
rect 2108 563 2118 597
rect 2152 563 2162 597
rect 1908 423 1918 457
rect 1952 423 1962 457
rect 1708 283 1718 317
rect 1752 283 1762 317
rect 1508 143 1518 177
rect 1552 143 1562 177
rect 1402 79 1468 80
rect 1402 27 1409 79
rect 1461 27 1468 79
rect 1402 26 1468 27
rect 1308 -67 1309 -15
rect 1361 -67 1362 -15
rect 1308 -79 1318 -67
rect 1352 -79 1362 -67
rect 1108 -132 1162 -131
rect 1108 -143 1118 -132
rect 1152 -143 1162 -132
rect 1108 -195 1109 -143
rect 1161 -195 1162 -143
rect 1108 -210 1162 -195
rect 1212 -133 1258 -81
rect 1212 -167 1218 -133
rect 1252 -167 1258 -133
rect 1118 -291 1125 -239
rect 1177 -291 1184 -239
rect 1012 -397 1018 -363
rect 1052 -397 1058 -363
rect 1012 -435 1058 -397
rect 1012 -469 1018 -435
rect 1052 -469 1058 -435
rect 1012 -512 1058 -469
rect 1109 -326 1161 -320
rect 1109 -390 1118 -378
rect 1152 -390 1161 -378
rect 1109 -454 1118 -442
rect 1152 -454 1161 -442
rect 1109 -555 1161 -506
rect 1212 -363 1258 -167
rect 1308 -131 1309 -79
rect 1361 -131 1362 -79
rect 1408 -22 1462 26
rect 1408 -74 1409 -22
rect 1461 -74 1462 -22
rect 1408 -81 1462 -74
rect 1508 -15 1562 143
rect 1608 177 1662 189
rect 1608 151 1618 177
rect 1652 151 1662 177
rect 1608 99 1609 151
rect 1661 99 1662 151
rect 1608 92 1662 99
rect 1708 177 1762 283
rect 1808 361 1862 368
rect 1808 309 1809 361
rect 1861 309 1862 361
rect 1808 283 1818 309
rect 1852 283 1862 309
rect 1808 271 1862 283
rect 1908 317 1962 423
rect 2008 457 2062 469
rect 2008 431 2018 457
rect 2052 431 2062 457
rect 2008 379 2009 431
rect 2061 379 2062 431
rect 2008 372 2062 379
rect 2108 457 2162 563
rect 2208 641 2262 648
rect 2208 589 2209 641
rect 2261 589 2262 641
rect 2208 563 2218 589
rect 2252 563 2262 589
rect 2208 551 2262 563
rect 2308 597 2362 703
rect 2408 737 2462 749
rect 2408 711 2418 737
rect 2452 711 2462 737
rect 2408 659 2409 711
rect 2461 659 2462 711
rect 2408 652 2462 659
rect 2508 737 2562 843
rect 2608 921 2662 928
rect 2608 869 2609 921
rect 2661 869 2662 921
rect 2608 843 2618 869
rect 2652 843 2662 869
rect 2608 831 2662 843
rect 2708 877 2762 983
rect 2808 1017 2862 1029
rect 2808 991 2818 1017
rect 2852 991 2862 1017
rect 2808 939 2809 991
rect 2861 939 2862 991
rect 2808 932 2862 939
rect 2908 1017 2962 1123
rect 3008 1201 3062 1208
rect 3008 1149 3009 1201
rect 3061 1149 3062 1201
rect 3008 1123 3018 1149
rect 3052 1123 3062 1149
rect 3008 1111 3062 1123
rect 3108 1157 3162 1353
rect 3208 1387 3262 1399
rect 3208 1361 3218 1387
rect 3252 1361 3262 1387
rect 3208 1309 3209 1361
rect 3261 1309 3262 1361
rect 3208 1302 3262 1309
rect 3308 1387 3362 1493
rect 3408 1571 3462 1578
rect 3408 1519 3409 1571
rect 3461 1519 3462 1571
rect 3408 1493 3418 1519
rect 3452 1493 3462 1519
rect 3408 1481 3462 1493
rect 3508 1527 3562 1633
rect 3608 1667 3662 1679
rect 3608 1641 3618 1667
rect 3652 1641 3662 1667
rect 3608 1589 3609 1641
rect 3661 1589 3662 1641
rect 3608 1582 3662 1589
rect 3708 1667 3762 1773
rect 3808 1851 3862 1858
rect 3808 1799 3809 1851
rect 3861 1799 3862 1851
rect 3808 1773 3818 1799
rect 3852 1773 3862 1799
rect 3808 1761 3862 1773
rect 3908 1807 3962 1913
rect 4008 1947 4062 1959
rect 4008 1921 4018 1947
rect 4052 1921 4062 1947
rect 4008 1869 4009 1921
rect 4061 1869 4062 1921
rect 4008 1862 4062 1869
rect 4108 1947 4162 2053
rect 4208 2131 4262 2138
rect 4208 2079 4209 2131
rect 4261 2079 4262 2131
rect 4208 2053 4218 2079
rect 4252 2053 4262 2079
rect 4208 2041 4262 2053
rect 4308 2087 4362 2193
rect 4408 2227 4462 2239
rect 4408 2201 4418 2227
rect 4452 2201 4462 2227
rect 4408 2149 4409 2201
rect 4461 2149 4462 2201
rect 4408 2142 4462 2149
rect 4508 2227 4562 2333
rect 4608 2411 4662 2418
rect 4608 2359 4609 2411
rect 4661 2359 4662 2411
rect 4608 2333 4618 2359
rect 4652 2333 4662 2359
rect 4608 2321 4662 2333
rect 4708 2367 4762 2563
rect 4808 2597 4862 2609
rect 4808 2571 4818 2597
rect 4852 2571 4862 2597
rect 4808 2519 4809 2571
rect 4861 2519 4862 2571
rect 4808 2512 4862 2519
rect 4908 2597 4962 2703
rect 5008 2781 5062 2788
rect 5008 2729 5009 2781
rect 5061 2729 5062 2781
rect 5008 2703 5018 2729
rect 5052 2703 5062 2729
rect 5008 2691 5062 2703
rect 5108 2737 5162 2843
rect 5208 2877 5262 2889
rect 5208 2851 5218 2877
rect 5252 2851 5262 2877
rect 5208 2799 5209 2851
rect 5261 2799 5262 2851
rect 5208 2792 5262 2799
rect 5308 2877 5362 2983
rect 5408 3061 5462 3068
rect 5408 3009 5409 3061
rect 5461 3009 5462 3061
rect 5408 2983 5418 3009
rect 5452 2983 5462 3009
rect 5408 2971 5462 2983
rect 5508 3017 5562 3123
rect 5608 3157 5662 3169
rect 5608 3131 5618 3157
rect 5652 3131 5662 3157
rect 5608 3079 5609 3131
rect 5661 3079 5662 3131
rect 5608 3072 5662 3079
rect 5708 3157 5762 3263
rect 5808 3341 5862 3348
rect 5808 3289 5809 3341
rect 5861 3289 5862 3341
rect 5808 3263 5818 3289
rect 5852 3263 5862 3289
rect 5808 3251 5862 3263
rect 5908 3297 5962 3403
rect 6008 3437 6062 3449
rect 6008 3411 6018 3437
rect 6052 3411 6062 3437
rect 6008 3359 6009 3411
rect 6061 3359 6062 3411
rect 6008 3352 6062 3359
rect 6108 3437 6162 3543
rect 6208 3621 6262 3628
rect 6208 3569 6209 3621
rect 6261 3569 6262 3621
rect 6208 3543 6218 3569
rect 6252 3543 6262 3569
rect 6208 3531 6262 3543
rect 6308 3577 6362 3773
rect 6408 3807 6462 3819
rect 6408 3781 6418 3807
rect 6452 3781 6462 3807
rect 6408 3729 6409 3781
rect 6461 3729 6462 3781
rect 6408 3722 6462 3729
rect 6508 3807 6562 3913
rect 6608 3991 6662 3998
rect 6608 3939 6609 3991
rect 6661 3939 6662 3991
rect 6608 3913 6618 3939
rect 6652 3913 6662 3939
rect 6608 3901 6662 3913
rect 6708 3947 6762 4053
rect 6808 4087 6862 4099
rect 6808 4061 6818 4087
rect 6852 4061 6862 4087
rect 6808 4009 6809 4061
rect 6861 4009 6862 4061
rect 6808 4002 6862 4009
rect 6908 4087 6962 4193
rect 7008 4271 7062 4278
rect 7008 4219 7009 4271
rect 7061 4219 7062 4271
rect 7008 4193 7018 4219
rect 7052 4193 7062 4219
rect 7008 4181 7062 4193
rect 7108 4227 7162 4333
rect 7208 4367 7262 4379
rect 7208 4341 7218 4367
rect 7252 4341 7262 4367
rect 7208 4289 7209 4341
rect 7261 4289 7262 4341
rect 7208 4282 7262 4289
rect 7308 4367 7362 4473
rect 7408 4551 7462 4558
rect 7408 4499 7409 4551
rect 7461 4499 7462 4551
rect 7408 4473 7418 4499
rect 7452 4473 7462 4499
rect 7408 4461 7462 4473
rect 7508 4507 7562 4613
rect 7608 4647 7662 4659
rect 7608 4621 7618 4647
rect 7652 4621 7662 4647
rect 7608 4569 7609 4621
rect 7661 4569 7662 4621
rect 7608 4562 7662 4569
rect 7708 4647 7762 4753
rect 7808 4831 7862 4838
rect 7808 4779 7809 4831
rect 7861 4779 7862 4831
rect 7808 4753 7818 4779
rect 7852 4753 7862 4779
rect 7808 4741 7862 4753
rect 7908 4787 7962 4960
rect 8002 4903 8068 4904
rect 8002 4851 8009 4903
rect 8061 4851 8068 4903
rect 8002 4850 8068 4851
rect 7908 4753 7918 4787
rect 7952 4753 7962 4787
rect 7708 4613 7718 4647
rect 7752 4613 7762 4647
rect 7508 4473 7518 4507
rect 7552 4473 7562 4507
rect 7308 4333 7318 4367
rect 7352 4333 7362 4367
rect 7108 4193 7118 4227
rect 7152 4193 7162 4227
rect 6908 4053 6918 4087
rect 6952 4053 6962 4087
rect 6708 3913 6718 3947
rect 6752 3913 6762 3947
rect 6508 3773 6518 3807
rect 6552 3773 6562 3807
rect 6402 3693 6468 3694
rect 6402 3641 6409 3693
rect 6461 3641 6468 3693
rect 6402 3640 6468 3641
rect 6308 3543 6318 3577
rect 6352 3543 6362 3577
rect 6108 3403 6118 3437
rect 6152 3403 6162 3437
rect 5908 3263 5918 3297
rect 5952 3263 5962 3297
rect 5708 3123 5718 3157
rect 5752 3123 5762 3157
rect 5508 2983 5518 3017
rect 5552 2983 5562 3017
rect 5308 2843 5318 2877
rect 5352 2843 5362 2877
rect 5108 2703 5118 2737
rect 5152 2703 5162 2737
rect 4908 2563 4918 2597
rect 4952 2563 4962 2597
rect 4802 2483 4868 2484
rect 4802 2431 4809 2483
rect 4861 2431 4868 2483
rect 4802 2430 4868 2431
rect 4708 2333 4718 2367
rect 4752 2333 4762 2367
rect 4508 2193 4518 2227
rect 4552 2193 4562 2227
rect 4308 2053 4318 2087
rect 4352 2053 4362 2087
rect 4108 1913 4118 1947
rect 4152 1913 4162 1947
rect 3908 1773 3918 1807
rect 3952 1773 3962 1807
rect 3708 1633 3718 1667
rect 3752 1633 3762 1667
rect 3508 1493 3518 1527
rect 3552 1493 3562 1527
rect 3308 1353 3318 1387
rect 3352 1353 3362 1387
rect 3202 1273 3268 1274
rect 3202 1221 3209 1273
rect 3261 1221 3268 1273
rect 3202 1220 3268 1221
rect 3108 1123 3118 1157
rect 3152 1123 3162 1157
rect 2908 983 2918 1017
rect 2952 983 2962 1017
rect 2708 843 2718 877
rect 2752 843 2762 877
rect 2508 703 2518 737
rect 2552 703 2562 737
rect 2308 563 2318 597
rect 2352 563 2362 597
rect 2108 423 2118 457
rect 2152 423 2162 457
rect 1908 283 1918 317
rect 1952 283 1962 317
rect 1708 143 1718 177
rect 1752 143 1762 177
rect 1602 63 1668 64
rect 1602 11 1609 63
rect 1661 11 1668 63
rect 1602 10 1668 11
rect 1508 -67 1509 -15
rect 1561 -67 1562 -15
rect 1508 -79 1518 -67
rect 1552 -79 1562 -67
rect 1308 -132 1362 -131
rect 1308 -143 1318 -132
rect 1352 -143 1362 -132
rect 1308 -195 1309 -143
rect 1361 -195 1362 -143
rect 1308 -210 1362 -195
rect 1412 -133 1458 -81
rect 1412 -167 1418 -133
rect 1452 -167 1458 -133
rect 1318 -291 1325 -239
rect 1377 -291 1384 -239
rect 1212 -397 1218 -363
rect 1252 -397 1258 -363
rect 1212 -435 1258 -397
rect 1212 -469 1218 -435
rect 1252 -469 1258 -435
rect 1212 -512 1258 -469
rect 1309 -326 1361 -320
rect 1309 -390 1318 -378
rect 1352 -390 1361 -378
rect 1309 -454 1318 -442
rect 1352 -454 1361 -442
rect 1309 -512 1361 -506
rect 1412 -363 1458 -167
rect 1508 -131 1509 -79
rect 1561 -131 1562 -79
rect 1608 -22 1662 10
rect 1608 -74 1609 -22
rect 1661 -74 1662 -22
rect 1608 -81 1662 -74
rect 1708 -15 1762 143
rect 1808 221 1862 228
rect 1808 169 1809 221
rect 1861 169 1862 221
rect 1808 143 1818 169
rect 1852 143 1862 169
rect 1808 131 1862 143
rect 1908 177 1962 283
rect 2008 317 2062 329
rect 2008 291 2018 317
rect 2052 291 2062 317
rect 2008 239 2009 291
rect 2061 239 2062 291
rect 2008 232 2062 239
rect 2108 317 2162 423
rect 2208 501 2262 508
rect 2208 449 2209 501
rect 2261 449 2262 501
rect 2208 423 2218 449
rect 2252 423 2262 449
rect 2208 411 2262 423
rect 2308 457 2362 563
rect 2408 597 2462 609
rect 2408 571 2418 597
rect 2452 571 2462 597
rect 2408 519 2409 571
rect 2461 519 2462 571
rect 2408 512 2462 519
rect 2508 597 2562 703
rect 2608 781 2662 788
rect 2608 729 2609 781
rect 2661 729 2662 781
rect 2608 703 2618 729
rect 2652 703 2662 729
rect 2608 691 2662 703
rect 2708 737 2762 843
rect 2808 877 2862 889
rect 2808 851 2818 877
rect 2852 851 2862 877
rect 2808 799 2809 851
rect 2861 799 2862 851
rect 2808 792 2862 799
rect 2908 877 2962 983
rect 3008 1061 3062 1068
rect 3008 1009 3009 1061
rect 3061 1009 3062 1061
rect 3008 983 3018 1009
rect 3052 983 3062 1009
rect 3008 971 3062 983
rect 3108 1017 3162 1123
rect 3208 1157 3262 1169
rect 3208 1131 3218 1157
rect 3252 1131 3262 1157
rect 3208 1079 3209 1131
rect 3261 1079 3262 1131
rect 3208 1072 3262 1079
rect 3308 1157 3362 1353
rect 3408 1431 3462 1438
rect 3408 1379 3409 1431
rect 3461 1379 3462 1431
rect 3408 1353 3418 1379
rect 3452 1353 3462 1379
rect 3408 1341 3462 1353
rect 3508 1387 3562 1493
rect 3608 1527 3662 1539
rect 3608 1501 3618 1527
rect 3652 1501 3662 1527
rect 3608 1449 3609 1501
rect 3661 1449 3662 1501
rect 3608 1442 3662 1449
rect 3708 1527 3762 1633
rect 3808 1711 3862 1718
rect 3808 1659 3809 1711
rect 3861 1659 3862 1711
rect 3808 1633 3818 1659
rect 3852 1633 3862 1659
rect 3808 1621 3862 1633
rect 3908 1667 3962 1773
rect 4008 1807 4062 1819
rect 4008 1781 4018 1807
rect 4052 1781 4062 1807
rect 4008 1729 4009 1781
rect 4061 1729 4062 1781
rect 4008 1722 4062 1729
rect 4108 1807 4162 1913
rect 4208 1991 4262 1998
rect 4208 1939 4209 1991
rect 4261 1939 4262 1991
rect 4208 1913 4218 1939
rect 4252 1913 4262 1939
rect 4208 1901 4262 1913
rect 4308 1947 4362 2053
rect 4408 2087 4462 2099
rect 4408 2061 4418 2087
rect 4452 2061 4462 2087
rect 4408 2009 4409 2061
rect 4461 2009 4462 2061
rect 4408 2002 4462 2009
rect 4508 2087 4562 2193
rect 4608 2271 4662 2278
rect 4608 2219 4609 2271
rect 4661 2219 4662 2271
rect 4608 2193 4618 2219
rect 4652 2193 4662 2219
rect 4608 2181 4662 2193
rect 4708 2227 4762 2333
rect 4808 2367 4862 2379
rect 4808 2341 4818 2367
rect 4852 2341 4862 2367
rect 4808 2289 4809 2341
rect 4861 2289 4862 2341
rect 4808 2282 4862 2289
rect 4908 2367 4962 2563
rect 5008 2641 5062 2648
rect 5008 2589 5009 2641
rect 5061 2589 5062 2641
rect 5008 2563 5018 2589
rect 5052 2563 5062 2589
rect 5008 2551 5062 2563
rect 5108 2597 5162 2703
rect 5208 2737 5262 2749
rect 5208 2711 5218 2737
rect 5252 2711 5262 2737
rect 5208 2659 5209 2711
rect 5261 2659 5262 2711
rect 5208 2652 5262 2659
rect 5308 2737 5362 2843
rect 5408 2921 5462 2928
rect 5408 2869 5409 2921
rect 5461 2869 5462 2921
rect 5408 2843 5418 2869
rect 5452 2843 5462 2869
rect 5408 2831 5462 2843
rect 5508 2877 5562 2983
rect 5608 3017 5662 3029
rect 5608 2991 5618 3017
rect 5652 2991 5662 3017
rect 5608 2939 5609 2991
rect 5661 2939 5662 2991
rect 5608 2932 5662 2939
rect 5708 3017 5762 3123
rect 5808 3201 5862 3208
rect 5808 3149 5809 3201
rect 5861 3149 5862 3201
rect 5808 3123 5818 3149
rect 5852 3123 5862 3149
rect 5808 3111 5862 3123
rect 5908 3157 5962 3263
rect 6008 3297 6062 3309
rect 6008 3271 6018 3297
rect 6052 3271 6062 3297
rect 6008 3219 6009 3271
rect 6061 3219 6062 3271
rect 6008 3212 6062 3219
rect 6108 3297 6162 3403
rect 6208 3481 6262 3488
rect 6208 3429 6209 3481
rect 6261 3429 6262 3481
rect 6208 3403 6218 3429
rect 6252 3403 6262 3429
rect 6208 3391 6262 3403
rect 6308 3437 6362 3543
rect 6408 3577 6462 3589
rect 6408 3551 6418 3577
rect 6452 3551 6462 3577
rect 6408 3499 6409 3551
rect 6461 3499 6462 3551
rect 6408 3492 6462 3499
rect 6508 3577 6562 3773
rect 6608 3851 6662 3858
rect 6608 3799 6609 3851
rect 6661 3799 6662 3851
rect 6608 3773 6618 3799
rect 6652 3773 6662 3799
rect 6608 3761 6662 3773
rect 6708 3807 6762 3913
rect 6808 3947 6862 3959
rect 6808 3921 6818 3947
rect 6852 3921 6862 3947
rect 6808 3869 6809 3921
rect 6861 3869 6862 3921
rect 6808 3862 6862 3869
rect 6908 3947 6962 4053
rect 7008 4131 7062 4138
rect 7008 4079 7009 4131
rect 7061 4079 7062 4131
rect 7008 4053 7018 4079
rect 7052 4053 7062 4079
rect 7008 4041 7062 4053
rect 7108 4087 7162 4193
rect 7208 4227 7262 4239
rect 7208 4201 7218 4227
rect 7252 4201 7262 4227
rect 7208 4149 7209 4201
rect 7261 4149 7262 4201
rect 7208 4142 7262 4149
rect 7308 4227 7362 4333
rect 7408 4411 7462 4418
rect 7408 4359 7409 4411
rect 7461 4359 7462 4411
rect 7408 4333 7418 4359
rect 7452 4333 7462 4359
rect 7408 4321 7462 4333
rect 7508 4367 7562 4473
rect 7608 4507 7662 4519
rect 7608 4481 7618 4507
rect 7652 4481 7662 4507
rect 7608 4429 7609 4481
rect 7661 4429 7662 4481
rect 7608 4422 7662 4429
rect 7708 4507 7762 4613
rect 7808 4691 7862 4698
rect 7808 4639 7809 4691
rect 7861 4639 7862 4691
rect 7808 4613 7818 4639
rect 7852 4613 7862 4639
rect 7808 4601 7862 4613
rect 7908 4647 7962 4753
rect 8008 4787 8062 4799
rect 8008 4761 8018 4787
rect 8052 4761 8062 4787
rect 8008 4709 8009 4761
rect 8061 4709 8062 4761
rect 8008 4702 8062 4709
rect 8108 4787 8162 4960
rect 8202 4919 8268 4920
rect 8202 4867 8209 4919
rect 8261 4867 8268 4919
rect 8202 4866 8268 4867
rect 8108 4753 8118 4787
rect 8152 4753 8162 4787
rect 7908 4613 7918 4647
rect 7952 4613 7962 4647
rect 7708 4473 7718 4507
rect 7752 4473 7762 4507
rect 7508 4333 7518 4367
rect 7552 4333 7562 4367
rect 7308 4193 7318 4227
rect 7352 4193 7362 4227
rect 7108 4053 7118 4087
rect 7152 4053 7162 4087
rect 6908 3913 6918 3947
rect 6952 3913 6962 3947
rect 6708 3773 6718 3807
rect 6752 3773 6762 3807
rect 6602 3709 6668 3710
rect 6602 3657 6609 3709
rect 6661 3657 6668 3709
rect 6602 3656 6668 3657
rect 6508 3543 6518 3577
rect 6552 3543 6562 3577
rect 6308 3403 6318 3437
rect 6352 3403 6362 3437
rect 6108 3263 6118 3297
rect 6152 3263 6162 3297
rect 5908 3123 5918 3157
rect 5952 3123 5962 3157
rect 5708 2983 5718 3017
rect 5752 2983 5762 3017
rect 5508 2843 5518 2877
rect 5552 2843 5562 2877
rect 5308 2703 5318 2737
rect 5352 2703 5362 2737
rect 5108 2563 5118 2597
rect 5152 2563 5162 2597
rect 5002 2499 5068 2500
rect 5002 2447 5009 2499
rect 5061 2447 5068 2499
rect 5002 2446 5068 2447
rect 4908 2333 4918 2367
rect 4952 2333 4962 2367
rect 4708 2193 4718 2227
rect 4752 2193 4762 2227
rect 4508 2053 4518 2087
rect 4552 2053 4562 2087
rect 4308 1913 4318 1947
rect 4352 1913 4362 1947
rect 4108 1773 4118 1807
rect 4152 1773 4162 1807
rect 3908 1633 3918 1667
rect 3952 1633 3962 1667
rect 3708 1493 3718 1527
rect 3752 1493 3762 1527
rect 3508 1353 3518 1387
rect 3552 1353 3562 1387
rect 3402 1289 3468 1290
rect 3402 1237 3409 1289
rect 3461 1237 3468 1289
rect 3402 1236 3468 1237
rect 3308 1123 3318 1157
rect 3352 1123 3362 1157
rect 3108 983 3118 1017
rect 3152 983 3162 1017
rect 2908 843 2918 877
rect 2952 843 2962 877
rect 2708 703 2718 737
rect 2752 703 2762 737
rect 2508 563 2518 597
rect 2552 563 2562 597
rect 2308 423 2318 457
rect 2352 423 2362 457
rect 2108 283 2118 317
rect 2152 283 2162 317
rect 1908 143 1918 177
rect 1952 143 1962 177
rect 1802 79 1868 80
rect 1802 27 1809 79
rect 1861 27 1868 79
rect 1802 26 1868 27
rect 1708 -67 1709 -15
rect 1761 -67 1762 -15
rect 1708 -79 1718 -67
rect 1752 -79 1762 -67
rect 1508 -132 1562 -131
rect 1508 -143 1518 -132
rect 1552 -143 1562 -132
rect 1508 -195 1509 -143
rect 1561 -195 1562 -143
rect 1508 -210 1562 -195
rect 1612 -133 1658 -81
rect 1612 -167 1618 -133
rect 1652 -167 1658 -133
rect 1518 -291 1525 -239
rect 1577 -291 1584 -239
rect 1412 -397 1418 -363
rect 1452 -397 1458 -363
rect 1412 -435 1458 -397
rect 1412 -469 1418 -435
rect 1452 -469 1458 -435
rect 1412 -512 1458 -469
rect 1509 -326 1561 -320
rect 1509 -390 1518 -378
rect 1552 -390 1561 -378
rect 1509 -454 1518 -442
rect 1552 -454 1561 -442
rect 1509 -555 1561 -506
rect 1612 -363 1658 -167
rect 1708 -131 1709 -79
rect 1761 -131 1762 -79
rect 1808 -22 1862 26
rect 1808 -74 1809 -22
rect 1861 -74 1862 -22
rect 1808 -81 1862 -74
rect 1908 -15 1962 143
rect 2008 177 2062 189
rect 2008 151 2018 177
rect 2052 151 2062 177
rect 2008 99 2009 151
rect 2061 99 2062 151
rect 2008 92 2062 99
rect 2108 177 2162 283
rect 2208 361 2262 368
rect 2208 309 2209 361
rect 2261 309 2262 361
rect 2208 283 2218 309
rect 2252 283 2262 309
rect 2208 271 2262 283
rect 2308 317 2362 423
rect 2408 457 2462 469
rect 2408 431 2418 457
rect 2452 431 2462 457
rect 2408 379 2409 431
rect 2461 379 2462 431
rect 2408 372 2462 379
rect 2508 457 2562 563
rect 2608 641 2662 648
rect 2608 589 2609 641
rect 2661 589 2662 641
rect 2608 563 2618 589
rect 2652 563 2662 589
rect 2608 551 2662 563
rect 2708 597 2762 703
rect 2808 737 2862 749
rect 2808 711 2818 737
rect 2852 711 2862 737
rect 2808 659 2809 711
rect 2861 659 2862 711
rect 2808 652 2862 659
rect 2908 737 2962 843
rect 3008 921 3062 928
rect 3008 869 3009 921
rect 3061 869 3062 921
rect 3008 843 3018 869
rect 3052 843 3062 869
rect 3008 831 3062 843
rect 3108 877 3162 983
rect 3208 1017 3262 1029
rect 3208 991 3218 1017
rect 3252 991 3262 1017
rect 3208 939 3209 991
rect 3261 939 3262 991
rect 3208 932 3262 939
rect 3308 1017 3362 1123
rect 3408 1201 3462 1208
rect 3408 1149 3409 1201
rect 3461 1149 3462 1201
rect 3408 1123 3418 1149
rect 3452 1123 3462 1149
rect 3408 1111 3462 1123
rect 3508 1157 3562 1353
rect 3608 1387 3662 1399
rect 3608 1361 3618 1387
rect 3652 1361 3662 1387
rect 3608 1309 3609 1361
rect 3661 1309 3662 1361
rect 3608 1302 3662 1309
rect 3708 1387 3762 1493
rect 3808 1571 3862 1578
rect 3808 1519 3809 1571
rect 3861 1519 3862 1571
rect 3808 1493 3818 1519
rect 3852 1493 3862 1519
rect 3808 1481 3862 1493
rect 3908 1527 3962 1633
rect 4008 1667 4062 1679
rect 4008 1641 4018 1667
rect 4052 1641 4062 1667
rect 4008 1589 4009 1641
rect 4061 1589 4062 1641
rect 4008 1582 4062 1589
rect 4108 1667 4162 1773
rect 4208 1851 4262 1858
rect 4208 1799 4209 1851
rect 4261 1799 4262 1851
rect 4208 1773 4218 1799
rect 4252 1773 4262 1799
rect 4208 1761 4262 1773
rect 4308 1807 4362 1913
rect 4408 1947 4462 1959
rect 4408 1921 4418 1947
rect 4452 1921 4462 1947
rect 4408 1869 4409 1921
rect 4461 1869 4462 1921
rect 4408 1862 4462 1869
rect 4508 1947 4562 2053
rect 4608 2131 4662 2138
rect 4608 2079 4609 2131
rect 4661 2079 4662 2131
rect 4608 2053 4618 2079
rect 4652 2053 4662 2079
rect 4608 2041 4662 2053
rect 4708 2087 4762 2193
rect 4808 2227 4862 2239
rect 4808 2201 4818 2227
rect 4852 2201 4862 2227
rect 4808 2149 4809 2201
rect 4861 2149 4862 2201
rect 4808 2142 4862 2149
rect 4908 2227 4962 2333
rect 5008 2411 5062 2418
rect 5008 2359 5009 2411
rect 5061 2359 5062 2411
rect 5008 2333 5018 2359
rect 5052 2333 5062 2359
rect 5008 2321 5062 2333
rect 5108 2367 5162 2563
rect 5208 2597 5262 2609
rect 5208 2571 5218 2597
rect 5252 2571 5262 2597
rect 5208 2519 5209 2571
rect 5261 2519 5262 2571
rect 5208 2512 5262 2519
rect 5308 2597 5362 2703
rect 5408 2781 5462 2788
rect 5408 2729 5409 2781
rect 5461 2729 5462 2781
rect 5408 2703 5418 2729
rect 5452 2703 5462 2729
rect 5408 2691 5462 2703
rect 5508 2737 5562 2843
rect 5608 2877 5662 2889
rect 5608 2851 5618 2877
rect 5652 2851 5662 2877
rect 5608 2799 5609 2851
rect 5661 2799 5662 2851
rect 5608 2792 5662 2799
rect 5708 2877 5762 2983
rect 5808 3061 5862 3068
rect 5808 3009 5809 3061
rect 5861 3009 5862 3061
rect 5808 2983 5818 3009
rect 5852 2983 5862 3009
rect 5808 2971 5862 2983
rect 5908 3017 5962 3123
rect 6008 3157 6062 3169
rect 6008 3131 6018 3157
rect 6052 3131 6062 3157
rect 6008 3079 6009 3131
rect 6061 3079 6062 3131
rect 6008 3072 6062 3079
rect 6108 3157 6162 3263
rect 6208 3341 6262 3348
rect 6208 3289 6209 3341
rect 6261 3289 6262 3341
rect 6208 3263 6218 3289
rect 6252 3263 6262 3289
rect 6208 3251 6262 3263
rect 6308 3297 6362 3403
rect 6408 3437 6462 3449
rect 6408 3411 6418 3437
rect 6452 3411 6462 3437
rect 6408 3359 6409 3411
rect 6461 3359 6462 3411
rect 6408 3352 6462 3359
rect 6508 3437 6562 3543
rect 6608 3621 6662 3628
rect 6608 3569 6609 3621
rect 6661 3569 6662 3621
rect 6608 3543 6618 3569
rect 6652 3543 6662 3569
rect 6608 3531 6662 3543
rect 6708 3577 6762 3773
rect 6808 3807 6862 3819
rect 6808 3781 6818 3807
rect 6852 3781 6862 3807
rect 6808 3729 6809 3781
rect 6861 3729 6862 3781
rect 6808 3722 6862 3729
rect 6908 3807 6962 3913
rect 7008 3991 7062 3998
rect 7008 3939 7009 3991
rect 7061 3939 7062 3991
rect 7008 3913 7018 3939
rect 7052 3913 7062 3939
rect 7008 3901 7062 3913
rect 7108 3947 7162 4053
rect 7208 4087 7262 4099
rect 7208 4061 7218 4087
rect 7252 4061 7262 4087
rect 7208 4009 7209 4061
rect 7261 4009 7262 4061
rect 7208 4002 7262 4009
rect 7308 4087 7362 4193
rect 7408 4271 7462 4278
rect 7408 4219 7409 4271
rect 7461 4219 7462 4271
rect 7408 4193 7418 4219
rect 7452 4193 7462 4219
rect 7408 4181 7462 4193
rect 7508 4227 7562 4333
rect 7608 4367 7662 4379
rect 7608 4341 7618 4367
rect 7652 4341 7662 4367
rect 7608 4289 7609 4341
rect 7661 4289 7662 4341
rect 7608 4282 7662 4289
rect 7708 4367 7762 4473
rect 7808 4551 7862 4558
rect 7808 4499 7809 4551
rect 7861 4499 7862 4551
rect 7808 4473 7818 4499
rect 7852 4473 7862 4499
rect 7808 4461 7862 4473
rect 7908 4507 7962 4613
rect 8008 4647 8062 4659
rect 8008 4621 8018 4647
rect 8052 4621 8062 4647
rect 8008 4569 8009 4621
rect 8061 4569 8062 4621
rect 8008 4562 8062 4569
rect 8108 4647 8162 4753
rect 8208 4831 8262 4838
rect 8208 4779 8209 4831
rect 8261 4779 8262 4831
rect 8208 4753 8218 4779
rect 8252 4753 8262 4779
rect 8208 4741 8262 4753
rect 8308 4787 8362 4960
rect 8402 4903 8468 4904
rect 8402 4851 8409 4903
rect 8461 4851 8468 4903
rect 8402 4850 8468 4851
rect 8308 4753 8318 4787
rect 8352 4753 8362 4787
rect 8108 4613 8118 4647
rect 8152 4613 8162 4647
rect 7908 4473 7918 4507
rect 7952 4473 7962 4507
rect 7708 4333 7718 4367
rect 7752 4333 7762 4367
rect 7508 4193 7518 4227
rect 7552 4193 7562 4227
rect 7308 4053 7318 4087
rect 7352 4053 7362 4087
rect 7108 3913 7118 3947
rect 7152 3913 7162 3947
rect 6908 3773 6918 3807
rect 6952 3773 6962 3807
rect 6802 3693 6868 3694
rect 6802 3641 6809 3693
rect 6861 3641 6868 3693
rect 6802 3640 6868 3641
rect 6708 3543 6718 3577
rect 6752 3543 6762 3577
rect 6508 3403 6518 3437
rect 6552 3403 6562 3437
rect 6308 3263 6318 3297
rect 6352 3263 6362 3297
rect 6108 3123 6118 3157
rect 6152 3123 6162 3157
rect 5908 2983 5918 3017
rect 5952 2983 5962 3017
rect 5708 2843 5718 2877
rect 5752 2843 5762 2877
rect 5508 2703 5518 2737
rect 5552 2703 5562 2737
rect 5308 2563 5318 2597
rect 5352 2563 5362 2597
rect 5202 2483 5268 2484
rect 5202 2431 5209 2483
rect 5261 2431 5268 2483
rect 5202 2430 5268 2431
rect 5108 2333 5118 2367
rect 5152 2333 5162 2367
rect 4908 2193 4918 2227
rect 4952 2193 4962 2227
rect 4708 2053 4718 2087
rect 4752 2053 4762 2087
rect 4508 1913 4518 1947
rect 4552 1913 4562 1947
rect 4308 1773 4318 1807
rect 4352 1773 4362 1807
rect 4108 1633 4118 1667
rect 4152 1633 4162 1667
rect 3908 1493 3918 1527
rect 3952 1493 3962 1527
rect 3708 1353 3718 1387
rect 3752 1353 3762 1387
rect 3602 1273 3668 1274
rect 3602 1221 3609 1273
rect 3661 1221 3668 1273
rect 3602 1220 3668 1221
rect 3508 1123 3518 1157
rect 3552 1123 3562 1157
rect 3308 983 3318 1017
rect 3352 983 3362 1017
rect 3108 843 3118 877
rect 3152 843 3162 877
rect 2908 703 2918 737
rect 2952 703 2962 737
rect 2708 563 2718 597
rect 2752 563 2762 597
rect 2508 423 2518 457
rect 2552 423 2562 457
rect 2308 283 2318 317
rect 2352 283 2362 317
rect 2108 143 2118 177
rect 2152 143 2162 177
rect 2002 63 2068 64
rect 2002 11 2009 63
rect 2061 11 2068 63
rect 2002 10 2068 11
rect 1908 -67 1909 -15
rect 1961 -67 1962 -15
rect 1908 -79 1918 -67
rect 1952 -79 1962 -67
rect 1708 -132 1762 -131
rect 1708 -143 1718 -132
rect 1752 -143 1762 -132
rect 1708 -195 1709 -143
rect 1761 -195 1762 -143
rect 1708 -210 1762 -195
rect 1812 -133 1858 -81
rect 1812 -167 1818 -133
rect 1852 -167 1858 -133
rect 1718 -291 1725 -239
rect 1777 -291 1784 -239
rect 1612 -397 1618 -363
rect 1652 -397 1658 -363
rect 1612 -435 1658 -397
rect 1612 -469 1618 -435
rect 1652 -469 1658 -435
rect 1612 -512 1658 -469
rect 1709 -326 1761 -320
rect 1709 -390 1718 -378
rect 1752 -390 1761 -378
rect 1709 -454 1718 -442
rect 1752 -454 1761 -442
rect 1709 -512 1761 -506
rect 1812 -363 1858 -167
rect 1908 -131 1909 -79
rect 1961 -131 1962 -79
rect 2008 -22 2062 10
rect 2008 -74 2009 -22
rect 2061 -74 2062 -22
rect 2008 -81 2062 -74
rect 2108 -15 2162 143
rect 2208 221 2262 228
rect 2208 169 2209 221
rect 2261 169 2262 221
rect 2208 143 2218 169
rect 2252 143 2262 169
rect 2208 131 2262 143
rect 2308 177 2362 283
rect 2408 317 2462 329
rect 2408 291 2418 317
rect 2452 291 2462 317
rect 2408 239 2409 291
rect 2461 239 2462 291
rect 2408 232 2462 239
rect 2508 317 2562 423
rect 2608 501 2662 508
rect 2608 449 2609 501
rect 2661 449 2662 501
rect 2608 423 2618 449
rect 2652 423 2662 449
rect 2608 411 2662 423
rect 2708 457 2762 563
rect 2808 597 2862 609
rect 2808 571 2818 597
rect 2852 571 2862 597
rect 2808 519 2809 571
rect 2861 519 2862 571
rect 2808 512 2862 519
rect 2908 597 2962 703
rect 3008 781 3062 788
rect 3008 729 3009 781
rect 3061 729 3062 781
rect 3008 703 3018 729
rect 3052 703 3062 729
rect 3008 691 3062 703
rect 3108 737 3162 843
rect 3208 877 3262 889
rect 3208 851 3218 877
rect 3252 851 3262 877
rect 3208 799 3209 851
rect 3261 799 3262 851
rect 3208 792 3262 799
rect 3308 877 3362 983
rect 3408 1061 3462 1068
rect 3408 1009 3409 1061
rect 3461 1009 3462 1061
rect 3408 983 3418 1009
rect 3452 983 3462 1009
rect 3408 971 3462 983
rect 3508 1017 3562 1123
rect 3608 1157 3662 1169
rect 3608 1131 3618 1157
rect 3652 1131 3662 1157
rect 3608 1079 3609 1131
rect 3661 1079 3662 1131
rect 3608 1072 3662 1079
rect 3708 1157 3762 1353
rect 3808 1431 3862 1438
rect 3808 1379 3809 1431
rect 3861 1379 3862 1431
rect 3808 1353 3818 1379
rect 3852 1353 3862 1379
rect 3808 1341 3862 1353
rect 3908 1387 3962 1493
rect 4008 1527 4062 1539
rect 4008 1501 4018 1527
rect 4052 1501 4062 1527
rect 4008 1449 4009 1501
rect 4061 1449 4062 1501
rect 4008 1442 4062 1449
rect 4108 1527 4162 1633
rect 4208 1711 4262 1718
rect 4208 1659 4209 1711
rect 4261 1659 4262 1711
rect 4208 1633 4218 1659
rect 4252 1633 4262 1659
rect 4208 1621 4262 1633
rect 4308 1667 4362 1773
rect 4408 1807 4462 1819
rect 4408 1781 4418 1807
rect 4452 1781 4462 1807
rect 4408 1729 4409 1781
rect 4461 1729 4462 1781
rect 4408 1722 4462 1729
rect 4508 1807 4562 1913
rect 4608 1991 4662 1998
rect 4608 1939 4609 1991
rect 4661 1939 4662 1991
rect 4608 1913 4618 1939
rect 4652 1913 4662 1939
rect 4608 1901 4662 1913
rect 4708 1947 4762 2053
rect 4808 2087 4862 2099
rect 4808 2061 4818 2087
rect 4852 2061 4862 2087
rect 4808 2009 4809 2061
rect 4861 2009 4862 2061
rect 4808 2002 4862 2009
rect 4908 2087 4962 2193
rect 5008 2271 5062 2278
rect 5008 2219 5009 2271
rect 5061 2219 5062 2271
rect 5008 2193 5018 2219
rect 5052 2193 5062 2219
rect 5008 2181 5062 2193
rect 5108 2227 5162 2333
rect 5208 2367 5262 2379
rect 5208 2341 5218 2367
rect 5252 2341 5262 2367
rect 5208 2289 5209 2341
rect 5261 2289 5262 2341
rect 5208 2282 5262 2289
rect 5308 2367 5362 2563
rect 5408 2641 5462 2648
rect 5408 2589 5409 2641
rect 5461 2589 5462 2641
rect 5408 2563 5418 2589
rect 5452 2563 5462 2589
rect 5408 2551 5462 2563
rect 5508 2597 5562 2703
rect 5608 2737 5662 2749
rect 5608 2711 5618 2737
rect 5652 2711 5662 2737
rect 5608 2659 5609 2711
rect 5661 2659 5662 2711
rect 5608 2652 5662 2659
rect 5708 2737 5762 2843
rect 5808 2921 5862 2928
rect 5808 2869 5809 2921
rect 5861 2869 5862 2921
rect 5808 2843 5818 2869
rect 5852 2843 5862 2869
rect 5808 2831 5862 2843
rect 5908 2877 5962 2983
rect 6008 3017 6062 3029
rect 6008 2991 6018 3017
rect 6052 2991 6062 3017
rect 6008 2939 6009 2991
rect 6061 2939 6062 2991
rect 6008 2932 6062 2939
rect 6108 3017 6162 3123
rect 6208 3201 6262 3208
rect 6208 3149 6209 3201
rect 6261 3149 6262 3201
rect 6208 3123 6218 3149
rect 6252 3123 6262 3149
rect 6208 3111 6262 3123
rect 6308 3157 6362 3263
rect 6408 3297 6462 3309
rect 6408 3271 6418 3297
rect 6452 3271 6462 3297
rect 6408 3219 6409 3271
rect 6461 3219 6462 3271
rect 6408 3212 6462 3219
rect 6508 3297 6562 3403
rect 6608 3481 6662 3488
rect 6608 3429 6609 3481
rect 6661 3429 6662 3481
rect 6608 3403 6618 3429
rect 6652 3403 6662 3429
rect 6608 3391 6662 3403
rect 6708 3437 6762 3543
rect 6808 3577 6862 3589
rect 6808 3551 6818 3577
rect 6852 3551 6862 3577
rect 6808 3499 6809 3551
rect 6861 3499 6862 3551
rect 6808 3492 6862 3499
rect 6908 3577 6962 3773
rect 7008 3851 7062 3858
rect 7008 3799 7009 3851
rect 7061 3799 7062 3851
rect 7008 3773 7018 3799
rect 7052 3773 7062 3799
rect 7008 3761 7062 3773
rect 7108 3807 7162 3913
rect 7208 3947 7262 3959
rect 7208 3921 7218 3947
rect 7252 3921 7262 3947
rect 7208 3869 7209 3921
rect 7261 3869 7262 3921
rect 7208 3862 7262 3869
rect 7308 3947 7362 4053
rect 7408 4131 7462 4138
rect 7408 4079 7409 4131
rect 7461 4079 7462 4131
rect 7408 4053 7418 4079
rect 7452 4053 7462 4079
rect 7408 4041 7462 4053
rect 7508 4087 7562 4193
rect 7608 4227 7662 4239
rect 7608 4201 7618 4227
rect 7652 4201 7662 4227
rect 7608 4149 7609 4201
rect 7661 4149 7662 4201
rect 7608 4142 7662 4149
rect 7708 4227 7762 4333
rect 7808 4411 7862 4418
rect 7808 4359 7809 4411
rect 7861 4359 7862 4411
rect 7808 4333 7818 4359
rect 7852 4333 7862 4359
rect 7808 4321 7862 4333
rect 7908 4367 7962 4473
rect 8008 4507 8062 4519
rect 8008 4481 8018 4507
rect 8052 4481 8062 4507
rect 8008 4429 8009 4481
rect 8061 4429 8062 4481
rect 8008 4422 8062 4429
rect 8108 4507 8162 4613
rect 8208 4691 8262 4698
rect 8208 4639 8209 4691
rect 8261 4639 8262 4691
rect 8208 4613 8218 4639
rect 8252 4613 8262 4639
rect 8208 4601 8262 4613
rect 8308 4647 8362 4753
rect 8408 4787 8462 4799
rect 8408 4761 8418 4787
rect 8452 4761 8462 4787
rect 8408 4709 8409 4761
rect 8461 4709 8462 4761
rect 8408 4702 8462 4709
rect 8508 4787 8562 4960
rect 8602 4919 8668 4920
rect 8602 4867 8609 4919
rect 8661 4867 8668 4919
rect 8602 4866 8668 4867
rect 8508 4753 8518 4787
rect 8552 4753 8562 4787
rect 8308 4613 8318 4647
rect 8352 4613 8362 4647
rect 8108 4473 8118 4507
rect 8152 4473 8162 4507
rect 7908 4333 7918 4367
rect 7952 4333 7962 4367
rect 7708 4193 7718 4227
rect 7752 4193 7762 4227
rect 7508 4053 7518 4087
rect 7552 4053 7562 4087
rect 7308 3913 7318 3947
rect 7352 3913 7362 3947
rect 7108 3773 7118 3807
rect 7152 3773 7162 3807
rect 7002 3709 7068 3710
rect 7002 3657 7009 3709
rect 7061 3657 7068 3709
rect 7002 3656 7068 3657
rect 6908 3543 6918 3577
rect 6952 3543 6962 3577
rect 6708 3403 6718 3437
rect 6752 3403 6762 3437
rect 6508 3263 6518 3297
rect 6552 3263 6562 3297
rect 6308 3123 6318 3157
rect 6352 3123 6362 3157
rect 6108 2983 6118 3017
rect 6152 2983 6162 3017
rect 5908 2843 5918 2877
rect 5952 2843 5962 2877
rect 5708 2703 5718 2737
rect 5752 2703 5762 2737
rect 5508 2563 5518 2597
rect 5552 2563 5562 2597
rect 5402 2499 5468 2500
rect 5402 2447 5409 2499
rect 5461 2447 5468 2499
rect 5402 2446 5468 2447
rect 5308 2333 5318 2367
rect 5352 2333 5362 2367
rect 5108 2193 5118 2227
rect 5152 2193 5162 2227
rect 4908 2053 4918 2087
rect 4952 2053 4962 2087
rect 4708 1913 4718 1947
rect 4752 1913 4762 1947
rect 4508 1773 4518 1807
rect 4552 1773 4562 1807
rect 4308 1633 4318 1667
rect 4352 1633 4362 1667
rect 4108 1493 4118 1527
rect 4152 1493 4162 1527
rect 3908 1353 3918 1387
rect 3952 1353 3962 1387
rect 3802 1289 3868 1290
rect 3802 1237 3809 1289
rect 3861 1237 3868 1289
rect 3802 1236 3868 1237
rect 3708 1123 3718 1157
rect 3752 1123 3762 1157
rect 3508 983 3518 1017
rect 3552 983 3562 1017
rect 3308 843 3318 877
rect 3352 843 3362 877
rect 3108 703 3118 737
rect 3152 703 3162 737
rect 2908 563 2918 597
rect 2952 563 2962 597
rect 2708 423 2718 457
rect 2752 423 2762 457
rect 2508 283 2518 317
rect 2552 283 2562 317
rect 2308 143 2318 177
rect 2352 143 2362 177
rect 2202 79 2268 80
rect 2202 27 2209 79
rect 2261 27 2268 79
rect 2202 26 2268 27
rect 2108 -67 2109 -15
rect 2161 -67 2162 -15
rect 2108 -79 2118 -67
rect 2152 -79 2162 -67
rect 1908 -132 1962 -131
rect 1908 -143 1918 -132
rect 1952 -143 1962 -132
rect 1908 -195 1909 -143
rect 1961 -195 1962 -143
rect 1908 -210 1962 -195
rect 2012 -133 2058 -81
rect 2012 -167 2018 -133
rect 2052 -167 2058 -133
rect 1918 -291 1925 -239
rect 1977 -291 1984 -239
rect 1812 -397 1818 -363
rect 1852 -397 1858 -363
rect 1812 -435 1858 -397
rect 1812 -469 1818 -435
rect 1852 -469 1858 -435
rect 1812 -512 1858 -469
rect 1909 -326 1961 -320
rect 1909 -390 1918 -378
rect 1952 -390 1961 -378
rect 1909 -454 1918 -442
rect 1952 -454 1961 -442
rect 1909 -555 1961 -506
rect 2012 -363 2058 -167
rect 2108 -131 2109 -79
rect 2161 -131 2162 -79
rect 2208 -22 2262 26
rect 2208 -74 2209 -22
rect 2261 -74 2262 -22
rect 2208 -81 2262 -74
rect 2308 -15 2362 143
rect 2408 177 2462 189
rect 2408 151 2418 177
rect 2452 151 2462 177
rect 2408 99 2409 151
rect 2461 99 2462 151
rect 2408 92 2462 99
rect 2508 177 2562 283
rect 2608 361 2662 368
rect 2608 309 2609 361
rect 2661 309 2662 361
rect 2608 283 2618 309
rect 2652 283 2662 309
rect 2608 271 2662 283
rect 2708 317 2762 423
rect 2808 457 2862 469
rect 2808 431 2818 457
rect 2852 431 2862 457
rect 2808 379 2809 431
rect 2861 379 2862 431
rect 2808 372 2862 379
rect 2908 457 2962 563
rect 3008 641 3062 648
rect 3008 589 3009 641
rect 3061 589 3062 641
rect 3008 563 3018 589
rect 3052 563 3062 589
rect 3008 551 3062 563
rect 3108 597 3162 703
rect 3208 737 3262 749
rect 3208 711 3218 737
rect 3252 711 3262 737
rect 3208 659 3209 711
rect 3261 659 3262 711
rect 3208 652 3262 659
rect 3308 737 3362 843
rect 3408 921 3462 928
rect 3408 869 3409 921
rect 3461 869 3462 921
rect 3408 843 3418 869
rect 3452 843 3462 869
rect 3408 831 3462 843
rect 3508 877 3562 983
rect 3608 1017 3662 1029
rect 3608 991 3618 1017
rect 3652 991 3662 1017
rect 3608 939 3609 991
rect 3661 939 3662 991
rect 3608 932 3662 939
rect 3708 1017 3762 1123
rect 3808 1201 3862 1208
rect 3808 1149 3809 1201
rect 3861 1149 3862 1201
rect 3808 1123 3818 1149
rect 3852 1123 3862 1149
rect 3808 1111 3862 1123
rect 3908 1157 3962 1353
rect 4008 1387 4062 1399
rect 4008 1361 4018 1387
rect 4052 1361 4062 1387
rect 4008 1309 4009 1361
rect 4061 1309 4062 1361
rect 4008 1302 4062 1309
rect 4108 1387 4162 1493
rect 4208 1571 4262 1578
rect 4208 1519 4209 1571
rect 4261 1519 4262 1571
rect 4208 1493 4218 1519
rect 4252 1493 4262 1519
rect 4208 1481 4262 1493
rect 4308 1527 4362 1633
rect 4408 1667 4462 1679
rect 4408 1641 4418 1667
rect 4452 1641 4462 1667
rect 4408 1589 4409 1641
rect 4461 1589 4462 1641
rect 4408 1582 4462 1589
rect 4508 1667 4562 1773
rect 4608 1851 4662 1858
rect 4608 1799 4609 1851
rect 4661 1799 4662 1851
rect 4608 1773 4618 1799
rect 4652 1773 4662 1799
rect 4608 1761 4662 1773
rect 4708 1807 4762 1913
rect 4808 1947 4862 1959
rect 4808 1921 4818 1947
rect 4852 1921 4862 1947
rect 4808 1869 4809 1921
rect 4861 1869 4862 1921
rect 4808 1862 4862 1869
rect 4908 1947 4962 2053
rect 5008 2131 5062 2138
rect 5008 2079 5009 2131
rect 5061 2079 5062 2131
rect 5008 2053 5018 2079
rect 5052 2053 5062 2079
rect 5008 2041 5062 2053
rect 5108 2087 5162 2193
rect 5208 2227 5262 2239
rect 5208 2201 5218 2227
rect 5252 2201 5262 2227
rect 5208 2149 5209 2201
rect 5261 2149 5262 2201
rect 5208 2142 5262 2149
rect 5308 2227 5362 2333
rect 5408 2411 5462 2418
rect 5408 2359 5409 2411
rect 5461 2359 5462 2411
rect 5408 2333 5418 2359
rect 5452 2333 5462 2359
rect 5408 2321 5462 2333
rect 5508 2367 5562 2563
rect 5608 2597 5662 2609
rect 5608 2571 5618 2597
rect 5652 2571 5662 2597
rect 5608 2519 5609 2571
rect 5661 2519 5662 2571
rect 5608 2512 5662 2519
rect 5708 2597 5762 2703
rect 5808 2781 5862 2788
rect 5808 2729 5809 2781
rect 5861 2729 5862 2781
rect 5808 2703 5818 2729
rect 5852 2703 5862 2729
rect 5808 2691 5862 2703
rect 5908 2737 5962 2843
rect 6008 2877 6062 2889
rect 6008 2851 6018 2877
rect 6052 2851 6062 2877
rect 6008 2799 6009 2851
rect 6061 2799 6062 2851
rect 6008 2792 6062 2799
rect 6108 2877 6162 2983
rect 6208 3061 6262 3068
rect 6208 3009 6209 3061
rect 6261 3009 6262 3061
rect 6208 2983 6218 3009
rect 6252 2983 6262 3009
rect 6208 2971 6262 2983
rect 6308 3017 6362 3123
rect 6408 3157 6462 3169
rect 6408 3131 6418 3157
rect 6452 3131 6462 3157
rect 6408 3079 6409 3131
rect 6461 3079 6462 3131
rect 6408 3072 6462 3079
rect 6508 3157 6562 3263
rect 6608 3341 6662 3348
rect 6608 3289 6609 3341
rect 6661 3289 6662 3341
rect 6608 3263 6618 3289
rect 6652 3263 6662 3289
rect 6608 3251 6662 3263
rect 6708 3297 6762 3403
rect 6808 3437 6862 3449
rect 6808 3411 6818 3437
rect 6852 3411 6862 3437
rect 6808 3359 6809 3411
rect 6861 3359 6862 3411
rect 6808 3352 6862 3359
rect 6908 3437 6962 3543
rect 7008 3621 7062 3628
rect 7008 3569 7009 3621
rect 7061 3569 7062 3621
rect 7008 3543 7018 3569
rect 7052 3543 7062 3569
rect 7008 3531 7062 3543
rect 7108 3577 7162 3773
rect 7208 3807 7262 3819
rect 7208 3781 7218 3807
rect 7252 3781 7262 3807
rect 7208 3729 7209 3781
rect 7261 3729 7262 3781
rect 7208 3722 7262 3729
rect 7308 3807 7362 3913
rect 7408 3991 7462 3998
rect 7408 3939 7409 3991
rect 7461 3939 7462 3991
rect 7408 3913 7418 3939
rect 7452 3913 7462 3939
rect 7408 3901 7462 3913
rect 7508 3947 7562 4053
rect 7608 4087 7662 4099
rect 7608 4061 7618 4087
rect 7652 4061 7662 4087
rect 7608 4009 7609 4061
rect 7661 4009 7662 4061
rect 7608 4002 7662 4009
rect 7708 4087 7762 4193
rect 7808 4271 7862 4278
rect 7808 4219 7809 4271
rect 7861 4219 7862 4271
rect 7808 4193 7818 4219
rect 7852 4193 7862 4219
rect 7808 4181 7862 4193
rect 7908 4227 7962 4333
rect 8008 4367 8062 4379
rect 8008 4341 8018 4367
rect 8052 4341 8062 4367
rect 8008 4289 8009 4341
rect 8061 4289 8062 4341
rect 8008 4282 8062 4289
rect 8108 4367 8162 4473
rect 8208 4551 8262 4558
rect 8208 4499 8209 4551
rect 8261 4499 8262 4551
rect 8208 4473 8218 4499
rect 8252 4473 8262 4499
rect 8208 4461 8262 4473
rect 8308 4507 8362 4613
rect 8408 4647 8462 4659
rect 8408 4621 8418 4647
rect 8452 4621 8462 4647
rect 8408 4569 8409 4621
rect 8461 4569 8462 4621
rect 8408 4562 8462 4569
rect 8508 4647 8562 4753
rect 8608 4831 8662 4838
rect 8608 4779 8609 4831
rect 8661 4779 8662 4831
rect 8608 4753 8618 4779
rect 8652 4753 8662 4779
rect 8608 4741 8662 4753
rect 8708 4787 8762 4960
rect 8802 4903 8868 4904
rect 8802 4851 8809 4903
rect 8861 4851 8868 4903
rect 8802 4850 8868 4851
rect 8708 4753 8718 4787
rect 8752 4753 8762 4787
rect 8508 4613 8518 4647
rect 8552 4613 8562 4647
rect 8308 4473 8318 4507
rect 8352 4473 8362 4507
rect 8108 4333 8118 4367
rect 8152 4333 8162 4367
rect 7908 4193 7918 4227
rect 7952 4193 7962 4227
rect 7708 4053 7718 4087
rect 7752 4053 7762 4087
rect 7508 3913 7518 3947
rect 7552 3913 7562 3947
rect 7308 3773 7318 3807
rect 7352 3773 7362 3807
rect 7202 3693 7268 3694
rect 7202 3641 7209 3693
rect 7261 3641 7268 3693
rect 7202 3640 7268 3641
rect 7108 3543 7118 3577
rect 7152 3543 7162 3577
rect 6908 3403 6918 3437
rect 6952 3403 6962 3437
rect 6708 3263 6718 3297
rect 6752 3263 6762 3297
rect 6508 3123 6518 3157
rect 6552 3123 6562 3157
rect 6308 2983 6318 3017
rect 6352 2983 6362 3017
rect 6108 2843 6118 2877
rect 6152 2843 6162 2877
rect 5908 2703 5918 2737
rect 5952 2703 5962 2737
rect 5708 2563 5718 2597
rect 5752 2563 5762 2597
rect 5602 2483 5668 2484
rect 5602 2431 5609 2483
rect 5661 2431 5668 2483
rect 5602 2430 5668 2431
rect 5508 2333 5518 2367
rect 5552 2333 5562 2367
rect 5308 2193 5318 2227
rect 5352 2193 5362 2227
rect 5108 2053 5118 2087
rect 5152 2053 5162 2087
rect 4908 1913 4918 1947
rect 4952 1913 4962 1947
rect 4708 1773 4718 1807
rect 4752 1773 4762 1807
rect 4508 1633 4518 1667
rect 4552 1633 4562 1667
rect 4308 1493 4318 1527
rect 4352 1493 4362 1527
rect 4108 1353 4118 1387
rect 4152 1353 4162 1387
rect 4002 1273 4068 1274
rect 4002 1221 4009 1273
rect 4061 1221 4068 1273
rect 4002 1220 4068 1221
rect 3908 1123 3918 1157
rect 3952 1123 3962 1157
rect 3708 983 3718 1017
rect 3752 983 3762 1017
rect 3508 843 3518 877
rect 3552 843 3562 877
rect 3308 703 3318 737
rect 3352 703 3362 737
rect 3108 563 3118 597
rect 3152 563 3162 597
rect 2908 423 2918 457
rect 2952 423 2962 457
rect 2708 283 2718 317
rect 2752 283 2762 317
rect 2508 143 2518 177
rect 2552 143 2562 177
rect 2402 63 2468 64
rect 2402 11 2409 63
rect 2461 11 2468 63
rect 2402 10 2468 11
rect 2308 -67 2309 -15
rect 2361 -67 2362 -15
rect 2308 -79 2318 -67
rect 2352 -79 2362 -67
rect 2108 -132 2162 -131
rect 2108 -143 2118 -132
rect 2152 -143 2162 -132
rect 2108 -195 2109 -143
rect 2161 -195 2162 -143
rect 2108 -210 2162 -195
rect 2212 -133 2258 -81
rect 2212 -167 2218 -133
rect 2252 -167 2258 -133
rect 2118 -291 2125 -239
rect 2177 -291 2184 -239
rect 2012 -397 2018 -363
rect 2052 -397 2058 -363
rect 2012 -435 2058 -397
rect 2012 -469 2018 -435
rect 2052 -469 2058 -435
rect 2012 -512 2058 -469
rect 2109 -326 2161 -320
rect 2109 -390 2118 -378
rect 2152 -390 2161 -378
rect 2109 -454 2118 -442
rect 2152 -454 2161 -442
rect 2109 -512 2161 -506
rect 2212 -363 2258 -167
rect 2308 -131 2309 -79
rect 2361 -131 2362 -79
rect 2408 -22 2462 10
rect 2408 -74 2409 -22
rect 2461 -74 2462 -22
rect 2408 -81 2462 -74
rect 2508 -15 2562 143
rect 2608 221 2662 228
rect 2608 169 2609 221
rect 2661 169 2662 221
rect 2608 143 2618 169
rect 2652 143 2662 169
rect 2608 131 2662 143
rect 2708 177 2762 283
rect 2808 317 2862 329
rect 2808 291 2818 317
rect 2852 291 2862 317
rect 2808 239 2809 291
rect 2861 239 2862 291
rect 2808 232 2862 239
rect 2908 317 2962 423
rect 3008 501 3062 508
rect 3008 449 3009 501
rect 3061 449 3062 501
rect 3008 423 3018 449
rect 3052 423 3062 449
rect 3008 411 3062 423
rect 3108 457 3162 563
rect 3208 597 3262 609
rect 3208 571 3218 597
rect 3252 571 3262 597
rect 3208 519 3209 571
rect 3261 519 3262 571
rect 3208 512 3262 519
rect 3308 597 3362 703
rect 3408 781 3462 788
rect 3408 729 3409 781
rect 3461 729 3462 781
rect 3408 703 3418 729
rect 3452 703 3462 729
rect 3408 691 3462 703
rect 3508 737 3562 843
rect 3608 877 3662 889
rect 3608 851 3618 877
rect 3652 851 3662 877
rect 3608 799 3609 851
rect 3661 799 3662 851
rect 3608 792 3662 799
rect 3708 877 3762 983
rect 3808 1061 3862 1068
rect 3808 1009 3809 1061
rect 3861 1009 3862 1061
rect 3808 983 3818 1009
rect 3852 983 3862 1009
rect 3808 971 3862 983
rect 3908 1017 3962 1123
rect 4008 1157 4062 1169
rect 4008 1131 4018 1157
rect 4052 1131 4062 1157
rect 4008 1079 4009 1131
rect 4061 1079 4062 1131
rect 4008 1072 4062 1079
rect 4108 1157 4162 1353
rect 4208 1431 4262 1438
rect 4208 1379 4209 1431
rect 4261 1379 4262 1431
rect 4208 1353 4218 1379
rect 4252 1353 4262 1379
rect 4208 1341 4262 1353
rect 4308 1387 4362 1493
rect 4408 1527 4462 1539
rect 4408 1501 4418 1527
rect 4452 1501 4462 1527
rect 4408 1449 4409 1501
rect 4461 1449 4462 1501
rect 4408 1442 4462 1449
rect 4508 1527 4562 1633
rect 4608 1711 4662 1718
rect 4608 1659 4609 1711
rect 4661 1659 4662 1711
rect 4608 1633 4618 1659
rect 4652 1633 4662 1659
rect 4608 1621 4662 1633
rect 4708 1667 4762 1773
rect 4808 1807 4862 1819
rect 4808 1781 4818 1807
rect 4852 1781 4862 1807
rect 4808 1729 4809 1781
rect 4861 1729 4862 1781
rect 4808 1722 4862 1729
rect 4908 1807 4962 1913
rect 5008 1991 5062 1998
rect 5008 1939 5009 1991
rect 5061 1939 5062 1991
rect 5008 1913 5018 1939
rect 5052 1913 5062 1939
rect 5008 1901 5062 1913
rect 5108 1947 5162 2053
rect 5208 2087 5262 2099
rect 5208 2061 5218 2087
rect 5252 2061 5262 2087
rect 5208 2009 5209 2061
rect 5261 2009 5262 2061
rect 5208 2002 5262 2009
rect 5308 2087 5362 2193
rect 5408 2271 5462 2278
rect 5408 2219 5409 2271
rect 5461 2219 5462 2271
rect 5408 2193 5418 2219
rect 5452 2193 5462 2219
rect 5408 2181 5462 2193
rect 5508 2227 5562 2333
rect 5608 2367 5662 2379
rect 5608 2341 5618 2367
rect 5652 2341 5662 2367
rect 5608 2289 5609 2341
rect 5661 2289 5662 2341
rect 5608 2282 5662 2289
rect 5708 2367 5762 2563
rect 5808 2641 5862 2648
rect 5808 2589 5809 2641
rect 5861 2589 5862 2641
rect 5808 2563 5818 2589
rect 5852 2563 5862 2589
rect 5808 2551 5862 2563
rect 5908 2597 5962 2703
rect 6008 2737 6062 2749
rect 6008 2711 6018 2737
rect 6052 2711 6062 2737
rect 6008 2659 6009 2711
rect 6061 2659 6062 2711
rect 6008 2652 6062 2659
rect 6108 2737 6162 2843
rect 6208 2921 6262 2928
rect 6208 2869 6209 2921
rect 6261 2869 6262 2921
rect 6208 2843 6218 2869
rect 6252 2843 6262 2869
rect 6208 2831 6262 2843
rect 6308 2877 6362 2983
rect 6408 3017 6462 3029
rect 6408 2991 6418 3017
rect 6452 2991 6462 3017
rect 6408 2939 6409 2991
rect 6461 2939 6462 2991
rect 6408 2932 6462 2939
rect 6508 3017 6562 3123
rect 6608 3201 6662 3208
rect 6608 3149 6609 3201
rect 6661 3149 6662 3201
rect 6608 3123 6618 3149
rect 6652 3123 6662 3149
rect 6608 3111 6662 3123
rect 6708 3157 6762 3263
rect 6808 3297 6862 3309
rect 6808 3271 6818 3297
rect 6852 3271 6862 3297
rect 6808 3219 6809 3271
rect 6861 3219 6862 3271
rect 6808 3212 6862 3219
rect 6908 3297 6962 3403
rect 7008 3481 7062 3488
rect 7008 3429 7009 3481
rect 7061 3429 7062 3481
rect 7008 3403 7018 3429
rect 7052 3403 7062 3429
rect 7008 3391 7062 3403
rect 7108 3437 7162 3543
rect 7208 3577 7262 3589
rect 7208 3551 7218 3577
rect 7252 3551 7262 3577
rect 7208 3499 7209 3551
rect 7261 3499 7262 3551
rect 7208 3492 7262 3499
rect 7308 3577 7362 3773
rect 7408 3851 7462 3858
rect 7408 3799 7409 3851
rect 7461 3799 7462 3851
rect 7408 3773 7418 3799
rect 7452 3773 7462 3799
rect 7408 3761 7462 3773
rect 7508 3807 7562 3913
rect 7608 3947 7662 3959
rect 7608 3921 7618 3947
rect 7652 3921 7662 3947
rect 7608 3869 7609 3921
rect 7661 3869 7662 3921
rect 7608 3862 7662 3869
rect 7708 3947 7762 4053
rect 7808 4131 7862 4138
rect 7808 4079 7809 4131
rect 7861 4079 7862 4131
rect 7808 4053 7818 4079
rect 7852 4053 7862 4079
rect 7808 4041 7862 4053
rect 7908 4087 7962 4193
rect 8008 4227 8062 4239
rect 8008 4201 8018 4227
rect 8052 4201 8062 4227
rect 8008 4149 8009 4201
rect 8061 4149 8062 4201
rect 8008 4142 8062 4149
rect 8108 4227 8162 4333
rect 8208 4411 8262 4418
rect 8208 4359 8209 4411
rect 8261 4359 8262 4411
rect 8208 4333 8218 4359
rect 8252 4333 8262 4359
rect 8208 4321 8262 4333
rect 8308 4367 8362 4473
rect 8408 4507 8462 4519
rect 8408 4481 8418 4507
rect 8452 4481 8462 4507
rect 8408 4429 8409 4481
rect 8461 4429 8462 4481
rect 8408 4422 8462 4429
rect 8508 4507 8562 4613
rect 8608 4691 8662 4698
rect 8608 4639 8609 4691
rect 8661 4639 8662 4691
rect 8608 4613 8618 4639
rect 8652 4613 8662 4639
rect 8608 4601 8662 4613
rect 8708 4647 8762 4753
rect 8808 4787 8862 4799
rect 8808 4761 8818 4787
rect 8852 4761 8862 4787
rect 8808 4709 8809 4761
rect 8861 4709 8862 4761
rect 8808 4702 8862 4709
rect 8908 4787 8962 4960
rect 9002 4919 9068 4920
rect 9002 4867 9009 4919
rect 9061 4867 9068 4919
rect 9002 4866 9068 4867
rect 8908 4753 8918 4787
rect 8952 4753 8962 4787
rect 8708 4613 8718 4647
rect 8752 4613 8762 4647
rect 8508 4473 8518 4507
rect 8552 4473 8562 4507
rect 8308 4333 8318 4367
rect 8352 4333 8362 4367
rect 8108 4193 8118 4227
rect 8152 4193 8162 4227
rect 7908 4053 7918 4087
rect 7952 4053 7962 4087
rect 7708 3913 7718 3947
rect 7752 3913 7762 3947
rect 7508 3773 7518 3807
rect 7552 3773 7562 3807
rect 7402 3709 7468 3710
rect 7402 3657 7409 3709
rect 7461 3657 7468 3709
rect 7402 3656 7468 3657
rect 7308 3543 7318 3577
rect 7352 3543 7362 3577
rect 7108 3403 7118 3437
rect 7152 3403 7162 3437
rect 6908 3263 6918 3297
rect 6952 3263 6962 3297
rect 6708 3123 6718 3157
rect 6752 3123 6762 3157
rect 6508 2983 6518 3017
rect 6552 2983 6562 3017
rect 6308 2843 6318 2877
rect 6352 2843 6362 2877
rect 6108 2703 6118 2737
rect 6152 2703 6162 2737
rect 5908 2563 5918 2597
rect 5952 2563 5962 2597
rect 5802 2499 5868 2500
rect 5802 2447 5809 2499
rect 5861 2447 5868 2499
rect 5802 2446 5868 2447
rect 5708 2333 5718 2367
rect 5752 2333 5762 2367
rect 5508 2193 5518 2227
rect 5552 2193 5562 2227
rect 5308 2053 5318 2087
rect 5352 2053 5362 2087
rect 5108 1913 5118 1947
rect 5152 1913 5162 1947
rect 4908 1773 4918 1807
rect 4952 1773 4962 1807
rect 4708 1633 4718 1667
rect 4752 1633 4762 1667
rect 4508 1493 4518 1527
rect 4552 1493 4562 1527
rect 4308 1353 4318 1387
rect 4352 1353 4362 1387
rect 4202 1289 4268 1290
rect 4202 1237 4209 1289
rect 4261 1237 4268 1289
rect 4202 1236 4268 1237
rect 4108 1123 4118 1157
rect 4152 1123 4162 1157
rect 3908 983 3918 1017
rect 3952 983 3962 1017
rect 3708 843 3718 877
rect 3752 843 3762 877
rect 3508 703 3518 737
rect 3552 703 3562 737
rect 3308 563 3318 597
rect 3352 563 3362 597
rect 3108 423 3118 457
rect 3152 423 3162 457
rect 2908 283 2918 317
rect 2952 283 2962 317
rect 2708 143 2718 177
rect 2752 143 2762 177
rect 2602 79 2668 80
rect 2602 27 2609 79
rect 2661 27 2668 79
rect 2602 26 2668 27
rect 2508 -67 2509 -15
rect 2561 -67 2562 -15
rect 2508 -79 2518 -67
rect 2552 -79 2562 -67
rect 2308 -132 2362 -131
rect 2308 -143 2318 -132
rect 2352 -143 2362 -132
rect 2308 -195 2309 -143
rect 2361 -195 2362 -143
rect 2308 -210 2362 -195
rect 2412 -133 2458 -81
rect 2412 -167 2418 -133
rect 2452 -167 2458 -133
rect 2318 -291 2325 -239
rect 2377 -291 2384 -239
rect 2212 -397 2218 -363
rect 2252 -397 2258 -363
rect 2212 -435 2258 -397
rect 2212 -469 2218 -435
rect 2252 -469 2258 -435
rect 2212 -512 2258 -469
rect 2309 -326 2361 -320
rect 2309 -390 2318 -378
rect 2352 -390 2361 -378
rect 2309 -454 2318 -442
rect 2352 -454 2361 -442
rect 2309 -555 2361 -506
rect 2412 -363 2458 -167
rect 2508 -131 2509 -79
rect 2561 -131 2562 -79
rect 2608 -22 2662 26
rect 2608 -74 2609 -22
rect 2661 -74 2662 -22
rect 2608 -81 2662 -74
rect 2708 -15 2762 143
rect 2808 177 2862 189
rect 2808 151 2818 177
rect 2852 151 2862 177
rect 2808 99 2809 151
rect 2861 99 2862 151
rect 2808 92 2862 99
rect 2908 177 2962 283
rect 3008 361 3062 368
rect 3008 309 3009 361
rect 3061 309 3062 361
rect 3008 283 3018 309
rect 3052 283 3062 309
rect 3008 271 3062 283
rect 3108 317 3162 423
rect 3208 457 3262 469
rect 3208 431 3218 457
rect 3252 431 3262 457
rect 3208 379 3209 431
rect 3261 379 3262 431
rect 3208 372 3262 379
rect 3308 457 3362 563
rect 3408 641 3462 648
rect 3408 589 3409 641
rect 3461 589 3462 641
rect 3408 563 3418 589
rect 3452 563 3462 589
rect 3408 551 3462 563
rect 3508 597 3562 703
rect 3608 737 3662 749
rect 3608 711 3618 737
rect 3652 711 3662 737
rect 3608 659 3609 711
rect 3661 659 3662 711
rect 3608 652 3662 659
rect 3708 737 3762 843
rect 3808 921 3862 928
rect 3808 869 3809 921
rect 3861 869 3862 921
rect 3808 843 3818 869
rect 3852 843 3862 869
rect 3808 831 3862 843
rect 3908 877 3962 983
rect 4008 1017 4062 1029
rect 4008 991 4018 1017
rect 4052 991 4062 1017
rect 4008 939 4009 991
rect 4061 939 4062 991
rect 4008 932 4062 939
rect 4108 1017 4162 1123
rect 4208 1201 4262 1208
rect 4208 1149 4209 1201
rect 4261 1149 4262 1201
rect 4208 1123 4218 1149
rect 4252 1123 4262 1149
rect 4208 1111 4262 1123
rect 4308 1157 4362 1353
rect 4408 1387 4462 1399
rect 4408 1361 4418 1387
rect 4452 1361 4462 1387
rect 4408 1309 4409 1361
rect 4461 1309 4462 1361
rect 4408 1302 4462 1309
rect 4508 1387 4562 1493
rect 4608 1571 4662 1578
rect 4608 1519 4609 1571
rect 4661 1519 4662 1571
rect 4608 1493 4618 1519
rect 4652 1493 4662 1519
rect 4608 1481 4662 1493
rect 4708 1527 4762 1633
rect 4808 1667 4862 1679
rect 4808 1641 4818 1667
rect 4852 1641 4862 1667
rect 4808 1589 4809 1641
rect 4861 1589 4862 1641
rect 4808 1582 4862 1589
rect 4908 1667 4962 1773
rect 5008 1851 5062 1858
rect 5008 1799 5009 1851
rect 5061 1799 5062 1851
rect 5008 1773 5018 1799
rect 5052 1773 5062 1799
rect 5008 1761 5062 1773
rect 5108 1807 5162 1913
rect 5208 1947 5262 1959
rect 5208 1921 5218 1947
rect 5252 1921 5262 1947
rect 5208 1869 5209 1921
rect 5261 1869 5262 1921
rect 5208 1862 5262 1869
rect 5308 1947 5362 2053
rect 5408 2131 5462 2138
rect 5408 2079 5409 2131
rect 5461 2079 5462 2131
rect 5408 2053 5418 2079
rect 5452 2053 5462 2079
rect 5408 2041 5462 2053
rect 5508 2087 5562 2193
rect 5608 2227 5662 2239
rect 5608 2201 5618 2227
rect 5652 2201 5662 2227
rect 5608 2149 5609 2201
rect 5661 2149 5662 2201
rect 5608 2142 5662 2149
rect 5708 2227 5762 2333
rect 5808 2411 5862 2418
rect 5808 2359 5809 2411
rect 5861 2359 5862 2411
rect 5808 2333 5818 2359
rect 5852 2333 5862 2359
rect 5808 2321 5862 2333
rect 5908 2367 5962 2563
rect 6008 2597 6062 2609
rect 6008 2571 6018 2597
rect 6052 2571 6062 2597
rect 6008 2519 6009 2571
rect 6061 2519 6062 2571
rect 6008 2512 6062 2519
rect 6108 2597 6162 2703
rect 6208 2781 6262 2788
rect 6208 2729 6209 2781
rect 6261 2729 6262 2781
rect 6208 2703 6218 2729
rect 6252 2703 6262 2729
rect 6208 2691 6262 2703
rect 6308 2737 6362 2843
rect 6408 2877 6462 2889
rect 6408 2851 6418 2877
rect 6452 2851 6462 2877
rect 6408 2799 6409 2851
rect 6461 2799 6462 2851
rect 6408 2792 6462 2799
rect 6508 2877 6562 2983
rect 6608 3061 6662 3068
rect 6608 3009 6609 3061
rect 6661 3009 6662 3061
rect 6608 2983 6618 3009
rect 6652 2983 6662 3009
rect 6608 2971 6662 2983
rect 6708 3017 6762 3123
rect 6808 3157 6862 3169
rect 6808 3131 6818 3157
rect 6852 3131 6862 3157
rect 6808 3079 6809 3131
rect 6861 3079 6862 3131
rect 6808 3072 6862 3079
rect 6908 3157 6962 3263
rect 7008 3341 7062 3348
rect 7008 3289 7009 3341
rect 7061 3289 7062 3341
rect 7008 3263 7018 3289
rect 7052 3263 7062 3289
rect 7008 3251 7062 3263
rect 7108 3297 7162 3403
rect 7208 3437 7262 3449
rect 7208 3411 7218 3437
rect 7252 3411 7262 3437
rect 7208 3359 7209 3411
rect 7261 3359 7262 3411
rect 7208 3352 7262 3359
rect 7308 3437 7362 3543
rect 7408 3621 7462 3628
rect 7408 3569 7409 3621
rect 7461 3569 7462 3621
rect 7408 3543 7418 3569
rect 7452 3543 7462 3569
rect 7408 3531 7462 3543
rect 7508 3577 7562 3773
rect 7608 3807 7662 3819
rect 7608 3781 7618 3807
rect 7652 3781 7662 3807
rect 7608 3729 7609 3781
rect 7661 3729 7662 3781
rect 7608 3722 7662 3729
rect 7708 3807 7762 3913
rect 7808 3991 7862 3998
rect 7808 3939 7809 3991
rect 7861 3939 7862 3991
rect 7808 3913 7818 3939
rect 7852 3913 7862 3939
rect 7808 3901 7862 3913
rect 7908 3947 7962 4053
rect 8008 4087 8062 4099
rect 8008 4061 8018 4087
rect 8052 4061 8062 4087
rect 8008 4009 8009 4061
rect 8061 4009 8062 4061
rect 8008 4002 8062 4009
rect 8108 4087 8162 4193
rect 8208 4271 8262 4278
rect 8208 4219 8209 4271
rect 8261 4219 8262 4271
rect 8208 4193 8218 4219
rect 8252 4193 8262 4219
rect 8208 4181 8262 4193
rect 8308 4227 8362 4333
rect 8408 4367 8462 4379
rect 8408 4341 8418 4367
rect 8452 4341 8462 4367
rect 8408 4289 8409 4341
rect 8461 4289 8462 4341
rect 8408 4282 8462 4289
rect 8508 4367 8562 4473
rect 8608 4551 8662 4558
rect 8608 4499 8609 4551
rect 8661 4499 8662 4551
rect 8608 4473 8618 4499
rect 8652 4473 8662 4499
rect 8608 4461 8662 4473
rect 8708 4507 8762 4613
rect 8808 4647 8862 4659
rect 8808 4621 8818 4647
rect 8852 4621 8862 4647
rect 8808 4569 8809 4621
rect 8861 4569 8862 4621
rect 8808 4562 8862 4569
rect 8908 4647 8962 4753
rect 9008 4831 9062 4838
rect 9008 4779 9009 4831
rect 9061 4779 9062 4831
rect 9008 4753 9018 4779
rect 9052 4753 9062 4779
rect 9008 4741 9062 4753
rect 9108 4787 9162 4960
rect 9202 4903 9268 4904
rect 9202 4851 9209 4903
rect 9261 4851 9268 4903
rect 9202 4850 9268 4851
rect 9108 4753 9118 4787
rect 9152 4753 9162 4787
rect 8908 4613 8918 4647
rect 8952 4613 8962 4647
rect 8708 4473 8718 4507
rect 8752 4473 8762 4507
rect 8508 4333 8518 4367
rect 8552 4333 8562 4367
rect 8308 4193 8318 4227
rect 8352 4193 8362 4227
rect 8108 4053 8118 4087
rect 8152 4053 8162 4087
rect 7908 3913 7918 3947
rect 7952 3913 7962 3947
rect 7708 3773 7718 3807
rect 7752 3773 7762 3807
rect 7602 3693 7668 3694
rect 7602 3641 7609 3693
rect 7661 3641 7668 3693
rect 7602 3640 7668 3641
rect 7508 3543 7518 3577
rect 7552 3543 7562 3577
rect 7308 3403 7318 3437
rect 7352 3403 7362 3437
rect 7108 3263 7118 3297
rect 7152 3263 7162 3297
rect 6908 3123 6918 3157
rect 6952 3123 6962 3157
rect 6708 2983 6718 3017
rect 6752 2983 6762 3017
rect 6508 2843 6518 2877
rect 6552 2843 6562 2877
rect 6308 2703 6318 2737
rect 6352 2703 6362 2737
rect 6108 2563 6118 2597
rect 6152 2563 6162 2597
rect 6002 2483 6068 2484
rect 6002 2431 6009 2483
rect 6061 2431 6068 2483
rect 6002 2430 6068 2431
rect 5908 2333 5918 2367
rect 5952 2333 5962 2367
rect 5708 2193 5718 2227
rect 5752 2193 5762 2227
rect 5508 2053 5518 2087
rect 5552 2053 5562 2087
rect 5308 1913 5318 1947
rect 5352 1913 5362 1947
rect 5108 1773 5118 1807
rect 5152 1773 5162 1807
rect 4908 1633 4918 1667
rect 4952 1633 4962 1667
rect 4708 1493 4718 1527
rect 4752 1493 4762 1527
rect 4508 1353 4518 1387
rect 4552 1353 4562 1387
rect 4402 1273 4468 1274
rect 4402 1221 4409 1273
rect 4461 1221 4468 1273
rect 4402 1220 4468 1221
rect 4308 1123 4318 1157
rect 4352 1123 4362 1157
rect 4108 983 4118 1017
rect 4152 983 4162 1017
rect 3908 843 3918 877
rect 3952 843 3962 877
rect 3708 703 3718 737
rect 3752 703 3762 737
rect 3508 563 3518 597
rect 3552 563 3562 597
rect 3308 423 3318 457
rect 3352 423 3362 457
rect 3108 283 3118 317
rect 3152 283 3162 317
rect 2908 143 2918 177
rect 2952 143 2962 177
rect 2802 63 2868 64
rect 2802 11 2809 63
rect 2861 11 2868 63
rect 2802 10 2868 11
rect 2708 -67 2709 -15
rect 2761 -67 2762 -15
rect 2708 -79 2718 -67
rect 2752 -79 2762 -67
rect 2508 -132 2562 -131
rect 2508 -143 2518 -132
rect 2552 -143 2562 -132
rect 2508 -195 2509 -143
rect 2561 -195 2562 -143
rect 2508 -210 2562 -195
rect 2612 -133 2658 -81
rect 2612 -167 2618 -133
rect 2652 -167 2658 -133
rect 2518 -291 2525 -239
rect 2577 -291 2584 -239
rect 2412 -397 2418 -363
rect 2452 -397 2458 -363
rect 2412 -435 2458 -397
rect 2412 -469 2418 -435
rect 2452 -469 2458 -435
rect 2412 -512 2458 -469
rect 2509 -326 2561 -320
rect 2509 -390 2518 -378
rect 2552 -390 2561 -378
rect 2509 -454 2518 -442
rect 2552 -454 2561 -442
rect 2509 -512 2561 -506
rect 2612 -363 2658 -167
rect 2708 -131 2709 -79
rect 2761 -131 2762 -79
rect 2808 -22 2862 10
rect 2808 -74 2809 -22
rect 2861 -74 2862 -22
rect 2808 -81 2862 -74
rect 2908 -15 2962 143
rect 3008 221 3062 228
rect 3008 169 3009 221
rect 3061 169 3062 221
rect 3008 143 3018 169
rect 3052 143 3062 169
rect 3008 131 3062 143
rect 3108 177 3162 283
rect 3208 317 3262 329
rect 3208 291 3218 317
rect 3252 291 3262 317
rect 3208 239 3209 291
rect 3261 239 3262 291
rect 3208 232 3262 239
rect 3308 317 3362 423
rect 3408 501 3462 508
rect 3408 449 3409 501
rect 3461 449 3462 501
rect 3408 423 3418 449
rect 3452 423 3462 449
rect 3408 411 3462 423
rect 3508 457 3562 563
rect 3608 597 3662 609
rect 3608 571 3618 597
rect 3652 571 3662 597
rect 3608 519 3609 571
rect 3661 519 3662 571
rect 3608 512 3662 519
rect 3708 597 3762 703
rect 3808 781 3862 788
rect 3808 729 3809 781
rect 3861 729 3862 781
rect 3808 703 3818 729
rect 3852 703 3862 729
rect 3808 691 3862 703
rect 3908 737 3962 843
rect 4008 877 4062 889
rect 4008 851 4018 877
rect 4052 851 4062 877
rect 4008 799 4009 851
rect 4061 799 4062 851
rect 4008 792 4062 799
rect 4108 877 4162 983
rect 4208 1061 4262 1068
rect 4208 1009 4209 1061
rect 4261 1009 4262 1061
rect 4208 983 4218 1009
rect 4252 983 4262 1009
rect 4208 971 4262 983
rect 4308 1017 4362 1123
rect 4408 1157 4462 1169
rect 4408 1131 4418 1157
rect 4452 1131 4462 1157
rect 4408 1079 4409 1131
rect 4461 1079 4462 1131
rect 4408 1072 4462 1079
rect 4508 1157 4562 1353
rect 4608 1431 4662 1438
rect 4608 1379 4609 1431
rect 4661 1379 4662 1431
rect 4608 1353 4618 1379
rect 4652 1353 4662 1379
rect 4608 1341 4662 1353
rect 4708 1387 4762 1493
rect 4808 1527 4862 1539
rect 4808 1501 4818 1527
rect 4852 1501 4862 1527
rect 4808 1449 4809 1501
rect 4861 1449 4862 1501
rect 4808 1442 4862 1449
rect 4908 1527 4962 1633
rect 5008 1711 5062 1718
rect 5008 1659 5009 1711
rect 5061 1659 5062 1711
rect 5008 1633 5018 1659
rect 5052 1633 5062 1659
rect 5008 1621 5062 1633
rect 5108 1667 5162 1773
rect 5208 1807 5262 1819
rect 5208 1781 5218 1807
rect 5252 1781 5262 1807
rect 5208 1729 5209 1781
rect 5261 1729 5262 1781
rect 5208 1722 5262 1729
rect 5308 1807 5362 1913
rect 5408 1991 5462 1998
rect 5408 1939 5409 1991
rect 5461 1939 5462 1991
rect 5408 1913 5418 1939
rect 5452 1913 5462 1939
rect 5408 1901 5462 1913
rect 5508 1947 5562 2053
rect 5608 2087 5662 2099
rect 5608 2061 5618 2087
rect 5652 2061 5662 2087
rect 5608 2009 5609 2061
rect 5661 2009 5662 2061
rect 5608 2002 5662 2009
rect 5708 2087 5762 2193
rect 5808 2271 5862 2278
rect 5808 2219 5809 2271
rect 5861 2219 5862 2271
rect 5808 2193 5818 2219
rect 5852 2193 5862 2219
rect 5808 2181 5862 2193
rect 5908 2227 5962 2333
rect 6008 2367 6062 2379
rect 6008 2341 6018 2367
rect 6052 2341 6062 2367
rect 6008 2289 6009 2341
rect 6061 2289 6062 2341
rect 6008 2282 6062 2289
rect 6108 2367 6162 2563
rect 6208 2641 6262 2648
rect 6208 2589 6209 2641
rect 6261 2589 6262 2641
rect 6208 2563 6218 2589
rect 6252 2563 6262 2589
rect 6208 2551 6262 2563
rect 6308 2597 6362 2703
rect 6408 2737 6462 2749
rect 6408 2711 6418 2737
rect 6452 2711 6462 2737
rect 6408 2659 6409 2711
rect 6461 2659 6462 2711
rect 6408 2652 6462 2659
rect 6508 2737 6562 2843
rect 6608 2921 6662 2928
rect 6608 2869 6609 2921
rect 6661 2869 6662 2921
rect 6608 2843 6618 2869
rect 6652 2843 6662 2869
rect 6608 2831 6662 2843
rect 6708 2877 6762 2983
rect 6808 3017 6862 3029
rect 6808 2991 6818 3017
rect 6852 2991 6862 3017
rect 6808 2939 6809 2991
rect 6861 2939 6862 2991
rect 6808 2932 6862 2939
rect 6908 3017 6962 3123
rect 7008 3201 7062 3208
rect 7008 3149 7009 3201
rect 7061 3149 7062 3201
rect 7008 3123 7018 3149
rect 7052 3123 7062 3149
rect 7008 3111 7062 3123
rect 7108 3157 7162 3263
rect 7208 3297 7262 3309
rect 7208 3271 7218 3297
rect 7252 3271 7262 3297
rect 7208 3219 7209 3271
rect 7261 3219 7262 3271
rect 7208 3212 7262 3219
rect 7308 3297 7362 3403
rect 7408 3481 7462 3488
rect 7408 3429 7409 3481
rect 7461 3429 7462 3481
rect 7408 3403 7418 3429
rect 7452 3403 7462 3429
rect 7408 3391 7462 3403
rect 7508 3437 7562 3543
rect 7608 3577 7662 3589
rect 7608 3551 7618 3577
rect 7652 3551 7662 3577
rect 7608 3499 7609 3551
rect 7661 3499 7662 3551
rect 7608 3492 7662 3499
rect 7708 3577 7762 3773
rect 7808 3851 7862 3858
rect 7808 3799 7809 3851
rect 7861 3799 7862 3851
rect 7808 3773 7818 3799
rect 7852 3773 7862 3799
rect 7808 3761 7862 3773
rect 7908 3807 7962 3913
rect 8008 3947 8062 3959
rect 8008 3921 8018 3947
rect 8052 3921 8062 3947
rect 8008 3869 8009 3921
rect 8061 3869 8062 3921
rect 8008 3862 8062 3869
rect 8108 3947 8162 4053
rect 8208 4131 8262 4138
rect 8208 4079 8209 4131
rect 8261 4079 8262 4131
rect 8208 4053 8218 4079
rect 8252 4053 8262 4079
rect 8208 4041 8262 4053
rect 8308 4087 8362 4193
rect 8408 4227 8462 4239
rect 8408 4201 8418 4227
rect 8452 4201 8462 4227
rect 8408 4149 8409 4201
rect 8461 4149 8462 4201
rect 8408 4142 8462 4149
rect 8508 4227 8562 4333
rect 8608 4411 8662 4418
rect 8608 4359 8609 4411
rect 8661 4359 8662 4411
rect 8608 4333 8618 4359
rect 8652 4333 8662 4359
rect 8608 4321 8662 4333
rect 8708 4367 8762 4473
rect 8808 4507 8862 4519
rect 8808 4481 8818 4507
rect 8852 4481 8862 4507
rect 8808 4429 8809 4481
rect 8861 4429 8862 4481
rect 8808 4422 8862 4429
rect 8908 4507 8962 4613
rect 9008 4691 9062 4698
rect 9008 4639 9009 4691
rect 9061 4639 9062 4691
rect 9008 4613 9018 4639
rect 9052 4613 9062 4639
rect 9008 4601 9062 4613
rect 9108 4647 9162 4753
rect 9208 4787 9262 4799
rect 9208 4761 9218 4787
rect 9252 4761 9262 4787
rect 9208 4709 9209 4761
rect 9261 4709 9262 4761
rect 9208 4702 9262 4709
rect 9308 4787 9362 4960
rect 9402 4919 9468 4920
rect 9402 4867 9409 4919
rect 9461 4867 9468 4919
rect 9402 4866 9468 4867
rect 9308 4753 9318 4787
rect 9352 4753 9362 4787
rect 9108 4613 9118 4647
rect 9152 4613 9162 4647
rect 8908 4473 8918 4507
rect 8952 4473 8962 4507
rect 8708 4333 8718 4367
rect 8752 4333 8762 4367
rect 8508 4193 8518 4227
rect 8552 4193 8562 4227
rect 8308 4053 8318 4087
rect 8352 4053 8362 4087
rect 8108 3913 8118 3947
rect 8152 3913 8162 3947
rect 7908 3773 7918 3807
rect 7952 3773 7962 3807
rect 7802 3709 7868 3710
rect 7802 3657 7809 3709
rect 7861 3657 7868 3709
rect 7802 3656 7868 3657
rect 7708 3543 7718 3577
rect 7752 3543 7762 3577
rect 7508 3403 7518 3437
rect 7552 3403 7562 3437
rect 7308 3263 7318 3297
rect 7352 3263 7362 3297
rect 7108 3123 7118 3157
rect 7152 3123 7162 3157
rect 6908 2983 6918 3017
rect 6952 2983 6962 3017
rect 6708 2843 6718 2877
rect 6752 2843 6762 2877
rect 6508 2703 6518 2737
rect 6552 2703 6562 2737
rect 6308 2563 6318 2597
rect 6352 2563 6362 2597
rect 6202 2499 6268 2500
rect 6202 2447 6209 2499
rect 6261 2447 6268 2499
rect 6202 2446 6268 2447
rect 6108 2333 6118 2367
rect 6152 2333 6162 2367
rect 5908 2193 5918 2227
rect 5952 2193 5962 2227
rect 5708 2053 5718 2087
rect 5752 2053 5762 2087
rect 5508 1913 5518 1947
rect 5552 1913 5562 1947
rect 5308 1773 5318 1807
rect 5352 1773 5362 1807
rect 5108 1633 5118 1667
rect 5152 1633 5162 1667
rect 4908 1493 4918 1527
rect 4952 1493 4962 1527
rect 4708 1353 4718 1387
rect 4752 1353 4762 1387
rect 4602 1289 4668 1290
rect 4602 1237 4609 1289
rect 4661 1237 4668 1289
rect 4602 1236 4668 1237
rect 4508 1123 4518 1157
rect 4552 1123 4562 1157
rect 4308 983 4318 1017
rect 4352 983 4362 1017
rect 4108 843 4118 877
rect 4152 843 4162 877
rect 3908 703 3918 737
rect 3952 703 3962 737
rect 3708 563 3718 597
rect 3752 563 3762 597
rect 3508 423 3518 457
rect 3552 423 3562 457
rect 3308 283 3318 317
rect 3352 283 3362 317
rect 3108 143 3118 177
rect 3152 143 3162 177
rect 3002 79 3068 80
rect 3002 27 3009 79
rect 3061 27 3068 79
rect 3002 26 3068 27
rect 2908 -67 2909 -15
rect 2961 -67 2962 -15
rect 2908 -79 2918 -67
rect 2952 -79 2962 -67
rect 2708 -132 2762 -131
rect 2708 -143 2718 -132
rect 2752 -143 2762 -132
rect 2708 -195 2709 -143
rect 2761 -195 2762 -143
rect 2708 -210 2762 -195
rect 2812 -133 2858 -81
rect 2812 -167 2818 -133
rect 2852 -167 2858 -133
rect 2718 -291 2725 -239
rect 2777 -291 2784 -239
rect 2612 -397 2618 -363
rect 2652 -397 2658 -363
rect 2612 -435 2658 -397
rect 2612 -469 2618 -435
rect 2652 -469 2658 -435
rect 2612 -512 2658 -469
rect 2709 -326 2761 -320
rect 2709 -390 2718 -378
rect 2752 -390 2761 -378
rect 2709 -454 2718 -442
rect 2752 -454 2761 -442
rect 2709 -555 2761 -506
rect 2812 -363 2858 -167
rect 2908 -131 2909 -79
rect 2961 -131 2962 -79
rect 3008 -22 3062 26
rect 3008 -74 3009 -22
rect 3061 -74 3062 -22
rect 3008 -81 3062 -74
rect 3108 -15 3162 143
rect 3208 177 3262 189
rect 3208 151 3218 177
rect 3252 151 3262 177
rect 3208 99 3209 151
rect 3261 99 3262 151
rect 3208 92 3262 99
rect 3308 177 3362 283
rect 3408 361 3462 368
rect 3408 309 3409 361
rect 3461 309 3462 361
rect 3408 283 3418 309
rect 3452 283 3462 309
rect 3408 271 3462 283
rect 3508 317 3562 423
rect 3608 457 3662 469
rect 3608 431 3618 457
rect 3652 431 3662 457
rect 3608 379 3609 431
rect 3661 379 3662 431
rect 3608 372 3662 379
rect 3708 457 3762 563
rect 3808 641 3862 648
rect 3808 589 3809 641
rect 3861 589 3862 641
rect 3808 563 3818 589
rect 3852 563 3862 589
rect 3808 551 3862 563
rect 3908 597 3962 703
rect 4008 737 4062 749
rect 4008 711 4018 737
rect 4052 711 4062 737
rect 4008 659 4009 711
rect 4061 659 4062 711
rect 4008 652 4062 659
rect 4108 737 4162 843
rect 4208 921 4262 928
rect 4208 869 4209 921
rect 4261 869 4262 921
rect 4208 843 4218 869
rect 4252 843 4262 869
rect 4208 831 4262 843
rect 4308 877 4362 983
rect 4408 1017 4462 1029
rect 4408 991 4418 1017
rect 4452 991 4462 1017
rect 4408 939 4409 991
rect 4461 939 4462 991
rect 4408 932 4462 939
rect 4508 1017 4562 1123
rect 4608 1201 4662 1208
rect 4608 1149 4609 1201
rect 4661 1149 4662 1201
rect 4608 1123 4618 1149
rect 4652 1123 4662 1149
rect 4608 1111 4662 1123
rect 4708 1157 4762 1353
rect 4808 1387 4862 1399
rect 4808 1361 4818 1387
rect 4852 1361 4862 1387
rect 4808 1309 4809 1361
rect 4861 1309 4862 1361
rect 4808 1302 4862 1309
rect 4908 1387 4962 1493
rect 5008 1571 5062 1578
rect 5008 1519 5009 1571
rect 5061 1519 5062 1571
rect 5008 1493 5018 1519
rect 5052 1493 5062 1519
rect 5008 1481 5062 1493
rect 5108 1527 5162 1633
rect 5208 1667 5262 1679
rect 5208 1641 5218 1667
rect 5252 1641 5262 1667
rect 5208 1589 5209 1641
rect 5261 1589 5262 1641
rect 5208 1582 5262 1589
rect 5308 1667 5362 1773
rect 5408 1851 5462 1858
rect 5408 1799 5409 1851
rect 5461 1799 5462 1851
rect 5408 1773 5418 1799
rect 5452 1773 5462 1799
rect 5408 1761 5462 1773
rect 5508 1807 5562 1913
rect 5608 1947 5662 1959
rect 5608 1921 5618 1947
rect 5652 1921 5662 1947
rect 5608 1869 5609 1921
rect 5661 1869 5662 1921
rect 5608 1862 5662 1869
rect 5708 1947 5762 2053
rect 5808 2131 5862 2138
rect 5808 2079 5809 2131
rect 5861 2079 5862 2131
rect 5808 2053 5818 2079
rect 5852 2053 5862 2079
rect 5808 2041 5862 2053
rect 5908 2087 5962 2193
rect 6008 2227 6062 2239
rect 6008 2201 6018 2227
rect 6052 2201 6062 2227
rect 6008 2149 6009 2201
rect 6061 2149 6062 2201
rect 6008 2142 6062 2149
rect 6108 2227 6162 2333
rect 6208 2411 6262 2418
rect 6208 2359 6209 2411
rect 6261 2359 6262 2411
rect 6208 2333 6218 2359
rect 6252 2333 6262 2359
rect 6208 2321 6262 2333
rect 6308 2367 6362 2563
rect 6408 2597 6462 2609
rect 6408 2571 6418 2597
rect 6452 2571 6462 2597
rect 6408 2519 6409 2571
rect 6461 2519 6462 2571
rect 6408 2512 6462 2519
rect 6508 2597 6562 2703
rect 6608 2781 6662 2788
rect 6608 2729 6609 2781
rect 6661 2729 6662 2781
rect 6608 2703 6618 2729
rect 6652 2703 6662 2729
rect 6608 2691 6662 2703
rect 6708 2737 6762 2843
rect 6808 2877 6862 2889
rect 6808 2851 6818 2877
rect 6852 2851 6862 2877
rect 6808 2799 6809 2851
rect 6861 2799 6862 2851
rect 6808 2792 6862 2799
rect 6908 2877 6962 2983
rect 7008 3061 7062 3068
rect 7008 3009 7009 3061
rect 7061 3009 7062 3061
rect 7008 2983 7018 3009
rect 7052 2983 7062 3009
rect 7008 2971 7062 2983
rect 7108 3017 7162 3123
rect 7208 3157 7262 3169
rect 7208 3131 7218 3157
rect 7252 3131 7262 3157
rect 7208 3079 7209 3131
rect 7261 3079 7262 3131
rect 7208 3072 7262 3079
rect 7308 3157 7362 3263
rect 7408 3341 7462 3348
rect 7408 3289 7409 3341
rect 7461 3289 7462 3341
rect 7408 3263 7418 3289
rect 7452 3263 7462 3289
rect 7408 3251 7462 3263
rect 7508 3297 7562 3403
rect 7608 3437 7662 3449
rect 7608 3411 7618 3437
rect 7652 3411 7662 3437
rect 7608 3359 7609 3411
rect 7661 3359 7662 3411
rect 7608 3352 7662 3359
rect 7708 3437 7762 3543
rect 7808 3621 7862 3628
rect 7808 3569 7809 3621
rect 7861 3569 7862 3621
rect 7808 3543 7818 3569
rect 7852 3543 7862 3569
rect 7808 3531 7862 3543
rect 7908 3577 7962 3773
rect 8008 3807 8062 3819
rect 8008 3781 8018 3807
rect 8052 3781 8062 3807
rect 8008 3729 8009 3781
rect 8061 3729 8062 3781
rect 8008 3722 8062 3729
rect 8108 3807 8162 3913
rect 8208 3991 8262 3998
rect 8208 3939 8209 3991
rect 8261 3939 8262 3991
rect 8208 3913 8218 3939
rect 8252 3913 8262 3939
rect 8208 3901 8262 3913
rect 8308 3947 8362 4053
rect 8408 4087 8462 4099
rect 8408 4061 8418 4087
rect 8452 4061 8462 4087
rect 8408 4009 8409 4061
rect 8461 4009 8462 4061
rect 8408 4002 8462 4009
rect 8508 4087 8562 4193
rect 8608 4271 8662 4278
rect 8608 4219 8609 4271
rect 8661 4219 8662 4271
rect 8608 4193 8618 4219
rect 8652 4193 8662 4219
rect 8608 4181 8662 4193
rect 8708 4227 8762 4333
rect 8808 4367 8862 4379
rect 8808 4341 8818 4367
rect 8852 4341 8862 4367
rect 8808 4289 8809 4341
rect 8861 4289 8862 4341
rect 8808 4282 8862 4289
rect 8908 4367 8962 4473
rect 9008 4551 9062 4558
rect 9008 4499 9009 4551
rect 9061 4499 9062 4551
rect 9008 4473 9018 4499
rect 9052 4473 9062 4499
rect 9008 4461 9062 4473
rect 9108 4507 9162 4613
rect 9208 4647 9262 4659
rect 9208 4621 9218 4647
rect 9252 4621 9262 4647
rect 9208 4569 9209 4621
rect 9261 4569 9262 4621
rect 9208 4562 9262 4569
rect 9308 4647 9362 4753
rect 9408 4831 9462 4838
rect 9408 4779 9409 4831
rect 9461 4779 9462 4831
rect 9408 4753 9418 4779
rect 9452 4753 9462 4779
rect 9408 4741 9462 4753
rect 9508 4787 9562 4960
rect 9602 4903 9668 4904
rect 9602 4851 9609 4903
rect 9661 4851 9668 4903
rect 9602 4850 9668 4851
rect 9508 4753 9518 4787
rect 9552 4753 9562 4787
rect 9308 4613 9318 4647
rect 9352 4613 9362 4647
rect 9108 4473 9118 4507
rect 9152 4473 9162 4507
rect 8908 4333 8918 4367
rect 8952 4333 8962 4367
rect 8708 4193 8718 4227
rect 8752 4193 8762 4227
rect 8508 4053 8518 4087
rect 8552 4053 8562 4087
rect 8308 3913 8318 3947
rect 8352 3913 8362 3947
rect 8108 3773 8118 3807
rect 8152 3773 8162 3807
rect 8002 3693 8068 3694
rect 8002 3641 8009 3693
rect 8061 3641 8068 3693
rect 8002 3640 8068 3641
rect 7908 3543 7918 3577
rect 7952 3543 7962 3577
rect 7708 3403 7718 3437
rect 7752 3403 7762 3437
rect 7508 3263 7518 3297
rect 7552 3263 7562 3297
rect 7308 3123 7318 3157
rect 7352 3123 7362 3157
rect 7108 2983 7118 3017
rect 7152 2983 7162 3017
rect 6908 2843 6918 2877
rect 6952 2843 6962 2877
rect 6708 2703 6718 2737
rect 6752 2703 6762 2737
rect 6508 2563 6518 2597
rect 6552 2563 6562 2597
rect 6402 2483 6468 2484
rect 6402 2431 6409 2483
rect 6461 2431 6468 2483
rect 6402 2430 6468 2431
rect 6308 2333 6318 2367
rect 6352 2333 6362 2367
rect 6108 2193 6118 2227
rect 6152 2193 6162 2227
rect 5908 2053 5918 2087
rect 5952 2053 5962 2087
rect 5708 1913 5718 1947
rect 5752 1913 5762 1947
rect 5508 1773 5518 1807
rect 5552 1773 5562 1807
rect 5308 1633 5318 1667
rect 5352 1633 5362 1667
rect 5108 1493 5118 1527
rect 5152 1493 5162 1527
rect 4908 1353 4918 1387
rect 4952 1353 4962 1387
rect 4802 1273 4868 1274
rect 4802 1221 4809 1273
rect 4861 1221 4868 1273
rect 4802 1220 4868 1221
rect 4708 1123 4718 1157
rect 4752 1123 4762 1157
rect 4508 983 4518 1017
rect 4552 983 4562 1017
rect 4308 843 4318 877
rect 4352 843 4362 877
rect 4108 703 4118 737
rect 4152 703 4162 737
rect 3908 563 3918 597
rect 3952 563 3962 597
rect 3708 423 3718 457
rect 3752 423 3762 457
rect 3508 283 3518 317
rect 3552 283 3562 317
rect 3308 143 3318 177
rect 3352 143 3362 177
rect 3202 63 3268 64
rect 3202 11 3209 63
rect 3261 11 3268 63
rect 3202 10 3268 11
rect 3108 -67 3109 -15
rect 3161 -67 3162 -15
rect 3108 -79 3118 -67
rect 3152 -79 3162 -67
rect 2908 -132 2962 -131
rect 2908 -143 2918 -132
rect 2952 -143 2962 -132
rect 2908 -195 2909 -143
rect 2961 -195 2962 -143
rect 2908 -210 2962 -195
rect 3012 -133 3058 -81
rect 3012 -167 3018 -133
rect 3052 -167 3058 -133
rect 2918 -291 2925 -239
rect 2977 -291 2984 -239
rect 2812 -397 2818 -363
rect 2852 -397 2858 -363
rect 2812 -435 2858 -397
rect 2812 -469 2818 -435
rect 2852 -469 2858 -435
rect 2812 -512 2858 -469
rect 2909 -326 2961 -320
rect 2909 -390 2918 -378
rect 2952 -390 2961 -378
rect 2909 -454 2918 -442
rect 2952 -454 2961 -442
rect 2909 -512 2961 -506
rect 3012 -363 3058 -167
rect 3108 -131 3109 -79
rect 3161 -131 3162 -79
rect 3208 -22 3262 10
rect 3208 -74 3209 -22
rect 3261 -74 3262 -22
rect 3208 -81 3262 -74
rect 3308 -15 3362 143
rect 3408 221 3462 228
rect 3408 169 3409 221
rect 3461 169 3462 221
rect 3408 143 3418 169
rect 3452 143 3462 169
rect 3408 131 3462 143
rect 3508 177 3562 283
rect 3608 317 3662 329
rect 3608 291 3618 317
rect 3652 291 3662 317
rect 3608 239 3609 291
rect 3661 239 3662 291
rect 3608 232 3662 239
rect 3708 317 3762 423
rect 3808 501 3862 508
rect 3808 449 3809 501
rect 3861 449 3862 501
rect 3808 423 3818 449
rect 3852 423 3862 449
rect 3808 411 3862 423
rect 3908 457 3962 563
rect 4008 597 4062 609
rect 4008 571 4018 597
rect 4052 571 4062 597
rect 4008 519 4009 571
rect 4061 519 4062 571
rect 4008 512 4062 519
rect 4108 597 4162 703
rect 4208 781 4262 788
rect 4208 729 4209 781
rect 4261 729 4262 781
rect 4208 703 4218 729
rect 4252 703 4262 729
rect 4208 691 4262 703
rect 4308 737 4362 843
rect 4408 877 4462 889
rect 4408 851 4418 877
rect 4452 851 4462 877
rect 4408 799 4409 851
rect 4461 799 4462 851
rect 4408 792 4462 799
rect 4508 877 4562 983
rect 4608 1061 4662 1068
rect 4608 1009 4609 1061
rect 4661 1009 4662 1061
rect 4608 983 4618 1009
rect 4652 983 4662 1009
rect 4608 971 4662 983
rect 4708 1017 4762 1123
rect 4808 1157 4862 1169
rect 4808 1131 4818 1157
rect 4852 1131 4862 1157
rect 4808 1079 4809 1131
rect 4861 1079 4862 1131
rect 4808 1072 4862 1079
rect 4908 1157 4962 1353
rect 5008 1431 5062 1438
rect 5008 1379 5009 1431
rect 5061 1379 5062 1431
rect 5008 1353 5018 1379
rect 5052 1353 5062 1379
rect 5008 1341 5062 1353
rect 5108 1387 5162 1493
rect 5208 1527 5262 1539
rect 5208 1501 5218 1527
rect 5252 1501 5262 1527
rect 5208 1449 5209 1501
rect 5261 1449 5262 1501
rect 5208 1442 5262 1449
rect 5308 1527 5362 1633
rect 5408 1711 5462 1718
rect 5408 1659 5409 1711
rect 5461 1659 5462 1711
rect 5408 1633 5418 1659
rect 5452 1633 5462 1659
rect 5408 1621 5462 1633
rect 5508 1667 5562 1773
rect 5608 1807 5662 1819
rect 5608 1781 5618 1807
rect 5652 1781 5662 1807
rect 5608 1729 5609 1781
rect 5661 1729 5662 1781
rect 5608 1722 5662 1729
rect 5708 1807 5762 1913
rect 5808 1991 5862 1998
rect 5808 1939 5809 1991
rect 5861 1939 5862 1991
rect 5808 1913 5818 1939
rect 5852 1913 5862 1939
rect 5808 1901 5862 1913
rect 5908 1947 5962 2053
rect 6008 2087 6062 2099
rect 6008 2061 6018 2087
rect 6052 2061 6062 2087
rect 6008 2009 6009 2061
rect 6061 2009 6062 2061
rect 6008 2002 6062 2009
rect 6108 2087 6162 2193
rect 6208 2271 6262 2278
rect 6208 2219 6209 2271
rect 6261 2219 6262 2271
rect 6208 2193 6218 2219
rect 6252 2193 6262 2219
rect 6208 2181 6262 2193
rect 6308 2227 6362 2333
rect 6408 2367 6462 2379
rect 6408 2341 6418 2367
rect 6452 2341 6462 2367
rect 6408 2289 6409 2341
rect 6461 2289 6462 2341
rect 6408 2282 6462 2289
rect 6508 2367 6562 2563
rect 6608 2641 6662 2648
rect 6608 2589 6609 2641
rect 6661 2589 6662 2641
rect 6608 2563 6618 2589
rect 6652 2563 6662 2589
rect 6608 2551 6662 2563
rect 6708 2597 6762 2703
rect 6808 2737 6862 2749
rect 6808 2711 6818 2737
rect 6852 2711 6862 2737
rect 6808 2659 6809 2711
rect 6861 2659 6862 2711
rect 6808 2652 6862 2659
rect 6908 2737 6962 2843
rect 7008 2921 7062 2928
rect 7008 2869 7009 2921
rect 7061 2869 7062 2921
rect 7008 2843 7018 2869
rect 7052 2843 7062 2869
rect 7008 2831 7062 2843
rect 7108 2877 7162 2983
rect 7208 3017 7262 3029
rect 7208 2991 7218 3017
rect 7252 2991 7262 3017
rect 7208 2939 7209 2991
rect 7261 2939 7262 2991
rect 7208 2932 7262 2939
rect 7308 3017 7362 3123
rect 7408 3201 7462 3208
rect 7408 3149 7409 3201
rect 7461 3149 7462 3201
rect 7408 3123 7418 3149
rect 7452 3123 7462 3149
rect 7408 3111 7462 3123
rect 7508 3157 7562 3263
rect 7608 3297 7662 3309
rect 7608 3271 7618 3297
rect 7652 3271 7662 3297
rect 7608 3219 7609 3271
rect 7661 3219 7662 3271
rect 7608 3212 7662 3219
rect 7708 3297 7762 3403
rect 7808 3481 7862 3488
rect 7808 3429 7809 3481
rect 7861 3429 7862 3481
rect 7808 3403 7818 3429
rect 7852 3403 7862 3429
rect 7808 3391 7862 3403
rect 7908 3437 7962 3543
rect 8008 3577 8062 3589
rect 8008 3551 8018 3577
rect 8052 3551 8062 3577
rect 8008 3499 8009 3551
rect 8061 3499 8062 3551
rect 8008 3492 8062 3499
rect 8108 3577 8162 3773
rect 8208 3851 8262 3858
rect 8208 3799 8209 3851
rect 8261 3799 8262 3851
rect 8208 3773 8218 3799
rect 8252 3773 8262 3799
rect 8208 3761 8262 3773
rect 8308 3807 8362 3913
rect 8408 3947 8462 3959
rect 8408 3921 8418 3947
rect 8452 3921 8462 3947
rect 8408 3869 8409 3921
rect 8461 3869 8462 3921
rect 8408 3862 8462 3869
rect 8508 3947 8562 4053
rect 8608 4131 8662 4138
rect 8608 4079 8609 4131
rect 8661 4079 8662 4131
rect 8608 4053 8618 4079
rect 8652 4053 8662 4079
rect 8608 4041 8662 4053
rect 8708 4087 8762 4193
rect 8808 4227 8862 4239
rect 8808 4201 8818 4227
rect 8852 4201 8862 4227
rect 8808 4149 8809 4201
rect 8861 4149 8862 4201
rect 8808 4142 8862 4149
rect 8908 4227 8962 4333
rect 9008 4411 9062 4418
rect 9008 4359 9009 4411
rect 9061 4359 9062 4411
rect 9008 4333 9018 4359
rect 9052 4333 9062 4359
rect 9008 4321 9062 4333
rect 9108 4367 9162 4473
rect 9208 4507 9262 4519
rect 9208 4481 9218 4507
rect 9252 4481 9262 4507
rect 9208 4429 9209 4481
rect 9261 4429 9262 4481
rect 9208 4422 9262 4429
rect 9308 4507 9362 4613
rect 9408 4691 9462 4698
rect 9408 4639 9409 4691
rect 9461 4639 9462 4691
rect 9408 4613 9418 4639
rect 9452 4613 9462 4639
rect 9408 4601 9462 4613
rect 9508 4647 9562 4753
rect 9608 4787 9662 4799
rect 9608 4761 9618 4787
rect 9652 4761 9662 4787
rect 9608 4709 9609 4761
rect 9661 4709 9662 4761
rect 9608 4702 9662 4709
rect 9708 4787 9762 4960
rect 9802 4919 9868 4920
rect 9802 4867 9809 4919
rect 9861 4867 9868 4919
rect 9802 4866 9868 4867
rect 9708 4753 9718 4787
rect 9752 4753 9762 4787
rect 9508 4613 9518 4647
rect 9552 4613 9562 4647
rect 9308 4473 9318 4507
rect 9352 4473 9362 4507
rect 9108 4333 9118 4367
rect 9152 4333 9162 4367
rect 8908 4193 8918 4227
rect 8952 4193 8962 4227
rect 8708 4053 8718 4087
rect 8752 4053 8762 4087
rect 8508 3913 8518 3947
rect 8552 3913 8562 3947
rect 8308 3773 8318 3807
rect 8352 3773 8362 3807
rect 8202 3709 8268 3710
rect 8202 3657 8209 3709
rect 8261 3657 8268 3709
rect 8202 3656 8268 3657
rect 8108 3543 8118 3577
rect 8152 3543 8162 3577
rect 7908 3403 7918 3437
rect 7952 3403 7962 3437
rect 7708 3263 7718 3297
rect 7752 3263 7762 3297
rect 7508 3123 7518 3157
rect 7552 3123 7562 3157
rect 7308 2983 7318 3017
rect 7352 2983 7362 3017
rect 7108 2843 7118 2877
rect 7152 2843 7162 2877
rect 6908 2703 6918 2737
rect 6952 2703 6962 2737
rect 6708 2563 6718 2597
rect 6752 2563 6762 2597
rect 6602 2499 6668 2500
rect 6602 2447 6609 2499
rect 6661 2447 6668 2499
rect 6602 2446 6668 2447
rect 6508 2333 6518 2367
rect 6552 2333 6562 2367
rect 6308 2193 6318 2227
rect 6352 2193 6362 2227
rect 6108 2053 6118 2087
rect 6152 2053 6162 2087
rect 5908 1913 5918 1947
rect 5952 1913 5962 1947
rect 5708 1773 5718 1807
rect 5752 1773 5762 1807
rect 5508 1633 5518 1667
rect 5552 1633 5562 1667
rect 5308 1493 5318 1527
rect 5352 1493 5362 1527
rect 5108 1353 5118 1387
rect 5152 1353 5162 1387
rect 5002 1289 5068 1290
rect 5002 1237 5009 1289
rect 5061 1237 5068 1289
rect 5002 1236 5068 1237
rect 4908 1123 4918 1157
rect 4952 1123 4962 1157
rect 4708 983 4718 1017
rect 4752 983 4762 1017
rect 4508 843 4518 877
rect 4552 843 4562 877
rect 4308 703 4318 737
rect 4352 703 4362 737
rect 4108 563 4118 597
rect 4152 563 4162 597
rect 3908 423 3918 457
rect 3952 423 3962 457
rect 3708 283 3718 317
rect 3752 283 3762 317
rect 3508 143 3518 177
rect 3552 143 3562 177
rect 3402 79 3468 80
rect 3402 27 3409 79
rect 3461 27 3468 79
rect 3402 26 3468 27
rect 3308 -67 3309 -15
rect 3361 -67 3362 -15
rect 3308 -79 3318 -67
rect 3352 -79 3362 -67
rect 3108 -132 3162 -131
rect 3108 -143 3118 -132
rect 3152 -143 3162 -132
rect 3108 -195 3109 -143
rect 3161 -195 3162 -143
rect 3108 -210 3162 -195
rect 3212 -133 3258 -81
rect 3212 -167 3218 -133
rect 3252 -167 3258 -133
rect 3118 -291 3125 -239
rect 3177 -291 3184 -239
rect 3012 -397 3018 -363
rect 3052 -397 3058 -363
rect 3012 -435 3058 -397
rect 3012 -469 3018 -435
rect 3052 -469 3058 -435
rect 3012 -512 3058 -469
rect 3109 -326 3161 -320
rect 3109 -390 3118 -378
rect 3152 -390 3161 -378
rect 3109 -454 3118 -442
rect 3152 -454 3161 -442
rect 3109 -555 3161 -506
rect 3212 -363 3258 -167
rect 3308 -131 3309 -79
rect 3361 -131 3362 -79
rect 3408 -22 3462 26
rect 3408 -74 3409 -22
rect 3461 -74 3462 -22
rect 3408 -81 3462 -74
rect 3508 -15 3562 143
rect 3608 177 3662 189
rect 3608 151 3618 177
rect 3652 151 3662 177
rect 3608 99 3609 151
rect 3661 99 3662 151
rect 3608 92 3662 99
rect 3708 177 3762 283
rect 3808 361 3862 368
rect 3808 309 3809 361
rect 3861 309 3862 361
rect 3808 283 3818 309
rect 3852 283 3862 309
rect 3808 271 3862 283
rect 3908 317 3962 423
rect 4008 457 4062 469
rect 4008 431 4018 457
rect 4052 431 4062 457
rect 4008 379 4009 431
rect 4061 379 4062 431
rect 4008 372 4062 379
rect 4108 457 4162 563
rect 4208 641 4262 648
rect 4208 589 4209 641
rect 4261 589 4262 641
rect 4208 563 4218 589
rect 4252 563 4262 589
rect 4208 551 4262 563
rect 4308 597 4362 703
rect 4408 737 4462 749
rect 4408 711 4418 737
rect 4452 711 4462 737
rect 4408 659 4409 711
rect 4461 659 4462 711
rect 4408 652 4462 659
rect 4508 737 4562 843
rect 4608 921 4662 928
rect 4608 869 4609 921
rect 4661 869 4662 921
rect 4608 843 4618 869
rect 4652 843 4662 869
rect 4608 831 4662 843
rect 4708 877 4762 983
rect 4808 1017 4862 1029
rect 4808 991 4818 1017
rect 4852 991 4862 1017
rect 4808 939 4809 991
rect 4861 939 4862 991
rect 4808 932 4862 939
rect 4908 1017 4962 1123
rect 5008 1201 5062 1208
rect 5008 1149 5009 1201
rect 5061 1149 5062 1201
rect 5008 1123 5018 1149
rect 5052 1123 5062 1149
rect 5008 1111 5062 1123
rect 5108 1157 5162 1353
rect 5208 1387 5262 1399
rect 5208 1361 5218 1387
rect 5252 1361 5262 1387
rect 5208 1309 5209 1361
rect 5261 1309 5262 1361
rect 5208 1302 5262 1309
rect 5308 1387 5362 1493
rect 5408 1571 5462 1578
rect 5408 1519 5409 1571
rect 5461 1519 5462 1571
rect 5408 1493 5418 1519
rect 5452 1493 5462 1519
rect 5408 1481 5462 1493
rect 5508 1527 5562 1633
rect 5608 1667 5662 1679
rect 5608 1641 5618 1667
rect 5652 1641 5662 1667
rect 5608 1589 5609 1641
rect 5661 1589 5662 1641
rect 5608 1582 5662 1589
rect 5708 1667 5762 1773
rect 5808 1851 5862 1858
rect 5808 1799 5809 1851
rect 5861 1799 5862 1851
rect 5808 1773 5818 1799
rect 5852 1773 5862 1799
rect 5808 1761 5862 1773
rect 5908 1807 5962 1913
rect 6008 1947 6062 1959
rect 6008 1921 6018 1947
rect 6052 1921 6062 1947
rect 6008 1869 6009 1921
rect 6061 1869 6062 1921
rect 6008 1862 6062 1869
rect 6108 1947 6162 2053
rect 6208 2131 6262 2138
rect 6208 2079 6209 2131
rect 6261 2079 6262 2131
rect 6208 2053 6218 2079
rect 6252 2053 6262 2079
rect 6208 2041 6262 2053
rect 6308 2087 6362 2193
rect 6408 2227 6462 2239
rect 6408 2201 6418 2227
rect 6452 2201 6462 2227
rect 6408 2149 6409 2201
rect 6461 2149 6462 2201
rect 6408 2142 6462 2149
rect 6508 2227 6562 2333
rect 6608 2411 6662 2418
rect 6608 2359 6609 2411
rect 6661 2359 6662 2411
rect 6608 2333 6618 2359
rect 6652 2333 6662 2359
rect 6608 2321 6662 2333
rect 6708 2367 6762 2563
rect 6808 2597 6862 2609
rect 6808 2571 6818 2597
rect 6852 2571 6862 2597
rect 6808 2519 6809 2571
rect 6861 2519 6862 2571
rect 6808 2512 6862 2519
rect 6908 2597 6962 2703
rect 7008 2781 7062 2788
rect 7008 2729 7009 2781
rect 7061 2729 7062 2781
rect 7008 2703 7018 2729
rect 7052 2703 7062 2729
rect 7008 2691 7062 2703
rect 7108 2737 7162 2843
rect 7208 2877 7262 2889
rect 7208 2851 7218 2877
rect 7252 2851 7262 2877
rect 7208 2799 7209 2851
rect 7261 2799 7262 2851
rect 7208 2792 7262 2799
rect 7308 2877 7362 2983
rect 7408 3061 7462 3068
rect 7408 3009 7409 3061
rect 7461 3009 7462 3061
rect 7408 2983 7418 3009
rect 7452 2983 7462 3009
rect 7408 2971 7462 2983
rect 7508 3017 7562 3123
rect 7608 3157 7662 3169
rect 7608 3131 7618 3157
rect 7652 3131 7662 3157
rect 7608 3079 7609 3131
rect 7661 3079 7662 3131
rect 7608 3072 7662 3079
rect 7708 3157 7762 3263
rect 7808 3341 7862 3348
rect 7808 3289 7809 3341
rect 7861 3289 7862 3341
rect 7808 3263 7818 3289
rect 7852 3263 7862 3289
rect 7808 3251 7862 3263
rect 7908 3297 7962 3403
rect 8008 3437 8062 3449
rect 8008 3411 8018 3437
rect 8052 3411 8062 3437
rect 8008 3359 8009 3411
rect 8061 3359 8062 3411
rect 8008 3352 8062 3359
rect 8108 3437 8162 3543
rect 8208 3621 8262 3628
rect 8208 3569 8209 3621
rect 8261 3569 8262 3621
rect 8208 3543 8218 3569
rect 8252 3543 8262 3569
rect 8208 3531 8262 3543
rect 8308 3577 8362 3773
rect 8408 3807 8462 3819
rect 8408 3781 8418 3807
rect 8452 3781 8462 3807
rect 8408 3729 8409 3781
rect 8461 3729 8462 3781
rect 8408 3722 8462 3729
rect 8508 3807 8562 3913
rect 8608 3991 8662 3998
rect 8608 3939 8609 3991
rect 8661 3939 8662 3991
rect 8608 3913 8618 3939
rect 8652 3913 8662 3939
rect 8608 3901 8662 3913
rect 8708 3947 8762 4053
rect 8808 4087 8862 4099
rect 8808 4061 8818 4087
rect 8852 4061 8862 4087
rect 8808 4009 8809 4061
rect 8861 4009 8862 4061
rect 8808 4002 8862 4009
rect 8908 4087 8962 4193
rect 9008 4271 9062 4278
rect 9008 4219 9009 4271
rect 9061 4219 9062 4271
rect 9008 4193 9018 4219
rect 9052 4193 9062 4219
rect 9008 4181 9062 4193
rect 9108 4227 9162 4333
rect 9208 4367 9262 4379
rect 9208 4341 9218 4367
rect 9252 4341 9262 4367
rect 9208 4289 9209 4341
rect 9261 4289 9262 4341
rect 9208 4282 9262 4289
rect 9308 4367 9362 4473
rect 9408 4551 9462 4558
rect 9408 4499 9409 4551
rect 9461 4499 9462 4551
rect 9408 4473 9418 4499
rect 9452 4473 9462 4499
rect 9408 4461 9462 4473
rect 9508 4507 9562 4613
rect 9608 4647 9662 4659
rect 9608 4621 9618 4647
rect 9652 4621 9662 4647
rect 9608 4569 9609 4621
rect 9661 4569 9662 4621
rect 9608 4562 9662 4569
rect 9708 4647 9762 4753
rect 9808 4831 9862 4838
rect 9808 4779 9809 4831
rect 9861 4779 9862 4831
rect 9808 4753 9818 4779
rect 9852 4753 9862 4779
rect 9808 4741 9862 4753
rect 9908 4787 9962 4960
rect 10002 4903 10068 4904
rect 10002 4851 10009 4903
rect 10061 4851 10068 4903
rect 10002 4850 10068 4851
rect 9908 4753 9918 4787
rect 9952 4753 9962 4787
rect 9708 4613 9718 4647
rect 9752 4613 9762 4647
rect 9508 4473 9518 4507
rect 9552 4473 9562 4507
rect 9308 4333 9318 4367
rect 9352 4333 9362 4367
rect 9108 4193 9118 4227
rect 9152 4193 9162 4227
rect 8908 4053 8918 4087
rect 8952 4053 8962 4087
rect 8708 3913 8718 3947
rect 8752 3913 8762 3947
rect 8508 3773 8518 3807
rect 8552 3773 8562 3807
rect 8402 3693 8468 3694
rect 8402 3641 8409 3693
rect 8461 3641 8468 3693
rect 8402 3640 8468 3641
rect 8308 3543 8318 3577
rect 8352 3543 8362 3577
rect 8108 3403 8118 3437
rect 8152 3403 8162 3437
rect 7908 3263 7918 3297
rect 7952 3263 7962 3297
rect 7708 3123 7718 3157
rect 7752 3123 7762 3157
rect 7508 2983 7518 3017
rect 7552 2983 7562 3017
rect 7308 2843 7318 2877
rect 7352 2843 7362 2877
rect 7108 2703 7118 2737
rect 7152 2703 7162 2737
rect 6908 2563 6918 2597
rect 6952 2563 6962 2597
rect 6802 2483 6868 2484
rect 6802 2431 6809 2483
rect 6861 2431 6868 2483
rect 6802 2430 6868 2431
rect 6708 2333 6718 2367
rect 6752 2333 6762 2367
rect 6508 2193 6518 2227
rect 6552 2193 6562 2227
rect 6308 2053 6318 2087
rect 6352 2053 6362 2087
rect 6108 1913 6118 1947
rect 6152 1913 6162 1947
rect 5908 1773 5918 1807
rect 5952 1773 5962 1807
rect 5708 1633 5718 1667
rect 5752 1633 5762 1667
rect 5508 1493 5518 1527
rect 5552 1493 5562 1527
rect 5308 1353 5318 1387
rect 5352 1353 5362 1387
rect 5202 1273 5268 1274
rect 5202 1221 5209 1273
rect 5261 1221 5268 1273
rect 5202 1220 5268 1221
rect 5108 1123 5118 1157
rect 5152 1123 5162 1157
rect 4908 983 4918 1017
rect 4952 983 4962 1017
rect 4708 843 4718 877
rect 4752 843 4762 877
rect 4508 703 4518 737
rect 4552 703 4562 737
rect 4308 563 4318 597
rect 4352 563 4362 597
rect 4108 423 4118 457
rect 4152 423 4162 457
rect 3908 283 3918 317
rect 3952 283 3962 317
rect 3708 143 3718 177
rect 3752 143 3762 177
rect 3602 63 3668 64
rect 3602 11 3609 63
rect 3661 11 3668 63
rect 3602 10 3668 11
rect 3508 -67 3509 -15
rect 3561 -67 3562 -15
rect 3508 -79 3518 -67
rect 3552 -79 3562 -67
rect 3308 -132 3362 -131
rect 3308 -143 3318 -132
rect 3352 -143 3362 -132
rect 3308 -195 3309 -143
rect 3361 -195 3362 -143
rect 3308 -210 3362 -195
rect 3412 -133 3458 -81
rect 3412 -167 3418 -133
rect 3452 -167 3458 -133
rect 3318 -291 3325 -239
rect 3377 -291 3384 -239
rect 3212 -397 3218 -363
rect 3252 -397 3258 -363
rect 3212 -435 3258 -397
rect 3212 -469 3218 -435
rect 3252 -469 3258 -435
rect 3212 -512 3258 -469
rect 3309 -326 3361 -320
rect 3309 -390 3318 -378
rect 3352 -390 3361 -378
rect 3309 -454 3318 -442
rect 3352 -454 3361 -442
rect 3309 -512 3361 -506
rect 3412 -363 3458 -167
rect 3508 -131 3509 -79
rect 3561 -131 3562 -79
rect 3608 -22 3662 10
rect 3608 -74 3609 -22
rect 3661 -74 3662 -22
rect 3608 -81 3662 -74
rect 3708 -15 3762 143
rect 3808 221 3862 228
rect 3808 169 3809 221
rect 3861 169 3862 221
rect 3808 143 3818 169
rect 3852 143 3862 169
rect 3808 131 3862 143
rect 3908 177 3962 283
rect 4008 317 4062 329
rect 4008 291 4018 317
rect 4052 291 4062 317
rect 4008 239 4009 291
rect 4061 239 4062 291
rect 4008 232 4062 239
rect 4108 317 4162 423
rect 4208 501 4262 508
rect 4208 449 4209 501
rect 4261 449 4262 501
rect 4208 423 4218 449
rect 4252 423 4262 449
rect 4208 411 4262 423
rect 4308 457 4362 563
rect 4408 597 4462 609
rect 4408 571 4418 597
rect 4452 571 4462 597
rect 4408 519 4409 571
rect 4461 519 4462 571
rect 4408 512 4462 519
rect 4508 597 4562 703
rect 4608 781 4662 788
rect 4608 729 4609 781
rect 4661 729 4662 781
rect 4608 703 4618 729
rect 4652 703 4662 729
rect 4608 691 4662 703
rect 4708 737 4762 843
rect 4808 877 4862 889
rect 4808 851 4818 877
rect 4852 851 4862 877
rect 4808 799 4809 851
rect 4861 799 4862 851
rect 4808 792 4862 799
rect 4908 877 4962 983
rect 5008 1061 5062 1068
rect 5008 1009 5009 1061
rect 5061 1009 5062 1061
rect 5008 983 5018 1009
rect 5052 983 5062 1009
rect 5008 971 5062 983
rect 5108 1017 5162 1123
rect 5208 1157 5262 1169
rect 5208 1131 5218 1157
rect 5252 1131 5262 1157
rect 5208 1079 5209 1131
rect 5261 1079 5262 1131
rect 5208 1072 5262 1079
rect 5308 1157 5362 1353
rect 5408 1431 5462 1438
rect 5408 1379 5409 1431
rect 5461 1379 5462 1431
rect 5408 1353 5418 1379
rect 5452 1353 5462 1379
rect 5408 1341 5462 1353
rect 5508 1387 5562 1493
rect 5608 1527 5662 1539
rect 5608 1501 5618 1527
rect 5652 1501 5662 1527
rect 5608 1449 5609 1501
rect 5661 1449 5662 1501
rect 5608 1442 5662 1449
rect 5708 1527 5762 1633
rect 5808 1711 5862 1718
rect 5808 1659 5809 1711
rect 5861 1659 5862 1711
rect 5808 1633 5818 1659
rect 5852 1633 5862 1659
rect 5808 1621 5862 1633
rect 5908 1667 5962 1773
rect 6008 1807 6062 1819
rect 6008 1781 6018 1807
rect 6052 1781 6062 1807
rect 6008 1729 6009 1781
rect 6061 1729 6062 1781
rect 6008 1722 6062 1729
rect 6108 1807 6162 1913
rect 6208 1991 6262 1998
rect 6208 1939 6209 1991
rect 6261 1939 6262 1991
rect 6208 1913 6218 1939
rect 6252 1913 6262 1939
rect 6208 1901 6262 1913
rect 6308 1947 6362 2053
rect 6408 2087 6462 2099
rect 6408 2061 6418 2087
rect 6452 2061 6462 2087
rect 6408 2009 6409 2061
rect 6461 2009 6462 2061
rect 6408 2002 6462 2009
rect 6508 2087 6562 2193
rect 6608 2271 6662 2278
rect 6608 2219 6609 2271
rect 6661 2219 6662 2271
rect 6608 2193 6618 2219
rect 6652 2193 6662 2219
rect 6608 2181 6662 2193
rect 6708 2227 6762 2333
rect 6808 2367 6862 2379
rect 6808 2341 6818 2367
rect 6852 2341 6862 2367
rect 6808 2289 6809 2341
rect 6861 2289 6862 2341
rect 6808 2282 6862 2289
rect 6908 2367 6962 2563
rect 7008 2641 7062 2648
rect 7008 2589 7009 2641
rect 7061 2589 7062 2641
rect 7008 2563 7018 2589
rect 7052 2563 7062 2589
rect 7008 2551 7062 2563
rect 7108 2597 7162 2703
rect 7208 2737 7262 2749
rect 7208 2711 7218 2737
rect 7252 2711 7262 2737
rect 7208 2659 7209 2711
rect 7261 2659 7262 2711
rect 7208 2652 7262 2659
rect 7308 2737 7362 2843
rect 7408 2921 7462 2928
rect 7408 2869 7409 2921
rect 7461 2869 7462 2921
rect 7408 2843 7418 2869
rect 7452 2843 7462 2869
rect 7408 2831 7462 2843
rect 7508 2877 7562 2983
rect 7608 3017 7662 3029
rect 7608 2991 7618 3017
rect 7652 2991 7662 3017
rect 7608 2939 7609 2991
rect 7661 2939 7662 2991
rect 7608 2932 7662 2939
rect 7708 3017 7762 3123
rect 7808 3201 7862 3208
rect 7808 3149 7809 3201
rect 7861 3149 7862 3201
rect 7808 3123 7818 3149
rect 7852 3123 7862 3149
rect 7808 3111 7862 3123
rect 7908 3157 7962 3263
rect 8008 3297 8062 3309
rect 8008 3271 8018 3297
rect 8052 3271 8062 3297
rect 8008 3219 8009 3271
rect 8061 3219 8062 3271
rect 8008 3212 8062 3219
rect 8108 3297 8162 3403
rect 8208 3481 8262 3488
rect 8208 3429 8209 3481
rect 8261 3429 8262 3481
rect 8208 3403 8218 3429
rect 8252 3403 8262 3429
rect 8208 3391 8262 3403
rect 8308 3437 8362 3543
rect 8408 3577 8462 3589
rect 8408 3551 8418 3577
rect 8452 3551 8462 3577
rect 8408 3499 8409 3551
rect 8461 3499 8462 3551
rect 8408 3492 8462 3499
rect 8508 3577 8562 3773
rect 8608 3851 8662 3858
rect 8608 3799 8609 3851
rect 8661 3799 8662 3851
rect 8608 3773 8618 3799
rect 8652 3773 8662 3799
rect 8608 3761 8662 3773
rect 8708 3807 8762 3913
rect 8808 3947 8862 3959
rect 8808 3921 8818 3947
rect 8852 3921 8862 3947
rect 8808 3869 8809 3921
rect 8861 3869 8862 3921
rect 8808 3862 8862 3869
rect 8908 3947 8962 4053
rect 9008 4131 9062 4138
rect 9008 4079 9009 4131
rect 9061 4079 9062 4131
rect 9008 4053 9018 4079
rect 9052 4053 9062 4079
rect 9008 4041 9062 4053
rect 9108 4087 9162 4193
rect 9208 4227 9262 4239
rect 9208 4201 9218 4227
rect 9252 4201 9262 4227
rect 9208 4149 9209 4201
rect 9261 4149 9262 4201
rect 9208 4142 9262 4149
rect 9308 4227 9362 4333
rect 9408 4411 9462 4418
rect 9408 4359 9409 4411
rect 9461 4359 9462 4411
rect 9408 4333 9418 4359
rect 9452 4333 9462 4359
rect 9408 4321 9462 4333
rect 9508 4367 9562 4473
rect 9608 4507 9662 4519
rect 9608 4481 9618 4507
rect 9652 4481 9662 4507
rect 9608 4429 9609 4481
rect 9661 4429 9662 4481
rect 9608 4422 9662 4429
rect 9708 4507 9762 4613
rect 9808 4691 9862 4698
rect 9808 4639 9809 4691
rect 9861 4639 9862 4691
rect 9808 4613 9818 4639
rect 9852 4613 9862 4639
rect 9808 4601 9862 4613
rect 9908 4647 9962 4753
rect 10008 4787 10062 4799
rect 10008 4761 10018 4787
rect 10052 4761 10062 4787
rect 10008 4709 10009 4761
rect 10061 4709 10062 4761
rect 10008 4702 10062 4709
rect 10108 4787 10162 4960
rect 10202 4919 10268 4920
rect 10202 4867 10209 4919
rect 10261 4867 10268 4919
rect 10202 4866 10268 4867
rect 10108 4753 10118 4787
rect 10152 4753 10162 4787
rect 9908 4613 9918 4647
rect 9952 4613 9962 4647
rect 9708 4473 9718 4507
rect 9752 4473 9762 4507
rect 9508 4333 9518 4367
rect 9552 4333 9562 4367
rect 9308 4193 9318 4227
rect 9352 4193 9362 4227
rect 9108 4053 9118 4087
rect 9152 4053 9162 4087
rect 8908 3913 8918 3947
rect 8952 3913 8962 3947
rect 8708 3773 8718 3807
rect 8752 3773 8762 3807
rect 8602 3709 8668 3710
rect 8602 3657 8609 3709
rect 8661 3657 8668 3709
rect 8602 3656 8668 3657
rect 8508 3543 8518 3577
rect 8552 3543 8562 3577
rect 8308 3403 8318 3437
rect 8352 3403 8362 3437
rect 8108 3263 8118 3297
rect 8152 3263 8162 3297
rect 7908 3123 7918 3157
rect 7952 3123 7962 3157
rect 7708 2983 7718 3017
rect 7752 2983 7762 3017
rect 7508 2843 7518 2877
rect 7552 2843 7562 2877
rect 7308 2703 7318 2737
rect 7352 2703 7362 2737
rect 7108 2563 7118 2597
rect 7152 2563 7162 2597
rect 7002 2499 7068 2500
rect 7002 2447 7009 2499
rect 7061 2447 7068 2499
rect 7002 2446 7068 2447
rect 6908 2333 6918 2367
rect 6952 2333 6962 2367
rect 6708 2193 6718 2227
rect 6752 2193 6762 2227
rect 6508 2053 6518 2087
rect 6552 2053 6562 2087
rect 6308 1913 6318 1947
rect 6352 1913 6362 1947
rect 6108 1773 6118 1807
rect 6152 1773 6162 1807
rect 5908 1633 5918 1667
rect 5952 1633 5962 1667
rect 5708 1493 5718 1527
rect 5752 1493 5762 1527
rect 5508 1353 5518 1387
rect 5552 1353 5562 1387
rect 5402 1289 5468 1290
rect 5402 1237 5409 1289
rect 5461 1237 5468 1289
rect 5402 1236 5468 1237
rect 5308 1123 5318 1157
rect 5352 1123 5362 1157
rect 5108 983 5118 1017
rect 5152 983 5162 1017
rect 4908 843 4918 877
rect 4952 843 4962 877
rect 4708 703 4718 737
rect 4752 703 4762 737
rect 4508 563 4518 597
rect 4552 563 4562 597
rect 4308 423 4318 457
rect 4352 423 4362 457
rect 4108 283 4118 317
rect 4152 283 4162 317
rect 3908 143 3918 177
rect 3952 143 3962 177
rect 3802 79 3868 80
rect 3802 27 3809 79
rect 3861 27 3868 79
rect 3802 26 3868 27
rect 3708 -67 3709 -15
rect 3761 -67 3762 -15
rect 3708 -79 3718 -67
rect 3752 -79 3762 -67
rect 3508 -132 3562 -131
rect 3508 -143 3518 -132
rect 3552 -143 3562 -132
rect 3508 -195 3509 -143
rect 3561 -195 3562 -143
rect 3508 -210 3562 -195
rect 3612 -133 3658 -81
rect 3612 -167 3618 -133
rect 3652 -167 3658 -133
rect 3518 -291 3525 -239
rect 3577 -291 3584 -239
rect 3412 -397 3418 -363
rect 3452 -397 3458 -363
rect 3412 -435 3458 -397
rect 3412 -469 3418 -435
rect 3452 -469 3458 -435
rect 3412 -512 3458 -469
rect 3509 -326 3561 -320
rect 3509 -390 3518 -378
rect 3552 -390 3561 -378
rect 3509 -454 3518 -442
rect 3552 -454 3561 -442
rect 3509 -555 3561 -506
rect 3612 -363 3658 -167
rect 3708 -131 3709 -79
rect 3761 -131 3762 -79
rect 3808 -22 3862 26
rect 3808 -74 3809 -22
rect 3861 -74 3862 -22
rect 3808 -81 3862 -74
rect 3908 -15 3962 143
rect 4008 177 4062 189
rect 4008 151 4018 177
rect 4052 151 4062 177
rect 4008 99 4009 151
rect 4061 99 4062 151
rect 4008 92 4062 99
rect 4108 177 4162 283
rect 4208 361 4262 368
rect 4208 309 4209 361
rect 4261 309 4262 361
rect 4208 283 4218 309
rect 4252 283 4262 309
rect 4208 271 4262 283
rect 4308 317 4362 423
rect 4408 457 4462 469
rect 4408 431 4418 457
rect 4452 431 4462 457
rect 4408 379 4409 431
rect 4461 379 4462 431
rect 4408 372 4462 379
rect 4508 457 4562 563
rect 4608 641 4662 648
rect 4608 589 4609 641
rect 4661 589 4662 641
rect 4608 563 4618 589
rect 4652 563 4662 589
rect 4608 551 4662 563
rect 4708 597 4762 703
rect 4808 737 4862 749
rect 4808 711 4818 737
rect 4852 711 4862 737
rect 4808 659 4809 711
rect 4861 659 4862 711
rect 4808 652 4862 659
rect 4908 737 4962 843
rect 5008 921 5062 928
rect 5008 869 5009 921
rect 5061 869 5062 921
rect 5008 843 5018 869
rect 5052 843 5062 869
rect 5008 831 5062 843
rect 5108 877 5162 983
rect 5208 1017 5262 1029
rect 5208 991 5218 1017
rect 5252 991 5262 1017
rect 5208 939 5209 991
rect 5261 939 5262 991
rect 5208 932 5262 939
rect 5308 1017 5362 1123
rect 5408 1201 5462 1208
rect 5408 1149 5409 1201
rect 5461 1149 5462 1201
rect 5408 1123 5418 1149
rect 5452 1123 5462 1149
rect 5408 1111 5462 1123
rect 5508 1157 5562 1353
rect 5608 1387 5662 1399
rect 5608 1361 5618 1387
rect 5652 1361 5662 1387
rect 5608 1309 5609 1361
rect 5661 1309 5662 1361
rect 5608 1302 5662 1309
rect 5708 1387 5762 1493
rect 5808 1571 5862 1578
rect 5808 1519 5809 1571
rect 5861 1519 5862 1571
rect 5808 1493 5818 1519
rect 5852 1493 5862 1519
rect 5808 1481 5862 1493
rect 5908 1527 5962 1633
rect 6008 1667 6062 1679
rect 6008 1641 6018 1667
rect 6052 1641 6062 1667
rect 6008 1589 6009 1641
rect 6061 1589 6062 1641
rect 6008 1582 6062 1589
rect 6108 1667 6162 1773
rect 6208 1851 6262 1858
rect 6208 1799 6209 1851
rect 6261 1799 6262 1851
rect 6208 1773 6218 1799
rect 6252 1773 6262 1799
rect 6208 1761 6262 1773
rect 6308 1807 6362 1913
rect 6408 1947 6462 1959
rect 6408 1921 6418 1947
rect 6452 1921 6462 1947
rect 6408 1869 6409 1921
rect 6461 1869 6462 1921
rect 6408 1862 6462 1869
rect 6508 1947 6562 2053
rect 6608 2131 6662 2138
rect 6608 2079 6609 2131
rect 6661 2079 6662 2131
rect 6608 2053 6618 2079
rect 6652 2053 6662 2079
rect 6608 2041 6662 2053
rect 6708 2087 6762 2193
rect 6808 2227 6862 2239
rect 6808 2201 6818 2227
rect 6852 2201 6862 2227
rect 6808 2149 6809 2201
rect 6861 2149 6862 2201
rect 6808 2142 6862 2149
rect 6908 2227 6962 2333
rect 7008 2411 7062 2418
rect 7008 2359 7009 2411
rect 7061 2359 7062 2411
rect 7008 2333 7018 2359
rect 7052 2333 7062 2359
rect 7008 2321 7062 2333
rect 7108 2367 7162 2563
rect 7208 2597 7262 2609
rect 7208 2571 7218 2597
rect 7252 2571 7262 2597
rect 7208 2519 7209 2571
rect 7261 2519 7262 2571
rect 7208 2512 7262 2519
rect 7308 2597 7362 2703
rect 7408 2781 7462 2788
rect 7408 2729 7409 2781
rect 7461 2729 7462 2781
rect 7408 2703 7418 2729
rect 7452 2703 7462 2729
rect 7408 2691 7462 2703
rect 7508 2737 7562 2843
rect 7608 2877 7662 2889
rect 7608 2851 7618 2877
rect 7652 2851 7662 2877
rect 7608 2799 7609 2851
rect 7661 2799 7662 2851
rect 7608 2792 7662 2799
rect 7708 2877 7762 2983
rect 7808 3061 7862 3068
rect 7808 3009 7809 3061
rect 7861 3009 7862 3061
rect 7808 2983 7818 3009
rect 7852 2983 7862 3009
rect 7808 2971 7862 2983
rect 7908 3017 7962 3123
rect 8008 3157 8062 3169
rect 8008 3131 8018 3157
rect 8052 3131 8062 3157
rect 8008 3079 8009 3131
rect 8061 3079 8062 3131
rect 8008 3072 8062 3079
rect 8108 3157 8162 3263
rect 8208 3341 8262 3348
rect 8208 3289 8209 3341
rect 8261 3289 8262 3341
rect 8208 3263 8218 3289
rect 8252 3263 8262 3289
rect 8208 3251 8262 3263
rect 8308 3297 8362 3403
rect 8408 3437 8462 3449
rect 8408 3411 8418 3437
rect 8452 3411 8462 3437
rect 8408 3359 8409 3411
rect 8461 3359 8462 3411
rect 8408 3352 8462 3359
rect 8508 3437 8562 3543
rect 8608 3621 8662 3628
rect 8608 3569 8609 3621
rect 8661 3569 8662 3621
rect 8608 3543 8618 3569
rect 8652 3543 8662 3569
rect 8608 3531 8662 3543
rect 8708 3577 8762 3773
rect 8808 3807 8862 3819
rect 8808 3781 8818 3807
rect 8852 3781 8862 3807
rect 8808 3729 8809 3781
rect 8861 3729 8862 3781
rect 8808 3722 8862 3729
rect 8908 3807 8962 3913
rect 9008 3991 9062 3998
rect 9008 3939 9009 3991
rect 9061 3939 9062 3991
rect 9008 3913 9018 3939
rect 9052 3913 9062 3939
rect 9008 3901 9062 3913
rect 9108 3947 9162 4053
rect 9208 4087 9262 4099
rect 9208 4061 9218 4087
rect 9252 4061 9262 4087
rect 9208 4009 9209 4061
rect 9261 4009 9262 4061
rect 9208 4002 9262 4009
rect 9308 4087 9362 4193
rect 9408 4271 9462 4278
rect 9408 4219 9409 4271
rect 9461 4219 9462 4271
rect 9408 4193 9418 4219
rect 9452 4193 9462 4219
rect 9408 4181 9462 4193
rect 9508 4227 9562 4333
rect 9608 4367 9662 4379
rect 9608 4341 9618 4367
rect 9652 4341 9662 4367
rect 9608 4289 9609 4341
rect 9661 4289 9662 4341
rect 9608 4282 9662 4289
rect 9708 4367 9762 4473
rect 9808 4551 9862 4558
rect 9808 4499 9809 4551
rect 9861 4499 9862 4551
rect 9808 4473 9818 4499
rect 9852 4473 9862 4499
rect 9808 4461 9862 4473
rect 9908 4507 9962 4613
rect 10008 4647 10062 4659
rect 10008 4621 10018 4647
rect 10052 4621 10062 4647
rect 10008 4569 10009 4621
rect 10061 4569 10062 4621
rect 10008 4562 10062 4569
rect 10108 4647 10162 4753
rect 10208 4831 10262 4838
rect 10208 4779 10209 4831
rect 10261 4779 10262 4831
rect 10208 4753 10218 4779
rect 10252 4753 10262 4779
rect 10208 4741 10262 4753
rect 10308 4787 10362 4960
rect 10402 4903 10468 4904
rect 10402 4851 10409 4903
rect 10461 4851 10468 4903
rect 10402 4850 10468 4851
rect 10308 4753 10318 4787
rect 10352 4753 10362 4787
rect 10108 4613 10118 4647
rect 10152 4613 10162 4647
rect 9908 4473 9918 4507
rect 9952 4473 9962 4507
rect 9708 4333 9718 4367
rect 9752 4333 9762 4367
rect 9508 4193 9518 4227
rect 9552 4193 9562 4227
rect 9308 4053 9318 4087
rect 9352 4053 9362 4087
rect 9108 3913 9118 3947
rect 9152 3913 9162 3947
rect 8908 3773 8918 3807
rect 8952 3773 8962 3807
rect 8802 3693 8868 3694
rect 8802 3641 8809 3693
rect 8861 3641 8868 3693
rect 8802 3640 8868 3641
rect 8708 3543 8718 3577
rect 8752 3543 8762 3577
rect 8508 3403 8518 3437
rect 8552 3403 8562 3437
rect 8308 3263 8318 3297
rect 8352 3263 8362 3297
rect 8108 3123 8118 3157
rect 8152 3123 8162 3157
rect 7908 2983 7918 3017
rect 7952 2983 7962 3017
rect 7708 2843 7718 2877
rect 7752 2843 7762 2877
rect 7508 2703 7518 2737
rect 7552 2703 7562 2737
rect 7308 2563 7318 2597
rect 7352 2563 7362 2597
rect 7202 2483 7268 2484
rect 7202 2431 7209 2483
rect 7261 2431 7268 2483
rect 7202 2430 7268 2431
rect 7108 2333 7118 2367
rect 7152 2333 7162 2367
rect 6908 2193 6918 2227
rect 6952 2193 6962 2227
rect 6708 2053 6718 2087
rect 6752 2053 6762 2087
rect 6508 1913 6518 1947
rect 6552 1913 6562 1947
rect 6308 1773 6318 1807
rect 6352 1773 6362 1807
rect 6108 1633 6118 1667
rect 6152 1633 6162 1667
rect 5908 1493 5918 1527
rect 5952 1493 5962 1527
rect 5708 1353 5718 1387
rect 5752 1353 5762 1387
rect 5602 1273 5668 1274
rect 5602 1221 5609 1273
rect 5661 1221 5668 1273
rect 5602 1220 5668 1221
rect 5508 1123 5518 1157
rect 5552 1123 5562 1157
rect 5308 983 5318 1017
rect 5352 983 5362 1017
rect 5108 843 5118 877
rect 5152 843 5162 877
rect 4908 703 4918 737
rect 4952 703 4962 737
rect 4708 563 4718 597
rect 4752 563 4762 597
rect 4508 423 4518 457
rect 4552 423 4562 457
rect 4308 283 4318 317
rect 4352 283 4362 317
rect 4108 143 4118 177
rect 4152 143 4162 177
rect 4002 63 4068 64
rect 4002 11 4009 63
rect 4061 11 4068 63
rect 4002 10 4068 11
rect 3908 -67 3909 -15
rect 3961 -67 3962 -15
rect 3908 -79 3918 -67
rect 3952 -79 3962 -67
rect 3708 -132 3762 -131
rect 3708 -143 3718 -132
rect 3752 -143 3762 -132
rect 3708 -195 3709 -143
rect 3761 -195 3762 -143
rect 3708 -210 3762 -195
rect 3812 -133 3858 -81
rect 3812 -167 3818 -133
rect 3852 -167 3858 -133
rect 3718 -291 3725 -239
rect 3777 -291 3784 -239
rect 3612 -397 3618 -363
rect 3652 -397 3658 -363
rect 3612 -435 3658 -397
rect 3612 -469 3618 -435
rect 3652 -469 3658 -435
rect 3612 -512 3658 -469
rect 3709 -326 3761 -320
rect 3709 -390 3718 -378
rect 3752 -390 3761 -378
rect 3709 -454 3718 -442
rect 3752 -454 3761 -442
rect 3709 -512 3761 -506
rect 3812 -363 3858 -167
rect 3908 -131 3909 -79
rect 3961 -131 3962 -79
rect 4008 -22 4062 10
rect 4008 -74 4009 -22
rect 4061 -74 4062 -22
rect 4008 -81 4062 -74
rect 4108 -15 4162 143
rect 4208 221 4262 228
rect 4208 169 4209 221
rect 4261 169 4262 221
rect 4208 143 4218 169
rect 4252 143 4262 169
rect 4208 131 4262 143
rect 4308 177 4362 283
rect 4408 317 4462 329
rect 4408 291 4418 317
rect 4452 291 4462 317
rect 4408 239 4409 291
rect 4461 239 4462 291
rect 4408 232 4462 239
rect 4508 317 4562 423
rect 4608 501 4662 508
rect 4608 449 4609 501
rect 4661 449 4662 501
rect 4608 423 4618 449
rect 4652 423 4662 449
rect 4608 411 4662 423
rect 4708 457 4762 563
rect 4808 597 4862 609
rect 4808 571 4818 597
rect 4852 571 4862 597
rect 4808 519 4809 571
rect 4861 519 4862 571
rect 4808 512 4862 519
rect 4908 597 4962 703
rect 5008 781 5062 788
rect 5008 729 5009 781
rect 5061 729 5062 781
rect 5008 703 5018 729
rect 5052 703 5062 729
rect 5008 691 5062 703
rect 5108 737 5162 843
rect 5208 877 5262 889
rect 5208 851 5218 877
rect 5252 851 5262 877
rect 5208 799 5209 851
rect 5261 799 5262 851
rect 5208 792 5262 799
rect 5308 877 5362 983
rect 5408 1061 5462 1068
rect 5408 1009 5409 1061
rect 5461 1009 5462 1061
rect 5408 983 5418 1009
rect 5452 983 5462 1009
rect 5408 971 5462 983
rect 5508 1017 5562 1123
rect 5608 1157 5662 1169
rect 5608 1131 5618 1157
rect 5652 1131 5662 1157
rect 5608 1079 5609 1131
rect 5661 1079 5662 1131
rect 5608 1072 5662 1079
rect 5708 1157 5762 1353
rect 5808 1431 5862 1438
rect 5808 1379 5809 1431
rect 5861 1379 5862 1431
rect 5808 1353 5818 1379
rect 5852 1353 5862 1379
rect 5808 1341 5862 1353
rect 5908 1387 5962 1493
rect 6008 1527 6062 1539
rect 6008 1501 6018 1527
rect 6052 1501 6062 1527
rect 6008 1449 6009 1501
rect 6061 1449 6062 1501
rect 6008 1442 6062 1449
rect 6108 1527 6162 1633
rect 6208 1711 6262 1718
rect 6208 1659 6209 1711
rect 6261 1659 6262 1711
rect 6208 1633 6218 1659
rect 6252 1633 6262 1659
rect 6208 1621 6262 1633
rect 6308 1667 6362 1773
rect 6408 1807 6462 1819
rect 6408 1781 6418 1807
rect 6452 1781 6462 1807
rect 6408 1729 6409 1781
rect 6461 1729 6462 1781
rect 6408 1722 6462 1729
rect 6508 1807 6562 1913
rect 6608 1991 6662 1998
rect 6608 1939 6609 1991
rect 6661 1939 6662 1991
rect 6608 1913 6618 1939
rect 6652 1913 6662 1939
rect 6608 1901 6662 1913
rect 6708 1947 6762 2053
rect 6808 2087 6862 2099
rect 6808 2061 6818 2087
rect 6852 2061 6862 2087
rect 6808 2009 6809 2061
rect 6861 2009 6862 2061
rect 6808 2002 6862 2009
rect 6908 2087 6962 2193
rect 7008 2271 7062 2278
rect 7008 2219 7009 2271
rect 7061 2219 7062 2271
rect 7008 2193 7018 2219
rect 7052 2193 7062 2219
rect 7008 2181 7062 2193
rect 7108 2227 7162 2333
rect 7208 2367 7262 2379
rect 7208 2341 7218 2367
rect 7252 2341 7262 2367
rect 7208 2289 7209 2341
rect 7261 2289 7262 2341
rect 7208 2282 7262 2289
rect 7308 2367 7362 2563
rect 7408 2641 7462 2648
rect 7408 2589 7409 2641
rect 7461 2589 7462 2641
rect 7408 2563 7418 2589
rect 7452 2563 7462 2589
rect 7408 2551 7462 2563
rect 7508 2597 7562 2703
rect 7608 2737 7662 2749
rect 7608 2711 7618 2737
rect 7652 2711 7662 2737
rect 7608 2659 7609 2711
rect 7661 2659 7662 2711
rect 7608 2652 7662 2659
rect 7708 2737 7762 2843
rect 7808 2921 7862 2928
rect 7808 2869 7809 2921
rect 7861 2869 7862 2921
rect 7808 2843 7818 2869
rect 7852 2843 7862 2869
rect 7808 2831 7862 2843
rect 7908 2877 7962 2983
rect 8008 3017 8062 3029
rect 8008 2991 8018 3017
rect 8052 2991 8062 3017
rect 8008 2939 8009 2991
rect 8061 2939 8062 2991
rect 8008 2932 8062 2939
rect 8108 3017 8162 3123
rect 8208 3201 8262 3208
rect 8208 3149 8209 3201
rect 8261 3149 8262 3201
rect 8208 3123 8218 3149
rect 8252 3123 8262 3149
rect 8208 3111 8262 3123
rect 8308 3157 8362 3263
rect 8408 3297 8462 3309
rect 8408 3271 8418 3297
rect 8452 3271 8462 3297
rect 8408 3219 8409 3271
rect 8461 3219 8462 3271
rect 8408 3212 8462 3219
rect 8508 3297 8562 3403
rect 8608 3481 8662 3488
rect 8608 3429 8609 3481
rect 8661 3429 8662 3481
rect 8608 3403 8618 3429
rect 8652 3403 8662 3429
rect 8608 3391 8662 3403
rect 8708 3437 8762 3543
rect 8808 3577 8862 3589
rect 8808 3551 8818 3577
rect 8852 3551 8862 3577
rect 8808 3499 8809 3551
rect 8861 3499 8862 3551
rect 8808 3492 8862 3499
rect 8908 3577 8962 3773
rect 9008 3851 9062 3858
rect 9008 3799 9009 3851
rect 9061 3799 9062 3851
rect 9008 3773 9018 3799
rect 9052 3773 9062 3799
rect 9008 3761 9062 3773
rect 9108 3807 9162 3913
rect 9208 3947 9262 3959
rect 9208 3921 9218 3947
rect 9252 3921 9262 3947
rect 9208 3869 9209 3921
rect 9261 3869 9262 3921
rect 9208 3862 9262 3869
rect 9308 3947 9362 4053
rect 9408 4131 9462 4138
rect 9408 4079 9409 4131
rect 9461 4079 9462 4131
rect 9408 4053 9418 4079
rect 9452 4053 9462 4079
rect 9408 4041 9462 4053
rect 9508 4087 9562 4193
rect 9608 4227 9662 4239
rect 9608 4201 9618 4227
rect 9652 4201 9662 4227
rect 9608 4149 9609 4201
rect 9661 4149 9662 4201
rect 9608 4142 9662 4149
rect 9708 4227 9762 4333
rect 9808 4411 9862 4418
rect 9808 4359 9809 4411
rect 9861 4359 9862 4411
rect 9808 4333 9818 4359
rect 9852 4333 9862 4359
rect 9808 4321 9862 4333
rect 9908 4367 9962 4473
rect 10008 4507 10062 4519
rect 10008 4481 10018 4507
rect 10052 4481 10062 4507
rect 10008 4429 10009 4481
rect 10061 4429 10062 4481
rect 10008 4422 10062 4429
rect 10108 4507 10162 4613
rect 10208 4691 10262 4698
rect 10208 4639 10209 4691
rect 10261 4639 10262 4691
rect 10208 4613 10218 4639
rect 10252 4613 10262 4639
rect 10208 4601 10262 4613
rect 10308 4647 10362 4753
rect 10408 4787 10462 4799
rect 10408 4761 10418 4787
rect 10452 4761 10462 4787
rect 10408 4709 10409 4761
rect 10461 4709 10462 4761
rect 10408 4702 10462 4709
rect 10508 4787 10562 4960
rect 10602 4919 10668 4920
rect 10602 4867 10609 4919
rect 10661 4867 10668 4919
rect 10602 4866 10668 4867
rect 10508 4753 10518 4787
rect 10552 4753 10562 4787
rect 10308 4613 10318 4647
rect 10352 4613 10362 4647
rect 10108 4473 10118 4507
rect 10152 4473 10162 4507
rect 9908 4333 9918 4367
rect 9952 4333 9962 4367
rect 9708 4193 9718 4227
rect 9752 4193 9762 4227
rect 9508 4053 9518 4087
rect 9552 4053 9562 4087
rect 9308 3913 9318 3947
rect 9352 3913 9362 3947
rect 9108 3773 9118 3807
rect 9152 3773 9162 3807
rect 9002 3709 9068 3710
rect 9002 3657 9009 3709
rect 9061 3657 9068 3709
rect 9002 3656 9068 3657
rect 8908 3543 8918 3577
rect 8952 3543 8962 3577
rect 8708 3403 8718 3437
rect 8752 3403 8762 3437
rect 8508 3263 8518 3297
rect 8552 3263 8562 3297
rect 8308 3123 8318 3157
rect 8352 3123 8362 3157
rect 8108 2983 8118 3017
rect 8152 2983 8162 3017
rect 7908 2843 7918 2877
rect 7952 2843 7962 2877
rect 7708 2703 7718 2737
rect 7752 2703 7762 2737
rect 7508 2563 7518 2597
rect 7552 2563 7562 2597
rect 7402 2499 7468 2500
rect 7402 2447 7409 2499
rect 7461 2447 7468 2499
rect 7402 2446 7468 2447
rect 7308 2333 7318 2367
rect 7352 2333 7362 2367
rect 7108 2193 7118 2227
rect 7152 2193 7162 2227
rect 6908 2053 6918 2087
rect 6952 2053 6962 2087
rect 6708 1913 6718 1947
rect 6752 1913 6762 1947
rect 6508 1773 6518 1807
rect 6552 1773 6562 1807
rect 6308 1633 6318 1667
rect 6352 1633 6362 1667
rect 6108 1493 6118 1527
rect 6152 1493 6162 1527
rect 5908 1353 5918 1387
rect 5952 1353 5962 1387
rect 5802 1289 5868 1290
rect 5802 1237 5809 1289
rect 5861 1237 5868 1289
rect 5802 1236 5868 1237
rect 5708 1123 5718 1157
rect 5752 1123 5762 1157
rect 5508 983 5518 1017
rect 5552 983 5562 1017
rect 5308 843 5318 877
rect 5352 843 5362 877
rect 5108 703 5118 737
rect 5152 703 5162 737
rect 4908 563 4918 597
rect 4952 563 4962 597
rect 4708 423 4718 457
rect 4752 423 4762 457
rect 4508 283 4518 317
rect 4552 283 4562 317
rect 4308 143 4318 177
rect 4352 143 4362 177
rect 4202 79 4268 80
rect 4202 27 4209 79
rect 4261 27 4268 79
rect 4202 26 4268 27
rect 4108 -67 4109 -15
rect 4161 -67 4162 -15
rect 4108 -79 4118 -67
rect 4152 -79 4162 -67
rect 3908 -132 3962 -131
rect 3908 -143 3918 -132
rect 3952 -143 3962 -132
rect 3908 -195 3909 -143
rect 3961 -195 3962 -143
rect 3908 -210 3962 -195
rect 4012 -133 4058 -81
rect 4012 -167 4018 -133
rect 4052 -167 4058 -133
rect 3918 -291 3925 -239
rect 3977 -291 3984 -239
rect 3812 -397 3818 -363
rect 3852 -397 3858 -363
rect 3812 -435 3858 -397
rect 3812 -469 3818 -435
rect 3852 -469 3858 -435
rect 3812 -512 3858 -469
rect 3909 -326 3961 -320
rect 3909 -390 3918 -378
rect 3952 -390 3961 -378
rect 3909 -454 3918 -442
rect 3952 -454 3961 -442
rect 3909 -555 3961 -506
rect 4012 -363 4058 -167
rect 4108 -131 4109 -79
rect 4161 -131 4162 -79
rect 4208 -22 4262 26
rect 4208 -74 4209 -22
rect 4261 -74 4262 -22
rect 4208 -81 4262 -74
rect 4308 -15 4362 143
rect 4408 177 4462 189
rect 4408 151 4418 177
rect 4452 151 4462 177
rect 4408 99 4409 151
rect 4461 99 4462 151
rect 4408 92 4462 99
rect 4508 177 4562 283
rect 4608 361 4662 368
rect 4608 309 4609 361
rect 4661 309 4662 361
rect 4608 283 4618 309
rect 4652 283 4662 309
rect 4608 271 4662 283
rect 4708 317 4762 423
rect 4808 457 4862 469
rect 4808 431 4818 457
rect 4852 431 4862 457
rect 4808 379 4809 431
rect 4861 379 4862 431
rect 4808 372 4862 379
rect 4908 457 4962 563
rect 5008 641 5062 648
rect 5008 589 5009 641
rect 5061 589 5062 641
rect 5008 563 5018 589
rect 5052 563 5062 589
rect 5008 551 5062 563
rect 5108 597 5162 703
rect 5208 737 5262 749
rect 5208 711 5218 737
rect 5252 711 5262 737
rect 5208 659 5209 711
rect 5261 659 5262 711
rect 5208 652 5262 659
rect 5308 737 5362 843
rect 5408 921 5462 928
rect 5408 869 5409 921
rect 5461 869 5462 921
rect 5408 843 5418 869
rect 5452 843 5462 869
rect 5408 831 5462 843
rect 5508 877 5562 983
rect 5608 1017 5662 1029
rect 5608 991 5618 1017
rect 5652 991 5662 1017
rect 5608 939 5609 991
rect 5661 939 5662 991
rect 5608 932 5662 939
rect 5708 1017 5762 1123
rect 5808 1201 5862 1208
rect 5808 1149 5809 1201
rect 5861 1149 5862 1201
rect 5808 1123 5818 1149
rect 5852 1123 5862 1149
rect 5808 1111 5862 1123
rect 5908 1157 5962 1353
rect 6008 1387 6062 1399
rect 6008 1361 6018 1387
rect 6052 1361 6062 1387
rect 6008 1309 6009 1361
rect 6061 1309 6062 1361
rect 6008 1302 6062 1309
rect 6108 1387 6162 1493
rect 6208 1571 6262 1578
rect 6208 1519 6209 1571
rect 6261 1519 6262 1571
rect 6208 1493 6218 1519
rect 6252 1493 6262 1519
rect 6208 1481 6262 1493
rect 6308 1527 6362 1633
rect 6408 1667 6462 1679
rect 6408 1641 6418 1667
rect 6452 1641 6462 1667
rect 6408 1589 6409 1641
rect 6461 1589 6462 1641
rect 6408 1582 6462 1589
rect 6508 1667 6562 1773
rect 6608 1851 6662 1858
rect 6608 1799 6609 1851
rect 6661 1799 6662 1851
rect 6608 1773 6618 1799
rect 6652 1773 6662 1799
rect 6608 1761 6662 1773
rect 6708 1807 6762 1913
rect 6808 1947 6862 1959
rect 6808 1921 6818 1947
rect 6852 1921 6862 1947
rect 6808 1869 6809 1921
rect 6861 1869 6862 1921
rect 6808 1862 6862 1869
rect 6908 1947 6962 2053
rect 7008 2131 7062 2138
rect 7008 2079 7009 2131
rect 7061 2079 7062 2131
rect 7008 2053 7018 2079
rect 7052 2053 7062 2079
rect 7008 2041 7062 2053
rect 7108 2087 7162 2193
rect 7208 2227 7262 2239
rect 7208 2201 7218 2227
rect 7252 2201 7262 2227
rect 7208 2149 7209 2201
rect 7261 2149 7262 2201
rect 7208 2142 7262 2149
rect 7308 2227 7362 2333
rect 7408 2411 7462 2418
rect 7408 2359 7409 2411
rect 7461 2359 7462 2411
rect 7408 2333 7418 2359
rect 7452 2333 7462 2359
rect 7408 2321 7462 2333
rect 7508 2367 7562 2563
rect 7608 2597 7662 2609
rect 7608 2571 7618 2597
rect 7652 2571 7662 2597
rect 7608 2519 7609 2571
rect 7661 2519 7662 2571
rect 7608 2512 7662 2519
rect 7708 2597 7762 2703
rect 7808 2781 7862 2788
rect 7808 2729 7809 2781
rect 7861 2729 7862 2781
rect 7808 2703 7818 2729
rect 7852 2703 7862 2729
rect 7808 2691 7862 2703
rect 7908 2737 7962 2843
rect 8008 2877 8062 2889
rect 8008 2851 8018 2877
rect 8052 2851 8062 2877
rect 8008 2799 8009 2851
rect 8061 2799 8062 2851
rect 8008 2792 8062 2799
rect 8108 2877 8162 2983
rect 8208 3061 8262 3068
rect 8208 3009 8209 3061
rect 8261 3009 8262 3061
rect 8208 2983 8218 3009
rect 8252 2983 8262 3009
rect 8208 2971 8262 2983
rect 8308 3017 8362 3123
rect 8408 3157 8462 3169
rect 8408 3131 8418 3157
rect 8452 3131 8462 3157
rect 8408 3079 8409 3131
rect 8461 3079 8462 3131
rect 8408 3072 8462 3079
rect 8508 3157 8562 3263
rect 8608 3341 8662 3348
rect 8608 3289 8609 3341
rect 8661 3289 8662 3341
rect 8608 3263 8618 3289
rect 8652 3263 8662 3289
rect 8608 3251 8662 3263
rect 8708 3297 8762 3403
rect 8808 3437 8862 3449
rect 8808 3411 8818 3437
rect 8852 3411 8862 3437
rect 8808 3359 8809 3411
rect 8861 3359 8862 3411
rect 8808 3352 8862 3359
rect 8908 3437 8962 3543
rect 9008 3621 9062 3628
rect 9008 3569 9009 3621
rect 9061 3569 9062 3621
rect 9008 3543 9018 3569
rect 9052 3543 9062 3569
rect 9008 3531 9062 3543
rect 9108 3577 9162 3773
rect 9208 3807 9262 3819
rect 9208 3781 9218 3807
rect 9252 3781 9262 3807
rect 9208 3729 9209 3781
rect 9261 3729 9262 3781
rect 9208 3722 9262 3729
rect 9308 3807 9362 3913
rect 9408 3991 9462 3998
rect 9408 3939 9409 3991
rect 9461 3939 9462 3991
rect 9408 3913 9418 3939
rect 9452 3913 9462 3939
rect 9408 3901 9462 3913
rect 9508 3947 9562 4053
rect 9608 4087 9662 4099
rect 9608 4061 9618 4087
rect 9652 4061 9662 4087
rect 9608 4009 9609 4061
rect 9661 4009 9662 4061
rect 9608 4002 9662 4009
rect 9708 4087 9762 4193
rect 9808 4271 9862 4278
rect 9808 4219 9809 4271
rect 9861 4219 9862 4271
rect 9808 4193 9818 4219
rect 9852 4193 9862 4219
rect 9808 4181 9862 4193
rect 9908 4227 9962 4333
rect 10008 4367 10062 4379
rect 10008 4341 10018 4367
rect 10052 4341 10062 4367
rect 10008 4289 10009 4341
rect 10061 4289 10062 4341
rect 10008 4282 10062 4289
rect 10108 4367 10162 4473
rect 10208 4551 10262 4558
rect 10208 4499 10209 4551
rect 10261 4499 10262 4551
rect 10208 4473 10218 4499
rect 10252 4473 10262 4499
rect 10208 4461 10262 4473
rect 10308 4507 10362 4613
rect 10408 4647 10462 4659
rect 10408 4621 10418 4647
rect 10452 4621 10462 4647
rect 10408 4569 10409 4621
rect 10461 4569 10462 4621
rect 10408 4562 10462 4569
rect 10508 4647 10562 4753
rect 10608 4831 10662 4838
rect 10608 4779 10609 4831
rect 10661 4779 10662 4831
rect 10608 4753 10618 4779
rect 10652 4753 10662 4779
rect 10608 4741 10662 4753
rect 10708 4787 10762 4960
rect 10802 4903 10868 4904
rect 10802 4851 10809 4903
rect 10861 4851 10868 4903
rect 10802 4850 10868 4851
rect 10708 4753 10718 4787
rect 10752 4753 10762 4787
rect 10508 4613 10518 4647
rect 10552 4613 10562 4647
rect 10308 4473 10318 4507
rect 10352 4473 10362 4507
rect 10108 4333 10118 4367
rect 10152 4333 10162 4367
rect 9908 4193 9918 4227
rect 9952 4193 9962 4227
rect 9708 4053 9718 4087
rect 9752 4053 9762 4087
rect 9508 3913 9518 3947
rect 9552 3913 9562 3947
rect 9308 3773 9318 3807
rect 9352 3773 9362 3807
rect 9202 3693 9268 3694
rect 9202 3641 9209 3693
rect 9261 3641 9268 3693
rect 9202 3640 9268 3641
rect 9108 3543 9118 3577
rect 9152 3543 9162 3577
rect 8908 3403 8918 3437
rect 8952 3403 8962 3437
rect 8708 3263 8718 3297
rect 8752 3263 8762 3297
rect 8508 3123 8518 3157
rect 8552 3123 8562 3157
rect 8308 2983 8318 3017
rect 8352 2983 8362 3017
rect 8108 2843 8118 2877
rect 8152 2843 8162 2877
rect 7908 2703 7918 2737
rect 7952 2703 7962 2737
rect 7708 2563 7718 2597
rect 7752 2563 7762 2597
rect 7602 2483 7668 2484
rect 7602 2431 7609 2483
rect 7661 2431 7668 2483
rect 7602 2430 7668 2431
rect 7508 2333 7518 2367
rect 7552 2333 7562 2367
rect 7308 2193 7318 2227
rect 7352 2193 7362 2227
rect 7108 2053 7118 2087
rect 7152 2053 7162 2087
rect 6908 1913 6918 1947
rect 6952 1913 6962 1947
rect 6708 1773 6718 1807
rect 6752 1773 6762 1807
rect 6508 1633 6518 1667
rect 6552 1633 6562 1667
rect 6308 1493 6318 1527
rect 6352 1493 6362 1527
rect 6108 1353 6118 1387
rect 6152 1353 6162 1387
rect 6002 1273 6068 1274
rect 6002 1221 6009 1273
rect 6061 1221 6068 1273
rect 6002 1220 6068 1221
rect 5908 1123 5918 1157
rect 5952 1123 5962 1157
rect 5708 983 5718 1017
rect 5752 983 5762 1017
rect 5508 843 5518 877
rect 5552 843 5562 877
rect 5308 703 5318 737
rect 5352 703 5362 737
rect 5108 563 5118 597
rect 5152 563 5162 597
rect 4908 423 4918 457
rect 4952 423 4962 457
rect 4708 283 4718 317
rect 4752 283 4762 317
rect 4508 143 4518 177
rect 4552 143 4562 177
rect 4402 63 4468 64
rect 4402 11 4409 63
rect 4461 11 4468 63
rect 4402 10 4468 11
rect 4308 -67 4309 -15
rect 4361 -67 4362 -15
rect 4308 -79 4318 -67
rect 4352 -79 4362 -67
rect 4108 -132 4162 -131
rect 4108 -143 4118 -132
rect 4152 -143 4162 -132
rect 4108 -195 4109 -143
rect 4161 -195 4162 -143
rect 4108 -210 4162 -195
rect 4212 -133 4258 -81
rect 4212 -167 4218 -133
rect 4252 -167 4258 -133
rect 4118 -291 4125 -239
rect 4177 -291 4184 -239
rect 4012 -397 4018 -363
rect 4052 -397 4058 -363
rect 4012 -435 4058 -397
rect 4012 -469 4018 -435
rect 4052 -469 4058 -435
rect 4012 -512 4058 -469
rect 4109 -326 4161 -320
rect 4109 -390 4118 -378
rect 4152 -390 4161 -378
rect 4109 -454 4118 -442
rect 4152 -454 4161 -442
rect 4109 -512 4161 -506
rect 4212 -363 4258 -167
rect 4308 -131 4309 -79
rect 4361 -131 4362 -79
rect 4408 -22 4462 10
rect 4408 -74 4409 -22
rect 4461 -74 4462 -22
rect 4408 -81 4462 -74
rect 4508 -15 4562 143
rect 4608 221 4662 228
rect 4608 169 4609 221
rect 4661 169 4662 221
rect 4608 143 4618 169
rect 4652 143 4662 169
rect 4608 131 4662 143
rect 4708 177 4762 283
rect 4808 317 4862 329
rect 4808 291 4818 317
rect 4852 291 4862 317
rect 4808 239 4809 291
rect 4861 239 4862 291
rect 4808 232 4862 239
rect 4908 317 4962 423
rect 5008 501 5062 508
rect 5008 449 5009 501
rect 5061 449 5062 501
rect 5008 423 5018 449
rect 5052 423 5062 449
rect 5008 411 5062 423
rect 5108 457 5162 563
rect 5208 597 5262 609
rect 5208 571 5218 597
rect 5252 571 5262 597
rect 5208 519 5209 571
rect 5261 519 5262 571
rect 5208 512 5262 519
rect 5308 597 5362 703
rect 5408 781 5462 788
rect 5408 729 5409 781
rect 5461 729 5462 781
rect 5408 703 5418 729
rect 5452 703 5462 729
rect 5408 691 5462 703
rect 5508 737 5562 843
rect 5608 877 5662 889
rect 5608 851 5618 877
rect 5652 851 5662 877
rect 5608 799 5609 851
rect 5661 799 5662 851
rect 5608 792 5662 799
rect 5708 877 5762 983
rect 5808 1061 5862 1068
rect 5808 1009 5809 1061
rect 5861 1009 5862 1061
rect 5808 983 5818 1009
rect 5852 983 5862 1009
rect 5808 971 5862 983
rect 5908 1017 5962 1123
rect 6008 1157 6062 1169
rect 6008 1131 6018 1157
rect 6052 1131 6062 1157
rect 6008 1079 6009 1131
rect 6061 1079 6062 1131
rect 6008 1072 6062 1079
rect 6108 1157 6162 1353
rect 6208 1431 6262 1438
rect 6208 1379 6209 1431
rect 6261 1379 6262 1431
rect 6208 1353 6218 1379
rect 6252 1353 6262 1379
rect 6208 1341 6262 1353
rect 6308 1387 6362 1493
rect 6408 1527 6462 1539
rect 6408 1501 6418 1527
rect 6452 1501 6462 1527
rect 6408 1449 6409 1501
rect 6461 1449 6462 1501
rect 6408 1442 6462 1449
rect 6508 1527 6562 1633
rect 6608 1711 6662 1718
rect 6608 1659 6609 1711
rect 6661 1659 6662 1711
rect 6608 1633 6618 1659
rect 6652 1633 6662 1659
rect 6608 1621 6662 1633
rect 6708 1667 6762 1773
rect 6808 1807 6862 1819
rect 6808 1781 6818 1807
rect 6852 1781 6862 1807
rect 6808 1729 6809 1781
rect 6861 1729 6862 1781
rect 6808 1722 6862 1729
rect 6908 1807 6962 1913
rect 7008 1991 7062 1998
rect 7008 1939 7009 1991
rect 7061 1939 7062 1991
rect 7008 1913 7018 1939
rect 7052 1913 7062 1939
rect 7008 1901 7062 1913
rect 7108 1947 7162 2053
rect 7208 2087 7262 2099
rect 7208 2061 7218 2087
rect 7252 2061 7262 2087
rect 7208 2009 7209 2061
rect 7261 2009 7262 2061
rect 7208 2002 7262 2009
rect 7308 2087 7362 2193
rect 7408 2271 7462 2278
rect 7408 2219 7409 2271
rect 7461 2219 7462 2271
rect 7408 2193 7418 2219
rect 7452 2193 7462 2219
rect 7408 2181 7462 2193
rect 7508 2227 7562 2333
rect 7608 2367 7662 2379
rect 7608 2341 7618 2367
rect 7652 2341 7662 2367
rect 7608 2289 7609 2341
rect 7661 2289 7662 2341
rect 7608 2282 7662 2289
rect 7708 2367 7762 2563
rect 7808 2641 7862 2648
rect 7808 2589 7809 2641
rect 7861 2589 7862 2641
rect 7808 2563 7818 2589
rect 7852 2563 7862 2589
rect 7808 2551 7862 2563
rect 7908 2597 7962 2703
rect 8008 2737 8062 2749
rect 8008 2711 8018 2737
rect 8052 2711 8062 2737
rect 8008 2659 8009 2711
rect 8061 2659 8062 2711
rect 8008 2652 8062 2659
rect 8108 2737 8162 2843
rect 8208 2921 8262 2928
rect 8208 2869 8209 2921
rect 8261 2869 8262 2921
rect 8208 2843 8218 2869
rect 8252 2843 8262 2869
rect 8208 2831 8262 2843
rect 8308 2877 8362 2983
rect 8408 3017 8462 3029
rect 8408 2991 8418 3017
rect 8452 2991 8462 3017
rect 8408 2939 8409 2991
rect 8461 2939 8462 2991
rect 8408 2932 8462 2939
rect 8508 3017 8562 3123
rect 8608 3201 8662 3208
rect 8608 3149 8609 3201
rect 8661 3149 8662 3201
rect 8608 3123 8618 3149
rect 8652 3123 8662 3149
rect 8608 3111 8662 3123
rect 8708 3157 8762 3263
rect 8808 3297 8862 3309
rect 8808 3271 8818 3297
rect 8852 3271 8862 3297
rect 8808 3219 8809 3271
rect 8861 3219 8862 3271
rect 8808 3212 8862 3219
rect 8908 3297 8962 3403
rect 9008 3481 9062 3488
rect 9008 3429 9009 3481
rect 9061 3429 9062 3481
rect 9008 3403 9018 3429
rect 9052 3403 9062 3429
rect 9008 3391 9062 3403
rect 9108 3437 9162 3543
rect 9208 3577 9262 3589
rect 9208 3551 9218 3577
rect 9252 3551 9262 3577
rect 9208 3499 9209 3551
rect 9261 3499 9262 3551
rect 9208 3492 9262 3499
rect 9308 3577 9362 3773
rect 9408 3851 9462 3858
rect 9408 3799 9409 3851
rect 9461 3799 9462 3851
rect 9408 3773 9418 3799
rect 9452 3773 9462 3799
rect 9408 3761 9462 3773
rect 9508 3807 9562 3913
rect 9608 3947 9662 3959
rect 9608 3921 9618 3947
rect 9652 3921 9662 3947
rect 9608 3869 9609 3921
rect 9661 3869 9662 3921
rect 9608 3862 9662 3869
rect 9708 3947 9762 4053
rect 9808 4131 9862 4138
rect 9808 4079 9809 4131
rect 9861 4079 9862 4131
rect 9808 4053 9818 4079
rect 9852 4053 9862 4079
rect 9808 4041 9862 4053
rect 9908 4087 9962 4193
rect 10008 4227 10062 4239
rect 10008 4201 10018 4227
rect 10052 4201 10062 4227
rect 10008 4149 10009 4201
rect 10061 4149 10062 4201
rect 10008 4142 10062 4149
rect 10108 4227 10162 4333
rect 10208 4411 10262 4418
rect 10208 4359 10209 4411
rect 10261 4359 10262 4411
rect 10208 4333 10218 4359
rect 10252 4333 10262 4359
rect 10208 4321 10262 4333
rect 10308 4367 10362 4473
rect 10408 4507 10462 4519
rect 10408 4481 10418 4507
rect 10452 4481 10462 4507
rect 10408 4429 10409 4481
rect 10461 4429 10462 4481
rect 10408 4422 10462 4429
rect 10508 4507 10562 4613
rect 10608 4691 10662 4698
rect 10608 4639 10609 4691
rect 10661 4639 10662 4691
rect 10608 4613 10618 4639
rect 10652 4613 10662 4639
rect 10608 4601 10662 4613
rect 10708 4647 10762 4753
rect 10808 4787 10862 4799
rect 10808 4761 10818 4787
rect 10852 4761 10862 4787
rect 10808 4709 10809 4761
rect 10861 4709 10862 4761
rect 10808 4702 10862 4709
rect 10908 4787 10962 4960
rect 11002 4919 11068 4920
rect 11002 4867 11009 4919
rect 11061 4867 11068 4919
rect 11002 4866 11068 4867
rect 10908 4753 10918 4787
rect 10952 4753 10962 4787
rect 10708 4613 10718 4647
rect 10752 4613 10762 4647
rect 10508 4473 10518 4507
rect 10552 4473 10562 4507
rect 10308 4333 10318 4367
rect 10352 4333 10362 4367
rect 10108 4193 10118 4227
rect 10152 4193 10162 4227
rect 9908 4053 9918 4087
rect 9952 4053 9962 4087
rect 9708 3913 9718 3947
rect 9752 3913 9762 3947
rect 9508 3773 9518 3807
rect 9552 3773 9562 3807
rect 9402 3709 9468 3710
rect 9402 3657 9409 3709
rect 9461 3657 9468 3709
rect 9402 3656 9468 3657
rect 9308 3543 9318 3577
rect 9352 3543 9362 3577
rect 9108 3403 9118 3437
rect 9152 3403 9162 3437
rect 8908 3263 8918 3297
rect 8952 3263 8962 3297
rect 8708 3123 8718 3157
rect 8752 3123 8762 3157
rect 8508 2983 8518 3017
rect 8552 2983 8562 3017
rect 8308 2843 8318 2877
rect 8352 2843 8362 2877
rect 8108 2703 8118 2737
rect 8152 2703 8162 2737
rect 7908 2563 7918 2597
rect 7952 2563 7962 2597
rect 7802 2499 7868 2500
rect 7802 2447 7809 2499
rect 7861 2447 7868 2499
rect 7802 2446 7868 2447
rect 7708 2333 7718 2367
rect 7752 2333 7762 2367
rect 7508 2193 7518 2227
rect 7552 2193 7562 2227
rect 7308 2053 7318 2087
rect 7352 2053 7362 2087
rect 7108 1913 7118 1947
rect 7152 1913 7162 1947
rect 6908 1773 6918 1807
rect 6952 1773 6962 1807
rect 6708 1633 6718 1667
rect 6752 1633 6762 1667
rect 6508 1493 6518 1527
rect 6552 1493 6562 1527
rect 6308 1353 6318 1387
rect 6352 1353 6362 1387
rect 6202 1289 6268 1290
rect 6202 1237 6209 1289
rect 6261 1237 6268 1289
rect 6202 1236 6268 1237
rect 6108 1123 6118 1157
rect 6152 1123 6162 1157
rect 5908 983 5918 1017
rect 5952 983 5962 1017
rect 5708 843 5718 877
rect 5752 843 5762 877
rect 5508 703 5518 737
rect 5552 703 5562 737
rect 5308 563 5318 597
rect 5352 563 5362 597
rect 5108 423 5118 457
rect 5152 423 5162 457
rect 4908 283 4918 317
rect 4952 283 4962 317
rect 4708 143 4718 177
rect 4752 143 4762 177
rect 4602 79 4668 80
rect 4602 27 4609 79
rect 4661 27 4668 79
rect 4602 26 4668 27
rect 4508 -67 4509 -15
rect 4561 -67 4562 -15
rect 4508 -79 4518 -67
rect 4552 -79 4562 -67
rect 4308 -132 4362 -131
rect 4308 -143 4318 -132
rect 4352 -143 4362 -132
rect 4308 -195 4309 -143
rect 4361 -195 4362 -143
rect 4308 -210 4362 -195
rect 4412 -133 4458 -81
rect 4412 -167 4418 -133
rect 4452 -167 4458 -133
rect 4318 -291 4325 -239
rect 4377 -291 4384 -239
rect 4212 -397 4218 -363
rect 4252 -397 4258 -363
rect 4212 -435 4258 -397
rect 4212 -469 4218 -435
rect 4252 -469 4258 -435
rect 4212 -512 4258 -469
rect 4309 -326 4361 -320
rect 4309 -390 4318 -378
rect 4352 -390 4361 -378
rect 4309 -454 4318 -442
rect 4352 -454 4361 -442
rect 4309 -555 4361 -506
rect 4412 -363 4458 -167
rect 4508 -131 4509 -79
rect 4561 -131 4562 -79
rect 4608 -22 4662 26
rect 4608 -74 4609 -22
rect 4661 -74 4662 -22
rect 4608 -81 4662 -74
rect 4708 -15 4762 143
rect 4808 177 4862 189
rect 4808 151 4818 177
rect 4852 151 4862 177
rect 4808 99 4809 151
rect 4861 99 4862 151
rect 4808 92 4862 99
rect 4908 177 4962 283
rect 5008 361 5062 368
rect 5008 309 5009 361
rect 5061 309 5062 361
rect 5008 283 5018 309
rect 5052 283 5062 309
rect 5008 271 5062 283
rect 5108 317 5162 423
rect 5208 457 5262 469
rect 5208 431 5218 457
rect 5252 431 5262 457
rect 5208 379 5209 431
rect 5261 379 5262 431
rect 5208 372 5262 379
rect 5308 457 5362 563
rect 5408 641 5462 648
rect 5408 589 5409 641
rect 5461 589 5462 641
rect 5408 563 5418 589
rect 5452 563 5462 589
rect 5408 551 5462 563
rect 5508 597 5562 703
rect 5608 737 5662 749
rect 5608 711 5618 737
rect 5652 711 5662 737
rect 5608 659 5609 711
rect 5661 659 5662 711
rect 5608 652 5662 659
rect 5708 737 5762 843
rect 5808 921 5862 928
rect 5808 869 5809 921
rect 5861 869 5862 921
rect 5808 843 5818 869
rect 5852 843 5862 869
rect 5808 831 5862 843
rect 5908 877 5962 983
rect 6008 1017 6062 1029
rect 6008 991 6018 1017
rect 6052 991 6062 1017
rect 6008 939 6009 991
rect 6061 939 6062 991
rect 6008 932 6062 939
rect 6108 1017 6162 1123
rect 6208 1201 6262 1208
rect 6208 1149 6209 1201
rect 6261 1149 6262 1201
rect 6208 1123 6218 1149
rect 6252 1123 6262 1149
rect 6208 1111 6262 1123
rect 6308 1157 6362 1353
rect 6408 1387 6462 1399
rect 6408 1361 6418 1387
rect 6452 1361 6462 1387
rect 6408 1309 6409 1361
rect 6461 1309 6462 1361
rect 6408 1302 6462 1309
rect 6508 1387 6562 1493
rect 6608 1571 6662 1578
rect 6608 1519 6609 1571
rect 6661 1519 6662 1571
rect 6608 1493 6618 1519
rect 6652 1493 6662 1519
rect 6608 1481 6662 1493
rect 6708 1527 6762 1633
rect 6808 1667 6862 1679
rect 6808 1641 6818 1667
rect 6852 1641 6862 1667
rect 6808 1589 6809 1641
rect 6861 1589 6862 1641
rect 6808 1582 6862 1589
rect 6908 1667 6962 1773
rect 7008 1851 7062 1858
rect 7008 1799 7009 1851
rect 7061 1799 7062 1851
rect 7008 1773 7018 1799
rect 7052 1773 7062 1799
rect 7008 1761 7062 1773
rect 7108 1807 7162 1913
rect 7208 1947 7262 1959
rect 7208 1921 7218 1947
rect 7252 1921 7262 1947
rect 7208 1869 7209 1921
rect 7261 1869 7262 1921
rect 7208 1862 7262 1869
rect 7308 1947 7362 2053
rect 7408 2131 7462 2138
rect 7408 2079 7409 2131
rect 7461 2079 7462 2131
rect 7408 2053 7418 2079
rect 7452 2053 7462 2079
rect 7408 2041 7462 2053
rect 7508 2087 7562 2193
rect 7608 2227 7662 2239
rect 7608 2201 7618 2227
rect 7652 2201 7662 2227
rect 7608 2149 7609 2201
rect 7661 2149 7662 2201
rect 7608 2142 7662 2149
rect 7708 2227 7762 2333
rect 7808 2411 7862 2418
rect 7808 2359 7809 2411
rect 7861 2359 7862 2411
rect 7808 2333 7818 2359
rect 7852 2333 7862 2359
rect 7808 2321 7862 2333
rect 7908 2367 7962 2563
rect 8008 2597 8062 2609
rect 8008 2571 8018 2597
rect 8052 2571 8062 2597
rect 8008 2519 8009 2571
rect 8061 2519 8062 2571
rect 8008 2512 8062 2519
rect 8108 2597 8162 2703
rect 8208 2781 8262 2788
rect 8208 2729 8209 2781
rect 8261 2729 8262 2781
rect 8208 2703 8218 2729
rect 8252 2703 8262 2729
rect 8208 2691 8262 2703
rect 8308 2737 8362 2843
rect 8408 2877 8462 2889
rect 8408 2851 8418 2877
rect 8452 2851 8462 2877
rect 8408 2799 8409 2851
rect 8461 2799 8462 2851
rect 8408 2792 8462 2799
rect 8508 2877 8562 2983
rect 8608 3061 8662 3068
rect 8608 3009 8609 3061
rect 8661 3009 8662 3061
rect 8608 2983 8618 3009
rect 8652 2983 8662 3009
rect 8608 2971 8662 2983
rect 8708 3017 8762 3123
rect 8808 3157 8862 3169
rect 8808 3131 8818 3157
rect 8852 3131 8862 3157
rect 8808 3079 8809 3131
rect 8861 3079 8862 3131
rect 8808 3072 8862 3079
rect 8908 3157 8962 3263
rect 9008 3341 9062 3348
rect 9008 3289 9009 3341
rect 9061 3289 9062 3341
rect 9008 3263 9018 3289
rect 9052 3263 9062 3289
rect 9008 3251 9062 3263
rect 9108 3297 9162 3403
rect 9208 3437 9262 3449
rect 9208 3411 9218 3437
rect 9252 3411 9262 3437
rect 9208 3359 9209 3411
rect 9261 3359 9262 3411
rect 9208 3352 9262 3359
rect 9308 3437 9362 3543
rect 9408 3621 9462 3628
rect 9408 3569 9409 3621
rect 9461 3569 9462 3621
rect 9408 3543 9418 3569
rect 9452 3543 9462 3569
rect 9408 3531 9462 3543
rect 9508 3577 9562 3773
rect 9608 3807 9662 3819
rect 9608 3781 9618 3807
rect 9652 3781 9662 3807
rect 9608 3729 9609 3781
rect 9661 3729 9662 3781
rect 9608 3722 9662 3729
rect 9708 3807 9762 3913
rect 9808 3991 9862 3998
rect 9808 3939 9809 3991
rect 9861 3939 9862 3991
rect 9808 3913 9818 3939
rect 9852 3913 9862 3939
rect 9808 3901 9862 3913
rect 9908 3947 9962 4053
rect 10008 4087 10062 4099
rect 10008 4061 10018 4087
rect 10052 4061 10062 4087
rect 10008 4009 10009 4061
rect 10061 4009 10062 4061
rect 10008 4002 10062 4009
rect 10108 4087 10162 4193
rect 10208 4271 10262 4278
rect 10208 4219 10209 4271
rect 10261 4219 10262 4271
rect 10208 4193 10218 4219
rect 10252 4193 10262 4219
rect 10208 4181 10262 4193
rect 10308 4227 10362 4333
rect 10408 4367 10462 4379
rect 10408 4341 10418 4367
rect 10452 4341 10462 4367
rect 10408 4289 10409 4341
rect 10461 4289 10462 4341
rect 10408 4282 10462 4289
rect 10508 4367 10562 4473
rect 10608 4551 10662 4558
rect 10608 4499 10609 4551
rect 10661 4499 10662 4551
rect 10608 4473 10618 4499
rect 10652 4473 10662 4499
rect 10608 4461 10662 4473
rect 10708 4507 10762 4613
rect 10808 4647 10862 4659
rect 10808 4621 10818 4647
rect 10852 4621 10862 4647
rect 10808 4569 10809 4621
rect 10861 4569 10862 4621
rect 10808 4562 10862 4569
rect 10908 4647 10962 4753
rect 11008 4831 11062 4838
rect 11008 4779 11009 4831
rect 11061 4779 11062 4831
rect 11008 4753 11018 4779
rect 11052 4753 11062 4779
rect 11008 4741 11062 4753
rect 11108 4787 11162 4960
rect 11202 4903 11268 4904
rect 11202 4851 11209 4903
rect 11261 4851 11268 4903
rect 11202 4850 11268 4851
rect 11108 4753 11118 4787
rect 11152 4753 11162 4787
rect 10908 4613 10918 4647
rect 10952 4613 10962 4647
rect 10708 4473 10718 4507
rect 10752 4473 10762 4507
rect 10508 4333 10518 4367
rect 10552 4333 10562 4367
rect 10308 4193 10318 4227
rect 10352 4193 10362 4227
rect 10108 4053 10118 4087
rect 10152 4053 10162 4087
rect 9908 3913 9918 3947
rect 9952 3913 9962 3947
rect 9708 3773 9718 3807
rect 9752 3773 9762 3807
rect 9602 3693 9668 3694
rect 9602 3641 9609 3693
rect 9661 3641 9668 3693
rect 9602 3640 9668 3641
rect 9508 3543 9518 3577
rect 9552 3543 9562 3577
rect 9308 3403 9318 3437
rect 9352 3403 9362 3437
rect 9108 3263 9118 3297
rect 9152 3263 9162 3297
rect 8908 3123 8918 3157
rect 8952 3123 8962 3157
rect 8708 2983 8718 3017
rect 8752 2983 8762 3017
rect 8508 2843 8518 2877
rect 8552 2843 8562 2877
rect 8308 2703 8318 2737
rect 8352 2703 8362 2737
rect 8108 2563 8118 2597
rect 8152 2563 8162 2597
rect 8002 2483 8068 2484
rect 8002 2431 8009 2483
rect 8061 2431 8068 2483
rect 8002 2430 8068 2431
rect 7908 2333 7918 2367
rect 7952 2333 7962 2367
rect 7708 2193 7718 2227
rect 7752 2193 7762 2227
rect 7508 2053 7518 2087
rect 7552 2053 7562 2087
rect 7308 1913 7318 1947
rect 7352 1913 7362 1947
rect 7108 1773 7118 1807
rect 7152 1773 7162 1807
rect 6908 1633 6918 1667
rect 6952 1633 6962 1667
rect 6708 1493 6718 1527
rect 6752 1493 6762 1527
rect 6508 1353 6518 1387
rect 6552 1353 6562 1387
rect 6402 1273 6468 1274
rect 6402 1221 6409 1273
rect 6461 1221 6468 1273
rect 6402 1220 6468 1221
rect 6308 1123 6318 1157
rect 6352 1123 6362 1157
rect 6108 983 6118 1017
rect 6152 983 6162 1017
rect 5908 843 5918 877
rect 5952 843 5962 877
rect 5708 703 5718 737
rect 5752 703 5762 737
rect 5508 563 5518 597
rect 5552 563 5562 597
rect 5308 423 5318 457
rect 5352 423 5362 457
rect 5108 283 5118 317
rect 5152 283 5162 317
rect 4908 143 4918 177
rect 4952 143 4962 177
rect 4802 63 4868 64
rect 4802 11 4809 63
rect 4861 11 4868 63
rect 4802 10 4868 11
rect 4708 -67 4709 -15
rect 4761 -67 4762 -15
rect 4708 -79 4718 -67
rect 4752 -79 4762 -67
rect 4508 -132 4562 -131
rect 4508 -143 4518 -132
rect 4552 -143 4562 -132
rect 4508 -195 4509 -143
rect 4561 -195 4562 -143
rect 4508 -210 4562 -195
rect 4612 -133 4658 -81
rect 4612 -167 4618 -133
rect 4652 -167 4658 -133
rect 4518 -291 4525 -239
rect 4577 -291 4584 -239
rect 4412 -397 4418 -363
rect 4452 -397 4458 -363
rect 4412 -435 4458 -397
rect 4412 -469 4418 -435
rect 4452 -469 4458 -435
rect 4412 -512 4458 -469
rect 4509 -326 4561 -320
rect 4509 -390 4518 -378
rect 4552 -390 4561 -378
rect 4509 -454 4518 -442
rect 4552 -454 4561 -442
rect 4509 -512 4561 -506
rect 4612 -363 4658 -167
rect 4708 -131 4709 -79
rect 4761 -131 4762 -79
rect 4808 -22 4862 10
rect 4808 -74 4809 -22
rect 4861 -74 4862 -22
rect 4808 -81 4862 -74
rect 4908 -15 4962 143
rect 5008 221 5062 228
rect 5008 169 5009 221
rect 5061 169 5062 221
rect 5008 143 5018 169
rect 5052 143 5062 169
rect 5008 131 5062 143
rect 5108 177 5162 283
rect 5208 317 5262 329
rect 5208 291 5218 317
rect 5252 291 5262 317
rect 5208 239 5209 291
rect 5261 239 5262 291
rect 5208 232 5262 239
rect 5308 317 5362 423
rect 5408 501 5462 508
rect 5408 449 5409 501
rect 5461 449 5462 501
rect 5408 423 5418 449
rect 5452 423 5462 449
rect 5408 411 5462 423
rect 5508 457 5562 563
rect 5608 597 5662 609
rect 5608 571 5618 597
rect 5652 571 5662 597
rect 5608 519 5609 571
rect 5661 519 5662 571
rect 5608 512 5662 519
rect 5708 597 5762 703
rect 5808 781 5862 788
rect 5808 729 5809 781
rect 5861 729 5862 781
rect 5808 703 5818 729
rect 5852 703 5862 729
rect 5808 691 5862 703
rect 5908 737 5962 843
rect 6008 877 6062 889
rect 6008 851 6018 877
rect 6052 851 6062 877
rect 6008 799 6009 851
rect 6061 799 6062 851
rect 6008 792 6062 799
rect 6108 877 6162 983
rect 6208 1061 6262 1068
rect 6208 1009 6209 1061
rect 6261 1009 6262 1061
rect 6208 983 6218 1009
rect 6252 983 6262 1009
rect 6208 971 6262 983
rect 6308 1017 6362 1123
rect 6408 1157 6462 1169
rect 6408 1131 6418 1157
rect 6452 1131 6462 1157
rect 6408 1079 6409 1131
rect 6461 1079 6462 1131
rect 6408 1072 6462 1079
rect 6508 1157 6562 1353
rect 6608 1431 6662 1438
rect 6608 1379 6609 1431
rect 6661 1379 6662 1431
rect 6608 1353 6618 1379
rect 6652 1353 6662 1379
rect 6608 1341 6662 1353
rect 6708 1387 6762 1493
rect 6808 1527 6862 1539
rect 6808 1501 6818 1527
rect 6852 1501 6862 1527
rect 6808 1449 6809 1501
rect 6861 1449 6862 1501
rect 6808 1442 6862 1449
rect 6908 1527 6962 1633
rect 7008 1711 7062 1718
rect 7008 1659 7009 1711
rect 7061 1659 7062 1711
rect 7008 1633 7018 1659
rect 7052 1633 7062 1659
rect 7008 1621 7062 1633
rect 7108 1667 7162 1773
rect 7208 1807 7262 1819
rect 7208 1781 7218 1807
rect 7252 1781 7262 1807
rect 7208 1729 7209 1781
rect 7261 1729 7262 1781
rect 7208 1722 7262 1729
rect 7308 1807 7362 1913
rect 7408 1991 7462 1998
rect 7408 1939 7409 1991
rect 7461 1939 7462 1991
rect 7408 1913 7418 1939
rect 7452 1913 7462 1939
rect 7408 1901 7462 1913
rect 7508 1947 7562 2053
rect 7608 2087 7662 2099
rect 7608 2061 7618 2087
rect 7652 2061 7662 2087
rect 7608 2009 7609 2061
rect 7661 2009 7662 2061
rect 7608 2002 7662 2009
rect 7708 2087 7762 2193
rect 7808 2271 7862 2278
rect 7808 2219 7809 2271
rect 7861 2219 7862 2271
rect 7808 2193 7818 2219
rect 7852 2193 7862 2219
rect 7808 2181 7862 2193
rect 7908 2227 7962 2333
rect 8008 2367 8062 2379
rect 8008 2341 8018 2367
rect 8052 2341 8062 2367
rect 8008 2289 8009 2341
rect 8061 2289 8062 2341
rect 8008 2282 8062 2289
rect 8108 2367 8162 2563
rect 8208 2641 8262 2648
rect 8208 2589 8209 2641
rect 8261 2589 8262 2641
rect 8208 2563 8218 2589
rect 8252 2563 8262 2589
rect 8208 2551 8262 2563
rect 8308 2597 8362 2703
rect 8408 2737 8462 2749
rect 8408 2711 8418 2737
rect 8452 2711 8462 2737
rect 8408 2659 8409 2711
rect 8461 2659 8462 2711
rect 8408 2652 8462 2659
rect 8508 2737 8562 2843
rect 8608 2921 8662 2928
rect 8608 2869 8609 2921
rect 8661 2869 8662 2921
rect 8608 2843 8618 2869
rect 8652 2843 8662 2869
rect 8608 2831 8662 2843
rect 8708 2877 8762 2983
rect 8808 3017 8862 3029
rect 8808 2991 8818 3017
rect 8852 2991 8862 3017
rect 8808 2939 8809 2991
rect 8861 2939 8862 2991
rect 8808 2932 8862 2939
rect 8908 3017 8962 3123
rect 9008 3201 9062 3208
rect 9008 3149 9009 3201
rect 9061 3149 9062 3201
rect 9008 3123 9018 3149
rect 9052 3123 9062 3149
rect 9008 3111 9062 3123
rect 9108 3157 9162 3263
rect 9208 3297 9262 3309
rect 9208 3271 9218 3297
rect 9252 3271 9262 3297
rect 9208 3219 9209 3271
rect 9261 3219 9262 3271
rect 9208 3212 9262 3219
rect 9308 3297 9362 3403
rect 9408 3481 9462 3488
rect 9408 3429 9409 3481
rect 9461 3429 9462 3481
rect 9408 3403 9418 3429
rect 9452 3403 9462 3429
rect 9408 3391 9462 3403
rect 9508 3437 9562 3543
rect 9608 3577 9662 3589
rect 9608 3551 9618 3577
rect 9652 3551 9662 3577
rect 9608 3499 9609 3551
rect 9661 3499 9662 3551
rect 9608 3492 9662 3499
rect 9708 3577 9762 3773
rect 9808 3851 9862 3858
rect 9808 3799 9809 3851
rect 9861 3799 9862 3851
rect 9808 3773 9818 3799
rect 9852 3773 9862 3799
rect 9808 3761 9862 3773
rect 9908 3807 9962 3913
rect 10008 3947 10062 3959
rect 10008 3921 10018 3947
rect 10052 3921 10062 3947
rect 10008 3869 10009 3921
rect 10061 3869 10062 3921
rect 10008 3862 10062 3869
rect 10108 3947 10162 4053
rect 10208 4131 10262 4138
rect 10208 4079 10209 4131
rect 10261 4079 10262 4131
rect 10208 4053 10218 4079
rect 10252 4053 10262 4079
rect 10208 4041 10262 4053
rect 10308 4087 10362 4193
rect 10408 4227 10462 4239
rect 10408 4201 10418 4227
rect 10452 4201 10462 4227
rect 10408 4149 10409 4201
rect 10461 4149 10462 4201
rect 10408 4142 10462 4149
rect 10508 4227 10562 4333
rect 10608 4411 10662 4418
rect 10608 4359 10609 4411
rect 10661 4359 10662 4411
rect 10608 4333 10618 4359
rect 10652 4333 10662 4359
rect 10608 4321 10662 4333
rect 10708 4367 10762 4473
rect 10808 4507 10862 4519
rect 10808 4481 10818 4507
rect 10852 4481 10862 4507
rect 10808 4429 10809 4481
rect 10861 4429 10862 4481
rect 10808 4422 10862 4429
rect 10908 4507 10962 4613
rect 11008 4691 11062 4698
rect 11008 4639 11009 4691
rect 11061 4639 11062 4691
rect 11008 4613 11018 4639
rect 11052 4613 11062 4639
rect 11008 4601 11062 4613
rect 11108 4647 11162 4753
rect 11208 4787 11262 4799
rect 11208 4761 11218 4787
rect 11252 4761 11262 4787
rect 11208 4709 11209 4761
rect 11261 4709 11262 4761
rect 11208 4702 11262 4709
rect 11308 4787 11362 4960
rect 11402 4919 11468 4920
rect 11402 4867 11409 4919
rect 11461 4867 11468 4919
rect 11402 4866 11468 4867
rect 11308 4753 11318 4787
rect 11352 4753 11362 4787
rect 11108 4613 11118 4647
rect 11152 4613 11162 4647
rect 10908 4473 10918 4507
rect 10952 4473 10962 4507
rect 10708 4333 10718 4367
rect 10752 4333 10762 4367
rect 10508 4193 10518 4227
rect 10552 4193 10562 4227
rect 10308 4053 10318 4087
rect 10352 4053 10362 4087
rect 10108 3913 10118 3947
rect 10152 3913 10162 3947
rect 9908 3773 9918 3807
rect 9952 3773 9962 3807
rect 9802 3709 9868 3710
rect 9802 3657 9809 3709
rect 9861 3657 9868 3709
rect 9802 3656 9868 3657
rect 9708 3543 9718 3577
rect 9752 3543 9762 3577
rect 9508 3403 9518 3437
rect 9552 3403 9562 3437
rect 9308 3263 9318 3297
rect 9352 3263 9362 3297
rect 9108 3123 9118 3157
rect 9152 3123 9162 3157
rect 8908 2983 8918 3017
rect 8952 2983 8962 3017
rect 8708 2843 8718 2877
rect 8752 2843 8762 2877
rect 8508 2703 8518 2737
rect 8552 2703 8562 2737
rect 8308 2563 8318 2597
rect 8352 2563 8362 2597
rect 8202 2499 8268 2500
rect 8202 2447 8209 2499
rect 8261 2447 8268 2499
rect 8202 2446 8268 2447
rect 8108 2333 8118 2367
rect 8152 2333 8162 2367
rect 7908 2193 7918 2227
rect 7952 2193 7962 2227
rect 7708 2053 7718 2087
rect 7752 2053 7762 2087
rect 7508 1913 7518 1947
rect 7552 1913 7562 1947
rect 7308 1773 7318 1807
rect 7352 1773 7362 1807
rect 7108 1633 7118 1667
rect 7152 1633 7162 1667
rect 6908 1493 6918 1527
rect 6952 1493 6962 1527
rect 6708 1353 6718 1387
rect 6752 1353 6762 1387
rect 6602 1289 6668 1290
rect 6602 1237 6609 1289
rect 6661 1237 6668 1289
rect 6602 1236 6668 1237
rect 6508 1123 6518 1157
rect 6552 1123 6562 1157
rect 6308 983 6318 1017
rect 6352 983 6362 1017
rect 6108 843 6118 877
rect 6152 843 6162 877
rect 5908 703 5918 737
rect 5952 703 5962 737
rect 5708 563 5718 597
rect 5752 563 5762 597
rect 5508 423 5518 457
rect 5552 423 5562 457
rect 5308 283 5318 317
rect 5352 283 5362 317
rect 5108 143 5118 177
rect 5152 143 5162 177
rect 5002 79 5068 80
rect 5002 27 5009 79
rect 5061 27 5068 79
rect 5002 26 5068 27
rect 4908 -67 4909 -15
rect 4961 -67 4962 -15
rect 4908 -79 4918 -67
rect 4952 -79 4962 -67
rect 4708 -132 4762 -131
rect 4708 -143 4718 -132
rect 4752 -143 4762 -132
rect 4708 -195 4709 -143
rect 4761 -195 4762 -143
rect 4708 -210 4762 -195
rect 4812 -133 4858 -81
rect 4812 -167 4818 -133
rect 4852 -167 4858 -133
rect 4718 -291 4725 -239
rect 4777 -291 4784 -239
rect 4612 -397 4618 -363
rect 4652 -397 4658 -363
rect 4612 -435 4658 -397
rect 4612 -469 4618 -435
rect 4652 -469 4658 -435
rect 4612 -512 4658 -469
rect 4709 -326 4761 -320
rect 4709 -390 4718 -378
rect 4752 -390 4761 -378
rect 4709 -454 4718 -442
rect 4752 -454 4761 -442
rect 4709 -555 4761 -506
rect 4812 -363 4858 -167
rect 4908 -131 4909 -79
rect 4961 -131 4962 -79
rect 5008 -22 5062 26
rect 5008 -74 5009 -22
rect 5061 -74 5062 -22
rect 5008 -81 5062 -74
rect 5108 -15 5162 143
rect 5208 177 5262 189
rect 5208 151 5218 177
rect 5252 151 5262 177
rect 5208 99 5209 151
rect 5261 99 5262 151
rect 5208 92 5262 99
rect 5308 177 5362 283
rect 5408 361 5462 368
rect 5408 309 5409 361
rect 5461 309 5462 361
rect 5408 283 5418 309
rect 5452 283 5462 309
rect 5408 271 5462 283
rect 5508 317 5562 423
rect 5608 457 5662 469
rect 5608 431 5618 457
rect 5652 431 5662 457
rect 5608 379 5609 431
rect 5661 379 5662 431
rect 5608 372 5662 379
rect 5708 457 5762 563
rect 5808 641 5862 648
rect 5808 589 5809 641
rect 5861 589 5862 641
rect 5808 563 5818 589
rect 5852 563 5862 589
rect 5808 551 5862 563
rect 5908 597 5962 703
rect 6008 737 6062 749
rect 6008 711 6018 737
rect 6052 711 6062 737
rect 6008 659 6009 711
rect 6061 659 6062 711
rect 6008 652 6062 659
rect 6108 737 6162 843
rect 6208 921 6262 928
rect 6208 869 6209 921
rect 6261 869 6262 921
rect 6208 843 6218 869
rect 6252 843 6262 869
rect 6208 831 6262 843
rect 6308 877 6362 983
rect 6408 1017 6462 1029
rect 6408 991 6418 1017
rect 6452 991 6462 1017
rect 6408 939 6409 991
rect 6461 939 6462 991
rect 6408 932 6462 939
rect 6508 1017 6562 1123
rect 6608 1201 6662 1208
rect 6608 1149 6609 1201
rect 6661 1149 6662 1201
rect 6608 1123 6618 1149
rect 6652 1123 6662 1149
rect 6608 1111 6662 1123
rect 6708 1157 6762 1353
rect 6808 1387 6862 1399
rect 6808 1361 6818 1387
rect 6852 1361 6862 1387
rect 6808 1309 6809 1361
rect 6861 1309 6862 1361
rect 6808 1302 6862 1309
rect 6908 1387 6962 1493
rect 7008 1571 7062 1578
rect 7008 1519 7009 1571
rect 7061 1519 7062 1571
rect 7008 1493 7018 1519
rect 7052 1493 7062 1519
rect 7008 1481 7062 1493
rect 7108 1527 7162 1633
rect 7208 1667 7262 1679
rect 7208 1641 7218 1667
rect 7252 1641 7262 1667
rect 7208 1589 7209 1641
rect 7261 1589 7262 1641
rect 7208 1582 7262 1589
rect 7308 1667 7362 1773
rect 7408 1851 7462 1858
rect 7408 1799 7409 1851
rect 7461 1799 7462 1851
rect 7408 1773 7418 1799
rect 7452 1773 7462 1799
rect 7408 1761 7462 1773
rect 7508 1807 7562 1913
rect 7608 1947 7662 1959
rect 7608 1921 7618 1947
rect 7652 1921 7662 1947
rect 7608 1869 7609 1921
rect 7661 1869 7662 1921
rect 7608 1862 7662 1869
rect 7708 1947 7762 2053
rect 7808 2131 7862 2138
rect 7808 2079 7809 2131
rect 7861 2079 7862 2131
rect 7808 2053 7818 2079
rect 7852 2053 7862 2079
rect 7808 2041 7862 2053
rect 7908 2087 7962 2193
rect 8008 2227 8062 2239
rect 8008 2201 8018 2227
rect 8052 2201 8062 2227
rect 8008 2149 8009 2201
rect 8061 2149 8062 2201
rect 8008 2142 8062 2149
rect 8108 2227 8162 2333
rect 8208 2411 8262 2418
rect 8208 2359 8209 2411
rect 8261 2359 8262 2411
rect 8208 2333 8218 2359
rect 8252 2333 8262 2359
rect 8208 2321 8262 2333
rect 8308 2367 8362 2563
rect 8408 2597 8462 2609
rect 8408 2571 8418 2597
rect 8452 2571 8462 2597
rect 8408 2519 8409 2571
rect 8461 2519 8462 2571
rect 8408 2512 8462 2519
rect 8508 2597 8562 2703
rect 8608 2781 8662 2788
rect 8608 2729 8609 2781
rect 8661 2729 8662 2781
rect 8608 2703 8618 2729
rect 8652 2703 8662 2729
rect 8608 2691 8662 2703
rect 8708 2737 8762 2843
rect 8808 2877 8862 2889
rect 8808 2851 8818 2877
rect 8852 2851 8862 2877
rect 8808 2799 8809 2851
rect 8861 2799 8862 2851
rect 8808 2792 8862 2799
rect 8908 2877 8962 2983
rect 9008 3061 9062 3068
rect 9008 3009 9009 3061
rect 9061 3009 9062 3061
rect 9008 2983 9018 3009
rect 9052 2983 9062 3009
rect 9008 2971 9062 2983
rect 9108 3017 9162 3123
rect 9208 3157 9262 3169
rect 9208 3131 9218 3157
rect 9252 3131 9262 3157
rect 9208 3079 9209 3131
rect 9261 3079 9262 3131
rect 9208 3072 9262 3079
rect 9308 3157 9362 3263
rect 9408 3341 9462 3348
rect 9408 3289 9409 3341
rect 9461 3289 9462 3341
rect 9408 3263 9418 3289
rect 9452 3263 9462 3289
rect 9408 3251 9462 3263
rect 9508 3297 9562 3403
rect 9608 3437 9662 3449
rect 9608 3411 9618 3437
rect 9652 3411 9662 3437
rect 9608 3359 9609 3411
rect 9661 3359 9662 3411
rect 9608 3352 9662 3359
rect 9708 3437 9762 3543
rect 9808 3621 9862 3628
rect 9808 3569 9809 3621
rect 9861 3569 9862 3621
rect 9808 3543 9818 3569
rect 9852 3543 9862 3569
rect 9808 3531 9862 3543
rect 9908 3577 9962 3773
rect 10008 3807 10062 3819
rect 10008 3781 10018 3807
rect 10052 3781 10062 3807
rect 10008 3729 10009 3781
rect 10061 3729 10062 3781
rect 10008 3722 10062 3729
rect 10108 3807 10162 3913
rect 10208 3991 10262 3998
rect 10208 3939 10209 3991
rect 10261 3939 10262 3991
rect 10208 3913 10218 3939
rect 10252 3913 10262 3939
rect 10208 3901 10262 3913
rect 10308 3947 10362 4053
rect 10408 4087 10462 4099
rect 10408 4061 10418 4087
rect 10452 4061 10462 4087
rect 10408 4009 10409 4061
rect 10461 4009 10462 4061
rect 10408 4002 10462 4009
rect 10508 4087 10562 4193
rect 10608 4271 10662 4278
rect 10608 4219 10609 4271
rect 10661 4219 10662 4271
rect 10608 4193 10618 4219
rect 10652 4193 10662 4219
rect 10608 4181 10662 4193
rect 10708 4227 10762 4333
rect 10808 4367 10862 4379
rect 10808 4341 10818 4367
rect 10852 4341 10862 4367
rect 10808 4289 10809 4341
rect 10861 4289 10862 4341
rect 10808 4282 10862 4289
rect 10908 4367 10962 4473
rect 11008 4551 11062 4558
rect 11008 4499 11009 4551
rect 11061 4499 11062 4551
rect 11008 4473 11018 4499
rect 11052 4473 11062 4499
rect 11008 4461 11062 4473
rect 11108 4507 11162 4613
rect 11208 4647 11262 4659
rect 11208 4621 11218 4647
rect 11252 4621 11262 4647
rect 11208 4569 11209 4621
rect 11261 4569 11262 4621
rect 11208 4562 11262 4569
rect 11308 4647 11362 4753
rect 11408 4831 11462 4838
rect 11408 4779 11409 4831
rect 11461 4779 11462 4831
rect 11408 4753 11418 4779
rect 11452 4753 11462 4779
rect 11408 4741 11462 4753
rect 11508 4787 11562 4960
rect 11602 4903 11668 4904
rect 11602 4851 11609 4903
rect 11661 4851 11668 4903
rect 11602 4850 11668 4851
rect 11508 4753 11518 4787
rect 11552 4753 11562 4787
rect 11308 4613 11318 4647
rect 11352 4613 11362 4647
rect 11108 4473 11118 4507
rect 11152 4473 11162 4507
rect 10908 4333 10918 4367
rect 10952 4333 10962 4367
rect 10708 4193 10718 4227
rect 10752 4193 10762 4227
rect 10508 4053 10518 4087
rect 10552 4053 10562 4087
rect 10308 3913 10318 3947
rect 10352 3913 10362 3947
rect 10108 3773 10118 3807
rect 10152 3773 10162 3807
rect 10002 3693 10068 3694
rect 10002 3641 10009 3693
rect 10061 3641 10068 3693
rect 10002 3640 10068 3641
rect 9908 3543 9918 3577
rect 9952 3543 9962 3577
rect 9708 3403 9718 3437
rect 9752 3403 9762 3437
rect 9508 3263 9518 3297
rect 9552 3263 9562 3297
rect 9308 3123 9318 3157
rect 9352 3123 9362 3157
rect 9108 2983 9118 3017
rect 9152 2983 9162 3017
rect 8908 2843 8918 2877
rect 8952 2843 8962 2877
rect 8708 2703 8718 2737
rect 8752 2703 8762 2737
rect 8508 2563 8518 2597
rect 8552 2563 8562 2597
rect 8402 2483 8468 2484
rect 8402 2431 8409 2483
rect 8461 2431 8468 2483
rect 8402 2430 8468 2431
rect 8308 2333 8318 2367
rect 8352 2333 8362 2367
rect 8108 2193 8118 2227
rect 8152 2193 8162 2227
rect 7908 2053 7918 2087
rect 7952 2053 7962 2087
rect 7708 1913 7718 1947
rect 7752 1913 7762 1947
rect 7508 1773 7518 1807
rect 7552 1773 7562 1807
rect 7308 1633 7318 1667
rect 7352 1633 7362 1667
rect 7108 1493 7118 1527
rect 7152 1493 7162 1527
rect 6908 1353 6918 1387
rect 6952 1353 6962 1387
rect 6802 1273 6868 1274
rect 6802 1221 6809 1273
rect 6861 1221 6868 1273
rect 6802 1220 6868 1221
rect 6708 1123 6718 1157
rect 6752 1123 6762 1157
rect 6508 983 6518 1017
rect 6552 983 6562 1017
rect 6308 843 6318 877
rect 6352 843 6362 877
rect 6108 703 6118 737
rect 6152 703 6162 737
rect 5908 563 5918 597
rect 5952 563 5962 597
rect 5708 423 5718 457
rect 5752 423 5762 457
rect 5508 283 5518 317
rect 5552 283 5562 317
rect 5308 143 5318 177
rect 5352 143 5362 177
rect 5202 63 5268 64
rect 5202 11 5209 63
rect 5261 11 5268 63
rect 5202 10 5268 11
rect 5108 -67 5109 -15
rect 5161 -67 5162 -15
rect 5108 -79 5118 -67
rect 5152 -79 5162 -67
rect 4908 -132 4962 -131
rect 4908 -143 4918 -132
rect 4952 -143 4962 -132
rect 4908 -195 4909 -143
rect 4961 -195 4962 -143
rect 4908 -210 4962 -195
rect 5012 -133 5058 -81
rect 5012 -167 5018 -133
rect 5052 -167 5058 -133
rect 4918 -291 4925 -239
rect 4977 -291 4984 -239
rect 4812 -397 4818 -363
rect 4852 -397 4858 -363
rect 4812 -435 4858 -397
rect 4812 -469 4818 -435
rect 4852 -469 4858 -435
rect 4812 -512 4858 -469
rect 4909 -326 4961 -320
rect 4909 -390 4918 -378
rect 4952 -390 4961 -378
rect 4909 -454 4918 -442
rect 4952 -454 4961 -442
rect 4909 -512 4961 -506
rect 5012 -363 5058 -167
rect 5108 -131 5109 -79
rect 5161 -131 5162 -79
rect 5208 -22 5262 10
rect 5208 -74 5209 -22
rect 5261 -74 5262 -22
rect 5208 -81 5262 -74
rect 5308 -15 5362 143
rect 5408 221 5462 228
rect 5408 169 5409 221
rect 5461 169 5462 221
rect 5408 143 5418 169
rect 5452 143 5462 169
rect 5408 131 5462 143
rect 5508 177 5562 283
rect 5608 317 5662 329
rect 5608 291 5618 317
rect 5652 291 5662 317
rect 5608 239 5609 291
rect 5661 239 5662 291
rect 5608 232 5662 239
rect 5708 317 5762 423
rect 5808 501 5862 508
rect 5808 449 5809 501
rect 5861 449 5862 501
rect 5808 423 5818 449
rect 5852 423 5862 449
rect 5808 411 5862 423
rect 5908 457 5962 563
rect 6008 597 6062 609
rect 6008 571 6018 597
rect 6052 571 6062 597
rect 6008 519 6009 571
rect 6061 519 6062 571
rect 6008 512 6062 519
rect 6108 597 6162 703
rect 6208 781 6262 788
rect 6208 729 6209 781
rect 6261 729 6262 781
rect 6208 703 6218 729
rect 6252 703 6262 729
rect 6208 691 6262 703
rect 6308 737 6362 843
rect 6408 877 6462 889
rect 6408 851 6418 877
rect 6452 851 6462 877
rect 6408 799 6409 851
rect 6461 799 6462 851
rect 6408 792 6462 799
rect 6508 877 6562 983
rect 6608 1061 6662 1068
rect 6608 1009 6609 1061
rect 6661 1009 6662 1061
rect 6608 983 6618 1009
rect 6652 983 6662 1009
rect 6608 971 6662 983
rect 6708 1017 6762 1123
rect 6808 1157 6862 1169
rect 6808 1131 6818 1157
rect 6852 1131 6862 1157
rect 6808 1079 6809 1131
rect 6861 1079 6862 1131
rect 6808 1072 6862 1079
rect 6908 1157 6962 1353
rect 7008 1431 7062 1438
rect 7008 1379 7009 1431
rect 7061 1379 7062 1431
rect 7008 1353 7018 1379
rect 7052 1353 7062 1379
rect 7008 1341 7062 1353
rect 7108 1387 7162 1493
rect 7208 1527 7262 1539
rect 7208 1501 7218 1527
rect 7252 1501 7262 1527
rect 7208 1449 7209 1501
rect 7261 1449 7262 1501
rect 7208 1442 7262 1449
rect 7308 1527 7362 1633
rect 7408 1711 7462 1718
rect 7408 1659 7409 1711
rect 7461 1659 7462 1711
rect 7408 1633 7418 1659
rect 7452 1633 7462 1659
rect 7408 1621 7462 1633
rect 7508 1667 7562 1773
rect 7608 1807 7662 1819
rect 7608 1781 7618 1807
rect 7652 1781 7662 1807
rect 7608 1729 7609 1781
rect 7661 1729 7662 1781
rect 7608 1722 7662 1729
rect 7708 1807 7762 1913
rect 7808 1991 7862 1998
rect 7808 1939 7809 1991
rect 7861 1939 7862 1991
rect 7808 1913 7818 1939
rect 7852 1913 7862 1939
rect 7808 1901 7862 1913
rect 7908 1947 7962 2053
rect 8008 2087 8062 2099
rect 8008 2061 8018 2087
rect 8052 2061 8062 2087
rect 8008 2009 8009 2061
rect 8061 2009 8062 2061
rect 8008 2002 8062 2009
rect 8108 2087 8162 2193
rect 8208 2271 8262 2278
rect 8208 2219 8209 2271
rect 8261 2219 8262 2271
rect 8208 2193 8218 2219
rect 8252 2193 8262 2219
rect 8208 2181 8262 2193
rect 8308 2227 8362 2333
rect 8408 2367 8462 2379
rect 8408 2341 8418 2367
rect 8452 2341 8462 2367
rect 8408 2289 8409 2341
rect 8461 2289 8462 2341
rect 8408 2282 8462 2289
rect 8508 2367 8562 2563
rect 8608 2641 8662 2648
rect 8608 2589 8609 2641
rect 8661 2589 8662 2641
rect 8608 2563 8618 2589
rect 8652 2563 8662 2589
rect 8608 2551 8662 2563
rect 8708 2597 8762 2703
rect 8808 2737 8862 2749
rect 8808 2711 8818 2737
rect 8852 2711 8862 2737
rect 8808 2659 8809 2711
rect 8861 2659 8862 2711
rect 8808 2652 8862 2659
rect 8908 2737 8962 2843
rect 9008 2921 9062 2928
rect 9008 2869 9009 2921
rect 9061 2869 9062 2921
rect 9008 2843 9018 2869
rect 9052 2843 9062 2869
rect 9008 2831 9062 2843
rect 9108 2877 9162 2983
rect 9208 3017 9262 3029
rect 9208 2991 9218 3017
rect 9252 2991 9262 3017
rect 9208 2939 9209 2991
rect 9261 2939 9262 2991
rect 9208 2932 9262 2939
rect 9308 3017 9362 3123
rect 9408 3201 9462 3208
rect 9408 3149 9409 3201
rect 9461 3149 9462 3201
rect 9408 3123 9418 3149
rect 9452 3123 9462 3149
rect 9408 3111 9462 3123
rect 9508 3157 9562 3263
rect 9608 3297 9662 3309
rect 9608 3271 9618 3297
rect 9652 3271 9662 3297
rect 9608 3219 9609 3271
rect 9661 3219 9662 3271
rect 9608 3212 9662 3219
rect 9708 3297 9762 3403
rect 9808 3481 9862 3488
rect 9808 3429 9809 3481
rect 9861 3429 9862 3481
rect 9808 3403 9818 3429
rect 9852 3403 9862 3429
rect 9808 3391 9862 3403
rect 9908 3437 9962 3543
rect 10008 3577 10062 3589
rect 10008 3551 10018 3577
rect 10052 3551 10062 3577
rect 10008 3499 10009 3551
rect 10061 3499 10062 3551
rect 10008 3492 10062 3499
rect 10108 3577 10162 3773
rect 10208 3851 10262 3858
rect 10208 3799 10209 3851
rect 10261 3799 10262 3851
rect 10208 3773 10218 3799
rect 10252 3773 10262 3799
rect 10208 3761 10262 3773
rect 10308 3807 10362 3913
rect 10408 3947 10462 3959
rect 10408 3921 10418 3947
rect 10452 3921 10462 3947
rect 10408 3869 10409 3921
rect 10461 3869 10462 3921
rect 10408 3862 10462 3869
rect 10508 3947 10562 4053
rect 10608 4131 10662 4138
rect 10608 4079 10609 4131
rect 10661 4079 10662 4131
rect 10608 4053 10618 4079
rect 10652 4053 10662 4079
rect 10608 4041 10662 4053
rect 10708 4087 10762 4193
rect 10808 4227 10862 4239
rect 10808 4201 10818 4227
rect 10852 4201 10862 4227
rect 10808 4149 10809 4201
rect 10861 4149 10862 4201
rect 10808 4142 10862 4149
rect 10908 4227 10962 4333
rect 11008 4411 11062 4418
rect 11008 4359 11009 4411
rect 11061 4359 11062 4411
rect 11008 4333 11018 4359
rect 11052 4333 11062 4359
rect 11008 4321 11062 4333
rect 11108 4367 11162 4473
rect 11208 4507 11262 4519
rect 11208 4481 11218 4507
rect 11252 4481 11262 4507
rect 11208 4429 11209 4481
rect 11261 4429 11262 4481
rect 11208 4422 11262 4429
rect 11308 4507 11362 4613
rect 11408 4691 11462 4698
rect 11408 4639 11409 4691
rect 11461 4639 11462 4691
rect 11408 4613 11418 4639
rect 11452 4613 11462 4639
rect 11408 4601 11462 4613
rect 11508 4647 11562 4753
rect 11608 4787 11662 4799
rect 11608 4761 11618 4787
rect 11652 4761 11662 4787
rect 11608 4709 11609 4761
rect 11661 4709 11662 4761
rect 11608 4702 11662 4709
rect 11708 4787 11762 4960
rect 11802 4919 11868 4920
rect 11802 4867 11809 4919
rect 11861 4867 11868 4919
rect 11802 4866 11868 4867
rect 11708 4753 11718 4787
rect 11752 4753 11762 4787
rect 11508 4613 11518 4647
rect 11552 4613 11562 4647
rect 11308 4473 11318 4507
rect 11352 4473 11362 4507
rect 11108 4333 11118 4367
rect 11152 4333 11162 4367
rect 10908 4193 10918 4227
rect 10952 4193 10962 4227
rect 10708 4053 10718 4087
rect 10752 4053 10762 4087
rect 10508 3913 10518 3947
rect 10552 3913 10562 3947
rect 10308 3773 10318 3807
rect 10352 3773 10362 3807
rect 10202 3709 10268 3710
rect 10202 3657 10209 3709
rect 10261 3657 10268 3709
rect 10202 3656 10268 3657
rect 10108 3543 10118 3577
rect 10152 3543 10162 3577
rect 9908 3403 9918 3437
rect 9952 3403 9962 3437
rect 9708 3263 9718 3297
rect 9752 3263 9762 3297
rect 9508 3123 9518 3157
rect 9552 3123 9562 3157
rect 9308 2983 9318 3017
rect 9352 2983 9362 3017
rect 9108 2843 9118 2877
rect 9152 2843 9162 2877
rect 8908 2703 8918 2737
rect 8952 2703 8962 2737
rect 8708 2563 8718 2597
rect 8752 2563 8762 2597
rect 8602 2499 8668 2500
rect 8602 2447 8609 2499
rect 8661 2447 8668 2499
rect 8602 2446 8668 2447
rect 8508 2333 8518 2367
rect 8552 2333 8562 2367
rect 8308 2193 8318 2227
rect 8352 2193 8362 2227
rect 8108 2053 8118 2087
rect 8152 2053 8162 2087
rect 7908 1913 7918 1947
rect 7952 1913 7962 1947
rect 7708 1773 7718 1807
rect 7752 1773 7762 1807
rect 7508 1633 7518 1667
rect 7552 1633 7562 1667
rect 7308 1493 7318 1527
rect 7352 1493 7362 1527
rect 7108 1353 7118 1387
rect 7152 1353 7162 1387
rect 7002 1289 7068 1290
rect 7002 1237 7009 1289
rect 7061 1237 7068 1289
rect 7002 1236 7068 1237
rect 6908 1123 6918 1157
rect 6952 1123 6962 1157
rect 6708 983 6718 1017
rect 6752 983 6762 1017
rect 6508 843 6518 877
rect 6552 843 6562 877
rect 6308 703 6318 737
rect 6352 703 6362 737
rect 6108 563 6118 597
rect 6152 563 6162 597
rect 5908 423 5918 457
rect 5952 423 5962 457
rect 5708 283 5718 317
rect 5752 283 5762 317
rect 5508 143 5518 177
rect 5552 143 5562 177
rect 5402 79 5468 80
rect 5402 27 5409 79
rect 5461 27 5468 79
rect 5402 26 5468 27
rect 5308 -67 5309 -15
rect 5361 -67 5362 -15
rect 5308 -79 5318 -67
rect 5352 -79 5362 -67
rect 5108 -132 5162 -131
rect 5108 -143 5118 -132
rect 5152 -143 5162 -132
rect 5108 -195 5109 -143
rect 5161 -195 5162 -143
rect 5108 -210 5162 -195
rect 5212 -133 5258 -81
rect 5212 -167 5218 -133
rect 5252 -167 5258 -133
rect 5118 -291 5125 -239
rect 5177 -291 5184 -239
rect 5012 -397 5018 -363
rect 5052 -397 5058 -363
rect 5012 -435 5058 -397
rect 5012 -469 5018 -435
rect 5052 -469 5058 -435
rect 5012 -512 5058 -469
rect 5109 -326 5161 -320
rect 5109 -390 5118 -378
rect 5152 -390 5161 -378
rect 5109 -454 5118 -442
rect 5152 -454 5161 -442
rect 5109 -555 5161 -506
rect 5212 -363 5258 -167
rect 5308 -131 5309 -79
rect 5361 -131 5362 -79
rect 5408 -22 5462 26
rect 5408 -74 5409 -22
rect 5461 -74 5462 -22
rect 5408 -81 5462 -74
rect 5508 -15 5562 143
rect 5608 177 5662 189
rect 5608 151 5618 177
rect 5652 151 5662 177
rect 5608 99 5609 151
rect 5661 99 5662 151
rect 5608 92 5662 99
rect 5708 177 5762 283
rect 5808 361 5862 368
rect 5808 309 5809 361
rect 5861 309 5862 361
rect 5808 283 5818 309
rect 5852 283 5862 309
rect 5808 271 5862 283
rect 5908 317 5962 423
rect 6008 457 6062 469
rect 6008 431 6018 457
rect 6052 431 6062 457
rect 6008 379 6009 431
rect 6061 379 6062 431
rect 6008 372 6062 379
rect 6108 457 6162 563
rect 6208 641 6262 648
rect 6208 589 6209 641
rect 6261 589 6262 641
rect 6208 563 6218 589
rect 6252 563 6262 589
rect 6208 551 6262 563
rect 6308 597 6362 703
rect 6408 737 6462 749
rect 6408 711 6418 737
rect 6452 711 6462 737
rect 6408 659 6409 711
rect 6461 659 6462 711
rect 6408 652 6462 659
rect 6508 737 6562 843
rect 6608 921 6662 928
rect 6608 869 6609 921
rect 6661 869 6662 921
rect 6608 843 6618 869
rect 6652 843 6662 869
rect 6608 831 6662 843
rect 6708 877 6762 983
rect 6808 1017 6862 1029
rect 6808 991 6818 1017
rect 6852 991 6862 1017
rect 6808 939 6809 991
rect 6861 939 6862 991
rect 6808 932 6862 939
rect 6908 1017 6962 1123
rect 7008 1201 7062 1208
rect 7008 1149 7009 1201
rect 7061 1149 7062 1201
rect 7008 1123 7018 1149
rect 7052 1123 7062 1149
rect 7008 1111 7062 1123
rect 7108 1157 7162 1353
rect 7208 1387 7262 1399
rect 7208 1361 7218 1387
rect 7252 1361 7262 1387
rect 7208 1309 7209 1361
rect 7261 1309 7262 1361
rect 7208 1302 7262 1309
rect 7308 1387 7362 1493
rect 7408 1571 7462 1578
rect 7408 1519 7409 1571
rect 7461 1519 7462 1571
rect 7408 1493 7418 1519
rect 7452 1493 7462 1519
rect 7408 1481 7462 1493
rect 7508 1527 7562 1633
rect 7608 1667 7662 1679
rect 7608 1641 7618 1667
rect 7652 1641 7662 1667
rect 7608 1589 7609 1641
rect 7661 1589 7662 1641
rect 7608 1582 7662 1589
rect 7708 1667 7762 1773
rect 7808 1851 7862 1858
rect 7808 1799 7809 1851
rect 7861 1799 7862 1851
rect 7808 1773 7818 1799
rect 7852 1773 7862 1799
rect 7808 1761 7862 1773
rect 7908 1807 7962 1913
rect 8008 1947 8062 1959
rect 8008 1921 8018 1947
rect 8052 1921 8062 1947
rect 8008 1869 8009 1921
rect 8061 1869 8062 1921
rect 8008 1862 8062 1869
rect 8108 1947 8162 2053
rect 8208 2131 8262 2138
rect 8208 2079 8209 2131
rect 8261 2079 8262 2131
rect 8208 2053 8218 2079
rect 8252 2053 8262 2079
rect 8208 2041 8262 2053
rect 8308 2087 8362 2193
rect 8408 2227 8462 2239
rect 8408 2201 8418 2227
rect 8452 2201 8462 2227
rect 8408 2149 8409 2201
rect 8461 2149 8462 2201
rect 8408 2142 8462 2149
rect 8508 2227 8562 2333
rect 8608 2411 8662 2418
rect 8608 2359 8609 2411
rect 8661 2359 8662 2411
rect 8608 2333 8618 2359
rect 8652 2333 8662 2359
rect 8608 2321 8662 2333
rect 8708 2367 8762 2563
rect 8808 2597 8862 2609
rect 8808 2571 8818 2597
rect 8852 2571 8862 2597
rect 8808 2519 8809 2571
rect 8861 2519 8862 2571
rect 8808 2512 8862 2519
rect 8908 2597 8962 2703
rect 9008 2781 9062 2788
rect 9008 2729 9009 2781
rect 9061 2729 9062 2781
rect 9008 2703 9018 2729
rect 9052 2703 9062 2729
rect 9008 2691 9062 2703
rect 9108 2737 9162 2843
rect 9208 2877 9262 2889
rect 9208 2851 9218 2877
rect 9252 2851 9262 2877
rect 9208 2799 9209 2851
rect 9261 2799 9262 2851
rect 9208 2792 9262 2799
rect 9308 2877 9362 2983
rect 9408 3061 9462 3068
rect 9408 3009 9409 3061
rect 9461 3009 9462 3061
rect 9408 2983 9418 3009
rect 9452 2983 9462 3009
rect 9408 2971 9462 2983
rect 9508 3017 9562 3123
rect 9608 3157 9662 3169
rect 9608 3131 9618 3157
rect 9652 3131 9662 3157
rect 9608 3079 9609 3131
rect 9661 3079 9662 3131
rect 9608 3072 9662 3079
rect 9708 3157 9762 3263
rect 9808 3341 9862 3348
rect 9808 3289 9809 3341
rect 9861 3289 9862 3341
rect 9808 3263 9818 3289
rect 9852 3263 9862 3289
rect 9808 3251 9862 3263
rect 9908 3297 9962 3403
rect 10008 3437 10062 3449
rect 10008 3411 10018 3437
rect 10052 3411 10062 3437
rect 10008 3359 10009 3411
rect 10061 3359 10062 3411
rect 10008 3352 10062 3359
rect 10108 3437 10162 3543
rect 10208 3621 10262 3628
rect 10208 3569 10209 3621
rect 10261 3569 10262 3621
rect 10208 3543 10218 3569
rect 10252 3543 10262 3569
rect 10208 3531 10262 3543
rect 10308 3577 10362 3773
rect 10408 3807 10462 3819
rect 10408 3781 10418 3807
rect 10452 3781 10462 3807
rect 10408 3729 10409 3781
rect 10461 3729 10462 3781
rect 10408 3722 10462 3729
rect 10508 3807 10562 3913
rect 10608 3991 10662 3998
rect 10608 3939 10609 3991
rect 10661 3939 10662 3991
rect 10608 3913 10618 3939
rect 10652 3913 10662 3939
rect 10608 3901 10662 3913
rect 10708 3947 10762 4053
rect 10808 4087 10862 4099
rect 10808 4061 10818 4087
rect 10852 4061 10862 4087
rect 10808 4009 10809 4061
rect 10861 4009 10862 4061
rect 10808 4002 10862 4009
rect 10908 4087 10962 4193
rect 11008 4271 11062 4278
rect 11008 4219 11009 4271
rect 11061 4219 11062 4271
rect 11008 4193 11018 4219
rect 11052 4193 11062 4219
rect 11008 4181 11062 4193
rect 11108 4227 11162 4333
rect 11208 4367 11262 4379
rect 11208 4341 11218 4367
rect 11252 4341 11262 4367
rect 11208 4289 11209 4341
rect 11261 4289 11262 4341
rect 11208 4282 11262 4289
rect 11308 4367 11362 4473
rect 11408 4551 11462 4558
rect 11408 4499 11409 4551
rect 11461 4499 11462 4551
rect 11408 4473 11418 4499
rect 11452 4473 11462 4499
rect 11408 4461 11462 4473
rect 11508 4507 11562 4613
rect 11608 4647 11662 4659
rect 11608 4621 11618 4647
rect 11652 4621 11662 4647
rect 11608 4569 11609 4621
rect 11661 4569 11662 4621
rect 11608 4562 11662 4569
rect 11708 4647 11762 4753
rect 11808 4831 11862 4838
rect 11808 4779 11809 4831
rect 11861 4779 11862 4831
rect 11808 4753 11818 4779
rect 11852 4753 11862 4779
rect 11808 4741 11862 4753
rect 11908 4787 11962 4960
rect 12002 4903 12068 4904
rect 12002 4851 12009 4903
rect 12061 4851 12068 4903
rect 12002 4850 12068 4851
rect 11908 4753 11918 4787
rect 11952 4753 11962 4787
rect 11708 4613 11718 4647
rect 11752 4613 11762 4647
rect 11508 4473 11518 4507
rect 11552 4473 11562 4507
rect 11308 4333 11318 4367
rect 11352 4333 11362 4367
rect 11108 4193 11118 4227
rect 11152 4193 11162 4227
rect 10908 4053 10918 4087
rect 10952 4053 10962 4087
rect 10708 3913 10718 3947
rect 10752 3913 10762 3947
rect 10508 3773 10518 3807
rect 10552 3773 10562 3807
rect 10402 3693 10468 3694
rect 10402 3641 10409 3693
rect 10461 3641 10468 3693
rect 10402 3640 10468 3641
rect 10308 3543 10318 3577
rect 10352 3543 10362 3577
rect 10108 3403 10118 3437
rect 10152 3403 10162 3437
rect 9908 3263 9918 3297
rect 9952 3263 9962 3297
rect 9708 3123 9718 3157
rect 9752 3123 9762 3157
rect 9508 2983 9518 3017
rect 9552 2983 9562 3017
rect 9308 2843 9318 2877
rect 9352 2843 9362 2877
rect 9108 2703 9118 2737
rect 9152 2703 9162 2737
rect 8908 2563 8918 2597
rect 8952 2563 8962 2597
rect 8802 2483 8868 2484
rect 8802 2431 8809 2483
rect 8861 2431 8868 2483
rect 8802 2430 8868 2431
rect 8708 2333 8718 2367
rect 8752 2333 8762 2367
rect 8508 2193 8518 2227
rect 8552 2193 8562 2227
rect 8308 2053 8318 2087
rect 8352 2053 8362 2087
rect 8108 1913 8118 1947
rect 8152 1913 8162 1947
rect 7908 1773 7918 1807
rect 7952 1773 7962 1807
rect 7708 1633 7718 1667
rect 7752 1633 7762 1667
rect 7508 1493 7518 1527
rect 7552 1493 7562 1527
rect 7308 1353 7318 1387
rect 7352 1353 7362 1387
rect 7202 1273 7268 1274
rect 7202 1221 7209 1273
rect 7261 1221 7268 1273
rect 7202 1220 7268 1221
rect 7108 1123 7118 1157
rect 7152 1123 7162 1157
rect 6908 983 6918 1017
rect 6952 983 6962 1017
rect 6708 843 6718 877
rect 6752 843 6762 877
rect 6508 703 6518 737
rect 6552 703 6562 737
rect 6308 563 6318 597
rect 6352 563 6362 597
rect 6108 423 6118 457
rect 6152 423 6162 457
rect 5908 283 5918 317
rect 5952 283 5962 317
rect 5708 143 5718 177
rect 5752 143 5762 177
rect 5602 63 5668 64
rect 5602 11 5609 63
rect 5661 11 5668 63
rect 5602 10 5668 11
rect 5508 -67 5509 -15
rect 5561 -67 5562 -15
rect 5508 -79 5518 -67
rect 5552 -79 5562 -67
rect 5308 -132 5362 -131
rect 5308 -143 5318 -132
rect 5352 -143 5362 -132
rect 5308 -195 5309 -143
rect 5361 -195 5362 -143
rect 5308 -210 5362 -195
rect 5412 -133 5458 -81
rect 5412 -167 5418 -133
rect 5452 -167 5458 -133
rect 5318 -291 5325 -239
rect 5377 -291 5384 -239
rect 5212 -397 5218 -363
rect 5252 -397 5258 -363
rect 5212 -435 5258 -397
rect 5212 -469 5218 -435
rect 5252 -469 5258 -435
rect 5212 -512 5258 -469
rect 5309 -326 5361 -320
rect 5309 -390 5318 -378
rect 5352 -390 5361 -378
rect 5309 -454 5318 -442
rect 5352 -454 5361 -442
rect 5309 -512 5361 -506
rect 5412 -363 5458 -167
rect 5508 -131 5509 -79
rect 5561 -131 5562 -79
rect 5608 -22 5662 10
rect 5608 -74 5609 -22
rect 5661 -74 5662 -22
rect 5608 -81 5662 -74
rect 5708 -15 5762 143
rect 5808 221 5862 228
rect 5808 169 5809 221
rect 5861 169 5862 221
rect 5808 143 5818 169
rect 5852 143 5862 169
rect 5808 131 5862 143
rect 5908 177 5962 283
rect 6008 317 6062 329
rect 6008 291 6018 317
rect 6052 291 6062 317
rect 6008 239 6009 291
rect 6061 239 6062 291
rect 6008 232 6062 239
rect 6108 317 6162 423
rect 6208 501 6262 508
rect 6208 449 6209 501
rect 6261 449 6262 501
rect 6208 423 6218 449
rect 6252 423 6262 449
rect 6208 411 6262 423
rect 6308 457 6362 563
rect 6408 597 6462 609
rect 6408 571 6418 597
rect 6452 571 6462 597
rect 6408 519 6409 571
rect 6461 519 6462 571
rect 6408 512 6462 519
rect 6508 597 6562 703
rect 6608 781 6662 788
rect 6608 729 6609 781
rect 6661 729 6662 781
rect 6608 703 6618 729
rect 6652 703 6662 729
rect 6608 691 6662 703
rect 6708 737 6762 843
rect 6808 877 6862 889
rect 6808 851 6818 877
rect 6852 851 6862 877
rect 6808 799 6809 851
rect 6861 799 6862 851
rect 6808 792 6862 799
rect 6908 877 6962 983
rect 7008 1061 7062 1068
rect 7008 1009 7009 1061
rect 7061 1009 7062 1061
rect 7008 983 7018 1009
rect 7052 983 7062 1009
rect 7008 971 7062 983
rect 7108 1017 7162 1123
rect 7208 1157 7262 1169
rect 7208 1131 7218 1157
rect 7252 1131 7262 1157
rect 7208 1079 7209 1131
rect 7261 1079 7262 1131
rect 7208 1072 7262 1079
rect 7308 1157 7362 1353
rect 7408 1431 7462 1438
rect 7408 1379 7409 1431
rect 7461 1379 7462 1431
rect 7408 1353 7418 1379
rect 7452 1353 7462 1379
rect 7408 1341 7462 1353
rect 7508 1387 7562 1493
rect 7608 1527 7662 1539
rect 7608 1501 7618 1527
rect 7652 1501 7662 1527
rect 7608 1449 7609 1501
rect 7661 1449 7662 1501
rect 7608 1442 7662 1449
rect 7708 1527 7762 1633
rect 7808 1711 7862 1718
rect 7808 1659 7809 1711
rect 7861 1659 7862 1711
rect 7808 1633 7818 1659
rect 7852 1633 7862 1659
rect 7808 1621 7862 1633
rect 7908 1667 7962 1773
rect 8008 1807 8062 1819
rect 8008 1781 8018 1807
rect 8052 1781 8062 1807
rect 8008 1729 8009 1781
rect 8061 1729 8062 1781
rect 8008 1722 8062 1729
rect 8108 1807 8162 1913
rect 8208 1991 8262 1998
rect 8208 1939 8209 1991
rect 8261 1939 8262 1991
rect 8208 1913 8218 1939
rect 8252 1913 8262 1939
rect 8208 1901 8262 1913
rect 8308 1947 8362 2053
rect 8408 2087 8462 2099
rect 8408 2061 8418 2087
rect 8452 2061 8462 2087
rect 8408 2009 8409 2061
rect 8461 2009 8462 2061
rect 8408 2002 8462 2009
rect 8508 2087 8562 2193
rect 8608 2271 8662 2278
rect 8608 2219 8609 2271
rect 8661 2219 8662 2271
rect 8608 2193 8618 2219
rect 8652 2193 8662 2219
rect 8608 2181 8662 2193
rect 8708 2227 8762 2333
rect 8808 2367 8862 2379
rect 8808 2341 8818 2367
rect 8852 2341 8862 2367
rect 8808 2289 8809 2341
rect 8861 2289 8862 2341
rect 8808 2282 8862 2289
rect 8908 2367 8962 2563
rect 9008 2641 9062 2648
rect 9008 2589 9009 2641
rect 9061 2589 9062 2641
rect 9008 2563 9018 2589
rect 9052 2563 9062 2589
rect 9008 2551 9062 2563
rect 9108 2597 9162 2703
rect 9208 2737 9262 2749
rect 9208 2711 9218 2737
rect 9252 2711 9262 2737
rect 9208 2659 9209 2711
rect 9261 2659 9262 2711
rect 9208 2652 9262 2659
rect 9308 2737 9362 2843
rect 9408 2921 9462 2928
rect 9408 2869 9409 2921
rect 9461 2869 9462 2921
rect 9408 2843 9418 2869
rect 9452 2843 9462 2869
rect 9408 2831 9462 2843
rect 9508 2877 9562 2983
rect 9608 3017 9662 3029
rect 9608 2991 9618 3017
rect 9652 2991 9662 3017
rect 9608 2939 9609 2991
rect 9661 2939 9662 2991
rect 9608 2932 9662 2939
rect 9708 3017 9762 3123
rect 9808 3201 9862 3208
rect 9808 3149 9809 3201
rect 9861 3149 9862 3201
rect 9808 3123 9818 3149
rect 9852 3123 9862 3149
rect 9808 3111 9862 3123
rect 9908 3157 9962 3263
rect 10008 3297 10062 3309
rect 10008 3271 10018 3297
rect 10052 3271 10062 3297
rect 10008 3219 10009 3271
rect 10061 3219 10062 3271
rect 10008 3212 10062 3219
rect 10108 3297 10162 3403
rect 10208 3481 10262 3488
rect 10208 3429 10209 3481
rect 10261 3429 10262 3481
rect 10208 3403 10218 3429
rect 10252 3403 10262 3429
rect 10208 3391 10262 3403
rect 10308 3437 10362 3543
rect 10408 3577 10462 3589
rect 10408 3551 10418 3577
rect 10452 3551 10462 3577
rect 10408 3499 10409 3551
rect 10461 3499 10462 3551
rect 10408 3492 10462 3499
rect 10508 3577 10562 3773
rect 10608 3851 10662 3858
rect 10608 3799 10609 3851
rect 10661 3799 10662 3851
rect 10608 3773 10618 3799
rect 10652 3773 10662 3799
rect 10608 3761 10662 3773
rect 10708 3807 10762 3913
rect 10808 3947 10862 3959
rect 10808 3921 10818 3947
rect 10852 3921 10862 3947
rect 10808 3869 10809 3921
rect 10861 3869 10862 3921
rect 10808 3862 10862 3869
rect 10908 3947 10962 4053
rect 11008 4131 11062 4138
rect 11008 4079 11009 4131
rect 11061 4079 11062 4131
rect 11008 4053 11018 4079
rect 11052 4053 11062 4079
rect 11008 4041 11062 4053
rect 11108 4087 11162 4193
rect 11208 4227 11262 4239
rect 11208 4201 11218 4227
rect 11252 4201 11262 4227
rect 11208 4149 11209 4201
rect 11261 4149 11262 4201
rect 11208 4142 11262 4149
rect 11308 4227 11362 4333
rect 11408 4411 11462 4418
rect 11408 4359 11409 4411
rect 11461 4359 11462 4411
rect 11408 4333 11418 4359
rect 11452 4333 11462 4359
rect 11408 4321 11462 4333
rect 11508 4367 11562 4473
rect 11608 4507 11662 4519
rect 11608 4481 11618 4507
rect 11652 4481 11662 4507
rect 11608 4429 11609 4481
rect 11661 4429 11662 4481
rect 11608 4422 11662 4429
rect 11708 4507 11762 4613
rect 11808 4691 11862 4698
rect 11808 4639 11809 4691
rect 11861 4639 11862 4691
rect 11808 4613 11818 4639
rect 11852 4613 11862 4639
rect 11808 4601 11862 4613
rect 11908 4647 11962 4753
rect 12008 4787 12062 4799
rect 12008 4761 12018 4787
rect 12052 4761 12062 4787
rect 12008 4709 12009 4761
rect 12061 4709 12062 4761
rect 12008 4702 12062 4709
rect 12108 4787 12162 4960
rect 12202 4919 12268 4920
rect 12202 4867 12209 4919
rect 12261 4867 12268 4919
rect 12202 4866 12268 4867
rect 12108 4753 12118 4787
rect 12152 4753 12162 4787
rect 11908 4613 11918 4647
rect 11952 4613 11962 4647
rect 11708 4473 11718 4507
rect 11752 4473 11762 4507
rect 11508 4333 11518 4367
rect 11552 4333 11562 4367
rect 11308 4193 11318 4227
rect 11352 4193 11362 4227
rect 11108 4053 11118 4087
rect 11152 4053 11162 4087
rect 10908 3913 10918 3947
rect 10952 3913 10962 3947
rect 10708 3773 10718 3807
rect 10752 3773 10762 3807
rect 10602 3709 10668 3710
rect 10602 3657 10609 3709
rect 10661 3657 10668 3709
rect 10602 3656 10668 3657
rect 10508 3543 10518 3577
rect 10552 3543 10562 3577
rect 10308 3403 10318 3437
rect 10352 3403 10362 3437
rect 10108 3263 10118 3297
rect 10152 3263 10162 3297
rect 9908 3123 9918 3157
rect 9952 3123 9962 3157
rect 9708 2983 9718 3017
rect 9752 2983 9762 3017
rect 9508 2843 9518 2877
rect 9552 2843 9562 2877
rect 9308 2703 9318 2737
rect 9352 2703 9362 2737
rect 9108 2563 9118 2597
rect 9152 2563 9162 2597
rect 9002 2499 9068 2500
rect 9002 2447 9009 2499
rect 9061 2447 9068 2499
rect 9002 2446 9068 2447
rect 8908 2333 8918 2367
rect 8952 2333 8962 2367
rect 8708 2193 8718 2227
rect 8752 2193 8762 2227
rect 8508 2053 8518 2087
rect 8552 2053 8562 2087
rect 8308 1913 8318 1947
rect 8352 1913 8362 1947
rect 8108 1773 8118 1807
rect 8152 1773 8162 1807
rect 7908 1633 7918 1667
rect 7952 1633 7962 1667
rect 7708 1493 7718 1527
rect 7752 1493 7762 1527
rect 7508 1353 7518 1387
rect 7552 1353 7562 1387
rect 7402 1289 7468 1290
rect 7402 1237 7409 1289
rect 7461 1237 7468 1289
rect 7402 1236 7468 1237
rect 7308 1123 7318 1157
rect 7352 1123 7362 1157
rect 7108 983 7118 1017
rect 7152 983 7162 1017
rect 6908 843 6918 877
rect 6952 843 6962 877
rect 6708 703 6718 737
rect 6752 703 6762 737
rect 6508 563 6518 597
rect 6552 563 6562 597
rect 6308 423 6318 457
rect 6352 423 6362 457
rect 6108 283 6118 317
rect 6152 283 6162 317
rect 5908 143 5918 177
rect 5952 143 5962 177
rect 5802 79 5868 80
rect 5802 27 5809 79
rect 5861 27 5868 79
rect 5802 26 5868 27
rect 5708 -67 5709 -15
rect 5761 -67 5762 -15
rect 5708 -79 5718 -67
rect 5752 -79 5762 -67
rect 5508 -132 5562 -131
rect 5508 -143 5518 -132
rect 5552 -143 5562 -132
rect 5508 -195 5509 -143
rect 5561 -195 5562 -143
rect 5508 -210 5562 -195
rect 5612 -133 5658 -81
rect 5612 -167 5618 -133
rect 5652 -167 5658 -133
rect 5518 -291 5525 -239
rect 5577 -291 5584 -239
rect 5412 -397 5418 -363
rect 5452 -397 5458 -363
rect 5412 -435 5458 -397
rect 5412 -469 5418 -435
rect 5452 -469 5458 -435
rect 5412 -512 5458 -469
rect 5509 -326 5561 -320
rect 5509 -390 5518 -378
rect 5552 -390 5561 -378
rect 5509 -454 5518 -442
rect 5552 -454 5561 -442
rect 5509 -555 5561 -506
rect 5612 -363 5658 -167
rect 5708 -131 5709 -79
rect 5761 -131 5762 -79
rect 5808 -22 5862 26
rect 5808 -74 5809 -22
rect 5861 -74 5862 -22
rect 5808 -81 5862 -74
rect 5908 -15 5962 143
rect 6008 177 6062 189
rect 6008 151 6018 177
rect 6052 151 6062 177
rect 6008 99 6009 151
rect 6061 99 6062 151
rect 6008 92 6062 99
rect 6108 177 6162 283
rect 6208 361 6262 368
rect 6208 309 6209 361
rect 6261 309 6262 361
rect 6208 283 6218 309
rect 6252 283 6262 309
rect 6208 271 6262 283
rect 6308 317 6362 423
rect 6408 457 6462 469
rect 6408 431 6418 457
rect 6452 431 6462 457
rect 6408 379 6409 431
rect 6461 379 6462 431
rect 6408 372 6462 379
rect 6508 457 6562 563
rect 6608 641 6662 648
rect 6608 589 6609 641
rect 6661 589 6662 641
rect 6608 563 6618 589
rect 6652 563 6662 589
rect 6608 551 6662 563
rect 6708 597 6762 703
rect 6808 737 6862 749
rect 6808 711 6818 737
rect 6852 711 6862 737
rect 6808 659 6809 711
rect 6861 659 6862 711
rect 6808 652 6862 659
rect 6908 737 6962 843
rect 7008 921 7062 928
rect 7008 869 7009 921
rect 7061 869 7062 921
rect 7008 843 7018 869
rect 7052 843 7062 869
rect 7008 831 7062 843
rect 7108 877 7162 983
rect 7208 1017 7262 1029
rect 7208 991 7218 1017
rect 7252 991 7262 1017
rect 7208 939 7209 991
rect 7261 939 7262 991
rect 7208 932 7262 939
rect 7308 1017 7362 1123
rect 7408 1201 7462 1208
rect 7408 1149 7409 1201
rect 7461 1149 7462 1201
rect 7408 1123 7418 1149
rect 7452 1123 7462 1149
rect 7408 1111 7462 1123
rect 7508 1157 7562 1353
rect 7608 1387 7662 1399
rect 7608 1361 7618 1387
rect 7652 1361 7662 1387
rect 7608 1309 7609 1361
rect 7661 1309 7662 1361
rect 7608 1302 7662 1309
rect 7708 1387 7762 1493
rect 7808 1571 7862 1578
rect 7808 1519 7809 1571
rect 7861 1519 7862 1571
rect 7808 1493 7818 1519
rect 7852 1493 7862 1519
rect 7808 1481 7862 1493
rect 7908 1527 7962 1633
rect 8008 1667 8062 1679
rect 8008 1641 8018 1667
rect 8052 1641 8062 1667
rect 8008 1589 8009 1641
rect 8061 1589 8062 1641
rect 8008 1582 8062 1589
rect 8108 1667 8162 1773
rect 8208 1851 8262 1858
rect 8208 1799 8209 1851
rect 8261 1799 8262 1851
rect 8208 1773 8218 1799
rect 8252 1773 8262 1799
rect 8208 1761 8262 1773
rect 8308 1807 8362 1913
rect 8408 1947 8462 1959
rect 8408 1921 8418 1947
rect 8452 1921 8462 1947
rect 8408 1869 8409 1921
rect 8461 1869 8462 1921
rect 8408 1862 8462 1869
rect 8508 1947 8562 2053
rect 8608 2131 8662 2138
rect 8608 2079 8609 2131
rect 8661 2079 8662 2131
rect 8608 2053 8618 2079
rect 8652 2053 8662 2079
rect 8608 2041 8662 2053
rect 8708 2087 8762 2193
rect 8808 2227 8862 2239
rect 8808 2201 8818 2227
rect 8852 2201 8862 2227
rect 8808 2149 8809 2201
rect 8861 2149 8862 2201
rect 8808 2142 8862 2149
rect 8908 2227 8962 2333
rect 9008 2411 9062 2418
rect 9008 2359 9009 2411
rect 9061 2359 9062 2411
rect 9008 2333 9018 2359
rect 9052 2333 9062 2359
rect 9008 2321 9062 2333
rect 9108 2367 9162 2563
rect 9208 2597 9262 2609
rect 9208 2571 9218 2597
rect 9252 2571 9262 2597
rect 9208 2519 9209 2571
rect 9261 2519 9262 2571
rect 9208 2512 9262 2519
rect 9308 2597 9362 2703
rect 9408 2781 9462 2788
rect 9408 2729 9409 2781
rect 9461 2729 9462 2781
rect 9408 2703 9418 2729
rect 9452 2703 9462 2729
rect 9408 2691 9462 2703
rect 9508 2737 9562 2843
rect 9608 2877 9662 2889
rect 9608 2851 9618 2877
rect 9652 2851 9662 2877
rect 9608 2799 9609 2851
rect 9661 2799 9662 2851
rect 9608 2792 9662 2799
rect 9708 2877 9762 2983
rect 9808 3061 9862 3068
rect 9808 3009 9809 3061
rect 9861 3009 9862 3061
rect 9808 2983 9818 3009
rect 9852 2983 9862 3009
rect 9808 2971 9862 2983
rect 9908 3017 9962 3123
rect 10008 3157 10062 3169
rect 10008 3131 10018 3157
rect 10052 3131 10062 3157
rect 10008 3079 10009 3131
rect 10061 3079 10062 3131
rect 10008 3072 10062 3079
rect 10108 3157 10162 3263
rect 10208 3341 10262 3348
rect 10208 3289 10209 3341
rect 10261 3289 10262 3341
rect 10208 3263 10218 3289
rect 10252 3263 10262 3289
rect 10208 3251 10262 3263
rect 10308 3297 10362 3403
rect 10408 3437 10462 3449
rect 10408 3411 10418 3437
rect 10452 3411 10462 3437
rect 10408 3359 10409 3411
rect 10461 3359 10462 3411
rect 10408 3352 10462 3359
rect 10508 3437 10562 3543
rect 10608 3621 10662 3628
rect 10608 3569 10609 3621
rect 10661 3569 10662 3621
rect 10608 3543 10618 3569
rect 10652 3543 10662 3569
rect 10608 3531 10662 3543
rect 10708 3577 10762 3773
rect 10808 3807 10862 3819
rect 10808 3781 10818 3807
rect 10852 3781 10862 3807
rect 10808 3729 10809 3781
rect 10861 3729 10862 3781
rect 10808 3722 10862 3729
rect 10908 3807 10962 3913
rect 11008 3991 11062 3998
rect 11008 3939 11009 3991
rect 11061 3939 11062 3991
rect 11008 3913 11018 3939
rect 11052 3913 11062 3939
rect 11008 3901 11062 3913
rect 11108 3947 11162 4053
rect 11208 4087 11262 4099
rect 11208 4061 11218 4087
rect 11252 4061 11262 4087
rect 11208 4009 11209 4061
rect 11261 4009 11262 4061
rect 11208 4002 11262 4009
rect 11308 4087 11362 4193
rect 11408 4271 11462 4278
rect 11408 4219 11409 4271
rect 11461 4219 11462 4271
rect 11408 4193 11418 4219
rect 11452 4193 11462 4219
rect 11408 4181 11462 4193
rect 11508 4227 11562 4333
rect 11608 4367 11662 4379
rect 11608 4341 11618 4367
rect 11652 4341 11662 4367
rect 11608 4289 11609 4341
rect 11661 4289 11662 4341
rect 11608 4282 11662 4289
rect 11708 4367 11762 4473
rect 11808 4551 11862 4558
rect 11808 4499 11809 4551
rect 11861 4499 11862 4551
rect 11808 4473 11818 4499
rect 11852 4473 11862 4499
rect 11808 4461 11862 4473
rect 11908 4507 11962 4613
rect 12008 4647 12062 4659
rect 12008 4621 12018 4647
rect 12052 4621 12062 4647
rect 12008 4569 12009 4621
rect 12061 4569 12062 4621
rect 12008 4562 12062 4569
rect 12108 4647 12162 4753
rect 12208 4831 12262 4838
rect 12208 4779 12209 4831
rect 12261 4779 12262 4831
rect 12208 4753 12218 4779
rect 12252 4753 12262 4779
rect 12208 4741 12262 4753
rect 12308 4787 12362 4960
rect 12402 4903 12468 4904
rect 12402 4851 12409 4903
rect 12461 4851 12468 4903
rect 12402 4850 12468 4851
rect 12308 4753 12318 4787
rect 12352 4753 12362 4787
rect 12108 4613 12118 4647
rect 12152 4613 12162 4647
rect 11908 4473 11918 4507
rect 11952 4473 11962 4507
rect 11708 4333 11718 4367
rect 11752 4333 11762 4367
rect 11508 4193 11518 4227
rect 11552 4193 11562 4227
rect 11308 4053 11318 4087
rect 11352 4053 11362 4087
rect 11108 3913 11118 3947
rect 11152 3913 11162 3947
rect 10908 3773 10918 3807
rect 10952 3773 10962 3807
rect 10802 3693 10868 3694
rect 10802 3641 10809 3693
rect 10861 3641 10868 3693
rect 10802 3640 10868 3641
rect 10708 3543 10718 3577
rect 10752 3543 10762 3577
rect 10508 3403 10518 3437
rect 10552 3403 10562 3437
rect 10308 3263 10318 3297
rect 10352 3263 10362 3297
rect 10108 3123 10118 3157
rect 10152 3123 10162 3157
rect 9908 2983 9918 3017
rect 9952 2983 9962 3017
rect 9708 2843 9718 2877
rect 9752 2843 9762 2877
rect 9508 2703 9518 2737
rect 9552 2703 9562 2737
rect 9308 2563 9318 2597
rect 9352 2563 9362 2597
rect 9202 2483 9268 2484
rect 9202 2431 9209 2483
rect 9261 2431 9268 2483
rect 9202 2430 9268 2431
rect 9108 2333 9118 2367
rect 9152 2333 9162 2367
rect 8908 2193 8918 2227
rect 8952 2193 8962 2227
rect 8708 2053 8718 2087
rect 8752 2053 8762 2087
rect 8508 1913 8518 1947
rect 8552 1913 8562 1947
rect 8308 1773 8318 1807
rect 8352 1773 8362 1807
rect 8108 1633 8118 1667
rect 8152 1633 8162 1667
rect 7908 1493 7918 1527
rect 7952 1493 7962 1527
rect 7708 1353 7718 1387
rect 7752 1353 7762 1387
rect 7602 1273 7668 1274
rect 7602 1221 7609 1273
rect 7661 1221 7668 1273
rect 7602 1220 7668 1221
rect 7508 1123 7518 1157
rect 7552 1123 7562 1157
rect 7308 983 7318 1017
rect 7352 983 7362 1017
rect 7108 843 7118 877
rect 7152 843 7162 877
rect 6908 703 6918 737
rect 6952 703 6962 737
rect 6708 563 6718 597
rect 6752 563 6762 597
rect 6508 423 6518 457
rect 6552 423 6562 457
rect 6308 283 6318 317
rect 6352 283 6362 317
rect 6108 143 6118 177
rect 6152 143 6162 177
rect 6002 63 6068 64
rect 6002 11 6009 63
rect 6061 11 6068 63
rect 6002 10 6068 11
rect 5908 -67 5909 -15
rect 5961 -67 5962 -15
rect 5908 -79 5918 -67
rect 5952 -79 5962 -67
rect 5708 -132 5762 -131
rect 5708 -143 5718 -132
rect 5752 -143 5762 -132
rect 5708 -195 5709 -143
rect 5761 -195 5762 -143
rect 5708 -210 5762 -195
rect 5812 -133 5858 -81
rect 5812 -167 5818 -133
rect 5852 -167 5858 -133
rect 5718 -291 5725 -239
rect 5777 -291 5784 -239
rect 5612 -397 5618 -363
rect 5652 -397 5658 -363
rect 5612 -435 5658 -397
rect 5612 -469 5618 -435
rect 5652 -469 5658 -435
rect 5612 -512 5658 -469
rect 5709 -326 5761 -320
rect 5709 -390 5718 -378
rect 5752 -390 5761 -378
rect 5709 -454 5718 -442
rect 5752 -454 5761 -442
rect 5709 -512 5761 -506
rect 5812 -363 5858 -167
rect 5908 -131 5909 -79
rect 5961 -131 5962 -79
rect 6008 -22 6062 10
rect 6008 -74 6009 -22
rect 6061 -74 6062 -22
rect 6008 -81 6062 -74
rect 6108 -15 6162 143
rect 6208 221 6262 228
rect 6208 169 6209 221
rect 6261 169 6262 221
rect 6208 143 6218 169
rect 6252 143 6262 169
rect 6208 131 6262 143
rect 6308 177 6362 283
rect 6408 317 6462 329
rect 6408 291 6418 317
rect 6452 291 6462 317
rect 6408 239 6409 291
rect 6461 239 6462 291
rect 6408 232 6462 239
rect 6508 317 6562 423
rect 6608 501 6662 508
rect 6608 449 6609 501
rect 6661 449 6662 501
rect 6608 423 6618 449
rect 6652 423 6662 449
rect 6608 411 6662 423
rect 6708 457 6762 563
rect 6808 597 6862 609
rect 6808 571 6818 597
rect 6852 571 6862 597
rect 6808 519 6809 571
rect 6861 519 6862 571
rect 6808 512 6862 519
rect 6908 597 6962 703
rect 7008 781 7062 788
rect 7008 729 7009 781
rect 7061 729 7062 781
rect 7008 703 7018 729
rect 7052 703 7062 729
rect 7008 691 7062 703
rect 7108 737 7162 843
rect 7208 877 7262 889
rect 7208 851 7218 877
rect 7252 851 7262 877
rect 7208 799 7209 851
rect 7261 799 7262 851
rect 7208 792 7262 799
rect 7308 877 7362 983
rect 7408 1061 7462 1068
rect 7408 1009 7409 1061
rect 7461 1009 7462 1061
rect 7408 983 7418 1009
rect 7452 983 7462 1009
rect 7408 971 7462 983
rect 7508 1017 7562 1123
rect 7608 1157 7662 1169
rect 7608 1131 7618 1157
rect 7652 1131 7662 1157
rect 7608 1079 7609 1131
rect 7661 1079 7662 1131
rect 7608 1072 7662 1079
rect 7708 1157 7762 1353
rect 7808 1431 7862 1438
rect 7808 1379 7809 1431
rect 7861 1379 7862 1431
rect 7808 1353 7818 1379
rect 7852 1353 7862 1379
rect 7808 1341 7862 1353
rect 7908 1387 7962 1493
rect 8008 1527 8062 1539
rect 8008 1501 8018 1527
rect 8052 1501 8062 1527
rect 8008 1449 8009 1501
rect 8061 1449 8062 1501
rect 8008 1442 8062 1449
rect 8108 1527 8162 1633
rect 8208 1711 8262 1718
rect 8208 1659 8209 1711
rect 8261 1659 8262 1711
rect 8208 1633 8218 1659
rect 8252 1633 8262 1659
rect 8208 1621 8262 1633
rect 8308 1667 8362 1773
rect 8408 1807 8462 1819
rect 8408 1781 8418 1807
rect 8452 1781 8462 1807
rect 8408 1729 8409 1781
rect 8461 1729 8462 1781
rect 8408 1722 8462 1729
rect 8508 1807 8562 1913
rect 8608 1991 8662 1998
rect 8608 1939 8609 1991
rect 8661 1939 8662 1991
rect 8608 1913 8618 1939
rect 8652 1913 8662 1939
rect 8608 1901 8662 1913
rect 8708 1947 8762 2053
rect 8808 2087 8862 2099
rect 8808 2061 8818 2087
rect 8852 2061 8862 2087
rect 8808 2009 8809 2061
rect 8861 2009 8862 2061
rect 8808 2002 8862 2009
rect 8908 2087 8962 2193
rect 9008 2271 9062 2278
rect 9008 2219 9009 2271
rect 9061 2219 9062 2271
rect 9008 2193 9018 2219
rect 9052 2193 9062 2219
rect 9008 2181 9062 2193
rect 9108 2227 9162 2333
rect 9208 2367 9262 2379
rect 9208 2341 9218 2367
rect 9252 2341 9262 2367
rect 9208 2289 9209 2341
rect 9261 2289 9262 2341
rect 9208 2282 9262 2289
rect 9308 2367 9362 2563
rect 9408 2641 9462 2648
rect 9408 2589 9409 2641
rect 9461 2589 9462 2641
rect 9408 2563 9418 2589
rect 9452 2563 9462 2589
rect 9408 2551 9462 2563
rect 9508 2597 9562 2703
rect 9608 2737 9662 2749
rect 9608 2711 9618 2737
rect 9652 2711 9662 2737
rect 9608 2659 9609 2711
rect 9661 2659 9662 2711
rect 9608 2652 9662 2659
rect 9708 2737 9762 2843
rect 9808 2921 9862 2928
rect 9808 2869 9809 2921
rect 9861 2869 9862 2921
rect 9808 2843 9818 2869
rect 9852 2843 9862 2869
rect 9808 2831 9862 2843
rect 9908 2877 9962 2983
rect 10008 3017 10062 3029
rect 10008 2991 10018 3017
rect 10052 2991 10062 3017
rect 10008 2939 10009 2991
rect 10061 2939 10062 2991
rect 10008 2932 10062 2939
rect 10108 3017 10162 3123
rect 10208 3201 10262 3208
rect 10208 3149 10209 3201
rect 10261 3149 10262 3201
rect 10208 3123 10218 3149
rect 10252 3123 10262 3149
rect 10208 3111 10262 3123
rect 10308 3157 10362 3263
rect 10408 3297 10462 3309
rect 10408 3271 10418 3297
rect 10452 3271 10462 3297
rect 10408 3219 10409 3271
rect 10461 3219 10462 3271
rect 10408 3212 10462 3219
rect 10508 3297 10562 3403
rect 10608 3481 10662 3488
rect 10608 3429 10609 3481
rect 10661 3429 10662 3481
rect 10608 3403 10618 3429
rect 10652 3403 10662 3429
rect 10608 3391 10662 3403
rect 10708 3437 10762 3543
rect 10808 3577 10862 3589
rect 10808 3551 10818 3577
rect 10852 3551 10862 3577
rect 10808 3499 10809 3551
rect 10861 3499 10862 3551
rect 10808 3492 10862 3499
rect 10908 3577 10962 3773
rect 11008 3851 11062 3858
rect 11008 3799 11009 3851
rect 11061 3799 11062 3851
rect 11008 3773 11018 3799
rect 11052 3773 11062 3799
rect 11008 3761 11062 3773
rect 11108 3807 11162 3913
rect 11208 3947 11262 3959
rect 11208 3921 11218 3947
rect 11252 3921 11262 3947
rect 11208 3869 11209 3921
rect 11261 3869 11262 3921
rect 11208 3862 11262 3869
rect 11308 3947 11362 4053
rect 11408 4131 11462 4138
rect 11408 4079 11409 4131
rect 11461 4079 11462 4131
rect 11408 4053 11418 4079
rect 11452 4053 11462 4079
rect 11408 4041 11462 4053
rect 11508 4087 11562 4193
rect 11608 4227 11662 4239
rect 11608 4201 11618 4227
rect 11652 4201 11662 4227
rect 11608 4149 11609 4201
rect 11661 4149 11662 4201
rect 11608 4142 11662 4149
rect 11708 4227 11762 4333
rect 11808 4411 11862 4418
rect 11808 4359 11809 4411
rect 11861 4359 11862 4411
rect 11808 4333 11818 4359
rect 11852 4333 11862 4359
rect 11808 4321 11862 4333
rect 11908 4367 11962 4473
rect 12008 4507 12062 4519
rect 12008 4481 12018 4507
rect 12052 4481 12062 4507
rect 12008 4429 12009 4481
rect 12061 4429 12062 4481
rect 12008 4422 12062 4429
rect 12108 4507 12162 4613
rect 12208 4691 12262 4698
rect 12208 4639 12209 4691
rect 12261 4639 12262 4691
rect 12208 4613 12218 4639
rect 12252 4613 12262 4639
rect 12208 4601 12262 4613
rect 12308 4647 12362 4753
rect 12408 4787 12462 4799
rect 12408 4761 12418 4787
rect 12452 4761 12462 4787
rect 12408 4709 12409 4761
rect 12461 4709 12462 4761
rect 12408 4702 12462 4709
rect 12508 4787 12562 4960
rect 12602 4919 12668 4920
rect 12602 4867 12609 4919
rect 12661 4867 12668 4919
rect 12602 4866 12668 4867
rect 12508 4753 12518 4787
rect 12552 4753 12562 4787
rect 12308 4613 12318 4647
rect 12352 4613 12362 4647
rect 12108 4473 12118 4507
rect 12152 4473 12162 4507
rect 11908 4333 11918 4367
rect 11952 4333 11962 4367
rect 11708 4193 11718 4227
rect 11752 4193 11762 4227
rect 11508 4053 11518 4087
rect 11552 4053 11562 4087
rect 11308 3913 11318 3947
rect 11352 3913 11362 3947
rect 11108 3773 11118 3807
rect 11152 3773 11162 3807
rect 11002 3709 11068 3710
rect 11002 3657 11009 3709
rect 11061 3657 11068 3709
rect 11002 3656 11068 3657
rect 10908 3543 10918 3577
rect 10952 3543 10962 3577
rect 10708 3403 10718 3437
rect 10752 3403 10762 3437
rect 10508 3263 10518 3297
rect 10552 3263 10562 3297
rect 10308 3123 10318 3157
rect 10352 3123 10362 3157
rect 10108 2983 10118 3017
rect 10152 2983 10162 3017
rect 9908 2843 9918 2877
rect 9952 2843 9962 2877
rect 9708 2703 9718 2737
rect 9752 2703 9762 2737
rect 9508 2563 9518 2597
rect 9552 2563 9562 2597
rect 9402 2499 9468 2500
rect 9402 2447 9409 2499
rect 9461 2447 9468 2499
rect 9402 2446 9468 2447
rect 9308 2333 9318 2367
rect 9352 2333 9362 2367
rect 9108 2193 9118 2227
rect 9152 2193 9162 2227
rect 8908 2053 8918 2087
rect 8952 2053 8962 2087
rect 8708 1913 8718 1947
rect 8752 1913 8762 1947
rect 8508 1773 8518 1807
rect 8552 1773 8562 1807
rect 8308 1633 8318 1667
rect 8352 1633 8362 1667
rect 8108 1493 8118 1527
rect 8152 1493 8162 1527
rect 7908 1353 7918 1387
rect 7952 1353 7962 1387
rect 7802 1289 7868 1290
rect 7802 1237 7809 1289
rect 7861 1237 7868 1289
rect 7802 1236 7868 1237
rect 7708 1123 7718 1157
rect 7752 1123 7762 1157
rect 7508 983 7518 1017
rect 7552 983 7562 1017
rect 7308 843 7318 877
rect 7352 843 7362 877
rect 7108 703 7118 737
rect 7152 703 7162 737
rect 6908 563 6918 597
rect 6952 563 6962 597
rect 6708 423 6718 457
rect 6752 423 6762 457
rect 6508 283 6518 317
rect 6552 283 6562 317
rect 6308 143 6318 177
rect 6352 143 6362 177
rect 6202 79 6268 80
rect 6202 27 6209 79
rect 6261 27 6268 79
rect 6202 26 6268 27
rect 6108 -67 6109 -15
rect 6161 -67 6162 -15
rect 6108 -79 6118 -67
rect 6152 -79 6162 -67
rect 5908 -132 5962 -131
rect 5908 -143 5918 -132
rect 5952 -143 5962 -132
rect 5908 -195 5909 -143
rect 5961 -195 5962 -143
rect 5908 -210 5962 -195
rect 6012 -133 6058 -81
rect 6012 -167 6018 -133
rect 6052 -167 6058 -133
rect 5918 -291 5925 -239
rect 5977 -291 5984 -239
rect 5812 -397 5818 -363
rect 5852 -397 5858 -363
rect 5812 -435 5858 -397
rect 5812 -469 5818 -435
rect 5852 -469 5858 -435
rect 5812 -512 5858 -469
rect 5909 -326 5961 -320
rect 5909 -390 5918 -378
rect 5952 -390 5961 -378
rect 5909 -454 5918 -442
rect 5952 -454 5961 -442
rect 5909 -555 5961 -506
rect 6012 -363 6058 -167
rect 6108 -131 6109 -79
rect 6161 -131 6162 -79
rect 6208 -22 6262 26
rect 6208 -74 6209 -22
rect 6261 -74 6262 -22
rect 6208 -81 6262 -74
rect 6308 -15 6362 143
rect 6408 177 6462 189
rect 6408 151 6418 177
rect 6452 151 6462 177
rect 6408 99 6409 151
rect 6461 99 6462 151
rect 6408 92 6462 99
rect 6508 177 6562 283
rect 6608 361 6662 368
rect 6608 309 6609 361
rect 6661 309 6662 361
rect 6608 283 6618 309
rect 6652 283 6662 309
rect 6608 271 6662 283
rect 6708 317 6762 423
rect 6808 457 6862 469
rect 6808 431 6818 457
rect 6852 431 6862 457
rect 6808 379 6809 431
rect 6861 379 6862 431
rect 6808 372 6862 379
rect 6908 457 6962 563
rect 7008 641 7062 648
rect 7008 589 7009 641
rect 7061 589 7062 641
rect 7008 563 7018 589
rect 7052 563 7062 589
rect 7008 551 7062 563
rect 7108 597 7162 703
rect 7208 737 7262 749
rect 7208 711 7218 737
rect 7252 711 7262 737
rect 7208 659 7209 711
rect 7261 659 7262 711
rect 7208 652 7262 659
rect 7308 737 7362 843
rect 7408 921 7462 928
rect 7408 869 7409 921
rect 7461 869 7462 921
rect 7408 843 7418 869
rect 7452 843 7462 869
rect 7408 831 7462 843
rect 7508 877 7562 983
rect 7608 1017 7662 1029
rect 7608 991 7618 1017
rect 7652 991 7662 1017
rect 7608 939 7609 991
rect 7661 939 7662 991
rect 7608 932 7662 939
rect 7708 1017 7762 1123
rect 7808 1201 7862 1208
rect 7808 1149 7809 1201
rect 7861 1149 7862 1201
rect 7808 1123 7818 1149
rect 7852 1123 7862 1149
rect 7808 1111 7862 1123
rect 7908 1157 7962 1353
rect 8008 1387 8062 1399
rect 8008 1361 8018 1387
rect 8052 1361 8062 1387
rect 8008 1309 8009 1361
rect 8061 1309 8062 1361
rect 8008 1302 8062 1309
rect 8108 1387 8162 1493
rect 8208 1571 8262 1578
rect 8208 1519 8209 1571
rect 8261 1519 8262 1571
rect 8208 1493 8218 1519
rect 8252 1493 8262 1519
rect 8208 1481 8262 1493
rect 8308 1527 8362 1633
rect 8408 1667 8462 1679
rect 8408 1641 8418 1667
rect 8452 1641 8462 1667
rect 8408 1589 8409 1641
rect 8461 1589 8462 1641
rect 8408 1582 8462 1589
rect 8508 1667 8562 1773
rect 8608 1851 8662 1858
rect 8608 1799 8609 1851
rect 8661 1799 8662 1851
rect 8608 1773 8618 1799
rect 8652 1773 8662 1799
rect 8608 1761 8662 1773
rect 8708 1807 8762 1913
rect 8808 1947 8862 1959
rect 8808 1921 8818 1947
rect 8852 1921 8862 1947
rect 8808 1869 8809 1921
rect 8861 1869 8862 1921
rect 8808 1862 8862 1869
rect 8908 1947 8962 2053
rect 9008 2131 9062 2138
rect 9008 2079 9009 2131
rect 9061 2079 9062 2131
rect 9008 2053 9018 2079
rect 9052 2053 9062 2079
rect 9008 2041 9062 2053
rect 9108 2087 9162 2193
rect 9208 2227 9262 2239
rect 9208 2201 9218 2227
rect 9252 2201 9262 2227
rect 9208 2149 9209 2201
rect 9261 2149 9262 2201
rect 9208 2142 9262 2149
rect 9308 2227 9362 2333
rect 9408 2411 9462 2418
rect 9408 2359 9409 2411
rect 9461 2359 9462 2411
rect 9408 2333 9418 2359
rect 9452 2333 9462 2359
rect 9408 2321 9462 2333
rect 9508 2367 9562 2563
rect 9608 2597 9662 2609
rect 9608 2571 9618 2597
rect 9652 2571 9662 2597
rect 9608 2519 9609 2571
rect 9661 2519 9662 2571
rect 9608 2512 9662 2519
rect 9708 2597 9762 2703
rect 9808 2781 9862 2788
rect 9808 2729 9809 2781
rect 9861 2729 9862 2781
rect 9808 2703 9818 2729
rect 9852 2703 9862 2729
rect 9808 2691 9862 2703
rect 9908 2737 9962 2843
rect 10008 2877 10062 2889
rect 10008 2851 10018 2877
rect 10052 2851 10062 2877
rect 10008 2799 10009 2851
rect 10061 2799 10062 2851
rect 10008 2792 10062 2799
rect 10108 2877 10162 2983
rect 10208 3061 10262 3068
rect 10208 3009 10209 3061
rect 10261 3009 10262 3061
rect 10208 2983 10218 3009
rect 10252 2983 10262 3009
rect 10208 2971 10262 2983
rect 10308 3017 10362 3123
rect 10408 3157 10462 3169
rect 10408 3131 10418 3157
rect 10452 3131 10462 3157
rect 10408 3079 10409 3131
rect 10461 3079 10462 3131
rect 10408 3072 10462 3079
rect 10508 3157 10562 3263
rect 10608 3341 10662 3348
rect 10608 3289 10609 3341
rect 10661 3289 10662 3341
rect 10608 3263 10618 3289
rect 10652 3263 10662 3289
rect 10608 3251 10662 3263
rect 10708 3297 10762 3403
rect 10808 3437 10862 3449
rect 10808 3411 10818 3437
rect 10852 3411 10862 3437
rect 10808 3359 10809 3411
rect 10861 3359 10862 3411
rect 10808 3352 10862 3359
rect 10908 3437 10962 3543
rect 11008 3621 11062 3628
rect 11008 3569 11009 3621
rect 11061 3569 11062 3621
rect 11008 3543 11018 3569
rect 11052 3543 11062 3569
rect 11008 3531 11062 3543
rect 11108 3577 11162 3773
rect 11208 3807 11262 3819
rect 11208 3781 11218 3807
rect 11252 3781 11262 3807
rect 11208 3729 11209 3781
rect 11261 3729 11262 3781
rect 11208 3722 11262 3729
rect 11308 3807 11362 3913
rect 11408 3991 11462 3998
rect 11408 3939 11409 3991
rect 11461 3939 11462 3991
rect 11408 3913 11418 3939
rect 11452 3913 11462 3939
rect 11408 3901 11462 3913
rect 11508 3947 11562 4053
rect 11608 4087 11662 4099
rect 11608 4061 11618 4087
rect 11652 4061 11662 4087
rect 11608 4009 11609 4061
rect 11661 4009 11662 4061
rect 11608 4002 11662 4009
rect 11708 4087 11762 4193
rect 11808 4271 11862 4278
rect 11808 4219 11809 4271
rect 11861 4219 11862 4271
rect 11808 4193 11818 4219
rect 11852 4193 11862 4219
rect 11808 4181 11862 4193
rect 11908 4227 11962 4333
rect 12008 4367 12062 4379
rect 12008 4341 12018 4367
rect 12052 4341 12062 4367
rect 12008 4289 12009 4341
rect 12061 4289 12062 4341
rect 12008 4282 12062 4289
rect 12108 4367 12162 4473
rect 12208 4551 12262 4558
rect 12208 4499 12209 4551
rect 12261 4499 12262 4551
rect 12208 4473 12218 4499
rect 12252 4473 12262 4499
rect 12208 4461 12262 4473
rect 12308 4507 12362 4613
rect 12408 4647 12462 4659
rect 12408 4621 12418 4647
rect 12452 4621 12462 4647
rect 12408 4569 12409 4621
rect 12461 4569 12462 4621
rect 12408 4562 12462 4569
rect 12508 4647 12562 4753
rect 12608 4831 12662 4838
rect 12608 4779 12609 4831
rect 12661 4779 12662 4831
rect 12608 4753 12618 4779
rect 12652 4753 12662 4779
rect 12608 4741 12662 4753
rect 12708 4787 12762 4960
rect 12990 4897 13020 5070
rect 12904 4891 13020 4897
rect 12904 4857 12916 4891
rect 12950 4857 13020 4891
rect 12904 4851 13020 4857
rect 12906 4802 12960 4814
rect 12708 4753 12718 4787
rect 12752 4753 12762 4787
rect 12508 4613 12518 4647
rect 12552 4613 12562 4647
rect 12308 4473 12318 4507
rect 12352 4473 12362 4507
rect 12108 4333 12118 4367
rect 12152 4333 12162 4367
rect 11908 4193 11918 4227
rect 11952 4193 11962 4227
rect 11708 4053 11718 4087
rect 11752 4053 11762 4087
rect 11508 3913 11518 3947
rect 11552 3913 11562 3947
rect 11308 3773 11318 3807
rect 11352 3773 11362 3807
rect 11202 3693 11268 3694
rect 11202 3641 11209 3693
rect 11261 3641 11268 3693
rect 11202 3640 11268 3641
rect 11108 3543 11118 3577
rect 11152 3543 11162 3577
rect 10908 3403 10918 3437
rect 10952 3403 10962 3437
rect 10708 3263 10718 3297
rect 10752 3263 10762 3297
rect 10508 3123 10518 3157
rect 10552 3123 10562 3157
rect 10308 2983 10318 3017
rect 10352 2983 10362 3017
rect 10108 2843 10118 2877
rect 10152 2843 10162 2877
rect 9908 2703 9918 2737
rect 9952 2703 9962 2737
rect 9708 2563 9718 2597
rect 9752 2563 9762 2597
rect 9602 2483 9668 2484
rect 9602 2431 9609 2483
rect 9661 2431 9668 2483
rect 9602 2430 9668 2431
rect 9508 2333 9518 2367
rect 9552 2333 9562 2367
rect 9308 2193 9318 2227
rect 9352 2193 9362 2227
rect 9108 2053 9118 2087
rect 9152 2053 9162 2087
rect 8908 1913 8918 1947
rect 8952 1913 8962 1947
rect 8708 1773 8718 1807
rect 8752 1773 8762 1807
rect 8508 1633 8518 1667
rect 8552 1633 8562 1667
rect 8308 1493 8318 1527
rect 8352 1493 8362 1527
rect 8108 1353 8118 1387
rect 8152 1353 8162 1387
rect 8002 1273 8068 1274
rect 8002 1221 8009 1273
rect 8061 1221 8068 1273
rect 8002 1220 8068 1221
rect 7908 1123 7918 1157
rect 7952 1123 7962 1157
rect 7708 983 7718 1017
rect 7752 983 7762 1017
rect 7508 843 7518 877
rect 7552 843 7562 877
rect 7308 703 7318 737
rect 7352 703 7362 737
rect 7108 563 7118 597
rect 7152 563 7162 597
rect 6908 423 6918 457
rect 6952 423 6962 457
rect 6708 283 6718 317
rect 6752 283 6762 317
rect 6508 143 6518 177
rect 6552 143 6562 177
rect 6402 63 6468 64
rect 6402 11 6409 63
rect 6461 11 6468 63
rect 6402 10 6468 11
rect 6308 -67 6309 -15
rect 6361 -67 6362 -15
rect 6308 -79 6318 -67
rect 6352 -79 6362 -67
rect 6108 -132 6162 -131
rect 6108 -143 6118 -132
rect 6152 -143 6162 -132
rect 6108 -195 6109 -143
rect 6161 -195 6162 -143
rect 6108 -210 6162 -195
rect 6212 -133 6258 -81
rect 6212 -167 6218 -133
rect 6252 -167 6258 -133
rect 6118 -291 6125 -239
rect 6177 -291 6184 -239
rect 6012 -397 6018 -363
rect 6052 -397 6058 -363
rect 6012 -435 6058 -397
rect 6012 -469 6018 -435
rect 6052 -469 6058 -435
rect 6012 -512 6058 -469
rect 6109 -326 6161 -320
rect 6109 -390 6118 -378
rect 6152 -390 6161 -378
rect 6109 -454 6118 -442
rect 6152 -454 6161 -442
rect 6109 -512 6161 -506
rect 6212 -363 6258 -167
rect 6308 -131 6309 -79
rect 6361 -131 6362 -79
rect 6408 -22 6462 10
rect 6408 -74 6409 -22
rect 6461 -74 6462 -22
rect 6408 -81 6462 -74
rect 6508 -15 6562 143
rect 6608 221 6662 228
rect 6608 169 6609 221
rect 6661 169 6662 221
rect 6608 143 6618 169
rect 6652 143 6662 169
rect 6608 131 6662 143
rect 6708 177 6762 283
rect 6808 317 6862 329
rect 6808 291 6818 317
rect 6852 291 6862 317
rect 6808 239 6809 291
rect 6861 239 6862 291
rect 6808 232 6862 239
rect 6908 317 6962 423
rect 7008 501 7062 508
rect 7008 449 7009 501
rect 7061 449 7062 501
rect 7008 423 7018 449
rect 7052 423 7062 449
rect 7008 411 7062 423
rect 7108 457 7162 563
rect 7208 597 7262 609
rect 7208 571 7218 597
rect 7252 571 7262 597
rect 7208 519 7209 571
rect 7261 519 7262 571
rect 7208 512 7262 519
rect 7308 597 7362 703
rect 7408 781 7462 788
rect 7408 729 7409 781
rect 7461 729 7462 781
rect 7408 703 7418 729
rect 7452 703 7462 729
rect 7408 691 7462 703
rect 7508 737 7562 843
rect 7608 877 7662 889
rect 7608 851 7618 877
rect 7652 851 7662 877
rect 7608 799 7609 851
rect 7661 799 7662 851
rect 7608 792 7662 799
rect 7708 877 7762 983
rect 7808 1061 7862 1068
rect 7808 1009 7809 1061
rect 7861 1009 7862 1061
rect 7808 983 7818 1009
rect 7852 983 7862 1009
rect 7808 971 7862 983
rect 7908 1017 7962 1123
rect 8008 1157 8062 1169
rect 8008 1131 8018 1157
rect 8052 1131 8062 1157
rect 8008 1079 8009 1131
rect 8061 1079 8062 1131
rect 8008 1072 8062 1079
rect 8108 1157 8162 1353
rect 8208 1431 8262 1438
rect 8208 1379 8209 1431
rect 8261 1379 8262 1431
rect 8208 1353 8218 1379
rect 8252 1353 8262 1379
rect 8208 1341 8262 1353
rect 8308 1387 8362 1493
rect 8408 1527 8462 1539
rect 8408 1501 8418 1527
rect 8452 1501 8462 1527
rect 8408 1449 8409 1501
rect 8461 1449 8462 1501
rect 8408 1442 8462 1449
rect 8508 1527 8562 1633
rect 8608 1711 8662 1718
rect 8608 1659 8609 1711
rect 8661 1659 8662 1711
rect 8608 1633 8618 1659
rect 8652 1633 8662 1659
rect 8608 1621 8662 1633
rect 8708 1667 8762 1773
rect 8808 1807 8862 1819
rect 8808 1781 8818 1807
rect 8852 1781 8862 1807
rect 8808 1729 8809 1781
rect 8861 1729 8862 1781
rect 8808 1722 8862 1729
rect 8908 1807 8962 1913
rect 9008 1991 9062 1998
rect 9008 1939 9009 1991
rect 9061 1939 9062 1991
rect 9008 1913 9018 1939
rect 9052 1913 9062 1939
rect 9008 1901 9062 1913
rect 9108 1947 9162 2053
rect 9208 2087 9262 2099
rect 9208 2061 9218 2087
rect 9252 2061 9262 2087
rect 9208 2009 9209 2061
rect 9261 2009 9262 2061
rect 9208 2002 9262 2009
rect 9308 2087 9362 2193
rect 9408 2271 9462 2278
rect 9408 2219 9409 2271
rect 9461 2219 9462 2271
rect 9408 2193 9418 2219
rect 9452 2193 9462 2219
rect 9408 2181 9462 2193
rect 9508 2227 9562 2333
rect 9608 2367 9662 2379
rect 9608 2341 9618 2367
rect 9652 2341 9662 2367
rect 9608 2289 9609 2341
rect 9661 2289 9662 2341
rect 9608 2282 9662 2289
rect 9708 2367 9762 2563
rect 9808 2641 9862 2648
rect 9808 2589 9809 2641
rect 9861 2589 9862 2641
rect 9808 2563 9818 2589
rect 9852 2563 9862 2589
rect 9808 2551 9862 2563
rect 9908 2597 9962 2703
rect 10008 2737 10062 2749
rect 10008 2711 10018 2737
rect 10052 2711 10062 2737
rect 10008 2659 10009 2711
rect 10061 2659 10062 2711
rect 10008 2652 10062 2659
rect 10108 2737 10162 2843
rect 10208 2921 10262 2928
rect 10208 2869 10209 2921
rect 10261 2869 10262 2921
rect 10208 2843 10218 2869
rect 10252 2843 10262 2869
rect 10208 2831 10262 2843
rect 10308 2877 10362 2983
rect 10408 3017 10462 3029
rect 10408 2991 10418 3017
rect 10452 2991 10462 3017
rect 10408 2939 10409 2991
rect 10461 2939 10462 2991
rect 10408 2932 10462 2939
rect 10508 3017 10562 3123
rect 10608 3201 10662 3208
rect 10608 3149 10609 3201
rect 10661 3149 10662 3201
rect 10608 3123 10618 3149
rect 10652 3123 10662 3149
rect 10608 3111 10662 3123
rect 10708 3157 10762 3263
rect 10808 3297 10862 3309
rect 10808 3271 10818 3297
rect 10852 3271 10862 3297
rect 10808 3219 10809 3271
rect 10861 3219 10862 3271
rect 10808 3212 10862 3219
rect 10908 3297 10962 3403
rect 11008 3481 11062 3488
rect 11008 3429 11009 3481
rect 11061 3429 11062 3481
rect 11008 3403 11018 3429
rect 11052 3403 11062 3429
rect 11008 3391 11062 3403
rect 11108 3437 11162 3543
rect 11208 3577 11262 3589
rect 11208 3551 11218 3577
rect 11252 3551 11262 3577
rect 11208 3499 11209 3551
rect 11261 3499 11262 3551
rect 11208 3492 11262 3499
rect 11308 3577 11362 3773
rect 11408 3851 11462 3858
rect 11408 3799 11409 3851
rect 11461 3799 11462 3851
rect 11408 3773 11418 3799
rect 11452 3773 11462 3799
rect 11408 3761 11462 3773
rect 11508 3807 11562 3913
rect 11608 3947 11662 3959
rect 11608 3921 11618 3947
rect 11652 3921 11662 3947
rect 11608 3869 11609 3921
rect 11661 3869 11662 3921
rect 11608 3862 11662 3869
rect 11708 3947 11762 4053
rect 11808 4131 11862 4138
rect 11808 4079 11809 4131
rect 11861 4079 11862 4131
rect 11808 4053 11818 4079
rect 11852 4053 11862 4079
rect 11808 4041 11862 4053
rect 11908 4087 11962 4193
rect 12008 4227 12062 4239
rect 12008 4201 12018 4227
rect 12052 4201 12062 4227
rect 12008 4149 12009 4201
rect 12061 4149 12062 4201
rect 12008 4142 12062 4149
rect 12108 4227 12162 4333
rect 12208 4411 12262 4418
rect 12208 4359 12209 4411
rect 12261 4359 12262 4411
rect 12208 4333 12218 4359
rect 12252 4333 12262 4359
rect 12208 4321 12262 4333
rect 12308 4367 12362 4473
rect 12408 4507 12462 4519
rect 12408 4481 12418 4507
rect 12452 4481 12462 4507
rect 12408 4429 12409 4481
rect 12461 4429 12462 4481
rect 12408 4422 12462 4429
rect 12508 4507 12562 4613
rect 12608 4691 12662 4698
rect 12608 4639 12609 4691
rect 12661 4639 12662 4691
rect 12608 4613 12618 4639
rect 12652 4613 12662 4639
rect 12608 4601 12662 4613
rect 12708 4647 12762 4753
rect 12808 4787 12862 4799
rect 12808 4761 12818 4787
rect 12852 4761 12862 4787
rect 12808 4709 12809 4761
rect 12861 4709 12862 4761
rect 12808 4702 12862 4709
rect 12906 4768 12916 4802
rect 12950 4768 12960 4802
rect 12906 4761 12960 4768
rect 12906 4709 12907 4761
rect 12959 4709 12960 4761
rect 12906 4702 12960 4709
rect 12906 4662 12960 4674
rect 12708 4613 12718 4647
rect 12752 4613 12762 4647
rect 12508 4473 12518 4507
rect 12552 4473 12562 4507
rect 12308 4333 12318 4367
rect 12352 4333 12362 4367
rect 12108 4193 12118 4227
rect 12152 4193 12162 4227
rect 11908 4053 11918 4087
rect 11952 4053 11962 4087
rect 11708 3913 11718 3947
rect 11752 3913 11762 3947
rect 11508 3773 11518 3807
rect 11552 3773 11562 3807
rect 11402 3709 11468 3710
rect 11402 3657 11409 3709
rect 11461 3657 11468 3709
rect 11402 3656 11468 3657
rect 11308 3543 11318 3577
rect 11352 3543 11362 3577
rect 11108 3403 11118 3437
rect 11152 3403 11162 3437
rect 10908 3263 10918 3297
rect 10952 3263 10962 3297
rect 10708 3123 10718 3157
rect 10752 3123 10762 3157
rect 10508 2983 10518 3017
rect 10552 2983 10562 3017
rect 10308 2843 10318 2877
rect 10352 2843 10362 2877
rect 10108 2703 10118 2737
rect 10152 2703 10162 2737
rect 9908 2563 9918 2597
rect 9952 2563 9962 2597
rect 9802 2499 9868 2500
rect 9802 2447 9809 2499
rect 9861 2447 9868 2499
rect 9802 2446 9868 2447
rect 9708 2333 9718 2367
rect 9752 2333 9762 2367
rect 9508 2193 9518 2227
rect 9552 2193 9562 2227
rect 9308 2053 9318 2087
rect 9352 2053 9362 2087
rect 9108 1913 9118 1947
rect 9152 1913 9162 1947
rect 8908 1773 8918 1807
rect 8952 1773 8962 1807
rect 8708 1633 8718 1667
rect 8752 1633 8762 1667
rect 8508 1493 8518 1527
rect 8552 1493 8562 1527
rect 8308 1353 8318 1387
rect 8352 1353 8362 1387
rect 8202 1289 8268 1290
rect 8202 1237 8209 1289
rect 8261 1237 8268 1289
rect 8202 1236 8268 1237
rect 8108 1123 8118 1157
rect 8152 1123 8162 1157
rect 7908 983 7918 1017
rect 7952 983 7962 1017
rect 7708 843 7718 877
rect 7752 843 7762 877
rect 7508 703 7518 737
rect 7552 703 7562 737
rect 7308 563 7318 597
rect 7352 563 7362 597
rect 7108 423 7118 457
rect 7152 423 7162 457
rect 6908 283 6918 317
rect 6952 283 6962 317
rect 6708 143 6718 177
rect 6752 143 6762 177
rect 6602 79 6668 80
rect 6602 27 6609 79
rect 6661 27 6668 79
rect 6602 26 6668 27
rect 6508 -67 6509 -15
rect 6561 -67 6562 -15
rect 6508 -79 6518 -67
rect 6552 -79 6562 -67
rect 6308 -132 6362 -131
rect 6308 -143 6318 -132
rect 6352 -143 6362 -132
rect 6308 -195 6309 -143
rect 6361 -195 6362 -143
rect 6308 -210 6362 -195
rect 6412 -133 6458 -81
rect 6412 -167 6418 -133
rect 6452 -167 6458 -133
rect 6318 -291 6325 -239
rect 6377 -291 6384 -239
rect 6212 -397 6218 -363
rect 6252 -397 6258 -363
rect 6212 -435 6258 -397
rect 6212 -469 6218 -435
rect 6252 -469 6258 -435
rect 6212 -512 6258 -469
rect 6309 -326 6361 -320
rect 6309 -390 6318 -378
rect 6352 -390 6361 -378
rect 6309 -454 6318 -442
rect 6352 -454 6361 -442
rect 6309 -555 6361 -506
rect 6412 -363 6458 -167
rect 6508 -131 6509 -79
rect 6561 -131 6562 -79
rect 6608 -22 6662 26
rect 6608 -74 6609 -22
rect 6661 -74 6662 -22
rect 6608 -81 6662 -74
rect 6708 -15 6762 143
rect 6808 177 6862 189
rect 6808 151 6818 177
rect 6852 151 6862 177
rect 6808 99 6809 151
rect 6861 99 6862 151
rect 6808 92 6862 99
rect 6908 177 6962 283
rect 7008 361 7062 368
rect 7008 309 7009 361
rect 7061 309 7062 361
rect 7008 283 7018 309
rect 7052 283 7062 309
rect 7008 271 7062 283
rect 7108 317 7162 423
rect 7208 457 7262 469
rect 7208 431 7218 457
rect 7252 431 7262 457
rect 7208 379 7209 431
rect 7261 379 7262 431
rect 7208 372 7262 379
rect 7308 457 7362 563
rect 7408 641 7462 648
rect 7408 589 7409 641
rect 7461 589 7462 641
rect 7408 563 7418 589
rect 7452 563 7462 589
rect 7408 551 7462 563
rect 7508 597 7562 703
rect 7608 737 7662 749
rect 7608 711 7618 737
rect 7652 711 7662 737
rect 7608 659 7609 711
rect 7661 659 7662 711
rect 7608 652 7662 659
rect 7708 737 7762 843
rect 7808 921 7862 928
rect 7808 869 7809 921
rect 7861 869 7862 921
rect 7808 843 7818 869
rect 7852 843 7862 869
rect 7808 831 7862 843
rect 7908 877 7962 983
rect 8008 1017 8062 1029
rect 8008 991 8018 1017
rect 8052 991 8062 1017
rect 8008 939 8009 991
rect 8061 939 8062 991
rect 8008 932 8062 939
rect 8108 1017 8162 1123
rect 8208 1201 8262 1208
rect 8208 1149 8209 1201
rect 8261 1149 8262 1201
rect 8208 1123 8218 1149
rect 8252 1123 8262 1149
rect 8208 1111 8262 1123
rect 8308 1157 8362 1353
rect 8408 1387 8462 1399
rect 8408 1361 8418 1387
rect 8452 1361 8462 1387
rect 8408 1309 8409 1361
rect 8461 1309 8462 1361
rect 8408 1302 8462 1309
rect 8508 1387 8562 1493
rect 8608 1571 8662 1578
rect 8608 1519 8609 1571
rect 8661 1519 8662 1571
rect 8608 1493 8618 1519
rect 8652 1493 8662 1519
rect 8608 1481 8662 1493
rect 8708 1527 8762 1633
rect 8808 1667 8862 1679
rect 8808 1641 8818 1667
rect 8852 1641 8862 1667
rect 8808 1589 8809 1641
rect 8861 1589 8862 1641
rect 8808 1582 8862 1589
rect 8908 1667 8962 1773
rect 9008 1851 9062 1858
rect 9008 1799 9009 1851
rect 9061 1799 9062 1851
rect 9008 1773 9018 1799
rect 9052 1773 9062 1799
rect 9008 1761 9062 1773
rect 9108 1807 9162 1913
rect 9208 1947 9262 1959
rect 9208 1921 9218 1947
rect 9252 1921 9262 1947
rect 9208 1869 9209 1921
rect 9261 1869 9262 1921
rect 9208 1862 9262 1869
rect 9308 1947 9362 2053
rect 9408 2131 9462 2138
rect 9408 2079 9409 2131
rect 9461 2079 9462 2131
rect 9408 2053 9418 2079
rect 9452 2053 9462 2079
rect 9408 2041 9462 2053
rect 9508 2087 9562 2193
rect 9608 2227 9662 2239
rect 9608 2201 9618 2227
rect 9652 2201 9662 2227
rect 9608 2149 9609 2201
rect 9661 2149 9662 2201
rect 9608 2142 9662 2149
rect 9708 2227 9762 2333
rect 9808 2411 9862 2418
rect 9808 2359 9809 2411
rect 9861 2359 9862 2411
rect 9808 2333 9818 2359
rect 9852 2333 9862 2359
rect 9808 2321 9862 2333
rect 9908 2367 9962 2563
rect 10008 2597 10062 2609
rect 10008 2571 10018 2597
rect 10052 2571 10062 2597
rect 10008 2519 10009 2571
rect 10061 2519 10062 2571
rect 10008 2512 10062 2519
rect 10108 2597 10162 2703
rect 10208 2781 10262 2788
rect 10208 2729 10209 2781
rect 10261 2729 10262 2781
rect 10208 2703 10218 2729
rect 10252 2703 10262 2729
rect 10208 2691 10262 2703
rect 10308 2737 10362 2843
rect 10408 2877 10462 2889
rect 10408 2851 10418 2877
rect 10452 2851 10462 2877
rect 10408 2799 10409 2851
rect 10461 2799 10462 2851
rect 10408 2792 10462 2799
rect 10508 2877 10562 2983
rect 10608 3061 10662 3068
rect 10608 3009 10609 3061
rect 10661 3009 10662 3061
rect 10608 2983 10618 3009
rect 10652 2983 10662 3009
rect 10608 2971 10662 2983
rect 10708 3017 10762 3123
rect 10808 3157 10862 3169
rect 10808 3131 10818 3157
rect 10852 3131 10862 3157
rect 10808 3079 10809 3131
rect 10861 3079 10862 3131
rect 10808 3072 10862 3079
rect 10908 3157 10962 3263
rect 11008 3341 11062 3348
rect 11008 3289 11009 3341
rect 11061 3289 11062 3341
rect 11008 3263 11018 3289
rect 11052 3263 11062 3289
rect 11008 3251 11062 3263
rect 11108 3297 11162 3403
rect 11208 3437 11262 3449
rect 11208 3411 11218 3437
rect 11252 3411 11262 3437
rect 11208 3359 11209 3411
rect 11261 3359 11262 3411
rect 11208 3352 11262 3359
rect 11308 3437 11362 3543
rect 11408 3621 11462 3628
rect 11408 3569 11409 3621
rect 11461 3569 11462 3621
rect 11408 3543 11418 3569
rect 11452 3543 11462 3569
rect 11408 3531 11462 3543
rect 11508 3577 11562 3773
rect 11608 3807 11662 3819
rect 11608 3781 11618 3807
rect 11652 3781 11662 3807
rect 11608 3729 11609 3781
rect 11661 3729 11662 3781
rect 11608 3722 11662 3729
rect 11708 3807 11762 3913
rect 11808 3991 11862 3998
rect 11808 3939 11809 3991
rect 11861 3939 11862 3991
rect 11808 3913 11818 3939
rect 11852 3913 11862 3939
rect 11808 3901 11862 3913
rect 11908 3947 11962 4053
rect 12008 4087 12062 4099
rect 12008 4061 12018 4087
rect 12052 4061 12062 4087
rect 12008 4009 12009 4061
rect 12061 4009 12062 4061
rect 12008 4002 12062 4009
rect 12108 4087 12162 4193
rect 12208 4271 12262 4278
rect 12208 4219 12209 4271
rect 12261 4219 12262 4271
rect 12208 4193 12218 4219
rect 12252 4193 12262 4219
rect 12208 4181 12262 4193
rect 12308 4227 12362 4333
rect 12408 4367 12462 4379
rect 12408 4341 12418 4367
rect 12452 4341 12462 4367
rect 12408 4289 12409 4341
rect 12461 4289 12462 4341
rect 12408 4282 12462 4289
rect 12508 4367 12562 4473
rect 12608 4551 12662 4558
rect 12608 4499 12609 4551
rect 12661 4499 12662 4551
rect 12608 4473 12618 4499
rect 12652 4473 12662 4499
rect 12608 4461 12662 4473
rect 12708 4507 12762 4613
rect 12808 4647 12862 4659
rect 12808 4621 12818 4647
rect 12852 4621 12862 4647
rect 12808 4569 12809 4621
rect 12861 4569 12862 4621
rect 12808 4562 12862 4569
rect 12906 4628 12916 4662
rect 12950 4628 12960 4662
rect 12906 4621 12960 4628
rect 12906 4569 12907 4621
rect 12959 4569 12960 4621
rect 12906 4562 12960 4569
rect 12906 4522 12960 4534
rect 12708 4473 12718 4507
rect 12752 4473 12762 4507
rect 12508 4333 12518 4367
rect 12552 4333 12562 4367
rect 12308 4193 12318 4227
rect 12352 4193 12362 4227
rect 12108 4053 12118 4087
rect 12152 4053 12162 4087
rect 11908 3913 11918 3947
rect 11952 3913 11962 3947
rect 11708 3773 11718 3807
rect 11752 3773 11762 3807
rect 11602 3693 11668 3694
rect 11602 3641 11609 3693
rect 11661 3641 11668 3693
rect 11602 3640 11668 3641
rect 11508 3543 11518 3577
rect 11552 3543 11562 3577
rect 11308 3403 11318 3437
rect 11352 3403 11362 3437
rect 11108 3263 11118 3297
rect 11152 3263 11162 3297
rect 10908 3123 10918 3157
rect 10952 3123 10962 3157
rect 10708 2983 10718 3017
rect 10752 2983 10762 3017
rect 10508 2843 10518 2877
rect 10552 2843 10562 2877
rect 10308 2703 10318 2737
rect 10352 2703 10362 2737
rect 10108 2563 10118 2597
rect 10152 2563 10162 2597
rect 10002 2483 10068 2484
rect 10002 2431 10009 2483
rect 10061 2431 10068 2483
rect 10002 2430 10068 2431
rect 9908 2333 9918 2367
rect 9952 2333 9962 2367
rect 9708 2193 9718 2227
rect 9752 2193 9762 2227
rect 9508 2053 9518 2087
rect 9552 2053 9562 2087
rect 9308 1913 9318 1947
rect 9352 1913 9362 1947
rect 9108 1773 9118 1807
rect 9152 1773 9162 1807
rect 8908 1633 8918 1667
rect 8952 1633 8962 1667
rect 8708 1493 8718 1527
rect 8752 1493 8762 1527
rect 8508 1353 8518 1387
rect 8552 1353 8562 1387
rect 8402 1273 8468 1274
rect 8402 1221 8409 1273
rect 8461 1221 8468 1273
rect 8402 1220 8468 1221
rect 8308 1123 8318 1157
rect 8352 1123 8362 1157
rect 8108 983 8118 1017
rect 8152 983 8162 1017
rect 7908 843 7918 877
rect 7952 843 7962 877
rect 7708 703 7718 737
rect 7752 703 7762 737
rect 7508 563 7518 597
rect 7552 563 7562 597
rect 7308 423 7318 457
rect 7352 423 7362 457
rect 7108 283 7118 317
rect 7152 283 7162 317
rect 6908 143 6918 177
rect 6952 143 6962 177
rect 6802 63 6868 64
rect 6802 11 6809 63
rect 6861 11 6868 63
rect 6802 10 6868 11
rect 6708 -67 6709 -15
rect 6761 -67 6762 -15
rect 6708 -79 6718 -67
rect 6752 -79 6762 -67
rect 6508 -132 6562 -131
rect 6508 -143 6518 -132
rect 6552 -143 6562 -132
rect 6508 -195 6509 -143
rect 6561 -195 6562 -143
rect 6508 -210 6562 -195
rect 6612 -133 6658 -81
rect 6612 -167 6618 -133
rect 6652 -167 6658 -133
rect 6518 -291 6525 -239
rect 6577 -291 6584 -239
rect 6412 -397 6418 -363
rect 6452 -397 6458 -363
rect 6412 -435 6458 -397
rect 6412 -469 6418 -435
rect 6452 -469 6458 -435
rect 6412 -512 6458 -469
rect 6509 -326 6561 -320
rect 6509 -390 6518 -378
rect 6552 -390 6561 -378
rect 6509 -454 6518 -442
rect 6552 -454 6561 -442
rect 6509 -512 6561 -506
rect 6612 -363 6658 -167
rect 6708 -131 6709 -79
rect 6761 -131 6762 -79
rect 6808 -22 6862 10
rect 6808 -74 6809 -22
rect 6861 -74 6862 -22
rect 6808 -81 6862 -74
rect 6908 -15 6962 143
rect 7008 221 7062 228
rect 7008 169 7009 221
rect 7061 169 7062 221
rect 7008 143 7018 169
rect 7052 143 7062 169
rect 7008 131 7062 143
rect 7108 177 7162 283
rect 7208 317 7262 329
rect 7208 291 7218 317
rect 7252 291 7262 317
rect 7208 239 7209 291
rect 7261 239 7262 291
rect 7208 232 7262 239
rect 7308 317 7362 423
rect 7408 501 7462 508
rect 7408 449 7409 501
rect 7461 449 7462 501
rect 7408 423 7418 449
rect 7452 423 7462 449
rect 7408 411 7462 423
rect 7508 457 7562 563
rect 7608 597 7662 609
rect 7608 571 7618 597
rect 7652 571 7662 597
rect 7608 519 7609 571
rect 7661 519 7662 571
rect 7608 512 7662 519
rect 7708 597 7762 703
rect 7808 781 7862 788
rect 7808 729 7809 781
rect 7861 729 7862 781
rect 7808 703 7818 729
rect 7852 703 7862 729
rect 7808 691 7862 703
rect 7908 737 7962 843
rect 8008 877 8062 889
rect 8008 851 8018 877
rect 8052 851 8062 877
rect 8008 799 8009 851
rect 8061 799 8062 851
rect 8008 792 8062 799
rect 8108 877 8162 983
rect 8208 1061 8262 1068
rect 8208 1009 8209 1061
rect 8261 1009 8262 1061
rect 8208 983 8218 1009
rect 8252 983 8262 1009
rect 8208 971 8262 983
rect 8308 1017 8362 1123
rect 8408 1157 8462 1169
rect 8408 1131 8418 1157
rect 8452 1131 8462 1157
rect 8408 1079 8409 1131
rect 8461 1079 8462 1131
rect 8408 1072 8462 1079
rect 8508 1157 8562 1353
rect 8608 1431 8662 1438
rect 8608 1379 8609 1431
rect 8661 1379 8662 1431
rect 8608 1353 8618 1379
rect 8652 1353 8662 1379
rect 8608 1341 8662 1353
rect 8708 1387 8762 1493
rect 8808 1527 8862 1539
rect 8808 1501 8818 1527
rect 8852 1501 8862 1527
rect 8808 1449 8809 1501
rect 8861 1449 8862 1501
rect 8808 1442 8862 1449
rect 8908 1527 8962 1633
rect 9008 1711 9062 1718
rect 9008 1659 9009 1711
rect 9061 1659 9062 1711
rect 9008 1633 9018 1659
rect 9052 1633 9062 1659
rect 9008 1621 9062 1633
rect 9108 1667 9162 1773
rect 9208 1807 9262 1819
rect 9208 1781 9218 1807
rect 9252 1781 9262 1807
rect 9208 1729 9209 1781
rect 9261 1729 9262 1781
rect 9208 1722 9262 1729
rect 9308 1807 9362 1913
rect 9408 1991 9462 1998
rect 9408 1939 9409 1991
rect 9461 1939 9462 1991
rect 9408 1913 9418 1939
rect 9452 1913 9462 1939
rect 9408 1901 9462 1913
rect 9508 1947 9562 2053
rect 9608 2087 9662 2099
rect 9608 2061 9618 2087
rect 9652 2061 9662 2087
rect 9608 2009 9609 2061
rect 9661 2009 9662 2061
rect 9608 2002 9662 2009
rect 9708 2087 9762 2193
rect 9808 2271 9862 2278
rect 9808 2219 9809 2271
rect 9861 2219 9862 2271
rect 9808 2193 9818 2219
rect 9852 2193 9862 2219
rect 9808 2181 9862 2193
rect 9908 2227 9962 2333
rect 10008 2367 10062 2379
rect 10008 2341 10018 2367
rect 10052 2341 10062 2367
rect 10008 2289 10009 2341
rect 10061 2289 10062 2341
rect 10008 2282 10062 2289
rect 10108 2367 10162 2563
rect 10208 2641 10262 2648
rect 10208 2589 10209 2641
rect 10261 2589 10262 2641
rect 10208 2563 10218 2589
rect 10252 2563 10262 2589
rect 10208 2551 10262 2563
rect 10308 2597 10362 2703
rect 10408 2737 10462 2749
rect 10408 2711 10418 2737
rect 10452 2711 10462 2737
rect 10408 2659 10409 2711
rect 10461 2659 10462 2711
rect 10408 2652 10462 2659
rect 10508 2737 10562 2843
rect 10608 2921 10662 2928
rect 10608 2869 10609 2921
rect 10661 2869 10662 2921
rect 10608 2843 10618 2869
rect 10652 2843 10662 2869
rect 10608 2831 10662 2843
rect 10708 2877 10762 2983
rect 10808 3017 10862 3029
rect 10808 2991 10818 3017
rect 10852 2991 10862 3017
rect 10808 2939 10809 2991
rect 10861 2939 10862 2991
rect 10808 2932 10862 2939
rect 10908 3017 10962 3123
rect 11008 3201 11062 3208
rect 11008 3149 11009 3201
rect 11061 3149 11062 3201
rect 11008 3123 11018 3149
rect 11052 3123 11062 3149
rect 11008 3111 11062 3123
rect 11108 3157 11162 3263
rect 11208 3297 11262 3309
rect 11208 3271 11218 3297
rect 11252 3271 11262 3297
rect 11208 3219 11209 3271
rect 11261 3219 11262 3271
rect 11208 3212 11262 3219
rect 11308 3297 11362 3403
rect 11408 3481 11462 3488
rect 11408 3429 11409 3481
rect 11461 3429 11462 3481
rect 11408 3403 11418 3429
rect 11452 3403 11462 3429
rect 11408 3391 11462 3403
rect 11508 3437 11562 3543
rect 11608 3577 11662 3589
rect 11608 3551 11618 3577
rect 11652 3551 11662 3577
rect 11608 3499 11609 3551
rect 11661 3499 11662 3551
rect 11608 3492 11662 3499
rect 11708 3577 11762 3773
rect 11808 3851 11862 3858
rect 11808 3799 11809 3851
rect 11861 3799 11862 3851
rect 11808 3773 11818 3799
rect 11852 3773 11862 3799
rect 11808 3761 11862 3773
rect 11908 3807 11962 3913
rect 12008 3947 12062 3959
rect 12008 3921 12018 3947
rect 12052 3921 12062 3947
rect 12008 3869 12009 3921
rect 12061 3869 12062 3921
rect 12008 3862 12062 3869
rect 12108 3947 12162 4053
rect 12208 4131 12262 4138
rect 12208 4079 12209 4131
rect 12261 4079 12262 4131
rect 12208 4053 12218 4079
rect 12252 4053 12262 4079
rect 12208 4041 12262 4053
rect 12308 4087 12362 4193
rect 12408 4227 12462 4239
rect 12408 4201 12418 4227
rect 12452 4201 12462 4227
rect 12408 4149 12409 4201
rect 12461 4149 12462 4201
rect 12408 4142 12462 4149
rect 12508 4227 12562 4333
rect 12608 4411 12662 4418
rect 12608 4359 12609 4411
rect 12661 4359 12662 4411
rect 12608 4333 12618 4359
rect 12652 4333 12662 4359
rect 12608 4321 12662 4333
rect 12708 4367 12762 4473
rect 12808 4507 12862 4519
rect 12808 4481 12818 4507
rect 12852 4481 12862 4507
rect 12808 4429 12809 4481
rect 12861 4429 12862 4481
rect 12808 4422 12862 4429
rect 12906 4488 12916 4522
rect 12950 4488 12960 4522
rect 12906 4481 12960 4488
rect 12906 4429 12907 4481
rect 12959 4429 12960 4481
rect 12906 4422 12960 4429
rect 12906 4382 12960 4394
rect 12708 4333 12718 4367
rect 12752 4333 12762 4367
rect 12508 4193 12518 4227
rect 12552 4193 12562 4227
rect 12308 4053 12318 4087
rect 12352 4053 12362 4087
rect 12108 3913 12118 3947
rect 12152 3913 12162 3947
rect 11908 3773 11918 3807
rect 11952 3773 11962 3807
rect 11802 3709 11868 3710
rect 11802 3657 11809 3709
rect 11861 3657 11868 3709
rect 11802 3656 11868 3657
rect 11708 3543 11718 3577
rect 11752 3543 11762 3577
rect 11508 3403 11518 3437
rect 11552 3403 11562 3437
rect 11308 3263 11318 3297
rect 11352 3263 11362 3297
rect 11108 3123 11118 3157
rect 11152 3123 11162 3157
rect 10908 2983 10918 3017
rect 10952 2983 10962 3017
rect 10708 2843 10718 2877
rect 10752 2843 10762 2877
rect 10508 2703 10518 2737
rect 10552 2703 10562 2737
rect 10308 2563 10318 2597
rect 10352 2563 10362 2597
rect 10202 2499 10268 2500
rect 10202 2447 10209 2499
rect 10261 2447 10268 2499
rect 10202 2446 10268 2447
rect 10108 2333 10118 2367
rect 10152 2333 10162 2367
rect 9908 2193 9918 2227
rect 9952 2193 9962 2227
rect 9708 2053 9718 2087
rect 9752 2053 9762 2087
rect 9508 1913 9518 1947
rect 9552 1913 9562 1947
rect 9308 1773 9318 1807
rect 9352 1773 9362 1807
rect 9108 1633 9118 1667
rect 9152 1633 9162 1667
rect 8908 1493 8918 1527
rect 8952 1493 8962 1527
rect 8708 1353 8718 1387
rect 8752 1353 8762 1387
rect 8602 1289 8668 1290
rect 8602 1237 8609 1289
rect 8661 1237 8668 1289
rect 8602 1236 8668 1237
rect 8508 1123 8518 1157
rect 8552 1123 8562 1157
rect 8308 983 8318 1017
rect 8352 983 8362 1017
rect 8108 843 8118 877
rect 8152 843 8162 877
rect 7908 703 7918 737
rect 7952 703 7962 737
rect 7708 563 7718 597
rect 7752 563 7762 597
rect 7508 423 7518 457
rect 7552 423 7562 457
rect 7308 283 7318 317
rect 7352 283 7362 317
rect 7108 143 7118 177
rect 7152 143 7162 177
rect 7002 79 7068 80
rect 7002 27 7009 79
rect 7061 27 7068 79
rect 7002 26 7068 27
rect 6908 -67 6909 -15
rect 6961 -67 6962 -15
rect 6908 -79 6918 -67
rect 6952 -79 6962 -67
rect 6708 -132 6762 -131
rect 6708 -143 6718 -132
rect 6752 -143 6762 -132
rect 6708 -195 6709 -143
rect 6761 -195 6762 -143
rect 6708 -210 6762 -195
rect 6812 -133 6858 -81
rect 6812 -167 6818 -133
rect 6852 -167 6858 -133
rect 6718 -291 6725 -239
rect 6777 -291 6784 -239
rect 6612 -397 6618 -363
rect 6652 -397 6658 -363
rect 6612 -435 6658 -397
rect 6612 -469 6618 -435
rect 6652 -469 6658 -435
rect 6612 -512 6658 -469
rect 6709 -326 6761 -320
rect 6709 -390 6718 -378
rect 6752 -390 6761 -378
rect 6709 -454 6718 -442
rect 6752 -454 6761 -442
rect 6709 -555 6761 -506
rect 6812 -363 6858 -167
rect 6908 -131 6909 -79
rect 6961 -131 6962 -79
rect 7008 -22 7062 26
rect 7008 -74 7009 -22
rect 7061 -74 7062 -22
rect 7008 -81 7062 -74
rect 7108 -15 7162 143
rect 7208 177 7262 189
rect 7208 151 7218 177
rect 7252 151 7262 177
rect 7208 99 7209 151
rect 7261 99 7262 151
rect 7208 92 7262 99
rect 7308 177 7362 283
rect 7408 361 7462 368
rect 7408 309 7409 361
rect 7461 309 7462 361
rect 7408 283 7418 309
rect 7452 283 7462 309
rect 7408 271 7462 283
rect 7508 317 7562 423
rect 7608 457 7662 469
rect 7608 431 7618 457
rect 7652 431 7662 457
rect 7608 379 7609 431
rect 7661 379 7662 431
rect 7608 372 7662 379
rect 7708 457 7762 563
rect 7808 641 7862 648
rect 7808 589 7809 641
rect 7861 589 7862 641
rect 7808 563 7818 589
rect 7852 563 7862 589
rect 7808 551 7862 563
rect 7908 597 7962 703
rect 8008 737 8062 749
rect 8008 711 8018 737
rect 8052 711 8062 737
rect 8008 659 8009 711
rect 8061 659 8062 711
rect 8008 652 8062 659
rect 8108 737 8162 843
rect 8208 921 8262 928
rect 8208 869 8209 921
rect 8261 869 8262 921
rect 8208 843 8218 869
rect 8252 843 8262 869
rect 8208 831 8262 843
rect 8308 877 8362 983
rect 8408 1017 8462 1029
rect 8408 991 8418 1017
rect 8452 991 8462 1017
rect 8408 939 8409 991
rect 8461 939 8462 991
rect 8408 932 8462 939
rect 8508 1017 8562 1123
rect 8608 1201 8662 1208
rect 8608 1149 8609 1201
rect 8661 1149 8662 1201
rect 8608 1123 8618 1149
rect 8652 1123 8662 1149
rect 8608 1111 8662 1123
rect 8708 1157 8762 1353
rect 8808 1387 8862 1399
rect 8808 1361 8818 1387
rect 8852 1361 8862 1387
rect 8808 1309 8809 1361
rect 8861 1309 8862 1361
rect 8808 1302 8862 1309
rect 8908 1387 8962 1493
rect 9008 1571 9062 1578
rect 9008 1519 9009 1571
rect 9061 1519 9062 1571
rect 9008 1493 9018 1519
rect 9052 1493 9062 1519
rect 9008 1481 9062 1493
rect 9108 1527 9162 1633
rect 9208 1667 9262 1679
rect 9208 1641 9218 1667
rect 9252 1641 9262 1667
rect 9208 1589 9209 1641
rect 9261 1589 9262 1641
rect 9208 1582 9262 1589
rect 9308 1667 9362 1773
rect 9408 1851 9462 1858
rect 9408 1799 9409 1851
rect 9461 1799 9462 1851
rect 9408 1773 9418 1799
rect 9452 1773 9462 1799
rect 9408 1761 9462 1773
rect 9508 1807 9562 1913
rect 9608 1947 9662 1959
rect 9608 1921 9618 1947
rect 9652 1921 9662 1947
rect 9608 1869 9609 1921
rect 9661 1869 9662 1921
rect 9608 1862 9662 1869
rect 9708 1947 9762 2053
rect 9808 2131 9862 2138
rect 9808 2079 9809 2131
rect 9861 2079 9862 2131
rect 9808 2053 9818 2079
rect 9852 2053 9862 2079
rect 9808 2041 9862 2053
rect 9908 2087 9962 2193
rect 10008 2227 10062 2239
rect 10008 2201 10018 2227
rect 10052 2201 10062 2227
rect 10008 2149 10009 2201
rect 10061 2149 10062 2201
rect 10008 2142 10062 2149
rect 10108 2227 10162 2333
rect 10208 2411 10262 2418
rect 10208 2359 10209 2411
rect 10261 2359 10262 2411
rect 10208 2333 10218 2359
rect 10252 2333 10262 2359
rect 10208 2321 10262 2333
rect 10308 2367 10362 2563
rect 10408 2597 10462 2609
rect 10408 2571 10418 2597
rect 10452 2571 10462 2597
rect 10408 2519 10409 2571
rect 10461 2519 10462 2571
rect 10408 2512 10462 2519
rect 10508 2597 10562 2703
rect 10608 2781 10662 2788
rect 10608 2729 10609 2781
rect 10661 2729 10662 2781
rect 10608 2703 10618 2729
rect 10652 2703 10662 2729
rect 10608 2691 10662 2703
rect 10708 2737 10762 2843
rect 10808 2877 10862 2889
rect 10808 2851 10818 2877
rect 10852 2851 10862 2877
rect 10808 2799 10809 2851
rect 10861 2799 10862 2851
rect 10808 2792 10862 2799
rect 10908 2877 10962 2983
rect 11008 3061 11062 3068
rect 11008 3009 11009 3061
rect 11061 3009 11062 3061
rect 11008 2983 11018 3009
rect 11052 2983 11062 3009
rect 11008 2971 11062 2983
rect 11108 3017 11162 3123
rect 11208 3157 11262 3169
rect 11208 3131 11218 3157
rect 11252 3131 11262 3157
rect 11208 3079 11209 3131
rect 11261 3079 11262 3131
rect 11208 3072 11262 3079
rect 11308 3157 11362 3263
rect 11408 3341 11462 3348
rect 11408 3289 11409 3341
rect 11461 3289 11462 3341
rect 11408 3263 11418 3289
rect 11452 3263 11462 3289
rect 11408 3251 11462 3263
rect 11508 3297 11562 3403
rect 11608 3437 11662 3449
rect 11608 3411 11618 3437
rect 11652 3411 11662 3437
rect 11608 3359 11609 3411
rect 11661 3359 11662 3411
rect 11608 3352 11662 3359
rect 11708 3437 11762 3543
rect 11808 3621 11862 3628
rect 11808 3569 11809 3621
rect 11861 3569 11862 3621
rect 11808 3543 11818 3569
rect 11852 3543 11862 3569
rect 11808 3531 11862 3543
rect 11908 3577 11962 3773
rect 12008 3807 12062 3819
rect 12008 3781 12018 3807
rect 12052 3781 12062 3807
rect 12008 3729 12009 3781
rect 12061 3729 12062 3781
rect 12008 3722 12062 3729
rect 12108 3807 12162 3913
rect 12208 3991 12262 3998
rect 12208 3939 12209 3991
rect 12261 3939 12262 3991
rect 12208 3913 12218 3939
rect 12252 3913 12262 3939
rect 12208 3901 12262 3913
rect 12308 3947 12362 4053
rect 12408 4087 12462 4099
rect 12408 4061 12418 4087
rect 12452 4061 12462 4087
rect 12408 4009 12409 4061
rect 12461 4009 12462 4061
rect 12408 4002 12462 4009
rect 12508 4087 12562 4193
rect 12608 4271 12662 4278
rect 12608 4219 12609 4271
rect 12661 4219 12662 4271
rect 12608 4193 12618 4219
rect 12652 4193 12662 4219
rect 12608 4181 12662 4193
rect 12708 4227 12762 4333
rect 12808 4367 12862 4379
rect 12808 4341 12818 4367
rect 12852 4341 12862 4367
rect 12808 4289 12809 4341
rect 12861 4289 12862 4341
rect 12808 4282 12862 4289
rect 12906 4348 12916 4382
rect 12950 4348 12960 4382
rect 12906 4341 12960 4348
rect 12906 4289 12907 4341
rect 12959 4289 12960 4341
rect 12906 4282 12960 4289
rect 12906 4242 12960 4254
rect 12708 4193 12718 4227
rect 12752 4193 12762 4227
rect 12508 4053 12518 4087
rect 12552 4053 12562 4087
rect 12308 3913 12318 3947
rect 12352 3913 12362 3947
rect 12108 3773 12118 3807
rect 12152 3773 12162 3807
rect 12002 3693 12068 3694
rect 12002 3641 12009 3693
rect 12061 3641 12068 3693
rect 12002 3640 12068 3641
rect 11908 3543 11918 3577
rect 11952 3543 11962 3577
rect 11708 3403 11718 3437
rect 11752 3403 11762 3437
rect 11508 3263 11518 3297
rect 11552 3263 11562 3297
rect 11308 3123 11318 3157
rect 11352 3123 11362 3157
rect 11108 2983 11118 3017
rect 11152 2983 11162 3017
rect 10908 2843 10918 2877
rect 10952 2843 10962 2877
rect 10708 2703 10718 2737
rect 10752 2703 10762 2737
rect 10508 2563 10518 2597
rect 10552 2563 10562 2597
rect 10402 2483 10468 2484
rect 10402 2431 10409 2483
rect 10461 2431 10468 2483
rect 10402 2430 10468 2431
rect 10308 2333 10318 2367
rect 10352 2333 10362 2367
rect 10108 2193 10118 2227
rect 10152 2193 10162 2227
rect 9908 2053 9918 2087
rect 9952 2053 9962 2087
rect 9708 1913 9718 1947
rect 9752 1913 9762 1947
rect 9508 1773 9518 1807
rect 9552 1773 9562 1807
rect 9308 1633 9318 1667
rect 9352 1633 9362 1667
rect 9108 1493 9118 1527
rect 9152 1493 9162 1527
rect 8908 1353 8918 1387
rect 8952 1353 8962 1387
rect 8802 1273 8868 1274
rect 8802 1221 8809 1273
rect 8861 1221 8868 1273
rect 8802 1220 8868 1221
rect 8708 1123 8718 1157
rect 8752 1123 8762 1157
rect 8508 983 8518 1017
rect 8552 983 8562 1017
rect 8308 843 8318 877
rect 8352 843 8362 877
rect 8108 703 8118 737
rect 8152 703 8162 737
rect 7908 563 7918 597
rect 7952 563 7962 597
rect 7708 423 7718 457
rect 7752 423 7762 457
rect 7508 283 7518 317
rect 7552 283 7562 317
rect 7308 143 7318 177
rect 7352 143 7362 177
rect 7202 63 7268 64
rect 7202 11 7209 63
rect 7261 11 7268 63
rect 7202 10 7268 11
rect 7108 -67 7109 -15
rect 7161 -67 7162 -15
rect 7108 -79 7118 -67
rect 7152 -79 7162 -67
rect 6908 -132 6962 -131
rect 6908 -143 6918 -132
rect 6952 -143 6962 -132
rect 6908 -195 6909 -143
rect 6961 -195 6962 -143
rect 6908 -210 6962 -195
rect 7012 -133 7058 -81
rect 7012 -167 7018 -133
rect 7052 -167 7058 -133
rect 6918 -291 6925 -239
rect 6977 -291 6984 -239
rect 6812 -397 6818 -363
rect 6852 -397 6858 -363
rect 6812 -435 6858 -397
rect 6812 -469 6818 -435
rect 6852 -469 6858 -435
rect 6812 -512 6858 -469
rect 6909 -326 6961 -320
rect 6909 -390 6918 -378
rect 6952 -390 6961 -378
rect 6909 -454 6918 -442
rect 6952 -454 6961 -442
rect 6909 -512 6961 -506
rect 7012 -363 7058 -167
rect 7108 -131 7109 -79
rect 7161 -131 7162 -79
rect 7208 -22 7262 10
rect 7208 -74 7209 -22
rect 7261 -74 7262 -22
rect 7208 -81 7262 -74
rect 7308 -15 7362 143
rect 7408 221 7462 228
rect 7408 169 7409 221
rect 7461 169 7462 221
rect 7408 143 7418 169
rect 7452 143 7462 169
rect 7408 131 7462 143
rect 7508 177 7562 283
rect 7608 317 7662 329
rect 7608 291 7618 317
rect 7652 291 7662 317
rect 7608 239 7609 291
rect 7661 239 7662 291
rect 7608 232 7662 239
rect 7708 317 7762 423
rect 7808 501 7862 508
rect 7808 449 7809 501
rect 7861 449 7862 501
rect 7808 423 7818 449
rect 7852 423 7862 449
rect 7808 411 7862 423
rect 7908 457 7962 563
rect 8008 597 8062 609
rect 8008 571 8018 597
rect 8052 571 8062 597
rect 8008 519 8009 571
rect 8061 519 8062 571
rect 8008 512 8062 519
rect 8108 597 8162 703
rect 8208 781 8262 788
rect 8208 729 8209 781
rect 8261 729 8262 781
rect 8208 703 8218 729
rect 8252 703 8262 729
rect 8208 691 8262 703
rect 8308 737 8362 843
rect 8408 877 8462 889
rect 8408 851 8418 877
rect 8452 851 8462 877
rect 8408 799 8409 851
rect 8461 799 8462 851
rect 8408 792 8462 799
rect 8508 877 8562 983
rect 8608 1061 8662 1068
rect 8608 1009 8609 1061
rect 8661 1009 8662 1061
rect 8608 983 8618 1009
rect 8652 983 8662 1009
rect 8608 971 8662 983
rect 8708 1017 8762 1123
rect 8808 1157 8862 1169
rect 8808 1131 8818 1157
rect 8852 1131 8862 1157
rect 8808 1079 8809 1131
rect 8861 1079 8862 1131
rect 8808 1072 8862 1079
rect 8908 1157 8962 1353
rect 9008 1431 9062 1438
rect 9008 1379 9009 1431
rect 9061 1379 9062 1431
rect 9008 1353 9018 1379
rect 9052 1353 9062 1379
rect 9008 1341 9062 1353
rect 9108 1387 9162 1493
rect 9208 1527 9262 1539
rect 9208 1501 9218 1527
rect 9252 1501 9262 1527
rect 9208 1449 9209 1501
rect 9261 1449 9262 1501
rect 9208 1442 9262 1449
rect 9308 1527 9362 1633
rect 9408 1711 9462 1718
rect 9408 1659 9409 1711
rect 9461 1659 9462 1711
rect 9408 1633 9418 1659
rect 9452 1633 9462 1659
rect 9408 1621 9462 1633
rect 9508 1667 9562 1773
rect 9608 1807 9662 1819
rect 9608 1781 9618 1807
rect 9652 1781 9662 1807
rect 9608 1729 9609 1781
rect 9661 1729 9662 1781
rect 9608 1722 9662 1729
rect 9708 1807 9762 1913
rect 9808 1991 9862 1998
rect 9808 1939 9809 1991
rect 9861 1939 9862 1991
rect 9808 1913 9818 1939
rect 9852 1913 9862 1939
rect 9808 1901 9862 1913
rect 9908 1947 9962 2053
rect 10008 2087 10062 2099
rect 10008 2061 10018 2087
rect 10052 2061 10062 2087
rect 10008 2009 10009 2061
rect 10061 2009 10062 2061
rect 10008 2002 10062 2009
rect 10108 2087 10162 2193
rect 10208 2271 10262 2278
rect 10208 2219 10209 2271
rect 10261 2219 10262 2271
rect 10208 2193 10218 2219
rect 10252 2193 10262 2219
rect 10208 2181 10262 2193
rect 10308 2227 10362 2333
rect 10408 2367 10462 2379
rect 10408 2341 10418 2367
rect 10452 2341 10462 2367
rect 10408 2289 10409 2341
rect 10461 2289 10462 2341
rect 10408 2282 10462 2289
rect 10508 2367 10562 2563
rect 10608 2641 10662 2648
rect 10608 2589 10609 2641
rect 10661 2589 10662 2641
rect 10608 2563 10618 2589
rect 10652 2563 10662 2589
rect 10608 2551 10662 2563
rect 10708 2597 10762 2703
rect 10808 2737 10862 2749
rect 10808 2711 10818 2737
rect 10852 2711 10862 2737
rect 10808 2659 10809 2711
rect 10861 2659 10862 2711
rect 10808 2652 10862 2659
rect 10908 2737 10962 2843
rect 11008 2921 11062 2928
rect 11008 2869 11009 2921
rect 11061 2869 11062 2921
rect 11008 2843 11018 2869
rect 11052 2843 11062 2869
rect 11008 2831 11062 2843
rect 11108 2877 11162 2983
rect 11208 3017 11262 3029
rect 11208 2991 11218 3017
rect 11252 2991 11262 3017
rect 11208 2939 11209 2991
rect 11261 2939 11262 2991
rect 11208 2932 11262 2939
rect 11308 3017 11362 3123
rect 11408 3201 11462 3208
rect 11408 3149 11409 3201
rect 11461 3149 11462 3201
rect 11408 3123 11418 3149
rect 11452 3123 11462 3149
rect 11408 3111 11462 3123
rect 11508 3157 11562 3263
rect 11608 3297 11662 3309
rect 11608 3271 11618 3297
rect 11652 3271 11662 3297
rect 11608 3219 11609 3271
rect 11661 3219 11662 3271
rect 11608 3212 11662 3219
rect 11708 3297 11762 3403
rect 11808 3481 11862 3488
rect 11808 3429 11809 3481
rect 11861 3429 11862 3481
rect 11808 3403 11818 3429
rect 11852 3403 11862 3429
rect 11808 3391 11862 3403
rect 11908 3437 11962 3543
rect 12008 3577 12062 3589
rect 12008 3551 12018 3577
rect 12052 3551 12062 3577
rect 12008 3499 12009 3551
rect 12061 3499 12062 3551
rect 12008 3492 12062 3499
rect 12108 3577 12162 3773
rect 12208 3851 12262 3858
rect 12208 3799 12209 3851
rect 12261 3799 12262 3851
rect 12208 3773 12218 3799
rect 12252 3773 12262 3799
rect 12208 3761 12262 3773
rect 12308 3807 12362 3913
rect 12408 3947 12462 3959
rect 12408 3921 12418 3947
rect 12452 3921 12462 3947
rect 12408 3869 12409 3921
rect 12461 3869 12462 3921
rect 12408 3862 12462 3869
rect 12508 3947 12562 4053
rect 12608 4131 12662 4138
rect 12608 4079 12609 4131
rect 12661 4079 12662 4131
rect 12608 4053 12618 4079
rect 12652 4053 12662 4079
rect 12608 4041 12662 4053
rect 12708 4087 12762 4193
rect 12808 4227 12862 4239
rect 12808 4201 12818 4227
rect 12852 4201 12862 4227
rect 12808 4149 12809 4201
rect 12861 4149 12862 4201
rect 12808 4142 12862 4149
rect 12906 4208 12916 4242
rect 12950 4208 12960 4242
rect 12906 4201 12960 4208
rect 12906 4149 12907 4201
rect 12959 4149 12960 4201
rect 12906 4142 12960 4149
rect 12906 4102 12960 4114
rect 12708 4053 12718 4087
rect 12752 4053 12762 4087
rect 12508 3913 12518 3947
rect 12552 3913 12562 3947
rect 12308 3773 12318 3807
rect 12352 3773 12362 3807
rect 12202 3709 12268 3710
rect 12202 3657 12209 3709
rect 12261 3657 12268 3709
rect 12202 3656 12268 3657
rect 12108 3543 12118 3577
rect 12152 3543 12162 3577
rect 11908 3403 11918 3437
rect 11952 3403 11962 3437
rect 11708 3263 11718 3297
rect 11752 3263 11762 3297
rect 11508 3123 11518 3157
rect 11552 3123 11562 3157
rect 11308 2983 11318 3017
rect 11352 2983 11362 3017
rect 11108 2843 11118 2877
rect 11152 2843 11162 2877
rect 10908 2703 10918 2737
rect 10952 2703 10962 2737
rect 10708 2563 10718 2597
rect 10752 2563 10762 2597
rect 10602 2499 10668 2500
rect 10602 2447 10609 2499
rect 10661 2447 10668 2499
rect 10602 2446 10668 2447
rect 10508 2333 10518 2367
rect 10552 2333 10562 2367
rect 10308 2193 10318 2227
rect 10352 2193 10362 2227
rect 10108 2053 10118 2087
rect 10152 2053 10162 2087
rect 9908 1913 9918 1947
rect 9952 1913 9962 1947
rect 9708 1773 9718 1807
rect 9752 1773 9762 1807
rect 9508 1633 9518 1667
rect 9552 1633 9562 1667
rect 9308 1493 9318 1527
rect 9352 1493 9362 1527
rect 9108 1353 9118 1387
rect 9152 1353 9162 1387
rect 9002 1289 9068 1290
rect 9002 1237 9009 1289
rect 9061 1237 9068 1289
rect 9002 1236 9068 1237
rect 8908 1123 8918 1157
rect 8952 1123 8962 1157
rect 8708 983 8718 1017
rect 8752 983 8762 1017
rect 8508 843 8518 877
rect 8552 843 8562 877
rect 8308 703 8318 737
rect 8352 703 8362 737
rect 8108 563 8118 597
rect 8152 563 8162 597
rect 7908 423 7918 457
rect 7952 423 7962 457
rect 7708 283 7718 317
rect 7752 283 7762 317
rect 7508 143 7518 177
rect 7552 143 7562 177
rect 7402 79 7468 80
rect 7402 27 7409 79
rect 7461 27 7468 79
rect 7402 26 7468 27
rect 7308 -67 7309 -15
rect 7361 -67 7362 -15
rect 7308 -79 7318 -67
rect 7352 -79 7362 -67
rect 7108 -132 7162 -131
rect 7108 -143 7118 -132
rect 7152 -143 7162 -132
rect 7108 -195 7109 -143
rect 7161 -195 7162 -143
rect 7108 -210 7162 -195
rect 7212 -133 7258 -81
rect 7212 -167 7218 -133
rect 7252 -167 7258 -133
rect 7118 -291 7125 -239
rect 7177 -291 7184 -239
rect 7012 -397 7018 -363
rect 7052 -397 7058 -363
rect 7012 -435 7058 -397
rect 7012 -469 7018 -435
rect 7052 -469 7058 -435
rect 7012 -512 7058 -469
rect 7109 -326 7161 -320
rect 7109 -390 7118 -378
rect 7152 -390 7161 -378
rect 7109 -454 7118 -442
rect 7152 -454 7161 -442
rect 7109 -555 7161 -506
rect 7212 -363 7258 -167
rect 7308 -131 7309 -79
rect 7361 -131 7362 -79
rect 7408 -22 7462 26
rect 7408 -74 7409 -22
rect 7461 -74 7462 -22
rect 7408 -81 7462 -74
rect 7508 -15 7562 143
rect 7608 177 7662 189
rect 7608 151 7618 177
rect 7652 151 7662 177
rect 7608 99 7609 151
rect 7661 99 7662 151
rect 7608 92 7662 99
rect 7708 177 7762 283
rect 7808 361 7862 368
rect 7808 309 7809 361
rect 7861 309 7862 361
rect 7808 283 7818 309
rect 7852 283 7862 309
rect 7808 271 7862 283
rect 7908 317 7962 423
rect 8008 457 8062 469
rect 8008 431 8018 457
rect 8052 431 8062 457
rect 8008 379 8009 431
rect 8061 379 8062 431
rect 8008 372 8062 379
rect 8108 457 8162 563
rect 8208 641 8262 648
rect 8208 589 8209 641
rect 8261 589 8262 641
rect 8208 563 8218 589
rect 8252 563 8262 589
rect 8208 551 8262 563
rect 8308 597 8362 703
rect 8408 737 8462 749
rect 8408 711 8418 737
rect 8452 711 8462 737
rect 8408 659 8409 711
rect 8461 659 8462 711
rect 8408 652 8462 659
rect 8508 737 8562 843
rect 8608 921 8662 928
rect 8608 869 8609 921
rect 8661 869 8662 921
rect 8608 843 8618 869
rect 8652 843 8662 869
rect 8608 831 8662 843
rect 8708 877 8762 983
rect 8808 1017 8862 1029
rect 8808 991 8818 1017
rect 8852 991 8862 1017
rect 8808 939 8809 991
rect 8861 939 8862 991
rect 8808 932 8862 939
rect 8908 1017 8962 1123
rect 9008 1201 9062 1208
rect 9008 1149 9009 1201
rect 9061 1149 9062 1201
rect 9008 1123 9018 1149
rect 9052 1123 9062 1149
rect 9008 1111 9062 1123
rect 9108 1157 9162 1353
rect 9208 1387 9262 1399
rect 9208 1361 9218 1387
rect 9252 1361 9262 1387
rect 9208 1309 9209 1361
rect 9261 1309 9262 1361
rect 9208 1302 9262 1309
rect 9308 1387 9362 1493
rect 9408 1571 9462 1578
rect 9408 1519 9409 1571
rect 9461 1519 9462 1571
rect 9408 1493 9418 1519
rect 9452 1493 9462 1519
rect 9408 1481 9462 1493
rect 9508 1527 9562 1633
rect 9608 1667 9662 1679
rect 9608 1641 9618 1667
rect 9652 1641 9662 1667
rect 9608 1589 9609 1641
rect 9661 1589 9662 1641
rect 9608 1582 9662 1589
rect 9708 1667 9762 1773
rect 9808 1851 9862 1858
rect 9808 1799 9809 1851
rect 9861 1799 9862 1851
rect 9808 1773 9818 1799
rect 9852 1773 9862 1799
rect 9808 1761 9862 1773
rect 9908 1807 9962 1913
rect 10008 1947 10062 1959
rect 10008 1921 10018 1947
rect 10052 1921 10062 1947
rect 10008 1869 10009 1921
rect 10061 1869 10062 1921
rect 10008 1862 10062 1869
rect 10108 1947 10162 2053
rect 10208 2131 10262 2138
rect 10208 2079 10209 2131
rect 10261 2079 10262 2131
rect 10208 2053 10218 2079
rect 10252 2053 10262 2079
rect 10208 2041 10262 2053
rect 10308 2087 10362 2193
rect 10408 2227 10462 2239
rect 10408 2201 10418 2227
rect 10452 2201 10462 2227
rect 10408 2149 10409 2201
rect 10461 2149 10462 2201
rect 10408 2142 10462 2149
rect 10508 2227 10562 2333
rect 10608 2411 10662 2418
rect 10608 2359 10609 2411
rect 10661 2359 10662 2411
rect 10608 2333 10618 2359
rect 10652 2333 10662 2359
rect 10608 2321 10662 2333
rect 10708 2367 10762 2563
rect 10808 2597 10862 2609
rect 10808 2571 10818 2597
rect 10852 2571 10862 2597
rect 10808 2519 10809 2571
rect 10861 2519 10862 2571
rect 10808 2512 10862 2519
rect 10908 2597 10962 2703
rect 11008 2781 11062 2788
rect 11008 2729 11009 2781
rect 11061 2729 11062 2781
rect 11008 2703 11018 2729
rect 11052 2703 11062 2729
rect 11008 2691 11062 2703
rect 11108 2737 11162 2843
rect 11208 2877 11262 2889
rect 11208 2851 11218 2877
rect 11252 2851 11262 2877
rect 11208 2799 11209 2851
rect 11261 2799 11262 2851
rect 11208 2792 11262 2799
rect 11308 2877 11362 2983
rect 11408 3061 11462 3068
rect 11408 3009 11409 3061
rect 11461 3009 11462 3061
rect 11408 2983 11418 3009
rect 11452 2983 11462 3009
rect 11408 2971 11462 2983
rect 11508 3017 11562 3123
rect 11608 3157 11662 3169
rect 11608 3131 11618 3157
rect 11652 3131 11662 3157
rect 11608 3079 11609 3131
rect 11661 3079 11662 3131
rect 11608 3072 11662 3079
rect 11708 3157 11762 3263
rect 11808 3341 11862 3348
rect 11808 3289 11809 3341
rect 11861 3289 11862 3341
rect 11808 3263 11818 3289
rect 11852 3263 11862 3289
rect 11808 3251 11862 3263
rect 11908 3297 11962 3403
rect 12008 3437 12062 3449
rect 12008 3411 12018 3437
rect 12052 3411 12062 3437
rect 12008 3359 12009 3411
rect 12061 3359 12062 3411
rect 12008 3352 12062 3359
rect 12108 3437 12162 3543
rect 12208 3621 12262 3628
rect 12208 3569 12209 3621
rect 12261 3569 12262 3621
rect 12208 3543 12218 3569
rect 12252 3543 12262 3569
rect 12208 3531 12262 3543
rect 12308 3577 12362 3773
rect 12408 3807 12462 3819
rect 12408 3781 12418 3807
rect 12452 3781 12462 3807
rect 12408 3729 12409 3781
rect 12461 3729 12462 3781
rect 12408 3722 12462 3729
rect 12508 3807 12562 3913
rect 12608 3991 12662 3998
rect 12608 3939 12609 3991
rect 12661 3939 12662 3991
rect 12608 3913 12618 3939
rect 12652 3913 12662 3939
rect 12608 3901 12662 3913
rect 12708 3947 12762 4053
rect 12808 4087 12862 4099
rect 12808 4061 12818 4087
rect 12852 4061 12862 4087
rect 12808 4009 12809 4061
rect 12861 4009 12862 4061
rect 12808 4002 12862 4009
rect 12906 4068 12916 4102
rect 12950 4068 12960 4102
rect 12906 4061 12960 4068
rect 12906 4009 12907 4061
rect 12959 4009 12960 4061
rect 12906 4002 12960 4009
rect 12906 3962 12960 3974
rect 12708 3913 12718 3947
rect 12752 3913 12762 3947
rect 12508 3773 12518 3807
rect 12552 3773 12562 3807
rect 12402 3693 12468 3694
rect 12402 3641 12409 3693
rect 12461 3641 12468 3693
rect 12402 3640 12468 3641
rect 12308 3543 12318 3577
rect 12352 3543 12362 3577
rect 12108 3403 12118 3437
rect 12152 3403 12162 3437
rect 11908 3263 11918 3297
rect 11952 3263 11962 3297
rect 11708 3123 11718 3157
rect 11752 3123 11762 3157
rect 11508 2983 11518 3017
rect 11552 2983 11562 3017
rect 11308 2843 11318 2877
rect 11352 2843 11362 2877
rect 11108 2703 11118 2737
rect 11152 2703 11162 2737
rect 10908 2563 10918 2597
rect 10952 2563 10962 2597
rect 10802 2483 10868 2484
rect 10802 2431 10809 2483
rect 10861 2431 10868 2483
rect 10802 2430 10868 2431
rect 10708 2333 10718 2367
rect 10752 2333 10762 2367
rect 10508 2193 10518 2227
rect 10552 2193 10562 2227
rect 10308 2053 10318 2087
rect 10352 2053 10362 2087
rect 10108 1913 10118 1947
rect 10152 1913 10162 1947
rect 9908 1773 9918 1807
rect 9952 1773 9962 1807
rect 9708 1633 9718 1667
rect 9752 1633 9762 1667
rect 9508 1493 9518 1527
rect 9552 1493 9562 1527
rect 9308 1353 9318 1387
rect 9352 1353 9362 1387
rect 9202 1273 9268 1274
rect 9202 1221 9209 1273
rect 9261 1221 9268 1273
rect 9202 1220 9268 1221
rect 9108 1123 9118 1157
rect 9152 1123 9162 1157
rect 8908 983 8918 1017
rect 8952 983 8962 1017
rect 8708 843 8718 877
rect 8752 843 8762 877
rect 8508 703 8518 737
rect 8552 703 8562 737
rect 8308 563 8318 597
rect 8352 563 8362 597
rect 8108 423 8118 457
rect 8152 423 8162 457
rect 7908 283 7918 317
rect 7952 283 7962 317
rect 7708 143 7718 177
rect 7752 143 7762 177
rect 7602 63 7668 64
rect 7602 11 7609 63
rect 7661 11 7668 63
rect 7602 10 7668 11
rect 7508 -67 7509 -15
rect 7561 -67 7562 -15
rect 7508 -79 7518 -67
rect 7552 -79 7562 -67
rect 7308 -132 7362 -131
rect 7308 -143 7318 -132
rect 7352 -143 7362 -132
rect 7308 -195 7309 -143
rect 7361 -195 7362 -143
rect 7308 -210 7362 -195
rect 7412 -133 7458 -81
rect 7412 -167 7418 -133
rect 7452 -167 7458 -133
rect 7318 -291 7325 -239
rect 7377 -291 7384 -239
rect 7212 -397 7218 -363
rect 7252 -397 7258 -363
rect 7212 -435 7258 -397
rect 7212 -469 7218 -435
rect 7252 -469 7258 -435
rect 7212 -512 7258 -469
rect 7309 -326 7361 -320
rect 7309 -390 7318 -378
rect 7352 -390 7361 -378
rect 7309 -454 7318 -442
rect 7352 -454 7361 -442
rect 7309 -512 7361 -506
rect 7412 -363 7458 -167
rect 7508 -131 7509 -79
rect 7561 -131 7562 -79
rect 7608 -22 7662 10
rect 7608 -74 7609 -22
rect 7661 -74 7662 -22
rect 7608 -81 7662 -74
rect 7708 -15 7762 143
rect 7808 221 7862 228
rect 7808 169 7809 221
rect 7861 169 7862 221
rect 7808 143 7818 169
rect 7852 143 7862 169
rect 7808 131 7862 143
rect 7908 177 7962 283
rect 8008 317 8062 329
rect 8008 291 8018 317
rect 8052 291 8062 317
rect 8008 239 8009 291
rect 8061 239 8062 291
rect 8008 232 8062 239
rect 8108 317 8162 423
rect 8208 501 8262 508
rect 8208 449 8209 501
rect 8261 449 8262 501
rect 8208 423 8218 449
rect 8252 423 8262 449
rect 8208 411 8262 423
rect 8308 457 8362 563
rect 8408 597 8462 609
rect 8408 571 8418 597
rect 8452 571 8462 597
rect 8408 519 8409 571
rect 8461 519 8462 571
rect 8408 512 8462 519
rect 8508 597 8562 703
rect 8608 781 8662 788
rect 8608 729 8609 781
rect 8661 729 8662 781
rect 8608 703 8618 729
rect 8652 703 8662 729
rect 8608 691 8662 703
rect 8708 737 8762 843
rect 8808 877 8862 889
rect 8808 851 8818 877
rect 8852 851 8862 877
rect 8808 799 8809 851
rect 8861 799 8862 851
rect 8808 792 8862 799
rect 8908 877 8962 983
rect 9008 1061 9062 1068
rect 9008 1009 9009 1061
rect 9061 1009 9062 1061
rect 9008 983 9018 1009
rect 9052 983 9062 1009
rect 9008 971 9062 983
rect 9108 1017 9162 1123
rect 9208 1157 9262 1169
rect 9208 1131 9218 1157
rect 9252 1131 9262 1157
rect 9208 1079 9209 1131
rect 9261 1079 9262 1131
rect 9208 1072 9262 1079
rect 9308 1157 9362 1353
rect 9408 1431 9462 1438
rect 9408 1379 9409 1431
rect 9461 1379 9462 1431
rect 9408 1353 9418 1379
rect 9452 1353 9462 1379
rect 9408 1341 9462 1353
rect 9508 1387 9562 1493
rect 9608 1527 9662 1539
rect 9608 1501 9618 1527
rect 9652 1501 9662 1527
rect 9608 1449 9609 1501
rect 9661 1449 9662 1501
rect 9608 1442 9662 1449
rect 9708 1527 9762 1633
rect 9808 1711 9862 1718
rect 9808 1659 9809 1711
rect 9861 1659 9862 1711
rect 9808 1633 9818 1659
rect 9852 1633 9862 1659
rect 9808 1621 9862 1633
rect 9908 1667 9962 1773
rect 10008 1807 10062 1819
rect 10008 1781 10018 1807
rect 10052 1781 10062 1807
rect 10008 1729 10009 1781
rect 10061 1729 10062 1781
rect 10008 1722 10062 1729
rect 10108 1807 10162 1913
rect 10208 1991 10262 1998
rect 10208 1939 10209 1991
rect 10261 1939 10262 1991
rect 10208 1913 10218 1939
rect 10252 1913 10262 1939
rect 10208 1901 10262 1913
rect 10308 1947 10362 2053
rect 10408 2087 10462 2099
rect 10408 2061 10418 2087
rect 10452 2061 10462 2087
rect 10408 2009 10409 2061
rect 10461 2009 10462 2061
rect 10408 2002 10462 2009
rect 10508 2087 10562 2193
rect 10608 2271 10662 2278
rect 10608 2219 10609 2271
rect 10661 2219 10662 2271
rect 10608 2193 10618 2219
rect 10652 2193 10662 2219
rect 10608 2181 10662 2193
rect 10708 2227 10762 2333
rect 10808 2367 10862 2379
rect 10808 2341 10818 2367
rect 10852 2341 10862 2367
rect 10808 2289 10809 2341
rect 10861 2289 10862 2341
rect 10808 2282 10862 2289
rect 10908 2367 10962 2563
rect 11008 2641 11062 2648
rect 11008 2589 11009 2641
rect 11061 2589 11062 2641
rect 11008 2563 11018 2589
rect 11052 2563 11062 2589
rect 11008 2551 11062 2563
rect 11108 2597 11162 2703
rect 11208 2737 11262 2749
rect 11208 2711 11218 2737
rect 11252 2711 11262 2737
rect 11208 2659 11209 2711
rect 11261 2659 11262 2711
rect 11208 2652 11262 2659
rect 11308 2737 11362 2843
rect 11408 2921 11462 2928
rect 11408 2869 11409 2921
rect 11461 2869 11462 2921
rect 11408 2843 11418 2869
rect 11452 2843 11462 2869
rect 11408 2831 11462 2843
rect 11508 2877 11562 2983
rect 11608 3017 11662 3029
rect 11608 2991 11618 3017
rect 11652 2991 11662 3017
rect 11608 2939 11609 2991
rect 11661 2939 11662 2991
rect 11608 2932 11662 2939
rect 11708 3017 11762 3123
rect 11808 3201 11862 3208
rect 11808 3149 11809 3201
rect 11861 3149 11862 3201
rect 11808 3123 11818 3149
rect 11852 3123 11862 3149
rect 11808 3111 11862 3123
rect 11908 3157 11962 3263
rect 12008 3297 12062 3309
rect 12008 3271 12018 3297
rect 12052 3271 12062 3297
rect 12008 3219 12009 3271
rect 12061 3219 12062 3271
rect 12008 3212 12062 3219
rect 12108 3297 12162 3403
rect 12208 3481 12262 3488
rect 12208 3429 12209 3481
rect 12261 3429 12262 3481
rect 12208 3403 12218 3429
rect 12252 3403 12262 3429
rect 12208 3391 12262 3403
rect 12308 3437 12362 3543
rect 12408 3577 12462 3589
rect 12408 3551 12418 3577
rect 12452 3551 12462 3577
rect 12408 3499 12409 3551
rect 12461 3499 12462 3551
rect 12408 3492 12462 3499
rect 12508 3577 12562 3773
rect 12608 3851 12662 3858
rect 12608 3799 12609 3851
rect 12661 3799 12662 3851
rect 12608 3773 12618 3799
rect 12652 3773 12662 3799
rect 12608 3761 12662 3773
rect 12708 3807 12762 3913
rect 12808 3947 12862 3959
rect 12808 3921 12818 3947
rect 12852 3921 12862 3947
rect 12808 3869 12809 3921
rect 12861 3869 12862 3921
rect 12808 3862 12862 3869
rect 12906 3928 12916 3962
rect 12950 3928 12960 3962
rect 12906 3921 12960 3928
rect 12906 3869 12907 3921
rect 12959 3869 12960 3921
rect 12906 3862 12960 3869
rect 12906 3822 12960 3834
rect 12708 3773 12718 3807
rect 12752 3773 12762 3807
rect 12602 3709 12668 3710
rect 12602 3657 12609 3709
rect 12661 3657 12668 3709
rect 12602 3656 12668 3657
rect 12508 3543 12518 3577
rect 12552 3543 12562 3577
rect 12308 3403 12318 3437
rect 12352 3403 12362 3437
rect 12108 3263 12118 3297
rect 12152 3263 12162 3297
rect 11908 3123 11918 3157
rect 11952 3123 11962 3157
rect 11708 2983 11718 3017
rect 11752 2983 11762 3017
rect 11508 2843 11518 2877
rect 11552 2843 11562 2877
rect 11308 2703 11318 2737
rect 11352 2703 11362 2737
rect 11108 2563 11118 2597
rect 11152 2563 11162 2597
rect 11002 2499 11068 2500
rect 11002 2447 11009 2499
rect 11061 2447 11068 2499
rect 11002 2446 11068 2447
rect 10908 2333 10918 2367
rect 10952 2333 10962 2367
rect 10708 2193 10718 2227
rect 10752 2193 10762 2227
rect 10508 2053 10518 2087
rect 10552 2053 10562 2087
rect 10308 1913 10318 1947
rect 10352 1913 10362 1947
rect 10108 1773 10118 1807
rect 10152 1773 10162 1807
rect 9908 1633 9918 1667
rect 9952 1633 9962 1667
rect 9708 1493 9718 1527
rect 9752 1493 9762 1527
rect 9508 1353 9518 1387
rect 9552 1353 9562 1387
rect 9402 1289 9468 1290
rect 9402 1237 9409 1289
rect 9461 1237 9468 1289
rect 9402 1236 9468 1237
rect 9308 1123 9318 1157
rect 9352 1123 9362 1157
rect 9108 983 9118 1017
rect 9152 983 9162 1017
rect 8908 843 8918 877
rect 8952 843 8962 877
rect 8708 703 8718 737
rect 8752 703 8762 737
rect 8508 563 8518 597
rect 8552 563 8562 597
rect 8308 423 8318 457
rect 8352 423 8362 457
rect 8108 283 8118 317
rect 8152 283 8162 317
rect 7908 143 7918 177
rect 7952 143 7962 177
rect 7802 79 7868 80
rect 7802 27 7809 79
rect 7861 27 7868 79
rect 7802 26 7868 27
rect 7708 -67 7709 -15
rect 7761 -67 7762 -15
rect 7708 -79 7718 -67
rect 7752 -79 7762 -67
rect 7508 -132 7562 -131
rect 7508 -143 7518 -132
rect 7552 -143 7562 -132
rect 7508 -195 7509 -143
rect 7561 -195 7562 -143
rect 7508 -210 7562 -195
rect 7612 -133 7658 -81
rect 7612 -167 7618 -133
rect 7652 -167 7658 -133
rect 7518 -291 7525 -239
rect 7577 -291 7584 -239
rect 7412 -397 7418 -363
rect 7452 -397 7458 -363
rect 7412 -435 7458 -397
rect 7412 -469 7418 -435
rect 7452 -469 7458 -435
rect 7412 -512 7458 -469
rect 7509 -326 7561 -320
rect 7509 -390 7518 -378
rect 7552 -390 7561 -378
rect 7509 -454 7518 -442
rect 7552 -454 7561 -442
rect 7509 -555 7561 -506
rect 7612 -363 7658 -167
rect 7708 -131 7709 -79
rect 7761 -131 7762 -79
rect 7808 -22 7862 26
rect 7808 -74 7809 -22
rect 7861 -74 7862 -22
rect 7808 -81 7862 -74
rect 7908 -15 7962 143
rect 8008 177 8062 189
rect 8008 151 8018 177
rect 8052 151 8062 177
rect 8008 99 8009 151
rect 8061 99 8062 151
rect 8008 92 8062 99
rect 8108 177 8162 283
rect 8208 361 8262 368
rect 8208 309 8209 361
rect 8261 309 8262 361
rect 8208 283 8218 309
rect 8252 283 8262 309
rect 8208 271 8262 283
rect 8308 317 8362 423
rect 8408 457 8462 469
rect 8408 431 8418 457
rect 8452 431 8462 457
rect 8408 379 8409 431
rect 8461 379 8462 431
rect 8408 372 8462 379
rect 8508 457 8562 563
rect 8608 641 8662 648
rect 8608 589 8609 641
rect 8661 589 8662 641
rect 8608 563 8618 589
rect 8652 563 8662 589
rect 8608 551 8662 563
rect 8708 597 8762 703
rect 8808 737 8862 749
rect 8808 711 8818 737
rect 8852 711 8862 737
rect 8808 659 8809 711
rect 8861 659 8862 711
rect 8808 652 8862 659
rect 8908 737 8962 843
rect 9008 921 9062 928
rect 9008 869 9009 921
rect 9061 869 9062 921
rect 9008 843 9018 869
rect 9052 843 9062 869
rect 9008 831 9062 843
rect 9108 877 9162 983
rect 9208 1017 9262 1029
rect 9208 991 9218 1017
rect 9252 991 9262 1017
rect 9208 939 9209 991
rect 9261 939 9262 991
rect 9208 932 9262 939
rect 9308 1017 9362 1123
rect 9408 1201 9462 1208
rect 9408 1149 9409 1201
rect 9461 1149 9462 1201
rect 9408 1123 9418 1149
rect 9452 1123 9462 1149
rect 9408 1111 9462 1123
rect 9508 1157 9562 1353
rect 9608 1387 9662 1399
rect 9608 1361 9618 1387
rect 9652 1361 9662 1387
rect 9608 1309 9609 1361
rect 9661 1309 9662 1361
rect 9608 1302 9662 1309
rect 9708 1387 9762 1493
rect 9808 1571 9862 1578
rect 9808 1519 9809 1571
rect 9861 1519 9862 1571
rect 9808 1493 9818 1519
rect 9852 1493 9862 1519
rect 9808 1481 9862 1493
rect 9908 1527 9962 1633
rect 10008 1667 10062 1679
rect 10008 1641 10018 1667
rect 10052 1641 10062 1667
rect 10008 1589 10009 1641
rect 10061 1589 10062 1641
rect 10008 1582 10062 1589
rect 10108 1667 10162 1773
rect 10208 1851 10262 1858
rect 10208 1799 10209 1851
rect 10261 1799 10262 1851
rect 10208 1773 10218 1799
rect 10252 1773 10262 1799
rect 10208 1761 10262 1773
rect 10308 1807 10362 1913
rect 10408 1947 10462 1959
rect 10408 1921 10418 1947
rect 10452 1921 10462 1947
rect 10408 1869 10409 1921
rect 10461 1869 10462 1921
rect 10408 1862 10462 1869
rect 10508 1947 10562 2053
rect 10608 2131 10662 2138
rect 10608 2079 10609 2131
rect 10661 2079 10662 2131
rect 10608 2053 10618 2079
rect 10652 2053 10662 2079
rect 10608 2041 10662 2053
rect 10708 2087 10762 2193
rect 10808 2227 10862 2239
rect 10808 2201 10818 2227
rect 10852 2201 10862 2227
rect 10808 2149 10809 2201
rect 10861 2149 10862 2201
rect 10808 2142 10862 2149
rect 10908 2227 10962 2333
rect 11008 2411 11062 2418
rect 11008 2359 11009 2411
rect 11061 2359 11062 2411
rect 11008 2333 11018 2359
rect 11052 2333 11062 2359
rect 11008 2321 11062 2333
rect 11108 2367 11162 2563
rect 11208 2597 11262 2609
rect 11208 2571 11218 2597
rect 11252 2571 11262 2597
rect 11208 2519 11209 2571
rect 11261 2519 11262 2571
rect 11208 2512 11262 2519
rect 11308 2597 11362 2703
rect 11408 2781 11462 2788
rect 11408 2729 11409 2781
rect 11461 2729 11462 2781
rect 11408 2703 11418 2729
rect 11452 2703 11462 2729
rect 11408 2691 11462 2703
rect 11508 2737 11562 2843
rect 11608 2877 11662 2889
rect 11608 2851 11618 2877
rect 11652 2851 11662 2877
rect 11608 2799 11609 2851
rect 11661 2799 11662 2851
rect 11608 2792 11662 2799
rect 11708 2877 11762 2983
rect 11808 3061 11862 3068
rect 11808 3009 11809 3061
rect 11861 3009 11862 3061
rect 11808 2983 11818 3009
rect 11852 2983 11862 3009
rect 11808 2971 11862 2983
rect 11908 3017 11962 3123
rect 12008 3157 12062 3169
rect 12008 3131 12018 3157
rect 12052 3131 12062 3157
rect 12008 3079 12009 3131
rect 12061 3079 12062 3131
rect 12008 3072 12062 3079
rect 12108 3157 12162 3263
rect 12208 3341 12262 3348
rect 12208 3289 12209 3341
rect 12261 3289 12262 3341
rect 12208 3263 12218 3289
rect 12252 3263 12262 3289
rect 12208 3251 12262 3263
rect 12308 3297 12362 3403
rect 12408 3437 12462 3449
rect 12408 3411 12418 3437
rect 12452 3411 12462 3437
rect 12408 3359 12409 3411
rect 12461 3359 12462 3411
rect 12408 3352 12462 3359
rect 12508 3437 12562 3543
rect 12608 3621 12662 3628
rect 12608 3569 12609 3621
rect 12661 3569 12662 3621
rect 12608 3543 12618 3569
rect 12652 3543 12662 3569
rect 12608 3531 12662 3543
rect 12708 3577 12762 3773
rect 12808 3807 12862 3819
rect 12808 3781 12818 3807
rect 12852 3781 12862 3807
rect 12808 3729 12809 3781
rect 12861 3729 12862 3781
rect 12808 3722 12862 3729
rect 12906 3788 12916 3822
rect 12950 3788 12960 3822
rect 12906 3781 12960 3788
rect 12906 3729 12907 3781
rect 12959 3729 12960 3781
rect 12906 3722 12960 3729
rect 12990 3687 13020 4851
rect 12904 3681 13020 3687
rect 12904 3647 12916 3681
rect 12950 3647 13020 3681
rect 12904 3641 13020 3647
rect 12906 3592 12960 3604
rect 12708 3543 12718 3577
rect 12752 3543 12762 3577
rect 12508 3403 12518 3437
rect 12552 3403 12562 3437
rect 12308 3263 12318 3297
rect 12352 3263 12362 3297
rect 12108 3123 12118 3157
rect 12152 3123 12162 3157
rect 11908 2983 11918 3017
rect 11952 2983 11962 3017
rect 11708 2843 11718 2877
rect 11752 2843 11762 2877
rect 11508 2703 11518 2737
rect 11552 2703 11562 2737
rect 11308 2563 11318 2597
rect 11352 2563 11362 2597
rect 11202 2483 11268 2484
rect 11202 2431 11209 2483
rect 11261 2431 11268 2483
rect 11202 2430 11268 2431
rect 11108 2333 11118 2367
rect 11152 2333 11162 2367
rect 10908 2193 10918 2227
rect 10952 2193 10962 2227
rect 10708 2053 10718 2087
rect 10752 2053 10762 2087
rect 10508 1913 10518 1947
rect 10552 1913 10562 1947
rect 10308 1773 10318 1807
rect 10352 1773 10362 1807
rect 10108 1633 10118 1667
rect 10152 1633 10162 1667
rect 9908 1493 9918 1527
rect 9952 1493 9962 1527
rect 9708 1353 9718 1387
rect 9752 1353 9762 1387
rect 9602 1273 9668 1274
rect 9602 1221 9609 1273
rect 9661 1221 9668 1273
rect 9602 1220 9668 1221
rect 9508 1123 9518 1157
rect 9552 1123 9562 1157
rect 9308 983 9318 1017
rect 9352 983 9362 1017
rect 9108 843 9118 877
rect 9152 843 9162 877
rect 8908 703 8918 737
rect 8952 703 8962 737
rect 8708 563 8718 597
rect 8752 563 8762 597
rect 8508 423 8518 457
rect 8552 423 8562 457
rect 8308 283 8318 317
rect 8352 283 8362 317
rect 8108 143 8118 177
rect 8152 143 8162 177
rect 8002 63 8068 64
rect 8002 11 8009 63
rect 8061 11 8068 63
rect 8002 10 8068 11
rect 7908 -67 7909 -15
rect 7961 -67 7962 -15
rect 7908 -79 7918 -67
rect 7952 -79 7962 -67
rect 7708 -132 7762 -131
rect 7708 -143 7718 -132
rect 7752 -143 7762 -132
rect 7708 -195 7709 -143
rect 7761 -195 7762 -143
rect 7708 -210 7762 -195
rect 7812 -133 7858 -81
rect 7812 -167 7818 -133
rect 7852 -167 7858 -133
rect 7718 -291 7725 -239
rect 7777 -291 7784 -239
rect 7612 -397 7618 -363
rect 7652 -397 7658 -363
rect 7612 -435 7658 -397
rect 7612 -469 7618 -435
rect 7652 -469 7658 -435
rect 7612 -512 7658 -469
rect 7709 -326 7761 -320
rect 7709 -390 7718 -378
rect 7752 -390 7761 -378
rect 7709 -454 7718 -442
rect 7752 -454 7761 -442
rect 7709 -512 7761 -506
rect 7812 -363 7858 -167
rect 7908 -131 7909 -79
rect 7961 -131 7962 -79
rect 8008 -22 8062 10
rect 8008 -74 8009 -22
rect 8061 -74 8062 -22
rect 8008 -81 8062 -74
rect 8108 -15 8162 143
rect 8208 221 8262 228
rect 8208 169 8209 221
rect 8261 169 8262 221
rect 8208 143 8218 169
rect 8252 143 8262 169
rect 8208 131 8262 143
rect 8308 177 8362 283
rect 8408 317 8462 329
rect 8408 291 8418 317
rect 8452 291 8462 317
rect 8408 239 8409 291
rect 8461 239 8462 291
rect 8408 232 8462 239
rect 8508 317 8562 423
rect 8608 501 8662 508
rect 8608 449 8609 501
rect 8661 449 8662 501
rect 8608 423 8618 449
rect 8652 423 8662 449
rect 8608 411 8662 423
rect 8708 457 8762 563
rect 8808 597 8862 609
rect 8808 571 8818 597
rect 8852 571 8862 597
rect 8808 519 8809 571
rect 8861 519 8862 571
rect 8808 512 8862 519
rect 8908 597 8962 703
rect 9008 781 9062 788
rect 9008 729 9009 781
rect 9061 729 9062 781
rect 9008 703 9018 729
rect 9052 703 9062 729
rect 9008 691 9062 703
rect 9108 737 9162 843
rect 9208 877 9262 889
rect 9208 851 9218 877
rect 9252 851 9262 877
rect 9208 799 9209 851
rect 9261 799 9262 851
rect 9208 792 9262 799
rect 9308 877 9362 983
rect 9408 1061 9462 1068
rect 9408 1009 9409 1061
rect 9461 1009 9462 1061
rect 9408 983 9418 1009
rect 9452 983 9462 1009
rect 9408 971 9462 983
rect 9508 1017 9562 1123
rect 9608 1157 9662 1169
rect 9608 1131 9618 1157
rect 9652 1131 9662 1157
rect 9608 1079 9609 1131
rect 9661 1079 9662 1131
rect 9608 1072 9662 1079
rect 9708 1157 9762 1353
rect 9808 1431 9862 1438
rect 9808 1379 9809 1431
rect 9861 1379 9862 1431
rect 9808 1353 9818 1379
rect 9852 1353 9862 1379
rect 9808 1341 9862 1353
rect 9908 1387 9962 1493
rect 10008 1527 10062 1539
rect 10008 1501 10018 1527
rect 10052 1501 10062 1527
rect 10008 1449 10009 1501
rect 10061 1449 10062 1501
rect 10008 1442 10062 1449
rect 10108 1527 10162 1633
rect 10208 1711 10262 1718
rect 10208 1659 10209 1711
rect 10261 1659 10262 1711
rect 10208 1633 10218 1659
rect 10252 1633 10262 1659
rect 10208 1621 10262 1633
rect 10308 1667 10362 1773
rect 10408 1807 10462 1819
rect 10408 1781 10418 1807
rect 10452 1781 10462 1807
rect 10408 1729 10409 1781
rect 10461 1729 10462 1781
rect 10408 1722 10462 1729
rect 10508 1807 10562 1913
rect 10608 1991 10662 1998
rect 10608 1939 10609 1991
rect 10661 1939 10662 1991
rect 10608 1913 10618 1939
rect 10652 1913 10662 1939
rect 10608 1901 10662 1913
rect 10708 1947 10762 2053
rect 10808 2087 10862 2099
rect 10808 2061 10818 2087
rect 10852 2061 10862 2087
rect 10808 2009 10809 2061
rect 10861 2009 10862 2061
rect 10808 2002 10862 2009
rect 10908 2087 10962 2193
rect 11008 2271 11062 2278
rect 11008 2219 11009 2271
rect 11061 2219 11062 2271
rect 11008 2193 11018 2219
rect 11052 2193 11062 2219
rect 11008 2181 11062 2193
rect 11108 2227 11162 2333
rect 11208 2367 11262 2379
rect 11208 2341 11218 2367
rect 11252 2341 11262 2367
rect 11208 2289 11209 2341
rect 11261 2289 11262 2341
rect 11208 2282 11262 2289
rect 11308 2367 11362 2563
rect 11408 2641 11462 2648
rect 11408 2589 11409 2641
rect 11461 2589 11462 2641
rect 11408 2563 11418 2589
rect 11452 2563 11462 2589
rect 11408 2551 11462 2563
rect 11508 2597 11562 2703
rect 11608 2737 11662 2749
rect 11608 2711 11618 2737
rect 11652 2711 11662 2737
rect 11608 2659 11609 2711
rect 11661 2659 11662 2711
rect 11608 2652 11662 2659
rect 11708 2737 11762 2843
rect 11808 2921 11862 2928
rect 11808 2869 11809 2921
rect 11861 2869 11862 2921
rect 11808 2843 11818 2869
rect 11852 2843 11862 2869
rect 11808 2831 11862 2843
rect 11908 2877 11962 2983
rect 12008 3017 12062 3029
rect 12008 2991 12018 3017
rect 12052 2991 12062 3017
rect 12008 2939 12009 2991
rect 12061 2939 12062 2991
rect 12008 2932 12062 2939
rect 12108 3017 12162 3123
rect 12208 3201 12262 3208
rect 12208 3149 12209 3201
rect 12261 3149 12262 3201
rect 12208 3123 12218 3149
rect 12252 3123 12262 3149
rect 12208 3111 12262 3123
rect 12308 3157 12362 3263
rect 12408 3297 12462 3309
rect 12408 3271 12418 3297
rect 12452 3271 12462 3297
rect 12408 3219 12409 3271
rect 12461 3219 12462 3271
rect 12408 3212 12462 3219
rect 12508 3297 12562 3403
rect 12608 3481 12662 3488
rect 12608 3429 12609 3481
rect 12661 3429 12662 3481
rect 12608 3403 12618 3429
rect 12652 3403 12662 3429
rect 12608 3391 12662 3403
rect 12708 3437 12762 3543
rect 12808 3577 12862 3589
rect 12808 3551 12818 3577
rect 12852 3551 12862 3577
rect 12808 3499 12809 3551
rect 12861 3499 12862 3551
rect 12808 3492 12862 3499
rect 12906 3558 12916 3592
rect 12950 3558 12960 3592
rect 12906 3551 12960 3558
rect 12906 3499 12907 3551
rect 12959 3499 12960 3551
rect 12906 3492 12960 3499
rect 12906 3452 12960 3464
rect 12708 3403 12718 3437
rect 12752 3403 12762 3437
rect 12508 3263 12518 3297
rect 12552 3263 12562 3297
rect 12308 3123 12318 3157
rect 12352 3123 12362 3157
rect 12108 2983 12118 3017
rect 12152 2983 12162 3017
rect 11908 2843 11918 2877
rect 11952 2843 11962 2877
rect 11708 2703 11718 2737
rect 11752 2703 11762 2737
rect 11508 2563 11518 2597
rect 11552 2563 11562 2597
rect 11402 2499 11468 2500
rect 11402 2447 11409 2499
rect 11461 2447 11468 2499
rect 11402 2446 11468 2447
rect 11308 2333 11318 2367
rect 11352 2333 11362 2367
rect 11108 2193 11118 2227
rect 11152 2193 11162 2227
rect 10908 2053 10918 2087
rect 10952 2053 10962 2087
rect 10708 1913 10718 1947
rect 10752 1913 10762 1947
rect 10508 1773 10518 1807
rect 10552 1773 10562 1807
rect 10308 1633 10318 1667
rect 10352 1633 10362 1667
rect 10108 1493 10118 1527
rect 10152 1493 10162 1527
rect 9908 1353 9918 1387
rect 9952 1353 9962 1387
rect 9802 1289 9868 1290
rect 9802 1237 9809 1289
rect 9861 1237 9868 1289
rect 9802 1236 9868 1237
rect 9708 1123 9718 1157
rect 9752 1123 9762 1157
rect 9508 983 9518 1017
rect 9552 983 9562 1017
rect 9308 843 9318 877
rect 9352 843 9362 877
rect 9108 703 9118 737
rect 9152 703 9162 737
rect 8908 563 8918 597
rect 8952 563 8962 597
rect 8708 423 8718 457
rect 8752 423 8762 457
rect 8508 283 8518 317
rect 8552 283 8562 317
rect 8308 143 8318 177
rect 8352 143 8362 177
rect 8202 79 8268 80
rect 8202 27 8209 79
rect 8261 27 8268 79
rect 8202 26 8268 27
rect 8108 -67 8109 -15
rect 8161 -67 8162 -15
rect 8108 -79 8118 -67
rect 8152 -79 8162 -67
rect 7908 -132 7962 -131
rect 7908 -143 7918 -132
rect 7952 -143 7962 -132
rect 7908 -195 7909 -143
rect 7961 -195 7962 -143
rect 7908 -210 7962 -195
rect 8012 -133 8058 -81
rect 8012 -167 8018 -133
rect 8052 -167 8058 -133
rect 7918 -291 7925 -239
rect 7977 -291 7984 -239
rect 7812 -397 7818 -363
rect 7852 -397 7858 -363
rect 7812 -435 7858 -397
rect 7812 -469 7818 -435
rect 7852 -469 7858 -435
rect 7812 -512 7858 -469
rect 7909 -326 7961 -320
rect 7909 -390 7918 -378
rect 7952 -390 7961 -378
rect 7909 -454 7918 -442
rect 7952 -454 7961 -442
rect 7909 -555 7961 -506
rect 8012 -363 8058 -167
rect 8108 -131 8109 -79
rect 8161 -131 8162 -79
rect 8208 -22 8262 26
rect 8208 -74 8209 -22
rect 8261 -74 8262 -22
rect 8208 -81 8262 -74
rect 8308 -15 8362 143
rect 8408 177 8462 189
rect 8408 151 8418 177
rect 8452 151 8462 177
rect 8408 99 8409 151
rect 8461 99 8462 151
rect 8408 92 8462 99
rect 8508 177 8562 283
rect 8608 361 8662 368
rect 8608 309 8609 361
rect 8661 309 8662 361
rect 8608 283 8618 309
rect 8652 283 8662 309
rect 8608 271 8662 283
rect 8708 317 8762 423
rect 8808 457 8862 469
rect 8808 431 8818 457
rect 8852 431 8862 457
rect 8808 379 8809 431
rect 8861 379 8862 431
rect 8808 372 8862 379
rect 8908 457 8962 563
rect 9008 641 9062 648
rect 9008 589 9009 641
rect 9061 589 9062 641
rect 9008 563 9018 589
rect 9052 563 9062 589
rect 9008 551 9062 563
rect 9108 597 9162 703
rect 9208 737 9262 749
rect 9208 711 9218 737
rect 9252 711 9262 737
rect 9208 659 9209 711
rect 9261 659 9262 711
rect 9208 652 9262 659
rect 9308 737 9362 843
rect 9408 921 9462 928
rect 9408 869 9409 921
rect 9461 869 9462 921
rect 9408 843 9418 869
rect 9452 843 9462 869
rect 9408 831 9462 843
rect 9508 877 9562 983
rect 9608 1017 9662 1029
rect 9608 991 9618 1017
rect 9652 991 9662 1017
rect 9608 939 9609 991
rect 9661 939 9662 991
rect 9608 932 9662 939
rect 9708 1017 9762 1123
rect 9808 1201 9862 1208
rect 9808 1149 9809 1201
rect 9861 1149 9862 1201
rect 9808 1123 9818 1149
rect 9852 1123 9862 1149
rect 9808 1111 9862 1123
rect 9908 1157 9962 1353
rect 10008 1387 10062 1399
rect 10008 1361 10018 1387
rect 10052 1361 10062 1387
rect 10008 1309 10009 1361
rect 10061 1309 10062 1361
rect 10008 1302 10062 1309
rect 10108 1387 10162 1493
rect 10208 1571 10262 1578
rect 10208 1519 10209 1571
rect 10261 1519 10262 1571
rect 10208 1493 10218 1519
rect 10252 1493 10262 1519
rect 10208 1481 10262 1493
rect 10308 1527 10362 1633
rect 10408 1667 10462 1679
rect 10408 1641 10418 1667
rect 10452 1641 10462 1667
rect 10408 1589 10409 1641
rect 10461 1589 10462 1641
rect 10408 1582 10462 1589
rect 10508 1667 10562 1773
rect 10608 1851 10662 1858
rect 10608 1799 10609 1851
rect 10661 1799 10662 1851
rect 10608 1773 10618 1799
rect 10652 1773 10662 1799
rect 10608 1761 10662 1773
rect 10708 1807 10762 1913
rect 10808 1947 10862 1959
rect 10808 1921 10818 1947
rect 10852 1921 10862 1947
rect 10808 1869 10809 1921
rect 10861 1869 10862 1921
rect 10808 1862 10862 1869
rect 10908 1947 10962 2053
rect 11008 2131 11062 2138
rect 11008 2079 11009 2131
rect 11061 2079 11062 2131
rect 11008 2053 11018 2079
rect 11052 2053 11062 2079
rect 11008 2041 11062 2053
rect 11108 2087 11162 2193
rect 11208 2227 11262 2239
rect 11208 2201 11218 2227
rect 11252 2201 11262 2227
rect 11208 2149 11209 2201
rect 11261 2149 11262 2201
rect 11208 2142 11262 2149
rect 11308 2227 11362 2333
rect 11408 2411 11462 2418
rect 11408 2359 11409 2411
rect 11461 2359 11462 2411
rect 11408 2333 11418 2359
rect 11452 2333 11462 2359
rect 11408 2321 11462 2333
rect 11508 2367 11562 2563
rect 11608 2597 11662 2609
rect 11608 2571 11618 2597
rect 11652 2571 11662 2597
rect 11608 2519 11609 2571
rect 11661 2519 11662 2571
rect 11608 2512 11662 2519
rect 11708 2597 11762 2703
rect 11808 2781 11862 2788
rect 11808 2729 11809 2781
rect 11861 2729 11862 2781
rect 11808 2703 11818 2729
rect 11852 2703 11862 2729
rect 11808 2691 11862 2703
rect 11908 2737 11962 2843
rect 12008 2877 12062 2889
rect 12008 2851 12018 2877
rect 12052 2851 12062 2877
rect 12008 2799 12009 2851
rect 12061 2799 12062 2851
rect 12008 2792 12062 2799
rect 12108 2877 12162 2983
rect 12208 3061 12262 3068
rect 12208 3009 12209 3061
rect 12261 3009 12262 3061
rect 12208 2983 12218 3009
rect 12252 2983 12262 3009
rect 12208 2971 12262 2983
rect 12308 3017 12362 3123
rect 12408 3157 12462 3169
rect 12408 3131 12418 3157
rect 12452 3131 12462 3157
rect 12408 3079 12409 3131
rect 12461 3079 12462 3131
rect 12408 3072 12462 3079
rect 12508 3157 12562 3263
rect 12608 3341 12662 3348
rect 12608 3289 12609 3341
rect 12661 3289 12662 3341
rect 12608 3263 12618 3289
rect 12652 3263 12662 3289
rect 12608 3251 12662 3263
rect 12708 3297 12762 3403
rect 12808 3437 12862 3449
rect 12808 3411 12818 3437
rect 12852 3411 12862 3437
rect 12808 3359 12809 3411
rect 12861 3359 12862 3411
rect 12808 3352 12862 3359
rect 12906 3418 12916 3452
rect 12950 3418 12960 3452
rect 12906 3411 12960 3418
rect 12906 3359 12907 3411
rect 12959 3359 12960 3411
rect 12906 3352 12960 3359
rect 12906 3312 12960 3324
rect 12708 3263 12718 3297
rect 12752 3263 12762 3297
rect 12508 3123 12518 3157
rect 12552 3123 12562 3157
rect 12308 2983 12318 3017
rect 12352 2983 12362 3017
rect 12108 2843 12118 2877
rect 12152 2843 12162 2877
rect 11908 2703 11918 2737
rect 11952 2703 11962 2737
rect 11708 2563 11718 2597
rect 11752 2563 11762 2597
rect 11602 2483 11668 2484
rect 11602 2431 11609 2483
rect 11661 2431 11668 2483
rect 11602 2430 11668 2431
rect 11508 2333 11518 2367
rect 11552 2333 11562 2367
rect 11308 2193 11318 2227
rect 11352 2193 11362 2227
rect 11108 2053 11118 2087
rect 11152 2053 11162 2087
rect 10908 1913 10918 1947
rect 10952 1913 10962 1947
rect 10708 1773 10718 1807
rect 10752 1773 10762 1807
rect 10508 1633 10518 1667
rect 10552 1633 10562 1667
rect 10308 1493 10318 1527
rect 10352 1493 10362 1527
rect 10108 1353 10118 1387
rect 10152 1353 10162 1387
rect 10002 1273 10068 1274
rect 10002 1221 10009 1273
rect 10061 1221 10068 1273
rect 10002 1220 10068 1221
rect 9908 1123 9918 1157
rect 9952 1123 9962 1157
rect 9708 983 9718 1017
rect 9752 983 9762 1017
rect 9508 843 9518 877
rect 9552 843 9562 877
rect 9308 703 9318 737
rect 9352 703 9362 737
rect 9108 563 9118 597
rect 9152 563 9162 597
rect 8908 423 8918 457
rect 8952 423 8962 457
rect 8708 283 8718 317
rect 8752 283 8762 317
rect 8508 143 8518 177
rect 8552 143 8562 177
rect 8402 63 8468 64
rect 8402 11 8409 63
rect 8461 11 8468 63
rect 8402 10 8468 11
rect 8308 -67 8309 -15
rect 8361 -67 8362 -15
rect 8308 -79 8318 -67
rect 8352 -79 8362 -67
rect 8108 -132 8162 -131
rect 8108 -143 8118 -132
rect 8152 -143 8162 -132
rect 8108 -195 8109 -143
rect 8161 -195 8162 -143
rect 8108 -210 8162 -195
rect 8212 -133 8258 -81
rect 8212 -167 8218 -133
rect 8252 -167 8258 -133
rect 8118 -291 8125 -239
rect 8177 -291 8184 -239
rect 8012 -397 8018 -363
rect 8052 -397 8058 -363
rect 8012 -435 8058 -397
rect 8012 -469 8018 -435
rect 8052 -469 8058 -435
rect 8012 -512 8058 -469
rect 8109 -326 8161 -320
rect 8109 -390 8118 -378
rect 8152 -390 8161 -378
rect 8109 -454 8118 -442
rect 8152 -454 8161 -442
rect 8109 -512 8161 -506
rect 8212 -363 8258 -167
rect 8308 -131 8309 -79
rect 8361 -131 8362 -79
rect 8408 -22 8462 10
rect 8408 -74 8409 -22
rect 8461 -74 8462 -22
rect 8408 -81 8462 -74
rect 8508 -15 8562 143
rect 8608 221 8662 228
rect 8608 169 8609 221
rect 8661 169 8662 221
rect 8608 143 8618 169
rect 8652 143 8662 169
rect 8608 131 8662 143
rect 8708 177 8762 283
rect 8808 317 8862 329
rect 8808 291 8818 317
rect 8852 291 8862 317
rect 8808 239 8809 291
rect 8861 239 8862 291
rect 8808 232 8862 239
rect 8908 317 8962 423
rect 9008 501 9062 508
rect 9008 449 9009 501
rect 9061 449 9062 501
rect 9008 423 9018 449
rect 9052 423 9062 449
rect 9008 411 9062 423
rect 9108 457 9162 563
rect 9208 597 9262 609
rect 9208 571 9218 597
rect 9252 571 9262 597
rect 9208 519 9209 571
rect 9261 519 9262 571
rect 9208 512 9262 519
rect 9308 597 9362 703
rect 9408 781 9462 788
rect 9408 729 9409 781
rect 9461 729 9462 781
rect 9408 703 9418 729
rect 9452 703 9462 729
rect 9408 691 9462 703
rect 9508 737 9562 843
rect 9608 877 9662 889
rect 9608 851 9618 877
rect 9652 851 9662 877
rect 9608 799 9609 851
rect 9661 799 9662 851
rect 9608 792 9662 799
rect 9708 877 9762 983
rect 9808 1061 9862 1068
rect 9808 1009 9809 1061
rect 9861 1009 9862 1061
rect 9808 983 9818 1009
rect 9852 983 9862 1009
rect 9808 971 9862 983
rect 9908 1017 9962 1123
rect 10008 1157 10062 1169
rect 10008 1131 10018 1157
rect 10052 1131 10062 1157
rect 10008 1079 10009 1131
rect 10061 1079 10062 1131
rect 10008 1072 10062 1079
rect 10108 1157 10162 1353
rect 10208 1431 10262 1438
rect 10208 1379 10209 1431
rect 10261 1379 10262 1431
rect 10208 1353 10218 1379
rect 10252 1353 10262 1379
rect 10208 1341 10262 1353
rect 10308 1387 10362 1493
rect 10408 1527 10462 1539
rect 10408 1501 10418 1527
rect 10452 1501 10462 1527
rect 10408 1449 10409 1501
rect 10461 1449 10462 1501
rect 10408 1442 10462 1449
rect 10508 1527 10562 1633
rect 10608 1711 10662 1718
rect 10608 1659 10609 1711
rect 10661 1659 10662 1711
rect 10608 1633 10618 1659
rect 10652 1633 10662 1659
rect 10608 1621 10662 1633
rect 10708 1667 10762 1773
rect 10808 1807 10862 1819
rect 10808 1781 10818 1807
rect 10852 1781 10862 1807
rect 10808 1729 10809 1781
rect 10861 1729 10862 1781
rect 10808 1722 10862 1729
rect 10908 1807 10962 1913
rect 11008 1991 11062 1998
rect 11008 1939 11009 1991
rect 11061 1939 11062 1991
rect 11008 1913 11018 1939
rect 11052 1913 11062 1939
rect 11008 1901 11062 1913
rect 11108 1947 11162 2053
rect 11208 2087 11262 2099
rect 11208 2061 11218 2087
rect 11252 2061 11262 2087
rect 11208 2009 11209 2061
rect 11261 2009 11262 2061
rect 11208 2002 11262 2009
rect 11308 2087 11362 2193
rect 11408 2271 11462 2278
rect 11408 2219 11409 2271
rect 11461 2219 11462 2271
rect 11408 2193 11418 2219
rect 11452 2193 11462 2219
rect 11408 2181 11462 2193
rect 11508 2227 11562 2333
rect 11608 2367 11662 2379
rect 11608 2341 11618 2367
rect 11652 2341 11662 2367
rect 11608 2289 11609 2341
rect 11661 2289 11662 2341
rect 11608 2282 11662 2289
rect 11708 2367 11762 2563
rect 11808 2641 11862 2648
rect 11808 2589 11809 2641
rect 11861 2589 11862 2641
rect 11808 2563 11818 2589
rect 11852 2563 11862 2589
rect 11808 2551 11862 2563
rect 11908 2597 11962 2703
rect 12008 2737 12062 2749
rect 12008 2711 12018 2737
rect 12052 2711 12062 2737
rect 12008 2659 12009 2711
rect 12061 2659 12062 2711
rect 12008 2652 12062 2659
rect 12108 2737 12162 2843
rect 12208 2921 12262 2928
rect 12208 2869 12209 2921
rect 12261 2869 12262 2921
rect 12208 2843 12218 2869
rect 12252 2843 12262 2869
rect 12208 2831 12262 2843
rect 12308 2877 12362 2983
rect 12408 3017 12462 3029
rect 12408 2991 12418 3017
rect 12452 2991 12462 3017
rect 12408 2939 12409 2991
rect 12461 2939 12462 2991
rect 12408 2932 12462 2939
rect 12508 3017 12562 3123
rect 12608 3201 12662 3208
rect 12608 3149 12609 3201
rect 12661 3149 12662 3201
rect 12608 3123 12618 3149
rect 12652 3123 12662 3149
rect 12608 3111 12662 3123
rect 12708 3157 12762 3263
rect 12808 3297 12862 3309
rect 12808 3271 12818 3297
rect 12852 3271 12862 3297
rect 12808 3219 12809 3271
rect 12861 3219 12862 3271
rect 12808 3212 12862 3219
rect 12906 3278 12916 3312
rect 12950 3278 12960 3312
rect 12906 3271 12960 3278
rect 12906 3219 12907 3271
rect 12959 3219 12960 3271
rect 12906 3212 12960 3219
rect 12906 3172 12960 3184
rect 12708 3123 12718 3157
rect 12752 3123 12762 3157
rect 12508 2983 12518 3017
rect 12552 2983 12562 3017
rect 12308 2843 12318 2877
rect 12352 2843 12362 2877
rect 12108 2703 12118 2737
rect 12152 2703 12162 2737
rect 11908 2563 11918 2597
rect 11952 2563 11962 2597
rect 11802 2499 11868 2500
rect 11802 2447 11809 2499
rect 11861 2447 11868 2499
rect 11802 2446 11868 2447
rect 11708 2333 11718 2367
rect 11752 2333 11762 2367
rect 11508 2193 11518 2227
rect 11552 2193 11562 2227
rect 11308 2053 11318 2087
rect 11352 2053 11362 2087
rect 11108 1913 11118 1947
rect 11152 1913 11162 1947
rect 10908 1773 10918 1807
rect 10952 1773 10962 1807
rect 10708 1633 10718 1667
rect 10752 1633 10762 1667
rect 10508 1493 10518 1527
rect 10552 1493 10562 1527
rect 10308 1353 10318 1387
rect 10352 1353 10362 1387
rect 10202 1289 10268 1290
rect 10202 1237 10209 1289
rect 10261 1237 10268 1289
rect 10202 1236 10268 1237
rect 10108 1123 10118 1157
rect 10152 1123 10162 1157
rect 9908 983 9918 1017
rect 9952 983 9962 1017
rect 9708 843 9718 877
rect 9752 843 9762 877
rect 9508 703 9518 737
rect 9552 703 9562 737
rect 9308 563 9318 597
rect 9352 563 9362 597
rect 9108 423 9118 457
rect 9152 423 9162 457
rect 8908 283 8918 317
rect 8952 283 8962 317
rect 8708 143 8718 177
rect 8752 143 8762 177
rect 8602 79 8668 80
rect 8602 27 8609 79
rect 8661 27 8668 79
rect 8602 26 8668 27
rect 8508 -67 8509 -15
rect 8561 -67 8562 -15
rect 8508 -79 8518 -67
rect 8552 -79 8562 -67
rect 8308 -132 8362 -131
rect 8308 -143 8318 -132
rect 8352 -143 8362 -132
rect 8308 -195 8309 -143
rect 8361 -195 8362 -143
rect 8308 -210 8362 -195
rect 8412 -133 8458 -81
rect 8412 -167 8418 -133
rect 8452 -167 8458 -133
rect 8318 -291 8325 -239
rect 8377 -291 8384 -239
rect 8212 -397 8218 -363
rect 8252 -397 8258 -363
rect 8212 -435 8258 -397
rect 8212 -469 8218 -435
rect 8252 -469 8258 -435
rect 8212 -512 8258 -469
rect 8309 -326 8361 -320
rect 8309 -390 8318 -378
rect 8352 -390 8361 -378
rect 8309 -454 8318 -442
rect 8352 -454 8361 -442
rect 8309 -555 8361 -506
rect 8412 -363 8458 -167
rect 8508 -131 8509 -79
rect 8561 -131 8562 -79
rect 8608 -22 8662 26
rect 8608 -74 8609 -22
rect 8661 -74 8662 -22
rect 8608 -81 8662 -74
rect 8708 -15 8762 143
rect 8808 177 8862 189
rect 8808 151 8818 177
rect 8852 151 8862 177
rect 8808 99 8809 151
rect 8861 99 8862 151
rect 8808 92 8862 99
rect 8908 177 8962 283
rect 9008 361 9062 368
rect 9008 309 9009 361
rect 9061 309 9062 361
rect 9008 283 9018 309
rect 9052 283 9062 309
rect 9008 271 9062 283
rect 9108 317 9162 423
rect 9208 457 9262 469
rect 9208 431 9218 457
rect 9252 431 9262 457
rect 9208 379 9209 431
rect 9261 379 9262 431
rect 9208 372 9262 379
rect 9308 457 9362 563
rect 9408 641 9462 648
rect 9408 589 9409 641
rect 9461 589 9462 641
rect 9408 563 9418 589
rect 9452 563 9462 589
rect 9408 551 9462 563
rect 9508 597 9562 703
rect 9608 737 9662 749
rect 9608 711 9618 737
rect 9652 711 9662 737
rect 9608 659 9609 711
rect 9661 659 9662 711
rect 9608 652 9662 659
rect 9708 737 9762 843
rect 9808 921 9862 928
rect 9808 869 9809 921
rect 9861 869 9862 921
rect 9808 843 9818 869
rect 9852 843 9862 869
rect 9808 831 9862 843
rect 9908 877 9962 983
rect 10008 1017 10062 1029
rect 10008 991 10018 1017
rect 10052 991 10062 1017
rect 10008 939 10009 991
rect 10061 939 10062 991
rect 10008 932 10062 939
rect 10108 1017 10162 1123
rect 10208 1201 10262 1208
rect 10208 1149 10209 1201
rect 10261 1149 10262 1201
rect 10208 1123 10218 1149
rect 10252 1123 10262 1149
rect 10208 1111 10262 1123
rect 10308 1157 10362 1353
rect 10408 1387 10462 1399
rect 10408 1361 10418 1387
rect 10452 1361 10462 1387
rect 10408 1309 10409 1361
rect 10461 1309 10462 1361
rect 10408 1302 10462 1309
rect 10508 1387 10562 1493
rect 10608 1571 10662 1578
rect 10608 1519 10609 1571
rect 10661 1519 10662 1571
rect 10608 1493 10618 1519
rect 10652 1493 10662 1519
rect 10608 1481 10662 1493
rect 10708 1527 10762 1633
rect 10808 1667 10862 1679
rect 10808 1641 10818 1667
rect 10852 1641 10862 1667
rect 10808 1589 10809 1641
rect 10861 1589 10862 1641
rect 10808 1582 10862 1589
rect 10908 1667 10962 1773
rect 11008 1851 11062 1858
rect 11008 1799 11009 1851
rect 11061 1799 11062 1851
rect 11008 1773 11018 1799
rect 11052 1773 11062 1799
rect 11008 1761 11062 1773
rect 11108 1807 11162 1913
rect 11208 1947 11262 1959
rect 11208 1921 11218 1947
rect 11252 1921 11262 1947
rect 11208 1869 11209 1921
rect 11261 1869 11262 1921
rect 11208 1862 11262 1869
rect 11308 1947 11362 2053
rect 11408 2131 11462 2138
rect 11408 2079 11409 2131
rect 11461 2079 11462 2131
rect 11408 2053 11418 2079
rect 11452 2053 11462 2079
rect 11408 2041 11462 2053
rect 11508 2087 11562 2193
rect 11608 2227 11662 2239
rect 11608 2201 11618 2227
rect 11652 2201 11662 2227
rect 11608 2149 11609 2201
rect 11661 2149 11662 2201
rect 11608 2142 11662 2149
rect 11708 2227 11762 2333
rect 11808 2411 11862 2418
rect 11808 2359 11809 2411
rect 11861 2359 11862 2411
rect 11808 2333 11818 2359
rect 11852 2333 11862 2359
rect 11808 2321 11862 2333
rect 11908 2367 11962 2563
rect 12008 2597 12062 2609
rect 12008 2571 12018 2597
rect 12052 2571 12062 2597
rect 12008 2519 12009 2571
rect 12061 2519 12062 2571
rect 12008 2512 12062 2519
rect 12108 2597 12162 2703
rect 12208 2781 12262 2788
rect 12208 2729 12209 2781
rect 12261 2729 12262 2781
rect 12208 2703 12218 2729
rect 12252 2703 12262 2729
rect 12208 2691 12262 2703
rect 12308 2737 12362 2843
rect 12408 2877 12462 2889
rect 12408 2851 12418 2877
rect 12452 2851 12462 2877
rect 12408 2799 12409 2851
rect 12461 2799 12462 2851
rect 12408 2792 12462 2799
rect 12508 2877 12562 2983
rect 12608 3061 12662 3068
rect 12608 3009 12609 3061
rect 12661 3009 12662 3061
rect 12608 2983 12618 3009
rect 12652 2983 12662 3009
rect 12608 2971 12662 2983
rect 12708 3017 12762 3123
rect 12808 3157 12862 3169
rect 12808 3131 12818 3157
rect 12852 3131 12862 3157
rect 12808 3079 12809 3131
rect 12861 3079 12862 3131
rect 12808 3072 12862 3079
rect 12906 3138 12916 3172
rect 12950 3138 12960 3172
rect 12906 3131 12960 3138
rect 12906 3079 12907 3131
rect 12959 3079 12960 3131
rect 12906 3072 12960 3079
rect 12906 3032 12960 3044
rect 12708 2983 12718 3017
rect 12752 2983 12762 3017
rect 12508 2843 12518 2877
rect 12552 2843 12562 2877
rect 12308 2703 12318 2737
rect 12352 2703 12362 2737
rect 12108 2563 12118 2597
rect 12152 2563 12162 2597
rect 12002 2483 12068 2484
rect 12002 2431 12009 2483
rect 12061 2431 12068 2483
rect 12002 2430 12068 2431
rect 11908 2333 11918 2367
rect 11952 2333 11962 2367
rect 11708 2193 11718 2227
rect 11752 2193 11762 2227
rect 11508 2053 11518 2087
rect 11552 2053 11562 2087
rect 11308 1913 11318 1947
rect 11352 1913 11362 1947
rect 11108 1773 11118 1807
rect 11152 1773 11162 1807
rect 10908 1633 10918 1667
rect 10952 1633 10962 1667
rect 10708 1493 10718 1527
rect 10752 1493 10762 1527
rect 10508 1353 10518 1387
rect 10552 1353 10562 1387
rect 10402 1273 10468 1274
rect 10402 1221 10409 1273
rect 10461 1221 10468 1273
rect 10402 1220 10468 1221
rect 10308 1123 10318 1157
rect 10352 1123 10362 1157
rect 10108 983 10118 1017
rect 10152 983 10162 1017
rect 9908 843 9918 877
rect 9952 843 9962 877
rect 9708 703 9718 737
rect 9752 703 9762 737
rect 9508 563 9518 597
rect 9552 563 9562 597
rect 9308 423 9318 457
rect 9352 423 9362 457
rect 9108 283 9118 317
rect 9152 283 9162 317
rect 8908 143 8918 177
rect 8952 143 8962 177
rect 8802 63 8868 64
rect 8802 11 8809 63
rect 8861 11 8868 63
rect 8802 10 8868 11
rect 8708 -67 8709 -15
rect 8761 -67 8762 -15
rect 8708 -79 8718 -67
rect 8752 -79 8762 -67
rect 8508 -132 8562 -131
rect 8508 -143 8518 -132
rect 8552 -143 8562 -132
rect 8508 -195 8509 -143
rect 8561 -195 8562 -143
rect 8508 -210 8562 -195
rect 8612 -133 8658 -81
rect 8612 -167 8618 -133
rect 8652 -167 8658 -133
rect 8518 -291 8525 -239
rect 8577 -291 8584 -239
rect 8412 -397 8418 -363
rect 8452 -397 8458 -363
rect 8412 -435 8458 -397
rect 8412 -469 8418 -435
rect 8452 -469 8458 -435
rect 8412 -512 8458 -469
rect 8509 -326 8561 -320
rect 8509 -390 8518 -378
rect 8552 -390 8561 -378
rect 8509 -454 8518 -442
rect 8552 -454 8561 -442
rect 8509 -512 8561 -506
rect 8612 -363 8658 -167
rect 8708 -131 8709 -79
rect 8761 -131 8762 -79
rect 8808 -22 8862 10
rect 8808 -74 8809 -22
rect 8861 -74 8862 -22
rect 8808 -81 8862 -74
rect 8908 -15 8962 143
rect 9008 221 9062 228
rect 9008 169 9009 221
rect 9061 169 9062 221
rect 9008 143 9018 169
rect 9052 143 9062 169
rect 9008 131 9062 143
rect 9108 177 9162 283
rect 9208 317 9262 329
rect 9208 291 9218 317
rect 9252 291 9262 317
rect 9208 239 9209 291
rect 9261 239 9262 291
rect 9208 232 9262 239
rect 9308 317 9362 423
rect 9408 501 9462 508
rect 9408 449 9409 501
rect 9461 449 9462 501
rect 9408 423 9418 449
rect 9452 423 9462 449
rect 9408 411 9462 423
rect 9508 457 9562 563
rect 9608 597 9662 609
rect 9608 571 9618 597
rect 9652 571 9662 597
rect 9608 519 9609 571
rect 9661 519 9662 571
rect 9608 512 9662 519
rect 9708 597 9762 703
rect 9808 781 9862 788
rect 9808 729 9809 781
rect 9861 729 9862 781
rect 9808 703 9818 729
rect 9852 703 9862 729
rect 9808 691 9862 703
rect 9908 737 9962 843
rect 10008 877 10062 889
rect 10008 851 10018 877
rect 10052 851 10062 877
rect 10008 799 10009 851
rect 10061 799 10062 851
rect 10008 792 10062 799
rect 10108 877 10162 983
rect 10208 1061 10262 1068
rect 10208 1009 10209 1061
rect 10261 1009 10262 1061
rect 10208 983 10218 1009
rect 10252 983 10262 1009
rect 10208 971 10262 983
rect 10308 1017 10362 1123
rect 10408 1157 10462 1169
rect 10408 1131 10418 1157
rect 10452 1131 10462 1157
rect 10408 1079 10409 1131
rect 10461 1079 10462 1131
rect 10408 1072 10462 1079
rect 10508 1157 10562 1353
rect 10608 1431 10662 1438
rect 10608 1379 10609 1431
rect 10661 1379 10662 1431
rect 10608 1353 10618 1379
rect 10652 1353 10662 1379
rect 10608 1341 10662 1353
rect 10708 1387 10762 1493
rect 10808 1527 10862 1539
rect 10808 1501 10818 1527
rect 10852 1501 10862 1527
rect 10808 1449 10809 1501
rect 10861 1449 10862 1501
rect 10808 1442 10862 1449
rect 10908 1527 10962 1633
rect 11008 1711 11062 1718
rect 11008 1659 11009 1711
rect 11061 1659 11062 1711
rect 11008 1633 11018 1659
rect 11052 1633 11062 1659
rect 11008 1621 11062 1633
rect 11108 1667 11162 1773
rect 11208 1807 11262 1819
rect 11208 1781 11218 1807
rect 11252 1781 11262 1807
rect 11208 1729 11209 1781
rect 11261 1729 11262 1781
rect 11208 1722 11262 1729
rect 11308 1807 11362 1913
rect 11408 1991 11462 1998
rect 11408 1939 11409 1991
rect 11461 1939 11462 1991
rect 11408 1913 11418 1939
rect 11452 1913 11462 1939
rect 11408 1901 11462 1913
rect 11508 1947 11562 2053
rect 11608 2087 11662 2099
rect 11608 2061 11618 2087
rect 11652 2061 11662 2087
rect 11608 2009 11609 2061
rect 11661 2009 11662 2061
rect 11608 2002 11662 2009
rect 11708 2087 11762 2193
rect 11808 2271 11862 2278
rect 11808 2219 11809 2271
rect 11861 2219 11862 2271
rect 11808 2193 11818 2219
rect 11852 2193 11862 2219
rect 11808 2181 11862 2193
rect 11908 2227 11962 2333
rect 12008 2367 12062 2379
rect 12008 2341 12018 2367
rect 12052 2341 12062 2367
rect 12008 2289 12009 2341
rect 12061 2289 12062 2341
rect 12008 2282 12062 2289
rect 12108 2367 12162 2563
rect 12208 2641 12262 2648
rect 12208 2589 12209 2641
rect 12261 2589 12262 2641
rect 12208 2563 12218 2589
rect 12252 2563 12262 2589
rect 12208 2551 12262 2563
rect 12308 2597 12362 2703
rect 12408 2737 12462 2749
rect 12408 2711 12418 2737
rect 12452 2711 12462 2737
rect 12408 2659 12409 2711
rect 12461 2659 12462 2711
rect 12408 2652 12462 2659
rect 12508 2737 12562 2843
rect 12608 2921 12662 2928
rect 12608 2869 12609 2921
rect 12661 2869 12662 2921
rect 12608 2843 12618 2869
rect 12652 2843 12662 2869
rect 12608 2831 12662 2843
rect 12708 2877 12762 2983
rect 12808 3017 12862 3029
rect 12808 2991 12818 3017
rect 12852 2991 12862 3017
rect 12808 2939 12809 2991
rect 12861 2939 12862 2991
rect 12808 2932 12862 2939
rect 12906 2998 12916 3032
rect 12950 2998 12960 3032
rect 12906 2991 12960 2998
rect 12906 2939 12907 2991
rect 12959 2939 12960 2991
rect 12906 2932 12960 2939
rect 12906 2892 12960 2904
rect 12708 2843 12718 2877
rect 12752 2843 12762 2877
rect 12508 2703 12518 2737
rect 12552 2703 12562 2737
rect 12308 2563 12318 2597
rect 12352 2563 12362 2597
rect 12202 2499 12268 2500
rect 12202 2447 12209 2499
rect 12261 2447 12268 2499
rect 12202 2446 12268 2447
rect 12108 2333 12118 2367
rect 12152 2333 12162 2367
rect 11908 2193 11918 2227
rect 11952 2193 11962 2227
rect 11708 2053 11718 2087
rect 11752 2053 11762 2087
rect 11508 1913 11518 1947
rect 11552 1913 11562 1947
rect 11308 1773 11318 1807
rect 11352 1773 11362 1807
rect 11108 1633 11118 1667
rect 11152 1633 11162 1667
rect 10908 1493 10918 1527
rect 10952 1493 10962 1527
rect 10708 1353 10718 1387
rect 10752 1353 10762 1387
rect 10602 1289 10668 1290
rect 10602 1237 10609 1289
rect 10661 1237 10668 1289
rect 10602 1236 10668 1237
rect 10508 1123 10518 1157
rect 10552 1123 10562 1157
rect 10308 983 10318 1017
rect 10352 983 10362 1017
rect 10108 843 10118 877
rect 10152 843 10162 877
rect 9908 703 9918 737
rect 9952 703 9962 737
rect 9708 563 9718 597
rect 9752 563 9762 597
rect 9508 423 9518 457
rect 9552 423 9562 457
rect 9308 283 9318 317
rect 9352 283 9362 317
rect 9108 143 9118 177
rect 9152 143 9162 177
rect 9002 79 9068 80
rect 9002 27 9009 79
rect 9061 27 9068 79
rect 9002 26 9068 27
rect 8908 -67 8909 -15
rect 8961 -67 8962 -15
rect 8908 -79 8918 -67
rect 8952 -79 8962 -67
rect 8708 -132 8762 -131
rect 8708 -143 8718 -132
rect 8752 -143 8762 -132
rect 8708 -195 8709 -143
rect 8761 -195 8762 -143
rect 8708 -210 8762 -195
rect 8812 -133 8858 -81
rect 8812 -167 8818 -133
rect 8852 -167 8858 -133
rect 8718 -291 8725 -239
rect 8777 -291 8784 -239
rect 8612 -397 8618 -363
rect 8652 -397 8658 -363
rect 8612 -435 8658 -397
rect 8612 -469 8618 -435
rect 8652 -469 8658 -435
rect 8612 -512 8658 -469
rect 8709 -326 8761 -320
rect 8709 -390 8718 -378
rect 8752 -390 8761 -378
rect 8709 -454 8718 -442
rect 8752 -454 8761 -442
rect 8709 -555 8761 -506
rect 8812 -363 8858 -167
rect 8908 -131 8909 -79
rect 8961 -131 8962 -79
rect 9008 -22 9062 26
rect 9008 -74 9009 -22
rect 9061 -74 9062 -22
rect 9008 -81 9062 -74
rect 9108 -15 9162 143
rect 9208 177 9262 189
rect 9208 151 9218 177
rect 9252 151 9262 177
rect 9208 99 9209 151
rect 9261 99 9262 151
rect 9208 92 9262 99
rect 9308 177 9362 283
rect 9408 361 9462 368
rect 9408 309 9409 361
rect 9461 309 9462 361
rect 9408 283 9418 309
rect 9452 283 9462 309
rect 9408 271 9462 283
rect 9508 317 9562 423
rect 9608 457 9662 469
rect 9608 431 9618 457
rect 9652 431 9662 457
rect 9608 379 9609 431
rect 9661 379 9662 431
rect 9608 372 9662 379
rect 9708 457 9762 563
rect 9808 641 9862 648
rect 9808 589 9809 641
rect 9861 589 9862 641
rect 9808 563 9818 589
rect 9852 563 9862 589
rect 9808 551 9862 563
rect 9908 597 9962 703
rect 10008 737 10062 749
rect 10008 711 10018 737
rect 10052 711 10062 737
rect 10008 659 10009 711
rect 10061 659 10062 711
rect 10008 652 10062 659
rect 10108 737 10162 843
rect 10208 921 10262 928
rect 10208 869 10209 921
rect 10261 869 10262 921
rect 10208 843 10218 869
rect 10252 843 10262 869
rect 10208 831 10262 843
rect 10308 877 10362 983
rect 10408 1017 10462 1029
rect 10408 991 10418 1017
rect 10452 991 10462 1017
rect 10408 939 10409 991
rect 10461 939 10462 991
rect 10408 932 10462 939
rect 10508 1017 10562 1123
rect 10608 1201 10662 1208
rect 10608 1149 10609 1201
rect 10661 1149 10662 1201
rect 10608 1123 10618 1149
rect 10652 1123 10662 1149
rect 10608 1111 10662 1123
rect 10708 1157 10762 1353
rect 10808 1387 10862 1399
rect 10808 1361 10818 1387
rect 10852 1361 10862 1387
rect 10808 1309 10809 1361
rect 10861 1309 10862 1361
rect 10808 1302 10862 1309
rect 10908 1387 10962 1493
rect 11008 1571 11062 1578
rect 11008 1519 11009 1571
rect 11061 1519 11062 1571
rect 11008 1493 11018 1519
rect 11052 1493 11062 1519
rect 11008 1481 11062 1493
rect 11108 1527 11162 1633
rect 11208 1667 11262 1679
rect 11208 1641 11218 1667
rect 11252 1641 11262 1667
rect 11208 1589 11209 1641
rect 11261 1589 11262 1641
rect 11208 1582 11262 1589
rect 11308 1667 11362 1773
rect 11408 1851 11462 1858
rect 11408 1799 11409 1851
rect 11461 1799 11462 1851
rect 11408 1773 11418 1799
rect 11452 1773 11462 1799
rect 11408 1761 11462 1773
rect 11508 1807 11562 1913
rect 11608 1947 11662 1959
rect 11608 1921 11618 1947
rect 11652 1921 11662 1947
rect 11608 1869 11609 1921
rect 11661 1869 11662 1921
rect 11608 1862 11662 1869
rect 11708 1947 11762 2053
rect 11808 2131 11862 2138
rect 11808 2079 11809 2131
rect 11861 2079 11862 2131
rect 11808 2053 11818 2079
rect 11852 2053 11862 2079
rect 11808 2041 11862 2053
rect 11908 2087 11962 2193
rect 12008 2227 12062 2239
rect 12008 2201 12018 2227
rect 12052 2201 12062 2227
rect 12008 2149 12009 2201
rect 12061 2149 12062 2201
rect 12008 2142 12062 2149
rect 12108 2227 12162 2333
rect 12208 2411 12262 2418
rect 12208 2359 12209 2411
rect 12261 2359 12262 2411
rect 12208 2333 12218 2359
rect 12252 2333 12262 2359
rect 12208 2321 12262 2333
rect 12308 2367 12362 2563
rect 12408 2597 12462 2609
rect 12408 2571 12418 2597
rect 12452 2571 12462 2597
rect 12408 2519 12409 2571
rect 12461 2519 12462 2571
rect 12408 2512 12462 2519
rect 12508 2597 12562 2703
rect 12608 2781 12662 2788
rect 12608 2729 12609 2781
rect 12661 2729 12662 2781
rect 12608 2703 12618 2729
rect 12652 2703 12662 2729
rect 12608 2691 12662 2703
rect 12708 2737 12762 2843
rect 12808 2877 12862 2889
rect 12808 2851 12818 2877
rect 12852 2851 12862 2877
rect 12808 2799 12809 2851
rect 12861 2799 12862 2851
rect 12808 2792 12862 2799
rect 12906 2858 12916 2892
rect 12950 2858 12960 2892
rect 12906 2851 12960 2858
rect 12906 2799 12907 2851
rect 12959 2799 12960 2851
rect 12906 2792 12960 2799
rect 12906 2752 12960 2764
rect 12708 2703 12718 2737
rect 12752 2703 12762 2737
rect 12508 2563 12518 2597
rect 12552 2563 12562 2597
rect 12402 2483 12468 2484
rect 12402 2431 12409 2483
rect 12461 2431 12468 2483
rect 12402 2430 12468 2431
rect 12308 2333 12318 2367
rect 12352 2333 12362 2367
rect 12108 2193 12118 2227
rect 12152 2193 12162 2227
rect 11908 2053 11918 2087
rect 11952 2053 11962 2087
rect 11708 1913 11718 1947
rect 11752 1913 11762 1947
rect 11508 1773 11518 1807
rect 11552 1773 11562 1807
rect 11308 1633 11318 1667
rect 11352 1633 11362 1667
rect 11108 1493 11118 1527
rect 11152 1493 11162 1527
rect 10908 1353 10918 1387
rect 10952 1353 10962 1387
rect 10802 1273 10868 1274
rect 10802 1221 10809 1273
rect 10861 1221 10868 1273
rect 10802 1220 10868 1221
rect 10708 1123 10718 1157
rect 10752 1123 10762 1157
rect 10508 983 10518 1017
rect 10552 983 10562 1017
rect 10308 843 10318 877
rect 10352 843 10362 877
rect 10108 703 10118 737
rect 10152 703 10162 737
rect 9908 563 9918 597
rect 9952 563 9962 597
rect 9708 423 9718 457
rect 9752 423 9762 457
rect 9508 283 9518 317
rect 9552 283 9562 317
rect 9308 143 9318 177
rect 9352 143 9362 177
rect 9202 63 9268 64
rect 9202 11 9209 63
rect 9261 11 9268 63
rect 9202 10 9268 11
rect 9108 -67 9109 -15
rect 9161 -67 9162 -15
rect 9108 -79 9118 -67
rect 9152 -79 9162 -67
rect 8908 -132 8962 -131
rect 8908 -143 8918 -132
rect 8952 -143 8962 -132
rect 8908 -195 8909 -143
rect 8961 -195 8962 -143
rect 8908 -210 8962 -195
rect 9012 -133 9058 -81
rect 9012 -167 9018 -133
rect 9052 -167 9058 -133
rect 8918 -291 8925 -239
rect 8977 -291 8984 -239
rect 8812 -397 8818 -363
rect 8852 -397 8858 -363
rect 8812 -435 8858 -397
rect 8812 -469 8818 -435
rect 8852 -469 8858 -435
rect 8812 -512 8858 -469
rect 8909 -326 8961 -320
rect 8909 -390 8918 -378
rect 8952 -390 8961 -378
rect 8909 -454 8918 -442
rect 8952 -454 8961 -442
rect 8909 -512 8961 -506
rect 9012 -363 9058 -167
rect 9108 -131 9109 -79
rect 9161 -131 9162 -79
rect 9208 -22 9262 10
rect 9208 -74 9209 -22
rect 9261 -74 9262 -22
rect 9208 -81 9262 -74
rect 9308 -15 9362 143
rect 9408 221 9462 228
rect 9408 169 9409 221
rect 9461 169 9462 221
rect 9408 143 9418 169
rect 9452 143 9462 169
rect 9408 131 9462 143
rect 9508 177 9562 283
rect 9608 317 9662 329
rect 9608 291 9618 317
rect 9652 291 9662 317
rect 9608 239 9609 291
rect 9661 239 9662 291
rect 9608 232 9662 239
rect 9708 317 9762 423
rect 9808 501 9862 508
rect 9808 449 9809 501
rect 9861 449 9862 501
rect 9808 423 9818 449
rect 9852 423 9862 449
rect 9808 411 9862 423
rect 9908 457 9962 563
rect 10008 597 10062 609
rect 10008 571 10018 597
rect 10052 571 10062 597
rect 10008 519 10009 571
rect 10061 519 10062 571
rect 10008 512 10062 519
rect 10108 597 10162 703
rect 10208 781 10262 788
rect 10208 729 10209 781
rect 10261 729 10262 781
rect 10208 703 10218 729
rect 10252 703 10262 729
rect 10208 691 10262 703
rect 10308 737 10362 843
rect 10408 877 10462 889
rect 10408 851 10418 877
rect 10452 851 10462 877
rect 10408 799 10409 851
rect 10461 799 10462 851
rect 10408 792 10462 799
rect 10508 877 10562 983
rect 10608 1061 10662 1068
rect 10608 1009 10609 1061
rect 10661 1009 10662 1061
rect 10608 983 10618 1009
rect 10652 983 10662 1009
rect 10608 971 10662 983
rect 10708 1017 10762 1123
rect 10808 1157 10862 1169
rect 10808 1131 10818 1157
rect 10852 1131 10862 1157
rect 10808 1079 10809 1131
rect 10861 1079 10862 1131
rect 10808 1072 10862 1079
rect 10908 1157 10962 1353
rect 11008 1431 11062 1438
rect 11008 1379 11009 1431
rect 11061 1379 11062 1431
rect 11008 1353 11018 1379
rect 11052 1353 11062 1379
rect 11008 1341 11062 1353
rect 11108 1387 11162 1493
rect 11208 1527 11262 1539
rect 11208 1501 11218 1527
rect 11252 1501 11262 1527
rect 11208 1449 11209 1501
rect 11261 1449 11262 1501
rect 11208 1442 11262 1449
rect 11308 1527 11362 1633
rect 11408 1711 11462 1718
rect 11408 1659 11409 1711
rect 11461 1659 11462 1711
rect 11408 1633 11418 1659
rect 11452 1633 11462 1659
rect 11408 1621 11462 1633
rect 11508 1667 11562 1773
rect 11608 1807 11662 1819
rect 11608 1781 11618 1807
rect 11652 1781 11662 1807
rect 11608 1729 11609 1781
rect 11661 1729 11662 1781
rect 11608 1722 11662 1729
rect 11708 1807 11762 1913
rect 11808 1991 11862 1998
rect 11808 1939 11809 1991
rect 11861 1939 11862 1991
rect 11808 1913 11818 1939
rect 11852 1913 11862 1939
rect 11808 1901 11862 1913
rect 11908 1947 11962 2053
rect 12008 2087 12062 2099
rect 12008 2061 12018 2087
rect 12052 2061 12062 2087
rect 12008 2009 12009 2061
rect 12061 2009 12062 2061
rect 12008 2002 12062 2009
rect 12108 2087 12162 2193
rect 12208 2271 12262 2278
rect 12208 2219 12209 2271
rect 12261 2219 12262 2271
rect 12208 2193 12218 2219
rect 12252 2193 12262 2219
rect 12208 2181 12262 2193
rect 12308 2227 12362 2333
rect 12408 2367 12462 2379
rect 12408 2341 12418 2367
rect 12452 2341 12462 2367
rect 12408 2289 12409 2341
rect 12461 2289 12462 2341
rect 12408 2282 12462 2289
rect 12508 2367 12562 2563
rect 12608 2641 12662 2648
rect 12608 2589 12609 2641
rect 12661 2589 12662 2641
rect 12608 2563 12618 2589
rect 12652 2563 12662 2589
rect 12608 2551 12662 2563
rect 12708 2597 12762 2703
rect 12808 2737 12862 2749
rect 12808 2711 12818 2737
rect 12852 2711 12862 2737
rect 12808 2659 12809 2711
rect 12861 2659 12862 2711
rect 12808 2652 12862 2659
rect 12906 2718 12916 2752
rect 12950 2718 12960 2752
rect 12906 2711 12960 2718
rect 12906 2659 12907 2711
rect 12959 2659 12960 2711
rect 12906 2652 12960 2659
rect 12906 2612 12960 2624
rect 12708 2563 12718 2597
rect 12752 2563 12762 2597
rect 12602 2499 12668 2500
rect 12602 2447 12609 2499
rect 12661 2447 12668 2499
rect 12602 2446 12668 2447
rect 12508 2333 12518 2367
rect 12552 2333 12562 2367
rect 12308 2193 12318 2227
rect 12352 2193 12362 2227
rect 12108 2053 12118 2087
rect 12152 2053 12162 2087
rect 11908 1913 11918 1947
rect 11952 1913 11962 1947
rect 11708 1773 11718 1807
rect 11752 1773 11762 1807
rect 11508 1633 11518 1667
rect 11552 1633 11562 1667
rect 11308 1493 11318 1527
rect 11352 1493 11362 1527
rect 11108 1353 11118 1387
rect 11152 1353 11162 1387
rect 11002 1289 11068 1290
rect 11002 1237 11009 1289
rect 11061 1237 11068 1289
rect 11002 1236 11068 1237
rect 10908 1123 10918 1157
rect 10952 1123 10962 1157
rect 10708 983 10718 1017
rect 10752 983 10762 1017
rect 10508 843 10518 877
rect 10552 843 10562 877
rect 10308 703 10318 737
rect 10352 703 10362 737
rect 10108 563 10118 597
rect 10152 563 10162 597
rect 9908 423 9918 457
rect 9952 423 9962 457
rect 9708 283 9718 317
rect 9752 283 9762 317
rect 9508 143 9518 177
rect 9552 143 9562 177
rect 9402 79 9468 80
rect 9402 27 9409 79
rect 9461 27 9468 79
rect 9402 26 9468 27
rect 9308 -67 9309 -15
rect 9361 -67 9362 -15
rect 9308 -79 9318 -67
rect 9352 -79 9362 -67
rect 9108 -132 9162 -131
rect 9108 -143 9118 -132
rect 9152 -143 9162 -132
rect 9108 -195 9109 -143
rect 9161 -195 9162 -143
rect 9108 -210 9162 -195
rect 9212 -133 9258 -81
rect 9212 -167 9218 -133
rect 9252 -167 9258 -133
rect 9118 -291 9125 -239
rect 9177 -291 9184 -239
rect 9012 -397 9018 -363
rect 9052 -397 9058 -363
rect 9012 -435 9058 -397
rect 9012 -469 9018 -435
rect 9052 -469 9058 -435
rect 9012 -512 9058 -469
rect 9109 -326 9161 -320
rect 9109 -390 9118 -378
rect 9152 -390 9161 -378
rect 9109 -454 9118 -442
rect 9152 -454 9161 -442
rect 9109 -555 9161 -506
rect 9212 -363 9258 -167
rect 9308 -131 9309 -79
rect 9361 -131 9362 -79
rect 9408 -22 9462 26
rect 9408 -74 9409 -22
rect 9461 -74 9462 -22
rect 9408 -81 9462 -74
rect 9508 -15 9562 143
rect 9608 177 9662 189
rect 9608 151 9618 177
rect 9652 151 9662 177
rect 9608 99 9609 151
rect 9661 99 9662 151
rect 9608 92 9662 99
rect 9708 177 9762 283
rect 9808 361 9862 368
rect 9808 309 9809 361
rect 9861 309 9862 361
rect 9808 283 9818 309
rect 9852 283 9862 309
rect 9808 271 9862 283
rect 9908 317 9962 423
rect 10008 457 10062 469
rect 10008 431 10018 457
rect 10052 431 10062 457
rect 10008 379 10009 431
rect 10061 379 10062 431
rect 10008 372 10062 379
rect 10108 457 10162 563
rect 10208 641 10262 648
rect 10208 589 10209 641
rect 10261 589 10262 641
rect 10208 563 10218 589
rect 10252 563 10262 589
rect 10208 551 10262 563
rect 10308 597 10362 703
rect 10408 737 10462 749
rect 10408 711 10418 737
rect 10452 711 10462 737
rect 10408 659 10409 711
rect 10461 659 10462 711
rect 10408 652 10462 659
rect 10508 737 10562 843
rect 10608 921 10662 928
rect 10608 869 10609 921
rect 10661 869 10662 921
rect 10608 843 10618 869
rect 10652 843 10662 869
rect 10608 831 10662 843
rect 10708 877 10762 983
rect 10808 1017 10862 1029
rect 10808 991 10818 1017
rect 10852 991 10862 1017
rect 10808 939 10809 991
rect 10861 939 10862 991
rect 10808 932 10862 939
rect 10908 1017 10962 1123
rect 11008 1201 11062 1208
rect 11008 1149 11009 1201
rect 11061 1149 11062 1201
rect 11008 1123 11018 1149
rect 11052 1123 11062 1149
rect 11008 1111 11062 1123
rect 11108 1157 11162 1353
rect 11208 1387 11262 1399
rect 11208 1361 11218 1387
rect 11252 1361 11262 1387
rect 11208 1309 11209 1361
rect 11261 1309 11262 1361
rect 11208 1302 11262 1309
rect 11308 1387 11362 1493
rect 11408 1571 11462 1578
rect 11408 1519 11409 1571
rect 11461 1519 11462 1571
rect 11408 1493 11418 1519
rect 11452 1493 11462 1519
rect 11408 1481 11462 1493
rect 11508 1527 11562 1633
rect 11608 1667 11662 1679
rect 11608 1641 11618 1667
rect 11652 1641 11662 1667
rect 11608 1589 11609 1641
rect 11661 1589 11662 1641
rect 11608 1582 11662 1589
rect 11708 1667 11762 1773
rect 11808 1851 11862 1858
rect 11808 1799 11809 1851
rect 11861 1799 11862 1851
rect 11808 1773 11818 1799
rect 11852 1773 11862 1799
rect 11808 1761 11862 1773
rect 11908 1807 11962 1913
rect 12008 1947 12062 1959
rect 12008 1921 12018 1947
rect 12052 1921 12062 1947
rect 12008 1869 12009 1921
rect 12061 1869 12062 1921
rect 12008 1862 12062 1869
rect 12108 1947 12162 2053
rect 12208 2131 12262 2138
rect 12208 2079 12209 2131
rect 12261 2079 12262 2131
rect 12208 2053 12218 2079
rect 12252 2053 12262 2079
rect 12208 2041 12262 2053
rect 12308 2087 12362 2193
rect 12408 2227 12462 2239
rect 12408 2201 12418 2227
rect 12452 2201 12462 2227
rect 12408 2149 12409 2201
rect 12461 2149 12462 2201
rect 12408 2142 12462 2149
rect 12508 2227 12562 2333
rect 12608 2411 12662 2418
rect 12608 2359 12609 2411
rect 12661 2359 12662 2411
rect 12608 2333 12618 2359
rect 12652 2333 12662 2359
rect 12608 2321 12662 2333
rect 12708 2367 12762 2563
rect 12808 2597 12862 2609
rect 12808 2571 12818 2597
rect 12852 2571 12862 2597
rect 12808 2519 12809 2571
rect 12861 2519 12862 2571
rect 12808 2512 12862 2519
rect 12906 2578 12916 2612
rect 12950 2578 12960 2612
rect 12906 2571 12960 2578
rect 12906 2519 12907 2571
rect 12959 2519 12960 2571
rect 12906 2512 12960 2519
rect 12990 2477 13020 3641
rect 12904 2471 13020 2477
rect 12904 2437 12916 2471
rect 12950 2437 13020 2471
rect 12904 2431 13020 2437
rect 12906 2382 12960 2394
rect 12708 2333 12718 2367
rect 12752 2333 12762 2367
rect 12508 2193 12518 2227
rect 12552 2193 12562 2227
rect 12308 2053 12318 2087
rect 12352 2053 12362 2087
rect 12108 1913 12118 1947
rect 12152 1913 12162 1947
rect 11908 1773 11918 1807
rect 11952 1773 11962 1807
rect 11708 1633 11718 1667
rect 11752 1633 11762 1667
rect 11508 1493 11518 1527
rect 11552 1493 11562 1527
rect 11308 1353 11318 1387
rect 11352 1353 11362 1387
rect 11202 1273 11268 1274
rect 11202 1221 11209 1273
rect 11261 1221 11268 1273
rect 11202 1220 11268 1221
rect 11108 1123 11118 1157
rect 11152 1123 11162 1157
rect 10908 983 10918 1017
rect 10952 983 10962 1017
rect 10708 843 10718 877
rect 10752 843 10762 877
rect 10508 703 10518 737
rect 10552 703 10562 737
rect 10308 563 10318 597
rect 10352 563 10362 597
rect 10108 423 10118 457
rect 10152 423 10162 457
rect 9908 283 9918 317
rect 9952 283 9962 317
rect 9708 143 9718 177
rect 9752 143 9762 177
rect 9602 63 9668 64
rect 9602 11 9609 63
rect 9661 11 9668 63
rect 9602 10 9668 11
rect 9508 -67 9509 -15
rect 9561 -67 9562 -15
rect 9508 -79 9518 -67
rect 9552 -79 9562 -67
rect 9308 -132 9362 -131
rect 9308 -143 9318 -132
rect 9352 -143 9362 -132
rect 9308 -195 9309 -143
rect 9361 -195 9362 -143
rect 9308 -210 9362 -195
rect 9412 -133 9458 -81
rect 9412 -167 9418 -133
rect 9452 -167 9458 -133
rect 9318 -291 9325 -239
rect 9377 -291 9384 -239
rect 9212 -397 9218 -363
rect 9252 -397 9258 -363
rect 9212 -435 9258 -397
rect 9212 -469 9218 -435
rect 9252 -469 9258 -435
rect 9212 -512 9258 -469
rect 9309 -326 9361 -320
rect 9309 -390 9318 -378
rect 9352 -390 9361 -378
rect 9309 -454 9318 -442
rect 9352 -454 9361 -442
rect 9309 -512 9361 -506
rect 9412 -363 9458 -167
rect 9508 -131 9509 -79
rect 9561 -131 9562 -79
rect 9608 -22 9662 10
rect 9608 -74 9609 -22
rect 9661 -74 9662 -22
rect 9608 -81 9662 -74
rect 9708 -15 9762 143
rect 9808 221 9862 228
rect 9808 169 9809 221
rect 9861 169 9862 221
rect 9808 143 9818 169
rect 9852 143 9862 169
rect 9808 131 9862 143
rect 9908 177 9962 283
rect 10008 317 10062 329
rect 10008 291 10018 317
rect 10052 291 10062 317
rect 10008 239 10009 291
rect 10061 239 10062 291
rect 10008 232 10062 239
rect 10108 317 10162 423
rect 10208 501 10262 508
rect 10208 449 10209 501
rect 10261 449 10262 501
rect 10208 423 10218 449
rect 10252 423 10262 449
rect 10208 411 10262 423
rect 10308 457 10362 563
rect 10408 597 10462 609
rect 10408 571 10418 597
rect 10452 571 10462 597
rect 10408 519 10409 571
rect 10461 519 10462 571
rect 10408 512 10462 519
rect 10508 597 10562 703
rect 10608 781 10662 788
rect 10608 729 10609 781
rect 10661 729 10662 781
rect 10608 703 10618 729
rect 10652 703 10662 729
rect 10608 691 10662 703
rect 10708 737 10762 843
rect 10808 877 10862 889
rect 10808 851 10818 877
rect 10852 851 10862 877
rect 10808 799 10809 851
rect 10861 799 10862 851
rect 10808 792 10862 799
rect 10908 877 10962 983
rect 11008 1061 11062 1068
rect 11008 1009 11009 1061
rect 11061 1009 11062 1061
rect 11008 983 11018 1009
rect 11052 983 11062 1009
rect 11008 971 11062 983
rect 11108 1017 11162 1123
rect 11208 1157 11262 1169
rect 11208 1131 11218 1157
rect 11252 1131 11262 1157
rect 11208 1079 11209 1131
rect 11261 1079 11262 1131
rect 11208 1072 11262 1079
rect 11308 1157 11362 1353
rect 11408 1431 11462 1438
rect 11408 1379 11409 1431
rect 11461 1379 11462 1431
rect 11408 1353 11418 1379
rect 11452 1353 11462 1379
rect 11408 1341 11462 1353
rect 11508 1387 11562 1493
rect 11608 1527 11662 1539
rect 11608 1501 11618 1527
rect 11652 1501 11662 1527
rect 11608 1449 11609 1501
rect 11661 1449 11662 1501
rect 11608 1442 11662 1449
rect 11708 1527 11762 1633
rect 11808 1711 11862 1718
rect 11808 1659 11809 1711
rect 11861 1659 11862 1711
rect 11808 1633 11818 1659
rect 11852 1633 11862 1659
rect 11808 1621 11862 1633
rect 11908 1667 11962 1773
rect 12008 1807 12062 1819
rect 12008 1781 12018 1807
rect 12052 1781 12062 1807
rect 12008 1729 12009 1781
rect 12061 1729 12062 1781
rect 12008 1722 12062 1729
rect 12108 1807 12162 1913
rect 12208 1991 12262 1998
rect 12208 1939 12209 1991
rect 12261 1939 12262 1991
rect 12208 1913 12218 1939
rect 12252 1913 12262 1939
rect 12208 1901 12262 1913
rect 12308 1947 12362 2053
rect 12408 2087 12462 2099
rect 12408 2061 12418 2087
rect 12452 2061 12462 2087
rect 12408 2009 12409 2061
rect 12461 2009 12462 2061
rect 12408 2002 12462 2009
rect 12508 2087 12562 2193
rect 12608 2271 12662 2278
rect 12608 2219 12609 2271
rect 12661 2219 12662 2271
rect 12608 2193 12618 2219
rect 12652 2193 12662 2219
rect 12608 2181 12662 2193
rect 12708 2227 12762 2333
rect 12808 2367 12862 2379
rect 12808 2341 12818 2367
rect 12852 2341 12862 2367
rect 12808 2289 12809 2341
rect 12861 2289 12862 2341
rect 12808 2282 12862 2289
rect 12906 2348 12916 2382
rect 12950 2348 12960 2382
rect 12906 2341 12960 2348
rect 12906 2289 12907 2341
rect 12959 2289 12960 2341
rect 12906 2282 12960 2289
rect 12906 2242 12960 2254
rect 12708 2193 12718 2227
rect 12752 2193 12762 2227
rect 12508 2053 12518 2087
rect 12552 2053 12562 2087
rect 12308 1913 12318 1947
rect 12352 1913 12362 1947
rect 12108 1773 12118 1807
rect 12152 1773 12162 1807
rect 11908 1633 11918 1667
rect 11952 1633 11962 1667
rect 11708 1493 11718 1527
rect 11752 1493 11762 1527
rect 11508 1353 11518 1387
rect 11552 1353 11562 1387
rect 11402 1289 11468 1290
rect 11402 1237 11409 1289
rect 11461 1237 11468 1289
rect 11402 1236 11468 1237
rect 11308 1123 11318 1157
rect 11352 1123 11362 1157
rect 11108 983 11118 1017
rect 11152 983 11162 1017
rect 10908 843 10918 877
rect 10952 843 10962 877
rect 10708 703 10718 737
rect 10752 703 10762 737
rect 10508 563 10518 597
rect 10552 563 10562 597
rect 10308 423 10318 457
rect 10352 423 10362 457
rect 10108 283 10118 317
rect 10152 283 10162 317
rect 9908 143 9918 177
rect 9952 143 9962 177
rect 9802 79 9868 80
rect 9802 27 9809 79
rect 9861 27 9868 79
rect 9802 26 9868 27
rect 9708 -67 9709 -15
rect 9761 -67 9762 -15
rect 9708 -79 9718 -67
rect 9752 -79 9762 -67
rect 9508 -132 9562 -131
rect 9508 -143 9518 -132
rect 9552 -143 9562 -132
rect 9508 -195 9509 -143
rect 9561 -195 9562 -143
rect 9508 -210 9562 -195
rect 9612 -133 9658 -81
rect 9612 -167 9618 -133
rect 9652 -167 9658 -133
rect 9518 -291 9525 -239
rect 9577 -291 9584 -239
rect 9412 -397 9418 -363
rect 9452 -397 9458 -363
rect 9412 -435 9458 -397
rect 9412 -469 9418 -435
rect 9452 -469 9458 -435
rect 9412 -512 9458 -469
rect 9509 -326 9561 -320
rect 9509 -390 9518 -378
rect 9552 -390 9561 -378
rect 9509 -454 9518 -442
rect 9552 -454 9561 -442
rect 9509 -555 9561 -506
rect 9612 -363 9658 -167
rect 9708 -131 9709 -79
rect 9761 -131 9762 -79
rect 9808 -22 9862 26
rect 9808 -74 9809 -22
rect 9861 -74 9862 -22
rect 9808 -81 9862 -74
rect 9908 -15 9962 143
rect 10008 177 10062 189
rect 10008 151 10018 177
rect 10052 151 10062 177
rect 10008 99 10009 151
rect 10061 99 10062 151
rect 10008 92 10062 99
rect 10108 177 10162 283
rect 10208 361 10262 368
rect 10208 309 10209 361
rect 10261 309 10262 361
rect 10208 283 10218 309
rect 10252 283 10262 309
rect 10208 271 10262 283
rect 10308 317 10362 423
rect 10408 457 10462 469
rect 10408 431 10418 457
rect 10452 431 10462 457
rect 10408 379 10409 431
rect 10461 379 10462 431
rect 10408 372 10462 379
rect 10508 457 10562 563
rect 10608 641 10662 648
rect 10608 589 10609 641
rect 10661 589 10662 641
rect 10608 563 10618 589
rect 10652 563 10662 589
rect 10608 551 10662 563
rect 10708 597 10762 703
rect 10808 737 10862 749
rect 10808 711 10818 737
rect 10852 711 10862 737
rect 10808 659 10809 711
rect 10861 659 10862 711
rect 10808 652 10862 659
rect 10908 737 10962 843
rect 11008 921 11062 928
rect 11008 869 11009 921
rect 11061 869 11062 921
rect 11008 843 11018 869
rect 11052 843 11062 869
rect 11008 831 11062 843
rect 11108 877 11162 983
rect 11208 1017 11262 1029
rect 11208 991 11218 1017
rect 11252 991 11262 1017
rect 11208 939 11209 991
rect 11261 939 11262 991
rect 11208 932 11262 939
rect 11308 1017 11362 1123
rect 11408 1201 11462 1208
rect 11408 1149 11409 1201
rect 11461 1149 11462 1201
rect 11408 1123 11418 1149
rect 11452 1123 11462 1149
rect 11408 1111 11462 1123
rect 11508 1157 11562 1353
rect 11608 1387 11662 1399
rect 11608 1361 11618 1387
rect 11652 1361 11662 1387
rect 11608 1309 11609 1361
rect 11661 1309 11662 1361
rect 11608 1302 11662 1309
rect 11708 1387 11762 1493
rect 11808 1571 11862 1578
rect 11808 1519 11809 1571
rect 11861 1519 11862 1571
rect 11808 1493 11818 1519
rect 11852 1493 11862 1519
rect 11808 1481 11862 1493
rect 11908 1527 11962 1633
rect 12008 1667 12062 1679
rect 12008 1641 12018 1667
rect 12052 1641 12062 1667
rect 12008 1589 12009 1641
rect 12061 1589 12062 1641
rect 12008 1582 12062 1589
rect 12108 1667 12162 1773
rect 12208 1851 12262 1858
rect 12208 1799 12209 1851
rect 12261 1799 12262 1851
rect 12208 1773 12218 1799
rect 12252 1773 12262 1799
rect 12208 1761 12262 1773
rect 12308 1807 12362 1913
rect 12408 1947 12462 1959
rect 12408 1921 12418 1947
rect 12452 1921 12462 1947
rect 12408 1869 12409 1921
rect 12461 1869 12462 1921
rect 12408 1862 12462 1869
rect 12508 1947 12562 2053
rect 12608 2131 12662 2138
rect 12608 2079 12609 2131
rect 12661 2079 12662 2131
rect 12608 2053 12618 2079
rect 12652 2053 12662 2079
rect 12608 2041 12662 2053
rect 12708 2087 12762 2193
rect 12808 2227 12862 2239
rect 12808 2201 12818 2227
rect 12852 2201 12862 2227
rect 12808 2149 12809 2201
rect 12861 2149 12862 2201
rect 12808 2142 12862 2149
rect 12906 2208 12916 2242
rect 12950 2208 12960 2242
rect 12906 2201 12960 2208
rect 12906 2149 12907 2201
rect 12959 2149 12960 2201
rect 12906 2142 12960 2149
rect 12906 2102 12960 2114
rect 12708 2053 12718 2087
rect 12752 2053 12762 2087
rect 12508 1913 12518 1947
rect 12552 1913 12562 1947
rect 12308 1773 12318 1807
rect 12352 1773 12362 1807
rect 12108 1633 12118 1667
rect 12152 1633 12162 1667
rect 11908 1493 11918 1527
rect 11952 1493 11962 1527
rect 11708 1353 11718 1387
rect 11752 1353 11762 1387
rect 11602 1273 11668 1274
rect 11602 1221 11609 1273
rect 11661 1221 11668 1273
rect 11602 1220 11668 1221
rect 11508 1123 11518 1157
rect 11552 1123 11562 1157
rect 11308 983 11318 1017
rect 11352 983 11362 1017
rect 11108 843 11118 877
rect 11152 843 11162 877
rect 10908 703 10918 737
rect 10952 703 10962 737
rect 10708 563 10718 597
rect 10752 563 10762 597
rect 10508 423 10518 457
rect 10552 423 10562 457
rect 10308 283 10318 317
rect 10352 283 10362 317
rect 10108 143 10118 177
rect 10152 143 10162 177
rect 10002 63 10068 64
rect 10002 11 10009 63
rect 10061 11 10068 63
rect 10002 10 10068 11
rect 9908 -67 9909 -15
rect 9961 -67 9962 -15
rect 9908 -79 9918 -67
rect 9952 -79 9962 -67
rect 9708 -132 9762 -131
rect 9708 -143 9718 -132
rect 9752 -143 9762 -132
rect 9708 -195 9709 -143
rect 9761 -195 9762 -143
rect 9708 -210 9762 -195
rect 9812 -133 9858 -81
rect 9812 -167 9818 -133
rect 9852 -167 9858 -133
rect 9718 -291 9725 -239
rect 9777 -291 9784 -239
rect 9612 -397 9618 -363
rect 9652 -397 9658 -363
rect 9612 -435 9658 -397
rect 9612 -469 9618 -435
rect 9652 -469 9658 -435
rect 9612 -512 9658 -469
rect 9709 -326 9761 -320
rect 9709 -390 9718 -378
rect 9752 -390 9761 -378
rect 9709 -454 9718 -442
rect 9752 -454 9761 -442
rect 9709 -512 9761 -506
rect 9812 -363 9858 -167
rect 9908 -131 9909 -79
rect 9961 -131 9962 -79
rect 10008 -22 10062 10
rect 10008 -74 10009 -22
rect 10061 -74 10062 -22
rect 10008 -81 10062 -74
rect 10108 -15 10162 143
rect 10208 221 10262 228
rect 10208 169 10209 221
rect 10261 169 10262 221
rect 10208 143 10218 169
rect 10252 143 10262 169
rect 10208 131 10262 143
rect 10308 177 10362 283
rect 10408 317 10462 329
rect 10408 291 10418 317
rect 10452 291 10462 317
rect 10408 239 10409 291
rect 10461 239 10462 291
rect 10408 232 10462 239
rect 10508 317 10562 423
rect 10608 501 10662 508
rect 10608 449 10609 501
rect 10661 449 10662 501
rect 10608 423 10618 449
rect 10652 423 10662 449
rect 10608 411 10662 423
rect 10708 457 10762 563
rect 10808 597 10862 609
rect 10808 571 10818 597
rect 10852 571 10862 597
rect 10808 519 10809 571
rect 10861 519 10862 571
rect 10808 512 10862 519
rect 10908 597 10962 703
rect 11008 781 11062 788
rect 11008 729 11009 781
rect 11061 729 11062 781
rect 11008 703 11018 729
rect 11052 703 11062 729
rect 11008 691 11062 703
rect 11108 737 11162 843
rect 11208 877 11262 889
rect 11208 851 11218 877
rect 11252 851 11262 877
rect 11208 799 11209 851
rect 11261 799 11262 851
rect 11208 792 11262 799
rect 11308 877 11362 983
rect 11408 1061 11462 1068
rect 11408 1009 11409 1061
rect 11461 1009 11462 1061
rect 11408 983 11418 1009
rect 11452 983 11462 1009
rect 11408 971 11462 983
rect 11508 1017 11562 1123
rect 11608 1157 11662 1169
rect 11608 1131 11618 1157
rect 11652 1131 11662 1157
rect 11608 1079 11609 1131
rect 11661 1079 11662 1131
rect 11608 1072 11662 1079
rect 11708 1157 11762 1353
rect 11808 1431 11862 1438
rect 11808 1379 11809 1431
rect 11861 1379 11862 1431
rect 11808 1353 11818 1379
rect 11852 1353 11862 1379
rect 11808 1341 11862 1353
rect 11908 1387 11962 1493
rect 12008 1527 12062 1539
rect 12008 1501 12018 1527
rect 12052 1501 12062 1527
rect 12008 1449 12009 1501
rect 12061 1449 12062 1501
rect 12008 1442 12062 1449
rect 12108 1527 12162 1633
rect 12208 1711 12262 1718
rect 12208 1659 12209 1711
rect 12261 1659 12262 1711
rect 12208 1633 12218 1659
rect 12252 1633 12262 1659
rect 12208 1621 12262 1633
rect 12308 1667 12362 1773
rect 12408 1807 12462 1819
rect 12408 1781 12418 1807
rect 12452 1781 12462 1807
rect 12408 1729 12409 1781
rect 12461 1729 12462 1781
rect 12408 1722 12462 1729
rect 12508 1807 12562 1913
rect 12608 1991 12662 1998
rect 12608 1939 12609 1991
rect 12661 1939 12662 1991
rect 12608 1913 12618 1939
rect 12652 1913 12662 1939
rect 12608 1901 12662 1913
rect 12708 1947 12762 2053
rect 12808 2087 12862 2099
rect 12808 2061 12818 2087
rect 12852 2061 12862 2087
rect 12808 2009 12809 2061
rect 12861 2009 12862 2061
rect 12808 2002 12862 2009
rect 12906 2068 12916 2102
rect 12950 2068 12960 2102
rect 12906 2061 12960 2068
rect 12906 2009 12907 2061
rect 12959 2009 12960 2061
rect 12906 2002 12960 2009
rect 12906 1962 12960 1974
rect 12708 1913 12718 1947
rect 12752 1913 12762 1947
rect 12508 1773 12518 1807
rect 12552 1773 12562 1807
rect 12308 1633 12318 1667
rect 12352 1633 12362 1667
rect 12108 1493 12118 1527
rect 12152 1493 12162 1527
rect 11908 1353 11918 1387
rect 11952 1353 11962 1387
rect 11802 1289 11868 1290
rect 11802 1237 11809 1289
rect 11861 1237 11868 1289
rect 11802 1236 11868 1237
rect 11708 1123 11718 1157
rect 11752 1123 11762 1157
rect 11508 983 11518 1017
rect 11552 983 11562 1017
rect 11308 843 11318 877
rect 11352 843 11362 877
rect 11108 703 11118 737
rect 11152 703 11162 737
rect 10908 563 10918 597
rect 10952 563 10962 597
rect 10708 423 10718 457
rect 10752 423 10762 457
rect 10508 283 10518 317
rect 10552 283 10562 317
rect 10308 143 10318 177
rect 10352 143 10362 177
rect 10202 79 10268 80
rect 10202 27 10209 79
rect 10261 27 10268 79
rect 10202 26 10268 27
rect 10108 -67 10109 -15
rect 10161 -67 10162 -15
rect 10108 -79 10118 -67
rect 10152 -79 10162 -67
rect 9908 -132 9962 -131
rect 9908 -143 9918 -132
rect 9952 -143 9962 -132
rect 9908 -195 9909 -143
rect 9961 -195 9962 -143
rect 9908 -210 9962 -195
rect 10012 -133 10058 -81
rect 10012 -167 10018 -133
rect 10052 -167 10058 -133
rect 9918 -291 9925 -239
rect 9977 -291 9984 -239
rect 9812 -397 9818 -363
rect 9852 -397 9858 -363
rect 9812 -435 9858 -397
rect 9812 -469 9818 -435
rect 9852 -469 9858 -435
rect 9812 -512 9858 -469
rect 9909 -326 9961 -320
rect 9909 -390 9918 -378
rect 9952 -390 9961 -378
rect 9909 -454 9918 -442
rect 9952 -454 9961 -442
rect 9909 -555 9961 -506
rect 10012 -363 10058 -167
rect 10108 -131 10109 -79
rect 10161 -131 10162 -79
rect 10208 -22 10262 26
rect 10208 -74 10209 -22
rect 10261 -74 10262 -22
rect 10208 -81 10262 -74
rect 10308 -15 10362 143
rect 10408 177 10462 189
rect 10408 151 10418 177
rect 10452 151 10462 177
rect 10408 99 10409 151
rect 10461 99 10462 151
rect 10408 92 10462 99
rect 10508 177 10562 283
rect 10608 361 10662 368
rect 10608 309 10609 361
rect 10661 309 10662 361
rect 10608 283 10618 309
rect 10652 283 10662 309
rect 10608 271 10662 283
rect 10708 317 10762 423
rect 10808 457 10862 469
rect 10808 431 10818 457
rect 10852 431 10862 457
rect 10808 379 10809 431
rect 10861 379 10862 431
rect 10808 372 10862 379
rect 10908 457 10962 563
rect 11008 641 11062 648
rect 11008 589 11009 641
rect 11061 589 11062 641
rect 11008 563 11018 589
rect 11052 563 11062 589
rect 11008 551 11062 563
rect 11108 597 11162 703
rect 11208 737 11262 749
rect 11208 711 11218 737
rect 11252 711 11262 737
rect 11208 659 11209 711
rect 11261 659 11262 711
rect 11208 652 11262 659
rect 11308 737 11362 843
rect 11408 921 11462 928
rect 11408 869 11409 921
rect 11461 869 11462 921
rect 11408 843 11418 869
rect 11452 843 11462 869
rect 11408 831 11462 843
rect 11508 877 11562 983
rect 11608 1017 11662 1029
rect 11608 991 11618 1017
rect 11652 991 11662 1017
rect 11608 939 11609 991
rect 11661 939 11662 991
rect 11608 932 11662 939
rect 11708 1017 11762 1123
rect 11808 1201 11862 1208
rect 11808 1149 11809 1201
rect 11861 1149 11862 1201
rect 11808 1123 11818 1149
rect 11852 1123 11862 1149
rect 11808 1111 11862 1123
rect 11908 1157 11962 1353
rect 12008 1387 12062 1399
rect 12008 1361 12018 1387
rect 12052 1361 12062 1387
rect 12008 1309 12009 1361
rect 12061 1309 12062 1361
rect 12008 1302 12062 1309
rect 12108 1387 12162 1493
rect 12208 1571 12262 1578
rect 12208 1519 12209 1571
rect 12261 1519 12262 1571
rect 12208 1493 12218 1519
rect 12252 1493 12262 1519
rect 12208 1481 12262 1493
rect 12308 1527 12362 1633
rect 12408 1667 12462 1679
rect 12408 1641 12418 1667
rect 12452 1641 12462 1667
rect 12408 1589 12409 1641
rect 12461 1589 12462 1641
rect 12408 1582 12462 1589
rect 12508 1667 12562 1773
rect 12608 1851 12662 1858
rect 12608 1799 12609 1851
rect 12661 1799 12662 1851
rect 12608 1773 12618 1799
rect 12652 1773 12662 1799
rect 12608 1761 12662 1773
rect 12708 1807 12762 1913
rect 12808 1947 12862 1959
rect 12808 1921 12818 1947
rect 12852 1921 12862 1947
rect 12808 1869 12809 1921
rect 12861 1869 12862 1921
rect 12808 1862 12862 1869
rect 12906 1928 12916 1962
rect 12950 1928 12960 1962
rect 12906 1921 12960 1928
rect 12906 1869 12907 1921
rect 12959 1869 12960 1921
rect 12906 1862 12960 1869
rect 12906 1822 12960 1834
rect 12708 1773 12718 1807
rect 12752 1773 12762 1807
rect 12508 1633 12518 1667
rect 12552 1633 12562 1667
rect 12308 1493 12318 1527
rect 12352 1493 12362 1527
rect 12108 1353 12118 1387
rect 12152 1353 12162 1387
rect 12002 1273 12068 1274
rect 12002 1221 12009 1273
rect 12061 1221 12068 1273
rect 12002 1220 12068 1221
rect 11908 1123 11918 1157
rect 11952 1123 11962 1157
rect 11708 983 11718 1017
rect 11752 983 11762 1017
rect 11508 843 11518 877
rect 11552 843 11562 877
rect 11308 703 11318 737
rect 11352 703 11362 737
rect 11108 563 11118 597
rect 11152 563 11162 597
rect 10908 423 10918 457
rect 10952 423 10962 457
rect 10708 283 10718 317
rect 10752 283 10762 317
rect 10508 143 10518 177
rect 10552 143 10562 177
rect 10402 63 10468 64
rect 10402 11 10409 63
rect 10461 11 10468 63
rect 10402 10 10468 11
rect 10308 -67 10309 -15
rect 10361 -67 10362 -15
rect 10308 -79 10318 -67
rect 10352 -79 10362 -67
rect 10108 -132 10162 -131
rect 10108 -143 10118 -132
rect 10152 -143 10162 -132
rect 10108 -195 10109 -143
rect 10161 -195 10162 -143
rect 10108 -210 10162 -195
rect 10212 -133 10258 -81
rect 10212 -167 10218 -133
rect 10252 -167 10258 -133
rect 10118 -291 10125 -239
rect 10177 -291 10184 -239
rect 10012 -397 10018 -363
rect 10052 -397 10058 -363
rect 10012 -435 10058 -397
rect 10012 -469 10018 -435
rect 10052 -469 10058 -435
rect 10012 -512 10058 -469
rect 10109 -326 10161 -320
rect 10109 -390 10118 -378
rect 10152 -390 10161 -378
rect 10109 -454 10118 -442
rect 10152 -454 10161 -442
rect 10109 -512 10161 -506
rect 10212 -363 10258 -167
rect 10308 -131 10309 -79
rect 10361 -131 10362 -79
rect 10408 -22 10462 10
rect 10408 -74 10409 -22
rect 10461 -74 10462 -22
rect 10408 -81 10462 -74
rect 10508 -15 10562 143
rect 10608 221 10662 228
rect 10608 169 10609 221
rect 10661 169 10662 221
rect 10608 143 10618 169
rect 10652 143 10662 169
rect 10608 131 10662 143
rect 10708 177 10762 283
rect 10808 317 10862 329
rect 10808 291 10818 317
rect 10852 291 10862 317
rect 10808 239 10809 291
rect 10861 239 10862 291
rect 10808 232 10862 239
rect 10908 317 10962 423
rect 11008 501 11062 508
rect 11008 449 11009 501
rect 11061 449 11062 501
rect 11008 423 11018 449
rect 11052 423 11062 449
rect 11008 411 11062 423
rect 11108 457 11162 563
rect 11208 597 11262 609
rect 11208 571 11218 597
rect 11252 571 11262 597
rect 11208 519 11209 571
rect 11261 519 11262 571
rect 11208 512 11262 519
rect 11308 597 11362 703
rect 11408 781 11462 788
rect 11408 729 11409 781
rect 11461 729 11462 781
rect 11408 703 11418 729
rect 11452 703 11462 729
rect 11408 691 11462 703
rect 11508 737 11562 843
rect 11608 877 11662 889
rect 11608 851 11618 877
rect 11652 851 11662 877
rect 11608 799 11609 851
rect 11661 799 11662 851
rect 11608 792 11662 799
rect 11708 877 11762 983
rect 11808 1061 11862 1068
rect 11808 1009 11809 1061
rect 11861 1009 11862 1061
rect 11808 983 11818 1009
rect 11852 983 11862 1009
rect 11808 971 11862 983
rect 11908 1017 11962 1123
rect 12008 1157 12062 1169
rect 12008 1131 12018 1157
rect 12052 1131 12062 1157
rect 12008 1079 12009 1131
rect 12061 1079 12062 1131
rect 12008 1072 12062 1079
rect 12108 1157 12162 1353
rect 12208 1431 12262 1438
rect 12208 1379 12209 1431
rect 12261 1379 12262 1431
rect 12208 1353 12218 1379
rect 12252 1353 12262 1379
rect 12208 1341 12262 1353
rect 12308 1387 12362 1493
rect 12408 1527 12462 1539
rect 12408 1501 12418 1527
rect 12452 1501 12462 1527
rect 12408 1449 12409 1501
rect 12461 1449 12462 1501
rect 12408 1442 12462 1449
rect 12508 1527 12562 1633
rect 12608 1711 12662 1718
rect 12608 1659 12609 1711
rect 12661 1659 12662 1711
rect 12608 1633 12618 1659
rect 12652 1633 12662 1659
rect 12608 1621 12662 1633
rect 12708 1667 12762 1773
rect 12808 1807 12862 1819
rect 12808 1781 12818 1807
rect 12852 1781 12862 1807
rect 12808 1729 12809 1781
rect 12861 1729 12862 1781
rect 12808 1722 12862 1729
rect 12906 1788 12916 1822
rect 12950 1788 12960 1822
rect 12906 1781 12960 1788
rect 12906 1729 12907 1781
rect 12959 1729 12960 1781
rect 12906 1722 12960 1729
rect 12906 1682 12960 1694
rect 12708 1633 12718 1667
rect 12752 1633 12762 1667
rect 12508 1493 12518 1527
rect 12552 1493 12562 1527
rect 12308 1353 12318 1387
rect 12352 1353 12362 1387
rect 12202 1289 12268 1290
rect 12202 1237 12209 1289
rect 12261 1237 12268 1289
rect 12202 1236 12268 1237
rect 12108 1123 12118 1157
rect 12152 1123 12162 1157
rect 11908 983 11918 1017
rect 11952 983 11962 1017
rect 11708 843 11718 877
rect 11752 843 11762 877
rect 11508 703 11518 737
rect 11552 703 11562 737
rect 11308 563 11318 597
rect 11352 563 11362 597
rect 11108 423 11118 457
rect 11152 423 11162 457
rect 10908 283 10918 317
rect 10952 283 10962 317
rect 10708 143 10718 177
rect 10752 143 10762 177
rect 10602 79 10668 80
rect 10602 27 10609 79
rect 10661 27 10668 79
rect 10602 26 10668 27
rect 10508 -67 10509 -15
rect 10561 -67 10562 -15
rect 10508 -79 10518 -67
rect 10552 -79 10562 -67
rect 10308 -132 10362 -131
rect 10308 -143 10318 -132
rect 10352 -143 10362 -132
rect 10308 -195 10309 -143
rect 10361 -195 10362 -143
rect 10308 -210 10362 -195
rect 10412 -133 10458 -81
rect 10412 -167 10418 -133
rect 10452 -167 10458 -133
rect 10318 -291 10325 -239
rect 10377 -291 10384 -239
rect 10212 -397 10218 -363
rect 10252 -397 10258 -363
rect 10212 -435 10258 -397
rect 10212 -469 10218 -435
rect 10252 -469 10258 -435
rect 10212 -512 10258 -469
rect 10309 -326 10361 -320
rect 10309 -390 10318 -378
rect 10352 -390 10361 -378
rect 10309 -454 10318 -442
rect 10352 -454 10361 -442
rect 10309 -555 10361 -506
rect 10412 -363 10458 -167
rect 10508 -131 10509 -79
rect 10561 -131 10562 -79
rect 10608 -22 10662 26
rect 10608 -74 10609 -22
rect 10661 -74 10662 -22
rect 10608 -81 10662 -74
rect 10708 -15 10762 143
rect 10808 177 10862 189
rect 10808 151 10818 177
rect 10852 151 10862 177
rect 10808 99 10809 151
rect 10861 99 10862 151
rect 10808 92 10862 99
rect 10908 177 10962 283
rect 11008 361 11062 368
rect 11008 309 11009 361
rect 11061 309 11062 361
rect 11008 283 11018 309
rect 11052 283 11062 309
rect 11008 271 11062 283
rect 11108 317 11162 423
rect 11208 457 11262 469
rect 11208 431 11218 457
rect 11252 431 11262 457
rect 11208 379 11209 431
rect 11261 379 11262 431
rect 11208 372 11262 379
rect 11308 457 11362 563
rect 11408 641 11462 648
rect 11408 589 11409 641
rect 11461 589 11462 641
rect 11408 563 11418 589
rect 11452 563 11462 589
rect 11408 551 11462 563
rect 11508 597 11562 703
rect 11608 737 11662 749
rect 11608 711 11618 737
rect 11652 711 11662 737
rect 11608 659 11609 711
rect 11661 659 11662 711
rect 11608 652 11662 659
rect 11708 737 11762 843
rect 11808 921 11862 928
rect 11808 869 11809 921
rect 11861 869 11862 921
rect 11808 843 11818 869
rect 11852 843 11862 869
rect 11808 831 11862 843
rect 11908 877 11962 983
rect 12008 1017 12062 1029
rect 12008 991 12018 1017
rect 12052 991 12062 1017
rect 12008 939 12009 991
rect 12061 939 12062 991
rect 12008 932 12062 939
rect 12108 1017 12162 1123
rect 12208 1201 12262 1208
rect 12208 1149 12209 1201
rect 12261 1149 12262 1201
rect 12208 1123 12218 1149
rect 12252 1123 12262 1149
rect 12208 1111 12262 1123
rect 12308 1157 12362 1353
rect 12408 1387 12462 1399
rect 12408 1361 12418 1387
rect 12452 1361 12462 1387
rect 12408 1309 12409 1361
rect 12461 1309 12462 1361
rect 12408 1302 12462 1309
rect 12508 1387 12562 1493
rect 12608 1571 12662 1578
rect 12608 1519 12609 1571
rect 12661 1519 12662 1571
rect 12608 1493 12618 1519
rect 12652 1493 12662 1519
rect 12608 1481 12662 1493
rect 12708 1527 12762 1633
rect 12808 1667 12862 1679
rect 12808 1641 12818 1667
rect 12852 1641 12862 1667
rect 12808 1589 12809 1641
rect 12861 1589 12862 1641
rect 12808 1582 12862 1589
rect 12906 1648 12916 1682
rect 12950 1648 12960 1682
rect 12906 1641 12960 1648
rect 12906 1589 12907 1641
rect 12959 1589 12960 1641
rect 12906 1582 12960 1589
rect 12906 1542 12960 1554
rect 12708 1493 12718 1527
rect 12752 1493 12762 1527
rect 12508 1353 12518 1387
rect 12552 1353 12562 1387
rect 12402 1273 12468 1274
rect 12402 1221 12409 1273
rect 12461 1221 12468 1273
rect 12402 1220 12468 1221
rect 12308 1123 12318 1157
rect 12352 1123 12362 1157
rect 12108 983 12118 1017
rect 12152 983 12162 1017
rect 11908 843 11918 877
rect 11952 843 11962 877
rect 11708 703 11718 737
rect 11752 703 11762 737
rect 11508 563 11518 597
rect 11552 563 11562 597
rect 11308 423 11318 457
rect 11352 423 11362 457
rect 11108 283 11118 317
rect 11152 283 11162 317
rect 10908 143 10918 177
rect 10952 143 10962 177
rect 10802 63 10868 64
rect 10802 11 10809 63
rect 10861 11 10868 63
rect 10802 10 10868 11
rect 10708 -67 10709 -15
rect 10761 -67 10762 -15
rect 10708 -79 10718 -67
rect 10752 -79 10762 -67
rect 10508 -132 10562 -131
rect 10508 -143 10518 -132
rect 10552 -143 10562 -132
rect 10508 -195 10509 -143
rect 10561 -195 10562 -143
rect 10508 -210 10562 -195
rect 10612 -133 10658 -81
rect 10612 -167 10618 -133
rect 10652 -167 10658 -133
rect 10518 -291 10525 -239
rect 10577 -291 10584 -239
rect 10412 -397 10418 -363
rect 10452 -397 10458 -363
rect 10412 -435 10458 -397
rect 10412 -469 10418 -435
rect 10452 -469 10458 -435
rect 10412 -512 10458 -469
rect 10509 -326 10561 -320
rect 10509 -390 10518 -378
rect 10552 -390 10561 -378
rect 10509 -454 10518 -442
rect 10552 -454 10561 -442
rect 10509 -512 10561 -506
rect 10612 -363 10658 -167
rect 10708 -131 10709 -79
rect 10761 -131 10762 -79
rect 10808 -22 10862 10
rect 10808 -74 10809 -22
rect 10861 -74 10862 -22
rect 10808 -81 10862 -74
rect 10908 -15 10962 143
rect 11008 221 11062 228
rect 11008 169 11009 221
rect 11061 169 11062 221
rect 11008 143 11018 169
rect 11052 143 11062 169
rect 11008 131 11062 143
rect 11108 177 11162 283
rect 11208 317 11262 329
rect 11208 291 11218 317
rect 11252 291 11262 317
rect 11208 239 11209 291
rect 11261 239 11262 291
rect 11208 232 11262 239
rect 11308 317 11362 423
rect 11408 501 11462 508
rect 11408 449 11409 501
rect 11461 449 11462 501
rect 11408 423 11418 449
rect 11452 423 11462 449
rect 11408 411 11462 423
rect 11508 457 11562 563
rect 11608 597 11662 609
rect 11608 571 11618 597
rect 11652 571 11662 597
rect 11608 519 11609 571
rect 11661 519 11662 571
rect 11608 512 11662 519
rect 11708 597 11762 703
rect 11808 781 11862 788
rect 11808 729 11809 781
rect 11861 729 11862 781
rect 11808 703 11818 729
rect 11852 703 11862 729
rect 11808 691 11862 703
rect 11908 737 11962 843
rect 12008 877 12062 889
rect 12008 851 12018 877
rect 12052 851 12062 877
rect 12008 799 12009 851
rect 12061 799 12062 851
rect 12008 792 12062 799
rect 12108 877 12162 983
rect 12208 1061 12262 1068
rect 12208 1009 12209 1061
rect 12261 1009 12262 1061
rect 12208 983 12218 1009
rect 12252 983 12262 1009
rect 12208 971 12262 983
rect 12308 1017 12362 1123
rect 12408 1157 12462 1169
rect 12408 1131 12418 1157
rect 12452 1131 12462 1157
rect 12408 1079 12409 1131
rect 12461 1079 12462 1131
rect 12408 1072 12462 1079
rect 12508 1157 12562 1353
rect 12608 1431 12662 1438
rect 12608 1379 12609 1431
rect 12661 1379 12662 1431
rect 12608 1353 12618 1379
rect 12652 1353 12662 1379
rect 12608 1341 12662 1353
rect 12708 1387 12762 1493
rect 12808 1527 12862 1539
rect 12808 1501 12818 1527
rect 12852 1501 12862 1527
rect 12808 1449 12809 1501
rect 12861 1449 12862 1501
rect 12808 1442 12862 1449
rect 12906 1508 12916 1542
rect 12950 1508 12960 1542
rect 12906 1501 12960 1508
rect 12906 1449 12907 1501
rect 12959 1449 12960 1501
rect 12906 1442 12960 1449
rect 12906 1402 12960 1414
rect 12708 1353 12718 1387
rect 12752 1353 12762 1387
rect 12602 1289 12668 1290
rect 12602 1237 12609 1289
rect 12661 1237 12668 1289
rect 12602 1236 12668 1237
rect 12508 1123 12518 1157
rect 12552 1123 12562 1157
rect 12308 983 12318 1017
rect 12352 983 12362 1017
rect 12108 843 12118 877
rect 12152 843 12162 877
rect 11908 703 11918 737
rect 11952 703 11962 737
rect 11708 563 11718 597
rect 11752 563 11762 597
rect 11508 423 11518 457
rect 11552 423 11562 457
rect 11308 283 11318 317
rect 11352 283 11362 317
rect 11108 143 11118 177
rect 11152 143 11162 177
rect 11002 79 11068 80
rect 11002 27 11009 79
rect 11061 27 11068 79
rect 11002 26 11068 27
rect 10908 -67 10909 -15
rect 10961 -67 10962 -15
rect 10908 -79 10918 -67
rect 10952 -79 10962 -67
rect 10708 -132 10762 -131
rect 10708 -143 10718 -132
rect 10752 -143 10762 -132
rect 10708 -195 10709 -143
rect 10761 -195 10762 -143
rect 10708 -210 10762 -195
rect 10812 -133 10858 -81
rect 10812 -167 10818 -133
rect 10852 -167 10858 -133
rect 10718 -291 10725 -239
rect 10777 -291 10784 -239
rect 10612 -397 10618 -363
rect 10652 -397 10658 -363
rect 10612 -435 10658 -397
rect 10612 -469 10618 -435
rect 10652 -469 10658 -435
rect 10612 -512 10658 -469
rect 10709 -326 10761 -320
rect 10709 -390 10718 -378
rect 10752 -390 10761 -378
rect 10709 -454 10718 -442
rect 10752 -454 10761 -442
rect 10709 -555 10761 -506
rect 10812 -363 10858 -167
rect 10908 -131 10909 -79
rect 10961 -131 10962 -79
rect 11008 -22 11062 26
rect 11008 -74 11009 -22
rect 11061 -74 11062 -22
rect 11008 -81 11062 -74
rect 11108 -15 11162 143
rect 11208 177 11262 189
rect 11208 151 11218 177
rect 11252 151 11262 177
rect 11208 99 11209 151
rect 11261 99 11262 151
rect 11208 92 11262 99
rect 11308 177 11362 283
rect 11408 361 11462 368
rect 11408 309 11409 361
rect 11461 309 11462 361
rect 11408 283 11418 309
rect 11452 283 11462 309
rect 11408 271 11462 283
rect 11508 317 11562 423
rect 11608 457 11662 469
rect 11608 431 11618 457
rect 11652 431 11662 457
rect 11608 379 11609 431
rect 11661 379 11662 431
rect 11608 372 11662 379
rect 11708 457 11762 563
rect 11808 641 11862 648
rect 11808 589 11809 641
rect 11861 589 11862 641
rect 11808 563 11818 589
rect 11852 563 11862 589
rect 11808 551 11862 563
rect 11908 597 11962 703
rect 12008 737 12062 749
rect 12008 711 12018 737
rect 12052 711 12062 737
rect 12008 659 12009 711
rect 12061 659 12062 711
rect 12008 652 12062 659
rect 12108 737 12162 843
rect 12208 921 12262 928
rect 12208 869 12209 921
rect 12261 869 12262 921
rect 12208 843 12218 869
rect 12252 843 12262 869
rect 12208 831 12262 843
rect 12308 877 12362 983
rect 12408 1017 12462 1029
rect 12408 991 12418 1017
rect 12452 991 12462 1017
rect 12408 939 12409 991
rect 12461 939 12462 991
rect 12408 932 12462 939
rect 12508 1017 12562 1123
rect 12608 1201 12662 1208
rect 12608 1149 12609 1201
rect 12661 1149 12662 1201
rect 12608 1123 12618 1149
rect 12652 1123 12662 1149
rect 12608 1111 12662 1123
rect 12708 1157 12762 1353
rect 12808 1387 12862 1399
rect 12808 1361 12818 1387
rect 12852 1361 12862 1387
rect 12808 1309 12809 1361
rect 12861 1309 12862 1361
rect 12808 1302 12862 1309
rect 12906 1368 12916 1402
rect 12950 1368 12960 1402
rect 12906 1361 12960 1368
rect 12906 1309 12907 1361
rect 12959 1309 12960 1361
rect 12906 1302 12960 1309
rect 12990 1267 13020 2431
rect 12904 1261 13020 1267
rect 12904 1227 12916 1261
rect 12950 1227 13020 1261
rect 12904 1221 13020 1227
rect 12906 1172 12960 1184
rect 12708 1123 12718 1157
rect 12752 1123 12762 1157
rect 12508 983 12518 1017
rect 12552 983 12562 1017
rect 12308 843 12318 877
rect 12352 843 12362 877
rect 12108 703 12118 737
rect 12152 703 12162 737
rect 11908 563 11918 597
rect 11952 563 11962 597
rect 11708 423 11718 457
rect 11752 423 11762 457
rect 11508 283 11518 317
rect 11552 283 11562 317
rect 11308 143 11318 177
rect 11352 143 11362 177
rect 11202 63 11268 64
rect 11202 11 11209 63
rect 11261 11 11268 63
rect 11202 10 11268 11
rect 11108 -67 11109 -15
rect 11161 -67 11162 -15
rect 11108 -79 11118 -67
rect 11152 -79 11162 -67
rect 10908 -132 10962 -131
rect 10908 -143 10918 -132
rect 10952 -143 10962 -132
rect 10908 -195 10909 -143
rect 10961 -195 10962 -143
rect 10908 -210 10962 -195
rect 11012 -133 11058 -81
rect 11012 -167 11018 -133
rect 11052 -167 11058 -133
rect 10918 -291 10925 -239
rect 10977 -291 10984 -239
rect 10812 -397 10818 -363
rect 10852 -397 10858 -363
rect 10812 -435 10858 -397
rect 10812 -469 10818 -435
rect 10852 -469 10858 -435
rect 10812 -512 10858 -469
rect 10909 -326 10961 -320
rect 10909 -390 10918 -378
rect 10952 -390 10961 -378
rect 10909 -454 10918 -442
rect 10952 -454 10961 -442
rect 10909 -512 10961 -506
rect 11012 -363 11058 -167
rect 11108 -131 11109 -79
rect 11161 -131 11162 -79
rect 11208 -22 11262 10
rect 11208 -74 11209 -22
rect 11261 -74 11262 -22
rect 11208 -81 11262 -74
rect 11308 -15 11362 143
rect 11408 221 11462 228
rect 11408 169 11409 221
rect 11461 169 11462 221
rect 11408 143 11418 169
rect 11452 143 11462 169
rect 11408 131 11462 143
rect 11508 177 11562 283
rect 11608 317 11662 329
rect 11608 291 11618 317
rect 11652 291 11662 317
rect 11608 239 11609 291
rect 11661 239 11662 291
rect 11608 232 11662 239
rect 11708 317 11762 423
rect 11808 501 11862 508
rect 11808 449 11809 501
rect 11861 449 11862 501
rect 11808 423 11818 449
rect 11852 423 11862 449
rect 11808 411 11862 423
rect 11908 457 11962 563
rect 12008 597 12062 609
rect 12008 571 12018 597
rect 12052 571 12062 597
rect 12008 519 12009 571
rect 12061 519 12062 571
rect 12008 512 12062 519
rect 12108 597 12162 703
rect 12208 781 12262 788
rect 12208 729 12209 781
rect 12261 729 12262 781
rect 12208 703 12218 729
rect 12252 703 12262 729
rect 12208 691 12262 703
rect 12308 737 12362 843
rect 12408 877 12462 889
rect 12408 851 12418 877
rect 12452 851 12462 877
rect 12408 799 12409 851
rect 12461 799 12462 851
rect 12408 792 12462 799
rect 12508 877 12562 983
rect 12608 1061 12662 1068
rect 12608 1009 12609 1061
rect 12661 1009 12662 1061
rect 12608 983 12618 1009
rect 12652 983 12662 1009
rect 12608 971 12662 983
rect 12708 1017 12762 1123
rect 12808 1157 12862 1169
rect 12808 1131 12818 1157
rect 12852 1131 12862 1157
rect 12808 1079 12809 1131
rect 12861 1079 12862 1131
rect 12808 1072 12862 1079
rect 12906 1138 12916 1172
rect 12950 1138 12960 1172
rect 12906 1131 12960 1138
rect 12906 1079 12907 1131
rect 12959 1079 12960 1131
rect 12906 1072 12960 1079
rect 12906 1032 12960 1044
rect 12708 983 12718 1017
rect 12752 983 12762 1017
rect 12508 843 12518 877
rect 12552 843 12562 877
rect 12308 703 12318 737
rect 12352 703 12362 737
rect 12108 563 12118 597
rect 12152 563 12162 597
rect 11908 423 11918 457
rect 11952 423 11962 457
rect 11708 283 11718 317
rect 11752 283 11762 317
rect 11508 143 11518 177
rect 11552 143 11562 177
rect 11402 79 11468 80
rect 11402 27 11409 79
rect 11461 27 11468 79
rect 11402 26 11468 27
rect 11308 -67 11309 -15
rect 11361 -67 11362 -15
rect 11308 -79 11318 -67
rect 11352 -79 11362 -67
rect 11108 -132 11162 -131
rect 11108 -143 11118 -132
rect 11152 -143 11162 -132
rect 11108 -195 11109 -143
rect 11161 -195 11162 -143
rect 11108 -210 11162 -195
rect 11212 -133 11258 -81
rect 11212 -167 11218 -133
rect 11252 -167 11258 -133
rect 11118 -291 11125 -239
rect 11177 -291 11184 -239
rect 11012 -397 11018 -363
rect 11052 -397 11058 -363
rect 11012 -435 11058 -397
rect 11012 -469 11018 -435
rect 11052 -469 11058 -435
rect 11012 -512 11058 -469
rect 11109 -326 11161 -320
rect 11109 -390 11118 -378
rect 11152 -390 11161 -378
rect 11109 -454 11118 -442
rect 11152 -454 11161 -442
rect 11109 -555 11161 -506
rect 11212 -363 11258 -167
rect 11308 -131 11309 -79
rect 11361 -131 11362 -79
rect 11408 -22 11462 26
rect 11408 -74 11409 -22
rect 11461 -74 11462 -22
rect 11408 -81 11462 -74
rect 11508 -15 11562 143
rect 11608 177 11662 189
rect 11608 151 11618 177
rect 11652 151 11662 177
rect 11608 99 11609 151
rect 11661 99 11662 151
rect 11608 92 11662 99
rect 11708 177 11762 283
rect 11808 361 11862 368
rect 11808 309 11809 361
rect 11861 309 11862 361
rect 11808 283 11818 309
rect 11852 283 11862 309
rect 11808 271 11862 283
rect 11908 317 11962 423
rect 12008 457 12062 469
rect 12008 431 12018 457
rect 12052 431 12062 457
rect 12008 379 12009 431
rect 12061 379 12062 431
rect 12008 372 12062 379
rect 12108 457 12162 563
rect 12208 641 12262 648
rect 12208 589 12209 641
rect 12261 589 12262 641
rect 12208 563 12218 589
rect 12252 563 12262 589
rect 12208 551 12262 563
rect 12308 597 12362 703
rect 12408 737 12462 749
rect 12408 711 12418 737
rect 12452 711 12462 737
rect 12408 659 12409 711
rect 12461 659 12462 711
rect 12408 652 12462 659
rect 12508 737 12562 843
rect 12608 921 12662 928
rect 12608 869 12609 921
rect 12661 869 12662 921
rect 12608 843 12618 869
rect 12652 843 12662 869
rect 12608 831 12662 843
rect 12708 877 12762 983
rect 12808 1017 12862 1029
rect 12808 991 12818 1017
rect 12852 991 12862 1017
rect 12808 939 12809 991
rect 12861 939 12862 991
rect 12808 932 12862 939
rect 12906 998 12916 1032
rect 12950 998 12960 1032
rect 12906 991 12960 998
rect 12906 939 12907 991
rect 12959 939 12960 991
rect 12906 932 12960 939
rect 12906 892 12960 904
rect 12708 843 12718 877
rect 12752 843 12762 877
rect 12508 703 12518 737
rect 12552 703 12562 737
rect 12308 563 12318 597
rect 12352 563 12362 597
rect 12108 423 12118 457
rect 12152 423 12162 457
rect 11908 283 11918 317
rect 11952 283 11962 317
rect 11708 143 11718 177
rect 11752 143 11762 177
rect 11602 63 11668 64
rect 11602 11 11609 63
rect 11661 11 11668 63
rect 11602 10 11668 11
rect 11508 -67 11509 -15
rect 11561 -67 11562 -15
rect 11508 -79 11518 -67
rect 11552 -79 11562 -67
rect 11308 -132 11362 -131
rect 11308 -143 11318 -132
rect 11352 -143 11362 -132
rect 11308 -195 11309 -143
rect 11361 -195 11362 -143
rect 11308 -210 11362 -195
rect 11412 -133 11458 -81
rect 11412 -167 11418 -133
rect 11452 -167 11458 -133
rect 11318 -291 11325 -239
rect 11377 -291 11384 -239
rect 11212 -397 11218 -363
rect 11252 -397 11258 -363
rect 11212 -435 11258 -397
rect 11212 -469 11218 -435
rect 11252 -469 11258 -435
rect 11212 -512 11258 -469
rect 11309 -326 11361 -320
rect 11309 -390 11318 -378
rect 11352 -390 11361 -378
rect 11309 -454 11318 -442
rect 11352 -454 11361 -442
rect 11309 -512 11361 -506
rect 11412 -363 11458 -167
rect 11508 -131 11509 -79
rect 11561 -131 11562 -79
rect 11608 -22 11662 10
rect 11608 -74 11609 -22
rect 11661 -74 11662 -22
rect 11608 -81 11662 -74
rect 11708 -15 11762 143
rect 11808 221 11862 228
rect 11808 169 11809 221
rect 11861 169 11862 221
rect 11808 143 11818 169
rect 11852 143 11862 169
rect 11808 131 11862 143
rect 11908 177 11962 283
rect 12008 317 12062 329
rect 12008 291 12018 317
rect 12052 291 12062 317
rect 12008 239 12009 291
rect 12061 239 12062 291
rect 12008 232 12062 239
rect 12108 317 12162 423
rect 12208 501 12262 508
rect 12208 449 12209 501
rect 12261 449 12262 501
rect 12208 423 12218 449
rect 12252 423 12262 449
rect 12208 411 12262 423
rect 12308 457 12362 563
rect 12408 597 12462 609
rect 12408 571 12418 597
rect 12452 571 12462 597
rect 12408 519 12409 571
rect 12461 519 12462 571
rect 12408 512 12462 519
rect 12508 597 12562 703
rect 12608 781 12662 788
rect 12608 729 12609 781
rect 12661 729 12662 781
rect 12608 703 12618 729
rect 12652 703 12662 729
rect 12608 691 12662 703
rect 12708 737 12762 843
rect 12808 877 12862 889
rect 12808 851 12818 877
rect 12852 851 12862 877
rect 12808 799 12809 851
rect 12861 799 12862 851
rect 12808 792 12862 799
rect 12906 858 12916 892
rect 12950 858 12960 892
rect 12906 851 12960 858
rect 12906 799 12907 851
rect 12959 799 12960 851
rect 12906 792 12960 799
rect 12906 752 12960 764
rect 12708 703 12718 737
rect 12752 703 12762 737
rect 12508 563 12518 597
rect 12552 563 12562 597
rect 12308 423 12318 457
rect 12352 423 12362 457
rect 12108 283 12118 317
rect 12152 283 12162 317
rect 11908 143 11918 177
rect 11952 143 11962 177
rect 11802 79 11868 80
rect 11802 27 11809 79
rect 11861 27 11868 79
rect 11802 26 11868 27
rect 11708 -67 11709 -15
rect 11761 -67 11762 -15
rect 11708 -79 11718 -67
rect 11752 -79 11762 -67
rect 11508 -132 11562 -131
rect 11508 -143 11518 -132
rect 11552 -143 11562 -132
rect 11508 -195 11509 -143
rect 11561 -195 11562 -143
rect 11508 -210 11562 -195
rect 11612 -133 11658 -81
rect 11612 -167 11618 -133
rect 11652 -167 11658 -133
rect 11518 -291 11525 -239
rect 11577 -291 11584 -239
rect 11412 -397 11418 -363
rect 11452 -397 11458 -363
rect 11412 -435 11458 -397
rect 11412 -469 11418 -435
rect 11452 -469 11458 -435
rect 11412 -512 11458 -469
rect 11509 -326 11561 -320
rect 11509 -390 11518 -378
rect 11552 -390 11561 -378
rect 11509 -454 11518 -442
rect 11552 -454 11561 -442
rect 11509 -555 11561 -506
rect 11612 -363 11658 -167
rect 11708 -131 11709 -79
rect 11761 -131 11762 -79
rect 11808 -22 11862 26
rect 11808 -74 11809 -22
rect 11861 -74 11862 -22
rect 11808 -81 11862 -74
rect 11908 -15 11962 143
rect 12008 177 12062 189
rect 12008 151 12018 177
rect 12052 151 12062 177
rect 12008 99 12009 151
rect 12061 99 12062 151
rect 12008 92 12062 99
rect 12108 177 12162 283
rect 12208 361 12262 368
rect 12208 309 12209 361
rect 12261 309 12262 361
rect 12208 283 12218 309
rect 12252 283 12262 309
rect 12208 271 12262 283
rect 12308 317 12362 423
rect 12408 457 12462 469
rect 12408 431 12418 457
rect 12452 431 12462 457
rect 12408 379 12409 431
rect 12461 379 12462 431
rect 12408 372 12462 379
rect 12508 457 12562 563
rect 12608 641 12662 648
rect 12608 589 12609 641
rect 12661 589 12662 641
rect 12608 563 12618 589
rect 12652 563 12662 589
rect 12608 551 12662 563
rect 12708 597 12762 703
rect 12808 737 12862 749
rect 12808 711 12818 737
rect 12852 711 12862 737
rect 12808 659 12809 711
rect 12861 659 12862 711
rect 12808 652 12862 659
rect 12906 718 12916 752
rect 12950 718 12960 752
rect 12906 711 12960 718
rect 12906 659 12907 711
rect 12959 659 12960 711
rect 12906 652 12960 659
rect 12906 612 12960 624
rect 12708 563 12718 597
rect 12752 563 12762 597
rect 12508 423 12518 457
rect 12552 423 12562 457
rect 12308 283 12318 317
rect 12352 283 12362 317
rect 12108 143 12118 177
rect 12152 143 12162 177
rect 12002 63 12068 64
rect 12002 11 12009 63
rect 12061 11 12068 63
rect 12002 10 12068 11
rect 11908 -67 11909 -15
rect 11961 -67 11962 -15
rect 11908 -79 11918 -67
rect 11952 -79 11962 -67
rect 11708 -132 11762 -131
rect 11708 -143 11718 -132
rect 11752 -143 11762 -132
rect 11708 -195 11709 -143
rect 11761 -195 11762 -143
rect 11708 -210 11762 -195
rect 11812 -133 11858 -81
rect 11812 -167 11818 -133
rect 11852 -167 11858 -133
rect 11718 -291 11725 -239
rect 11777 -291 11784 -239
rect 11612 -397 11618 -363
rect 11652 -397 11658 -363
rect 11612 -435 11658 -397
rect 11612 -469 11618 -435
rect 11652 -469 11658 -435
rect 11612 -512 11658 -469
rect 11709 -326 11761 -320
rect 11709 -390 11718 -378
rect 11752 -390 11761 -378
rect 11709 -454 11718 -442
rect 11752 -454 11761 -442
rect 11709 -512 11761 -506
rect 11812 -363 11858 -167
rect 11908 -131 11909 -79
rect 11961 -131 11962 -79
rect 12008 -22 12062 10
rect 12008 -74 12009 -22
rect 12061 -74 12062 -22
rect 12008 -81 12062 -74
rect 12108 -15 12162 143
rect 12208 221 12262 228
rect 12208 169 12209 221
rect 12261 169 12262 221
rect 12208 143 12218 169
rect 12252 143 12262 169
rect 12208 131 12262 143
rect 12308 177 12362 283
rect 12408 317 12462 329
rect 12408 291 12418 317
rect 12452 291 12462 317
rect 12408 239 12409 291
rect 12461 239 12462 291
rect 12408 232 12462 239
rect 12508 317 12562 423
rect 12608 501 12662 508
rect 12608 449 12609 501
rect 12661 449 12662 501
rect 12608 423 12618 449
rect 12652 423 12662 449
rect 12608 411 12662 423
rect 12708 457 12762 563
rect 12808 597 12862 609
rect 12808 571 12818 597
rect 12852 571 12862 597
rect 12808 519 12809 571
rect 12861 519 12862 571
rect 12808 512 12862 519
rect 12906 578 12916 612
rect 12950 578 12960 612
rect 12906 571 12960 578
rect 12906 519 12907 571
rect 12959 519 12960 571
rect 12906 512 12960 519
rect 12906 472 12960 484
rect 12708 423 12718 457
rect 12752 423 12762 457
rect 12508 283 12518 317
rect 12552 283 12562 317
rect 12308 143 12318 177
rect 12352 143 12362 177
rect 12202 79 12268 80
rect 12202 27 12209 79
rect 12261 27 12268 79
rect 12202 26 12268 27
rect 12108 -67 12109 -15
rect 12161 -67 12162 -15
rect 12108 -79 12118 -67
rect 12152 -79 12162 -67
rect 11908 -132 11962 -131
rect 11908 -143 11918 -132
rect 11952 -143 11962 -132
rect 11908 -195 11909 -143
rect 11961 -195 11962 -143
rect 11908 -210 11962 -195
rect 12012 -133 12058 -81
rect 12012 -167 12018 -133
rect 12052 -167 12058 -133
rect 11918 -291 11925 -239
rect 11977 -291 11984 -239
rect 11812 -397 11818 -363
rect 11852 -397 11858 -363
rect 11812 -435 11858 -397
rect 11812 -469 11818 -435
rect 11852 -469 11858 -435
rect 11812 -512 11858 -469
rect 11909 -326 11961 -320
rect 11909 -390 11918 -378
rect 11952 -390 11961 -378
rect 11909 -454 11918 -442
rect 11952 -454 11961 -442
rect 11909 -555 11961 -506
rect 12012 -363 12058 -167
rect 12108 -131 12109 -79
rect 12161 -131 12162 -79
rect 12208 -22 12262 26
rect 12208 -74 12209 -22
rect 12261 -74 12262 -22
rect 12208 -81 12262 -74
rect 12308 -15 12362 143
rect 12408 177 12462 189
rect 12408 151 12418 177
rect 12452 151 12462 177
rect 12408 99 12409 151
rect 12461 99 12462 151
rect 12408 92 12462 99
rect 12508 177 12562 283
rect 12608 361 12662 368
rect 12608 309 12609 361
rect 12661 309 12662 361
rect 12608 283 12618 309
rect 12652 283 12662 309
rect 12608 271 12662 283
rect 12708 317 12762 423
rect 12808 457 12862 469
rect 12808 431 12818 457
rect 12852 431 12862 457
rect 12808 379 12809 431
rect 12861 379 12862 431
rect 12808 372 12862 379
rect 12906 438 12916 472
rect 12950 438 12960 472
rect 12906 431 12960 438
rect 12906 379 12907 431
rect 12959 379 12960 431
rect 12906 372 12960 379
rect 12906 332 12960 344
rect 12708 283 12718 317
rect 12752 283 12762 317
rect 12508 143 12518 177
rect 12552 143 12562 177
rect 12402 63 12468 64
rect 12402 11 12409 63
rect 12461 11 12468 63
rect 12402 10 12468 11
rect 12308 -67 12309 -15
rect 12361 -67 12362 -15
rect 12308 -79 12318 -67
rect 12352 -79 12362 -67
rect 12108 -132 12162 -131
rect 12108 -143 12118 -132
rect 12152 -143 12162 -132
rect 12108 -195 12109 -143
rect 12161 -195 12162 -143
rect 12108 -210 12162 -195
rect 12212 -133 12258 -81
rect 12212 -167 12218 -133
rect 12252 -167 12258 -133
rect 12118 -291 12125 -239
rect 12177 -291 12184 -239
rect 12012 -397 12018 -363
rect 12052 -397 12058 -363
rect 12012 -435 12058 -397
rect 12012 -469 12018 -435
rect 12052 -469 12058 -435
rect 12012 -512 12058 -469
rect 12109 -326 12161 -320
rect 12109 -390 12118 -378
rect 12152 -390 12161 -378
rect 12109 -454 12118 -442
rect 12152 -454 12161 -442
rect 12109 -512 12161 -506
rect 12212 -363 12258 -167
rect 12308 -131 12309 -79
rect 12361 -131 12362 -79
rect 12408 -22 12462 10
rect 12408 -74 12409 -22
rect 12461 -74 12462 -22
rect 12408 -81 12462 -74
rect 12508 -15 12562 143
rect 12608 221 12662 228
rect 12608 169 12609 221
rect 12661 169 12662 221
rect 12608 143 12618 169
rect 12652 143 12662 169
rect 12608 131 12662 143
rect 12708 177 12762 283
rect 12808 317 12862 329
rect 12808 291 12818 317
rect 12852 291 12862 317
rect 12808 239 12809 291
rect 12861 239 12862 291
rect 12808 232 12862 239
rect 12906 298 12916 332
rect 12950 298 12960 332
rect 12906 291 12960 298
rect 12906 239 12907 291
rect 12959 239 12960 291
rect 12906 232 12960 239
rect 12906 192 12960 204
rect 12708 143 12718 177
rect 12752 143 12762 177
rect 12602 79 12668 80
rect 12602 27 12609 79
rect 12661 27 12668 79
rect 12602 26 12668 27
rect 12508 -67 12509 -15
rect 12561 -67 12562 -15
rect 12508 -79 12518 -67
rect 12552 -79 12562 -67
rect 12308 -132 12362 -131
rect 12308 -143 12318 -132
rect 12352 -143 12362 -132
rect 12308 -195 12309 -143
rect 12361 -195 12362 -143
rect 12308 -210 12362 -195
rect 12412 -133 12458 -81
rect 12412 -167 12418 -133
rect 12452 -167 12458 -133
rect 12318 -291 12325 -239
rect 12377 -291 12384 -239
rect 12212 -397 12218 -363
rect 12252 -397 12258 -363
rect 12212 -435 12258 -397
rect 12212 -469 12218 -435
rect 12252 -469 12258 -435
rect 12212 -512 12258 -469
rect 12309 -326 12361 -320
rect 12309 -390 12318 -378
rect 12352 -390 12361 -378
rect 12309 -454 12318 -442
rect 12352 -454 12361 -442
rect 12309 -555 12361 -506
rect 12412 -363 12458 -167
rect 12508 -131 12509 -79
rect 12561 -131 12562 -79
rect 12608 -22 12662 26
rect 12608 -74 12609 -22
rect 12661 -74 12662 -22
rect 12608 -81 12662 -74
rect 12708 -15 12762 143
rect 12808 177 12862 189
rect 12808 151 12818 177
rect 12852 151 12862 177
rect 12808 99 12809 151
rect 12861 99 12862 151
rect 12808 92 12862 99
rect 12906 158 12916 192
rect 12950 158 12960 192
rect 12906 151 12960 158
rect 12906 99 12907 151
rect 12959 99 12960 151
rect 12906 92 12960 99
rect 12990 57 13020 1221
rect 12904 51 13020 57
rect 12904 17 12916 51
rect 12950 17 13020 51
rect 12904 11 13020 17
rect 12990 0 13020 11
rect 13050 4919 13080 5070
rect 13280 4920 13310 5070
rect 13380 4920 13410 5070
rect 13480 4920 13510 5070
rect 13580 4920 13610 5070
rect 13050 4913 13166 4919
rect 13050 4879 13120 4913
rect 13154 4879 13166 4913
rect 13050 4873 13166 4879
rect 13272 4908 13318 4920
rect 13272 4874 13278 4908
rect 13312 4874 13318 4908
rect 13050 3709 13080 4873
rect 13272 4862 13318 4874
rect 13372 4908 13418 4920
rect 13372 4874 13378 4908
rect 13412 4874 13418 4908
rect 13372 4862 13418 4874
rect 13472 4908 13518 4920
rect 13472 4874 13478 4908
rect 13512 4874 13518 4908
rect 13472 4862 13518 4874
rect 13572 4908 13618 4920
rect 13572 4874 13578 4908
rect 13612 4874 13618 4908
rect 13572 4862 13618 4874
rect 13110 4831 13164 4838
rect 13110 4779 13111 4831
rect 13163 4779 13164 4831
rect 13110 4772 13164 4779
rect 13110 4738 13120 4772
rect 13154 4738 13164 4772
rect 13110 4726 13164 4738
rect 13110 4691 13164 4698
rect 13110 4639 13111 4691
rect 13163 4639 13164 4691
rect 13110 4632 13164 4639
rect 13110 4598 13120 4632
rect 13154 4598 13164 4632
rect 13110 4586 13164 4598
rect 13110 4551 13164 4558
rect 13110 4499 13111 4551
rect 13163 4499 13164 4551
rect 13110 4492 13164 4499
rect 13110 4458 13120 4492
rect 13154 4458 13164 4492
rect 13110 4446 13164 4458
rect 13110 4411 13164 4418
rect 13110 4359 13111 4411
rect 13163 4359 13164 4411
rect 13110 4352 13164 4359
rect 13110 4318 13120 4352
rect 13154 4318 13164 4352
rect 13110 4306 13164 4318
rect 13110 4271 13164 4278
rect 13110 4219 13111 4271
rect 13163 4219 13164 4271
rect 13110 4212 13164 4219
rect 13110 4178 13120 4212
rect 13154 4178 13164 4212
rect 13110 4166 13164 4178
rect 13110 4131 13164 4138
rect 13110 4079 13111 4131
rect 13163 4079 13164 4131
rect 13110 4072 13164 4079
rect 13110 4038 13120 4072
rect 13154 4038 13164 4072
rect 13110 4026 13164 4038
rect 13110 3991 13164 3998
rect 13110 3939 13111 3991
rect 13163 3939 13164 3991
rect 13110 3932 13164 3939
rect 13110 3898 13120 3932
rect 13154 3898 13164 3932
rect 13110 3886 13164 3898
rect 13110 3851 13164 3858
rect 13110 3799 13111 3851
rect 13163 3799 13164 3851
rect 13110 3792 13164 3799
rect 13110 3758 13120 3792
rect 13154 3758 13164 3792
rect 13110 3746 13164 3758
rect 13280 3710 13310 4862
rect 13380 3710 13410 4862
rect 13480 3710 13510 4862
rect 13580 3710 13610 4862
rect 13050 3703 13166 3709
rect 13050 3669 13120 3703
rect 13154 3669 13166 3703
rect 13050 3663 13166 3669
rect 13272 3698 13318 3710
rect 13272 3664 13278 3698
rect 13312 3664 13318 3698
rect 13050 2499 13080 3663
rect 13272 3652 13318 3664
rect 13372 3698 13418 3710
rect 13372 3664 13378 3698
rect 13412 3664 13418 3698
rect 13372 3652 13418 3664
rect 13472 3698 13518 3710
rect 13472 3664 13478 3698
rect 13512 3664 13518 3698
rect 13472 3652 13518 3664
rect 13572 3698 13618 3710
rect 13572 3664 13578 3698
rect 13612 3664 13618 3698
rect 13572 3652 13618 3664
rect 13110 3621 13164 3628
rect 13110 3569 13111 3621
rect 13163 3569 13164 3621
rect 13110 3562 13164 3569
rect 13110 3528 13120 3562
rect 13154 3528 13164 3562
rect 13110 3516 13164 3528
rect 13110 3481 13164 3488
rect 13110 3429 13111 3481
rect 13163 3429 13164 3481
rect 13110 3422 13164 3429
rect 13110 3388 13120 3422
rect 13154 3388 13164 3422
rect 13110 3376 13164 3388
rect 13110 3341 13164 3348
rect 13110 3289 13111 3341
rect 13163 3289 13164 3341
rect 13110 3282 13164 3289
rect 13110 3248 13120 3282
rect 13154 3248 13164 3282
rect 13110 3236 13164 3248
rect 13110 3201 13164 3208
rect 13110 3149 13111 3201
rect 13163 3149 13164 3201
rect 13110 3142 13164 3149
rect 13110 3108 13120 3142
rect 13154 3108 13164 3142
rect 13110 3096 13164 3108
rect 13110 3061 13164 3068
rect 13110 3009 13111 3061
rect 13163 3009 13164 3061
rect 13110 3002 13164 3009
rect 13110 2968 13120 3002
rect 13154 2968 13164 3002
rect 13110 2956 13164 2968
rect 13110 2921 13164 2928
rect 13110 2869 13111 2921
rect 13163 2869 13164 2921
rect 13110 2862 13164 2869
rect 13110 2828 13120 2862
rect 13154 2828 13164 2862
rect 13110 2816 13164 2828
rect 13110 2781 13164 2788
rect 13110 2729 13111 2781
rect 13163 2729 13164 2781
rect 13110 2722 13164 2729
rect 13110 2688 13120 2722
rect 13154 2688 13164 2722
rect 13110 2676 13164 2688
rect 13110 2641 13164 2648
rect 13110 2589 13111 2641
rect 13163 2589 13164 2641
rect 13110 2582 13164 2589
rect 13110 2548 13120 2582
rect 13154 2548 13164 2582
rect 13110 2536 13164 2548
rect 13280 2500 13310 3652
rect 13380 2500 13410 3652
rect 13480 2500 13510 3652
rect 13580 2500 13610 3652
rect 13050 2493 13166 2499
rect 13050 2459 13120 2493
rect 13154 2459 13166 2493
rect 13050 2453 13166 2459
rect 13272 2488 13318 2500
rect 13272 2454 13278 2488
rect 13312 2454 13318 2488
rect 13050 1289 13080 2453
rect 13272 2442 13318 2454
rect 13372 2488 13418 2500
rect 13372 2454 13378 2488
rect 13412 2454 13418 2488
rect 13372 2442 13418 2454
rect 13472 2488 13518 2500
rect 13472 2454 13478 2488
rect 13512 2454 13518 2488
rect 13472 2442 13518 2454
rect 13572 2488 13618 2500
rect 13572 2454 13578 2488
rect 13612 2454 13618 2488
rect 13572 2442 13618 2454
rect 13110 2411 13164 2418
rect 13110 2359 13111 2411
rect 13163 2359 13164 2411
rect 13110 2352 13164 2359
rect 13110 2318 13120 2352
rect 13154 2318 13164 2352
rect 13110 2306 13164 2318
rect 13110 2271 13164 2278
rect 13110 2219 13111 2271
rect 13163 2219 13164 2271
rect 13110 2212 13164 2219
rect 13110 2178 13120 2212
rect 13154 2178 13164 2212
rect 13110 2166 13164 2178
rect 13110 2131 13164 2138
rect 13110 2079 13111 2131
rect 13163 2079 13164 2131
rect 13110 2072 13164 2079
rect 13110 2038 13120 2072
rect 13154 2038 13164 2072
rect 13110 2026 13164 2038
rect 13110 1991 13164 1998
rect 13110 1939 13111 1991
rect 13163 1939 13164 1991
rect 13110 1932 13164 1939
rect 13110 1898 13120 1932
rect 13154 1898 13164 1932
rect 13110 1886 13164 1898
rect 13110 1851 13164 1858
rect 13110 1799 13111 1851
rect 13163 1799 13164 1851
rect 13110 1792 13164 1799
rect 13110 1758 13120 1792
rect 13154 1758 13164 1792
rect 13110 1746 13164 1758
rect 13110 1711 13164 1718
rect 13110 1659 13111 1711
rect 13163 1659 13164 1711
rect 13110 1652 13164 1659
rect 13110 1618 13120 1652
rect 13154 1618 13164 1652
rect 13110 1606 13164 1618
rect 13110 1571 13164 1578
rect 13110 1519 13111 1571
rect 13163 1519 13164 1571
rect 13110 1512 13164 1519
rect 13110 1478 13120 1512
rect 13154 1478 13164 1512
rect 13110 1466 13164 1478
rect 13110 1431 13164 1438
rect 13110 1379 13111 1431
rect 13163 1379 13164 1431
rect 13110 1372 13164 1379
rect 13110 1338 13120 1372
rect 13154 1338 13164 1372
rect 13110 1326 13164 1338
rect 13280 1290 13310 2442
rect 13380 1290 13410 2442
rect 13480 1290 13510 2442
rect 13580 1290 13610 2442
rect 13050 1283 13166 1289
rect 13050 1249 13120 1283
rect 13154 1249 13166 1283
rect 13050 1243 13166 1249
rect 13272 1278 13318 1290
rect 13272 1244 13278 1278
rect 13312 1244 13318 1278
rect 13050 79 13080 1243
rect 13272 1232 13318 1244
rect 13372 1278 13418 1290
rect 13372 1244 13378 1278
rect 13412 1244 13418 1278
rect 13372 1232 13418 1244
rect 13472 1278 13518 1290
rect 13472 1244 13478 1278
rect 13512 1244 13518 1278
rect 13472 1232 13518 1244
rect 13572 1278 13618 1290
rect 13572 1244 13578 1278
rect 13612 1244 13618 1278
rect 13572 1232 13618 1244
rect 13110 1201 13164 1208
rect 13110 1149 13111 1201
rect 13163 1149 13164 1201
rect 13110 1142 13164 1149
rect 13110 1108 13120 1142
rect 13154 1108 13164 1142
rect 13110 1096 13164 1108
rect 13110 1061 13164 1068
rect 13110 1009 13111 1061
rect 13163 1009 13164 1061
rect 13110 1002 13164 1009
rect 13110 968 13120 1002
rect 13154 968 13164 1002
rect 13110 956 13164 968
rect 13110 921 13164 928
rect 13110 869 13111 921
rect 13163 869 13164 921
rect 13110 862 13164 869
rect 13110 828 13120 862
rect 13154 828 13164 862
rect 13110 816 13164 828
rect 13110 781 13164 788
rect 13110 729 13111 781
rect 13163 729 13164 781
rect 13110 722 13164 729
rect 13110 688 13120 722
rect 13154 688 13164 722
rect 13110 676 13164 688
rect 13110 641 13164 648
rect 13110 589 13111 641
rect 13163 589 13164 641
rect 13110 582 13164 589
rect 13110 548 13120 582
rect 13154 548 13164 582
rect 13110 536 13164 548
rect 13110 501 13164 508
rect 13110 449 13111 501
rect 13163 449 13164 501
rect 13110 442 13164 449
rect 13110 408 13120 442
rect 13154 408 13164 442
rect 13110 396 13164 408
rect 13110 361 13164 368
rect 13110 309 13111 361
rect 13163 309 13164 361
rect 13110 302 13164 309
rect 13110 268 13120 302
rect 13154 268 13164 302
rect 13110 256 13164 268
rect 13110 221 13164 228
rect 13110 169 13111 221
rect 13163 169 13164 221
rect 13110 162 13164 169
rect 13110 128 13120 162
rect 13154 128 13164 162
rect 13110 116 13164 128
rect 13280 80 13310 1232
rect 13380 80 13410 1232
rect 13480 80 13510 1232
rect 13580 80 13610 1232
rect 13050 73 13166 79
rect 13050 39 13120 73
rect 13154 39 13166 73
rect 13050 33 13166 39
rect 13272 68 13318 80
rect 13272 34 13278 68
rect 13312 34 13318 68
rect 13050 0 13080 33
rect 13272 22 13318 34
rect 13372 68 13418 80
rect 13372 34 13378 68
rect 13412 34 13418 68
rect 13372 22 13418 34
rect 13472 68 13518 80
rect 13472 34 13478 68
rect 13512 34 13518 68
rect 13472 22 13518 34
rect 13572 68 13618 80
rect 13572 34 13578 68
rect 13612 34 13618 68
rect 13572 22 13618 34
rect 13280 0 13310 22
rect 13380 0 13410 22
rect 13480 0 13510 22
rect 13580 0 13610 22
rect 12708 -67 12709 -15
rect 12761 -67 12762 -15
rect 12708 -79 12718 -67
rect 12752 -79 12762 -67
rect 12508 -132 12562 -131
rect 12508 -143 12518 -132
rect 12552 -143 12562 -132
rect 12508 -195 12509 -143
rect 12561 -195 12562 -143
rect 12508 -210 12562 -195
rect 12612 -133 12658 -81
rect 12612 -167 12618 -133
rect 12652 -167 12658 -133
rect 12518 -291 12525 -239
rect 12577 -291 12584 -239
rect 12412 -397 12418 -363
rect 12452 -397 12458 -363
rect 12412 -435 12458 -397
rect 12412 -469 12418 -435
rect 12452 -469 12458 -435
rect 12412 -512 12458 -469
rect 12509 -326 12561 -320
rect 12509 -390 12518 -378
rect 12552 -390 12561 -378
rect 12509 -454 12518 -442
rect 12552 -454 12561 -442
rect 12509 -512 12561 -506
rect 12612 -363 12658 -167
rect 12708 -131 12709 -79
rect 12761 -131 12762 -79
rect 12708 -132 12762 -131
rect 12708 -143 12718 -132
rect 12752 -143 12762 -132
rect 12708 -195 12709 -143
rect 12761 -195 12762 -143
rect 12708 -210 12762 -195
rect 14526 -199 14697 -193
rect 14526 -251 14553 -199
rect 14605 -251 14617 -199
rect 14669 -251 14697 -199
rect 14526 -257 14697 -251
rect 14805 -199 15136 -193
rect 14805 -251 14816 -199
rect 14868 -208 14880 -199
rect 14932 -208 14944 -199
rect 14996 -208 15008 -199
rect 15060 -208 15072 -199
rect 14876 -242 14880 -208
rect 14868 -251 14880 -242
rect 14932 -251 14944 -242
rect 14996 -251 15008 -242
rect 15060 -251 15072 -242
rect 15124 -251 15136 -199
rect 14805 -257 15136 -251
rect 15206 -199 15537 -193
rect 15206 -251 15217 -199
rect 15269 -208 15281 -199
rect 15333 -208 15345 -199
rect 15397 -208 15409 -199
rect 15461 -208 15473 -199
rect 15461 -242 15465 -208
rect 15269 -251 15281 -242
rect 15333 -251 15345 -242
rect 15397 -251 15409 -242
rect 15461 -251 15473 -242
rect 15525 -251 15537 -199
rect 15206 -257 15537 -251
rect 15645 -199 15816 -193
rect 15645 -251 15672 -199
rect 15724 -251 15736 -199
rect 15788 -251 15816 -199
rect 15645 -257 15816 -251
rect 14520 -308 15136 -302
rect 14520 -310 14560 -308
rect 12612 -397 12618 -363
rect 12652 -397 12658 -363
rect 12612 -435 12658 -397
rect 12612 -469 12618 -435
rect 12652 -469 12658 -435
rect 12612 -512 12658 -469
rect 12709 -326 12761 -320
rect 14400 -340 14560 -310
rect 14520 -342 14560 -340
rect 14594 -342 14632 -308
rect 14666 -342 14841 -308
rect 14875 -342 14913 -308
rect 14947 -342 14985 -308
rect 15019 -342 15057 -308
rect 15091 -342 15136 -308
rect 14520 -348 15136 -342
rect 15206 -351 15212 -299
rect 15264 -302 15270 -299
rect 15264 -308 15822 -302
rect 15285 -342 15323 -308
rect 15357 -342 15395 -308
rect 15429 -342 15467 -308
rect 15501 -342 15676 -308
rect 15710 -342 15748 -308
rect 15782 -342 15822 -308
rect 15264 -348 15822 -342
rect 15264 -351 15270 -348
rect 12709 -390 12718 -378
rect 12752 -390 12761 -378
rect 14526 -399 14697 -393
rect 14434 -410 14440 -399
rect 14400 -440 14440 -410
rect 12709 -454 12718 -442
rect 12752 -454 12761 -442
rect 14434 -451 14440 -440
rect 14492 -451 14498 -399
rect 14526 -451 14553 -399
rect 14605 -451 14617 -399
rect 14669 -451 14697 -399
rect 14526 -457 14697 -451
rect 14725 -399 14777 -393
rect 14725 -457 14777 -451
rect 14805 -399 15136 -393
rect 14805 -451 14816 -399
rect 14868 -408 14880 -399
rect 14932 -408 14944 -399
rect 14996 -408 15008 -399
rect 15060 -408 15072 -399
rect 14876 -442 14880 -408
rect 14868 -451 14880 -442
rect 14932 -451 14944 -442
rect 14996 -451 15008 -442
rect 15060 -451 15072 -442
rect 15124 -451 15136 -399
rect 14805 -457 15136 -451
rect 15206 -399 15537 -393
rect 15206 -451 15217 -399
rect 15269 -408 15281 -399
rect 15333 -408 15345 -399
rect 15397 -408 15409 -399
rect 15461 -408 15473 -399
rect 15461 -442 15465 -408
rect 15269 -451 15281 -442
rect 15333 -451 15345 -442
rect 15397 -451 15409 -442
rect 15461 -451 15473 -442
rect 15525 -451 15537 -399
rect 15206 -457 15537 -451
rect 15565 -399 15617 -393
rect 15565 -457 15617 -451
rect 15645 -399 15816 -393
rect 15645 -451 15672 -399
rect 15724 -451 15736 -399
rect 15788 -451 15816 -399
rect 15645 -457 15816 -451
rect 12709 -555 12761 -506
rect 14520 -508 15136 -502
rect 14520 -510 14560 -508
rect 14400 -540 14560 -510
rect 14520 -542 14560 -540
rect 14594 -542 14632 -508
rect 14666 -542 14841 -508
rect 14875 -542 14913 -508
rect 14947 -542 14985 -508
rect 15019 -542 15057 -508
rect 15091 -542 15136 -508
rect 14520 -548 15136 -542
rect 15206 -551 15212 -499
rect 15264 -502 15270 -499
rect 15264 -508 15822 -502
rect 15285 -542 15323 -508
rect 15357 -542 15395 -508
rect 15429 -542 15467 -508
rect 15501 -542 15676 -508
rect 15710 -542 15748 -508
rect 15782 -542 15822 -508
rect 15264 -548 15822 -542
rect 15264 -551 15270 -548
rect -137 -561 7 -555
rect -137 -595 -118 -561
rect -84 -595 -46 -561
rect -12 -595 7 -561
rect -137 -601 7 -595
rect 263 -561 407 -555
rect 263 -595 282 -561
rect 316 -595 354 -561
rect 388 -595 407 -561
rect 263 -601 407 -595
rect 663 -561 807 -555
rect 663 -595 682 -561
rect 716 -595 754 -561
rect 788 -595 807 -561
rect 663 -601 807 -595
rect 1063 -561 1207 -555
rect 1063 -595 1082 -561
rect 1116 -595 1154 -561
rect 1188 -595 1207 -561
rect 1063 -601 1207 -595
rect 1463 -561 1607 -555
rect 1463 -595 1482 -561
rect 1516 -595 1554 -561
rect 1588 -595 1607 -561
rect 1463 -601 1607 -595
rect 1863 -561 2007 -555
rect 1863 -595 1882 -561
rect 1916 -595 1954 -561
rect 1988 -595 2007 -561
rect 1863 -601 2007 -595
rect 2263 -561 2407 -555
rect 2263 -595 2282 -561
rect 2316 -595 2354 -561
rect 2388 -595 2407 -561
rect 2263 -601 2407 -595
rect 2663 -561 2807 -555
rect 2663 -595 2682 -561
rect 2716 -595 2754 -561
rect 2788 -595 2807 -561
rect 2663 -601 2807 -595
rect 3063 -561 3207 -555
rect 3063 -595 3082 -561
rect 3116 -595 3154 -561
rect 3188 -595 3207 -561
rect 3063 -601 3207 -595
rect 3463 -561 3607 -555
rect 3463 -595 3482 -561
rect 3516 -595 3554 -561
rect 3588 -595 3607 -561
rect 3463 -601 3607 -595
rect 3863 -561 4007 -555
rect 3863 -595 3882 -561
rect 3916 -595 3954 -561
rect 3988 -595 4007 -561
rect 3863 -601 4007 -595
rect 4263 -561 4407 -555
rect 4263 -595 4282 -561
rect 4316 -595 4354 -561
rect 4388 -595 4407 -561
rect 4263 -601 4407 -595
rect 4663 -561 4807 -555
rect 4663 -595 4682 -561
rect 4716 -595 4754 -561
rect 4788 -595 4807 -561
rect 4663 -601 4807 -595
rect 5063 -561 5207 -555
rect 5063 -595 5082 -561
rect 5116 -595 5154 -561
rect 5188 -595 5207 -561
rect 5063 -601 5207 -595
rect 5463 -561 5607 -555
rect 5463 -595 5482 -561
rect 5516 -595 5554 -561
rect 5588 -595 5607 -561
rect 5463 -601 5607 -595
rect 5863 -561 6007 -555
rect 5863 -595 5882 -561
rect 5916 -595 5954 -561
rect 5988 -595 6007 -561
rect 5863 -601 6007 -595
rect 6263 -561 6407 -555
rect 6263 -595 6282 -561
rect 6316 -595 6354 -561
rect 6388 -595 6407 -561
rect 6263 -601 6407 -595
rect 6663 -561 6807 -555
rect 6663 -595 6682 -561
rect 6716 -595 6754 -561
rect 6788 -595 6807 -561
rect 6663 -601 6807 -595
rect 7063 -561 7207 -555
rect 7063 -595 7082 -561
rect 7116 -595 7154 -561
rect 7188 -595 7207 -561
rect 7063 -601 7207 -595
rect 7463 -561 7607 -555
rect 7463 -595 7482 -561
rect 7516 -595 7554 -561
rect 7588 -595 7607 -561
rect 7463 -601 7607 -595
rect 7863 -561 8007 -555
rect 7863 -595 7882 -561
rect 7916 -595 7954 -561
rect 7988 -595 8007 -561
rect 7863 -601 8007 -595
rect 8263 -561 8407 -555
rect 8263 -595 8282 -561
rect 8316 -595 8354 -561
rect 8388 -595 8407 -561
rect 8263 -601 8407 -595
rect 8663 -561 8807 -555
rect 8663 -595 8682 -561
rect 8716 -595 8754 -561
rect 8788 -595 8807 -561
rect 8663 -601 8807 -595
rect 9063 -561 9207 -555
rect 9063 -595 9082 -561
rect 9116 -595 9154 -561
rect 9188 -595 9207 -561
rect 9063 -601 9207 -595
rect 9463 -561 9607 -555
rect 9463 -595 9482 -561
rect 9516 -595 9554 -561
rect 9588 -595 9607 -561
rect 9463 -601 9607 -595
rect 9863 -561 10007 -555
rect 9863 -595 9882 -561
rect 9916 -595 9954 -561
rect 9988 -595 10007 -561
rect 9863 -601 10007 -595
rect 10263 -561 10407 -555
rect 10263 -595 10282 -561
rect 10316 -595 10354 -561
rect 10388 -595 10407 -561
rect 10263 -601 10407 -595
rect 10663 -561 10807 -555
rect 10663 -595 10682 -561
rect 10716 -595 10754 -561
rect 10788 -595 10807 -561
rect 10663 -601 10807 -595
rect 11063 -561 11207 -555
rect 11063 -595 11082 -561
rect 11116 -595 11154 -561
rect 11188 -595 11207 -561
rect 11063 -601 11207 -595
rect 11463 -561 11607 -555
rect 11463 -595 11482 -561
rect 11516 -595 11554 -561
rect 11588 -595 11607 -561
rect 11463 -601 11607 -595
rect 11863 -561 12007 -555
rect 11863 -595 11882 -561
rect 11916 -595 11954 -561
rect 11988 -595 12007 -561
rect 11863 -601 12007 -595
rect 12263 -561 12407 -555
rect 12263 -595 12282 -561
rect 12316 -595 12354 -561
rect 12388 -595 12407 -561
rect 12263 -601 12407 -595
rect 12663 -561 12807 -555
rect 12663 -595 12682 -561
rect 12716 -595 12754 -561
rect 12788 -595 12807 -561
rect 12663 -601 12807 -595
rect 14526 -599 14697 -593
rect 14434 -610 14440 -599
rect 32 -630 90 -624
rect 32 -632 44 -630
rect -148 -662 44 -632
rect 32 -664 44 -662
rect 78 -632 90 -630
rect 180 -630 238 -624
rect 180 -632 192 -630
rect 78 -662 192 -632
rect 78 -664 90 -662
rect 32 -670 90 -664
rect 180 -664 192 -662
rect 226 -632 238 -630
rect 432 -630 490 -624
rect 432 -632 444 -630
rect 226 -662 444 -632
rect 226 -664 238 -662
rect 180 -670 238 -664
rect 432 -664 444 -662
rect 478 -632 490 -630
rect 580 -630 638 -624
rect 580 -632 592 -630
rect 478 -662 592 -632
rect 478 -664 490 -662
rect 432 -670 490 -664
rect 580 -664 592 -662
rect 626 -632 638 -630
rect 832 -630 890 -624
rect 832 -632 844 -630
rect 626 -662 844 -632
rect 626 -664 638 -662
rect 580 -670 638 -664
rect 832 -664 844 -662
rect 878 -632 890 -630
rect 980 -630 1038 -624
rect 980 -632 992 -630
rect 878 -662 992 -632
rect 878 -664 890 -662
rect 832 -670 890 -664
rect 980 -664 992 -662
rect 1026 -632 1038 -630
rect 1232 -630 1290 -624
rect 1232 -632 1244 -630
rect 1026 -662 1244 -632
rect 1026 -664 1038 -662
rect 980 -670 1038 -664
rect 1232 -664 1244 -662
rect 1278 -632 1290 -630
rect 1380 -630 1438 -624
rect 1380 -632 1392 -630
rect 1278 -662 1392 -632
rect 1278 -664 1290 -662
rect 1232 -670 1290 -664
rect 1380 -664 1392 -662
rect 1426 -632 1438 -630
rect 1632 -630 1690 -624
rect 1632 -632 1644 -630
rect 1426 -662 1644 -632
rect 1426 -664 1438 -662
rect 1380 -670 1438 -664
rect 1632 -664 1644 -662
rect 1678 -632 1690 -630
rect 1780 -630 1838 -624
rect 1780 -632 1792 -630
rect 1678 -662 1792 -632
rect 1678 -664 1690 -662
rect 1632 -670 1690 -664
rect 1780 -664 1792 -662
rect 1826 -632 1838 -630
rect 2032 -630 2090 -624
rect 2032 -632 2044 -630
rect 1826 -662 2044 -632
rect 1826 -664 1838 -662
rect 1780 -670 1838 -664
rect 2032 -664 2044 -662
rect 2078 -632 2090 -630
rect 2180 -630 2238 -624
rect 2180 -632 2192 -630
rect 2078 -662 2192 -632
rect 2078 -664 2090 -662
rect 2032 -670 2090 -664
rect 2180 -664 2192 -662
rect 2226 -632 2238 -630
rect 2432 -630 2490 -624
rect 2432 -632 2444 -630
rect 2226 -662 2444 -632
rect 2226 -664 2238 -662
rect 2180 -670 2238 -664
rect 2432 -664 2444 -662
rect 2478 -632 2490 -630
rect 2580 -630 2638 -624
rect 2580 -632 2592 -630
rect 2478 -662 2592 -632
rect 2478 -664 2490 -662
rect 2432 -670 2490 -664
rect 2580 -664 2592 -662
rect 2626 -632 2638 -630
rect 2832 -630 2890 -624
rect 2832 -632 2844 -630
rect 2626 -662 2844 -632
rect 2626 -664 2638 -662
rect 2580 -670 2638 -664
rect 2832 -664 2844 -662
rect 2878 -632 2890 -630
rect 2980 -630 3038 -624
rect 2980 -632 2992 -630
rect 2878 -662 2992 -632
rect 2878 -664 2890 -662
rect 2832 -670 2890 -664
rect 2980 -664 2992 -662
rect 3026 -632 3038 -630
rect 3232 -630 3290 -624
rect 3232 -632 3244 -630
rect 3026 -662 3244 -632
rect 3026 -664 3038 -662
rect 2980 -670 3038 -664
rect 3232 -664 3244 -662
rect 3278 -632 3290 -630
rect 3380 -630 3438 -624
rect 3380 -632 3392 -630
rect 3278 -662 3392 -632
rect 3278 -664 3290 -662
rect 3232 -670 3290 -664
rect 3380 -664 3392 -662
rect 3426 -632 3438 -630
rect 3632 -630 3690 -624
rect 3632 -632 3644 -630
rect 3426 -662 3644 -632
rect 3426 -664 3438 -662
rect 3380 -670 3438 -664
rect 3632 -664 3644 -662
rect 3678 -632 3690 -630
rect 3780 -630 3838 -624
rect 3780 -632 3792 -630
rect 3678 -662 3792 -632
rect 3678 -664 3690 -662
rect 3632 -670 3690 -664
rect 3780 -664 3792 -662
rect 3826 -632 3838 -630
rect 4032 -630 4090 -624
rect 4032 -632 4044 -630
rect 3826 -662 4044 -632
rect 3826 -664 3838 -662
rect 3780 -670 3838 -664
rect 4032 -664 4044 -662
rect 4078 -632 4090 -630
rect 4180 -630 4238 -624
rect 4180 -632 4192 -630
rect 4078 -662 4192 -632
rect 4078 -664 4090 -662
rect 4032 -670 4090 -664
rect 4180 -664 4192 -662
rect 4226 -632 4238 -630
rect 4432 -630 4490 -624
rect 4432 -632 4444 -630
rect 4226 -662 4444 -632
rect 4226 -664 4238 -662
rect 4180 -670 4238 -664
rect 4432 -664 4444 -662
rect 4478 -632 4490 -630
rect 4580 -630 4638 -624
rect 4580 -632 4592 -630
rect 4478 -662 4592 -632
rect 4478 -664 4490 -662
rect 4432 -670 4490 -664
rect 4580 -664 4592 -662
rect 4626 -632 4638 -630
rect 4832 -630 4890 -624
rect 4832 -632 4844 -630
rect 4626 -662 4844 -632
rect 4626 -664 4638 -662
rect 4580 -670 4638 -664
rect 4832 -664 4844 -662
rect 4878 -632 4890 -630
rect 4980 -630 5038 -624
rect 4980 -632 4992 -630
rect 4878 -662 4992 -632
rect 4878 -664 4890 -662
rect 4832 -670 4890 -664
rect 4980 -664 4992 -662
rect 5026 -632 5038 -630
rect 5232 -630 5290 -624
rect 5232 -632 5244 -630
rect 5026 -662 5244 -632
rect 5026 -664 5038 -662
rect 4980 -670 5038 -664
rect 5232 -664 5244 -662
rect 5278 -632 5290 -630
rect 5380 -630 5438 -624
rect 5380 -632 5392 -630
rect 5278 -662 5392 -632
rect 5278 -664 5290 -662
rect 5232 -670 5290 -664
rect 5380 -664 5392 -662
rect 5426 -632 5438 -630
rect 5632 -630 5690 -624
rect 5632 -632 5644 -630
rect 5426 -662 5644 -632
rect 5426 -664 5438 -662
rect 5380 -670 5438 -664
rect 5632 -664 5644 -662
rect 5678 -632 5690 -630
rect 5780 -630 5838 -624
rect 5780 -632 5792 -630
rect 5678 -662 5792 -632
rect 5678 -664 5690 -662
rect 5632 -670 5690 -664
rect 5780 -664 5792 -662
rect 5826 -632 5838 -630
rect 6032 -630 6090 -624
rect 6032 -632 6044 -630
rect 5826 -662 6044 -632
rect 5826 -664 5838 -662
rect 5780 -670 5838 -664
rect 6032 -664 6044 -662
rect 6078 -632 6090 -630
rect 6180 -630 6238 -624
rect 6180 -632 6192 -630
rect 6078 -662 6192 -632
rect 6078 -664 6090 -662
rect 6032 -670 6090 -664
rect 6180 -664 6192 -662
rect 6226 -632 6238 -630
rect 6432 -630 6490 -624
rect 6432 -632 6444 -630
rect 6226 -662 6444 -632
rect 6226 -664 6238 -662
rect 6180 -670 6238 -664
rect 6432 -664 6444 -662
rect 6478 -632 6490 -630
rect 6580 -630 6638 -624
rect 6580 -632 6592 -630
rect 6478 -662 6592 -632
rect 6478 -664 6490 -662
rect 6432 -670 6490 -664
rect 6580 -664 6592 -662
rect 6626 -632 6638 -630
rect 6832 -630 6890 -624
rect 6832 -632 6844 -630
rect 6626 -662 6844 -632
rect 6626 -664 6638 -662
rect 6580 -670 6638 -664
rect 6832 -664 6844 -662
rect 6878 -632 6890 -630
rect 6980 -630 7038 -624
rect 6980 -632 6992 -630
rect 6878 -662 6992 -632
rect 6878 -664 6890 -662
rect 6832 -670 6890 -664
rect 6980 -664 6992 -662
rect 7026 -632 7038 -630
rect 7232 -630 7290 -624
rect 7232 -632 7244 -630
rect 7026 -662 7244 -632
rect 7026 -664 7038 -662
rect 6980 -670 7038 -664
rect 7232 -664 7244 -662
rect 7278 -632 7290 -630
rect 7380 -630 7438 -624
rect 7380 -632 7392 -630
rect 7278 -662 7392 -632
rect 7278 -664 7290 -662
rect 7232 -670 7290 -664
rect 7380 -664 7392 -662
rect 7426 -632 7438 -630
rect 7632 -630 7690 -624
rect 7632 -632 7644 -630
rect 7426 -662 7644 -632
rect 7426 -664 7438 -662
rect 7380 -670 7438 -664
rect 7632 -664 7644 -662
rect 7678 -632 7690 -630
rect 7780 -630 7838 -624
rect 7780 -632 7792 -630
rect 7678 -662 7792 -632
rect 7678 -664 7690 -662
rect 7632 -670 7690 -664
rect 7780 -664 7792 -662
rect 7826 -632 7838 -630
rect 8032 -630 8090 -624
rect 8032 -632 8044 -630
rect 7826 -662 8044 -632
rect 7826 -664 7838 -662
rect 7780 -670 7838 -664
rect 8032 -664 8044 -662
rect 8078 -632 8090 -630
rect 8180 -630 8238 -624
rect 8180 -632 8192 -630
rect 8078 -662 8192 -632
rect 8078 -664 8090 -662
rect 8032 -670 8090 -664
rect 8180 -664 8192 -662
rect 8226 -632 8238 -630
rect 8432 -630 8490 -624
rect 8432 -632 8444 -630
rect 8226 -662 8444 -632
rect 8226 -664 8238 -662
rect 8180 -670 8238 -664
rect 8432 -664 8444 -662
rect 8478 -632 8490 -630
rect 8580 -630 8638 -624
rect 8580 -632 8592 -630
rect 8478 -662 8592 -632
rect 8478 -664 8490 -662
rect 8432 -670 8490 -664
rect 8580 -664 8592 -662
rect 8626 -632 8638 -630
rect 8832 -630 8890 -624
rect 8832 -632 8844 -630
rect 8626 -662 8844 -632
rect 8626 -664 8638 -662
rect 8580 -670 8638 -664
rect 8832 -664 8844 -662
rect 8878 -632 8890 -630
rect 8980 -630 9038 -624
rect 8980 -632 8992 -630
rect 8878 -662 8992 -632
rect 8878 -664 8890 -662
rect 8832 -670 8890 -664
rect 8980 -664 8992 -662
rect 9026 -632 9038 -630
rect 9232 -630 9290 -624
rect 9232 -632 9244 -630
rect 9026 -662 9244 -632
rect 9026 -664 9038 -662
rect 8980 -670 9038 -664
rect 9232 -664 9244 -662
rect 9278 -632 9290 -630
rect 9380 -630 9438 -624
rect 9380 -632 9392 -630
rect 9278 -662 9392 -632
rect 9278 -664 9290 -662
rect 9232 -670 9290 -664
rect 9380 -664 9392 -662
rect 9426 -632 9438 -630
rect 9632 -630 9690 -624
rect 9632 -632 9644 -630
rect 9426 -662 9644 -632
rect 9426 -664 9438 -662
rect 9380 -670 9438 -664
rect 9632 -664 9644 -662
rect 9678 -632 9690 -630
rect 9780 -630 9838 -624
rect 9780 -632 9792 -630
rect 9678 -662 9792 -632
rect 9678 -664 9690 -662
rect 9632 -670 9690 -664
rect 9780 -664 9792 -662
rect 9826 -632 9838 -630
rect 10032 -630 10090 -624
rect 10032 -632 10044 -630
rect 9826 -662 10044 -632
rect 9826 -664 9838 -662
rect 9780 -670 9838 -664
rect 10032 -664 10044 -662
rect 10078 -632 10090 -630
rect 10180 -630 10238 -624
rect 10180 -632 10192 -630
rect 10078 -662 10192 -632
rect 10078 -664 10090 -662
rect 10032 -670 10090 -664
rect 10180 -664 10192 -662
rect 10226 -632 10238 -630
rect 10432 -630 10490 -624
rect 10432 -632 10444 -630
rect 10226 -662 10444 -632
rect 10226 -664 10238 -662
rect 10180 -670 10238 -664
rect 10432 -664 10444 -662
rect 10478 -632 10490 -630
rect 10580 -630 10638 -624
rect 10580 -632 10592 -630
rect 10478 -662 10592 -632
rect 10478 -664 10490 -662
rect 10432 -670 10490 -664
rect 10580 -664 10592 -662
rect 10626 -632 10638 -630
rect 10832 -630 10890 -624
rect 10832 -632 10844 -630
rect 10626 -662 10844 -632
rect 10626 -664 10638 -662
rect 10580 -670 10638 -664
rect 10832 -664 10844 -662
rect 10878 -632 10890 -630
rect 10980 -630 11038 -624
rect 10980 -632 10992 -630
rect 10878 -662 10992 -632
rect 10878 -664 10890 -662
rect 10832 -670 10890 -664
rect 10980 -664 10992 -662
rect 11026 -632 11038 -630
rect 11232 -630 11290 -624
rect 11232 -632 11244 -630
rect 11026 -662 11244 -632
rect 11026 -664 11038 -662
rect 10980 -670 11038 -664
rect 11232 -664 11244 -662
rect 11278 -632 11290 -630
rect 11380 -630 11438 -624
rect 11380 -632 11392 -630
rect 11278 -662 11392 -632
rect 11278 -664 11290 -662
rect 11232 -670 11290 -664
rect 11380 -664 11392 -662
rect 11426 -632 11438 -630
rect 11632 -630 11690 -624
rect 11632 -632 11644 -630
rect 11426 -662 11644 -632
rect 11426 -664 11438 -662
rect 11380 -670 11438 -664
rect 11632 -664 11644 -662
rect 11678 -632 11690 -630
rect 11780 -630 11838 -624
rect 11780 -632 11792 -630
rect 11678 -662 11792 -632
rect 11678 -664 11690 -662
rect 11632 -670 11690 -664
rect 11780 -664 11792 -662
rect 11826 -632 11838 -630
rect 12032 -630 12090 -624
rect 12032 -632 12044 -630
rect 11826 -662 12044 -632
rect 11826 -664 11838 -662
rect 11780 -670 11838 -664
rect 12032 -664 12044 -662
rect 12078 -632 12090 -630
rect 12180 -630 12238 -624
rect 12180 -632 12192 -630
rect 12078 -662 12192 -632
rect 12078 -664 12090 -662
rect 12032 -670 12090 -664
rect 12180 -664 12192 -662
rect 12226 -632 12238 -630
rect 12432 -630 12490 -624
rect 12432 -632 12444 -630
rect 12226 -662 12444 -632
rect 12226 -664 12238 -662
rect 12180 -670 12238 -664
rect 12432 -664 12444 -662
rect 12478 -632 12490 -630
rect 12580 -630 12638 -624
rect 12580 -632 12592 -630
rect 12478 -662 12592 -632
rect 12478 -664 12490 -662
rect 12432 -670 12490 -664
rect 12580 -664 12592 -662
rect 12626 -632 12638 -630
rect 12626 -662 12818 -632
rect 14400 -640 14440 -610
rect 14434 -651 14440 -640
rect 14492 -651 14498 -599
rect 14526 -651 14553 -599
rect 14605 -651 14617 -599
rect 14669 -651 14697 -599
rect 14526 -657 14697 -651
rect 14725 -599 14777 -593
rect 14725 -657 14777 -651
rect 14805 -599 15136 -593
rect 14805 -651 14816 -599
rect 14868 -608 14880 -599
rect 14932 -608 14944 -599
rect 14996 -608 15008 -599
rect 15060 -608 15072 -599
rect 14876 -642 14880 -608
rect 14868 -651 14880 -642
rect 14932 -651 14944 -642
rect 14996 -651 15008 -642
rect 15060 -651 15072 -642
rect 15124 -651 15136 -599
rect 14805 -657 15136 -651
rect 15206 -599 15537 -593
rect 15206 -651 15217 -599
rect 15269 -608 15281 -599
rect 15333 -608 15345 -599
rect 15397 -608 15409 -599
rect 15461 -608 15473 -599
rect 15461 -642 15465 -608
rect 15269 -651 15281 -642
rect 15333 -651 15345 -642
rect 15397 -651 15409 -642
rect 15461 -651 15473 -642
rect 15525 -651 15537 -599
rect 15206 -657 15537 -651
rect 15565 -599 15617 -593
rect 15565 -657 15617 -651
rect 15645 -599 15816 -593
rect 15645 -651 15672 -599
rect 15724 -651 15736 -599
rect 15788 -651 15816 -599
rect 15645 -657 15816 -651
rect 12626 -664 12638 -662
rect 12580 -670 12638 -664
rect 14520 -708 15136 -702
rect 14520 -710 14560 -708
rect 14400 -740 14560 -710
rect 14520 -742 14560 -740
rect 14594 -742 14632 -708
rect 14666 -742 14841 -708
rect 14875 -742 14913 -708
rect 14947 -742 14985 -708
rect 15019 -742 15057 -708
rect 15091 -742 15136 -708
rect 14520 -748 15136 -742
rect 15206 -751 15212 -699
rect 15264 -702 15270 -699
rect 15264 -708 15822 -702
rect 15285 -742 15323 -708
rect 15357 -742 15395 -708
rect 15429 -742 15467 -708
rect 15501 -742 15676 -708
rect 15710 -742 15748 -708
rect 15782 -742 15822 -708
rect 15264 -748 15822 -742
rect 15264 -751 15270 -748
rect 14526 -799 14697 -793
rect 14434 -810 14440 -799
rect -18 -880 -9 -828
rect 43 -880 55 -828
rect 107 -880 116 -828
rect 154 -880 163 -828
rect 215 -880 227 -828
rect 279 -880 288 -828
rect 382 -880 391 -828
rect 443 -880 455 -828
rect 507 -880 516 -828
rect 554 -880 563 -828
rect 615 -880 627 -828
rect 679 -880 688 -828
rect 782 -880 791 -828
rect 843 -880 855 -828
rect 907 -880 916 -828
rect 954 -880 963 -828
rect 1015 -880 1027 -828
rect 1079 -880 1088 -828
rect 1182 -880 1191 -828
rect 1243 -880 1255 -828
rect 1307 -880 1316 -828
rect 1354 -880 1363 -828
rect 1415 -880 1427 -828
rect 1479 -880 1488 -828
rect 1582 -880 1591 -828
rect 1643 -880 1655 -828
rect 1707 -880 1716 -828
rect 1754 -880 1763 -828
rect 1815 -880 1827 -828
rect 1879 -880 1888 -828
rect 1982 -880 1991 -828
rect 2043 -880 2055 -828
rect 2107 -880 2116 -828
rect 2154 -880 2163 -828
rect 2215 -880 2227 -828
rect 2279 -880 2288 -828
rect 2382 -880 2391 -828
rect 2443 -880 2455 -828
rect 2507 -880 2516 -828
rect 2554 -880 2563 -828
rect 2615 -880 2627 -828
rect 2679 -880 2688 -828
rect 2782 -880 2791 -828
rect 2843 -880 2855 -828
rect 2907 -880 2916 -828
rect 2954 -880 2963 -828
rect 3015 -880 3027 -828
rect 3079 -880 3088 -828
rect 3182 -880 3191 -828
rect 3243 -880 3255 -828
rect 3307 -880 3316 -828
rect 3354 -880 3363 -828
rect 3415 -880 3427 -828
rect 3479 -880 3488 -828
rect 3582 -880 3591 -828
rect 3643 -880 3655 -828
rect 3707 -880 3716 -828
rect 3754 -880 3763 -828
rect 3815 -880 3827 -828
rect 3879 -880 3888 -828
rect 3982 -880 3991 -828
rect 4043 -880 4055 -828
rect 4107 -880 4116 -828
rect 4154 -880 4163 -828
rect 4215 -880 4227 -828
rect 4279 -880 4288 -828
rect 4382 -880 4391 -828
rect 4443 -880 4455 -828
rect 4507 -880 4516 -828
rect 4554 -880 4563 -828
rect 4615 -880 4627 -828
rect 4679 -880 4688 -828
rect 4782 -880 4791 -828
rect 4843 -880 4855 -828
rect 4907 -880 4916 -828
rect 4954 -880 4963 -828
rect 5015 -880 5027 -828
rect 5079 -880 5088 -828
rect 5182 -880 5191 -828
rect 5243 -880 5255 -828
rect 5307 -880 5316 -828
rect 5354 -880 5363 -828
rect 5415 -880 5427 -828
rect 5479 -880 5488 -828
rect 5582 -880 5591 -828
rect 5643 -880 5655 -828
rect 5707 -880 5716 -828
rect 5754 -880 5763 -828
rect 5815 -880 5827 -828
rect 5879 -880 5888 -828
rect 5982 -880 5991 -828
rect 6043 -880 6055 -828
rect 6107 -880 6116 -828
rect 6154 -880 6163 -828
rect 6215 -880 6227 -828
rect 6279 -880 6288 -828
rect 6382 -880 6391 -828
rect 6443 -880 6455 -828
rect 6507 -880 6516 -828
rect 6554 -880 6563 -828
rect 6615 -880 6627 -828
rect 6679 -880 6688 -828
rect 6782 -880 6791 -828
rect 6843 -880 6855 -828
rect 6907 -880 6916 -828
rect 6954 -880 6963 -828
rect 7015 -880 7027 -828
rect 7079 -880 7088 -828
rect 7182 -880 7191 -828
rect 7243 -880 7255 -828
rect 7307 -880 7316 -828
rect 7354 -880 7363 -828
rect 7415 -880 7427 -828
rect 7479 -880 7488 -828
rect 7582 -880 7591 -828
rect 7643 -880 7655 -828
rect 7707 -880 7716 -828
rect 7754 -880 7763 -828
rect 7815 -880 7827 -828
rect 7879 -880 7888 -828
rect 7982 -880 7991 -828
rect 8043 -880 8055 -828
rect 8107 -880 8116 -828
rect 8154 -880 8163 -828
rect 8215 -880 8227 -828
rect 8279 -880 8288 -828
rect 8382 -880 8391 -828
rect 8443 -880 8455 -828
rect 8507 -880 8516 -828
rect 8554 -880 8563 -828
rect 8615 -880 8627 -828
rect 8679 -880 8688 -828
rect 8782 -880 8791 -828
rect 8843 -880 8855 -828
rect 8907 -880 8916 -828
rect 8954 -880 8963 -828
rect 9015 -880 9027 -828
rect 9079 -880 9088 -828
rect 9182 -880 9191 -828
rect 9243 -880 9255 -828
rect 9307 -880 9316 -828
rect 9354 -880 9363 -828
rect 9415 -880 9427 -828
rect 9479 -880 9488 -828
rect 9582 -880 9591 -828
rect 9643 -880 9655 -828
rect 9707 -880 9716 -828
rect 9754 -880 9763 -828
rect 9815 -880 9827 -828
rect 9879 -880 9888 -828
rect 9982 -880 9991 -828
rect 10043 -880 10055 -828
rect 10107 -880 10116 -828
rect 10154 -880 10163 -828
rect 10215 -880 10227 -828
rect 10279 -880 10288 -828
rect 10382 -880 10391 -828
rect 10443 -880 10455 -828
rect 10507 -880 10516 -828
rect 10554 -880 10563 -828
rect 10615 -880 10627 -828
rect 10679 -880 10688 -828
rect 10782 -880 10791 -828
rect 10843 -880 10855 -828
rect 10907 -880 10916 -828
rect 10954 -880 10963 -828
rect 11015 -880 11027 -828
rect 11079 -880 11088 -828
rect 11182 -880 11191 -828
rect 11243 -880 11255 -828
rect 11307 -880 11316 -828
rect 11354 -880 11363 -828
rect 11415 -880 11427 -828
rect 11479 -880 11488 -828
rect 11582 -880 11591 -828
rect 11643 -880 11655 -828
rect 11707 -880 11716 -828
rect 11754 -880 11763 -828
rect 11815 -880 11827 -828
rect 11879 -880 11888 -828
rect 11982 -880 11991 -828
rect 12043 -880 12055 -828
rect 12107 -880 12116 -828
rect 12154 -880 12163 -828
rect 12215 -880 12227 -828
rect 12279 -880 12288 -828
rect 12382 -880 12391 -828
rect 12443 -880 12455 -828
rect 12507 -880 12516 -828
rect 12554 -880 12563 -828
rect 12615 -880 12627 -828
rect 12679 -880 12688 -828
rect 14400 -840 14440 -810
rect 14434 -851 14440 -840
rect 14492 -851 14498 -799
rect 14526 -851 14553 -799
rect 14605 -851 14617 -799
rect 14669 -851 14697 -799
rect 14526 -857 14697 -851
rect 14725 -799 14777 -793
rect 14725 -857 14777 -851
rect 14805 -799 15136 -793
rect 14805 -851 14816 -799
rect 14868 -808 14880 -799
rect 14932 -808 14944 -799
rect 14996 -808 15008 -799
rect 15060 -808 15072 -799
rect 14876 -842 14880 -808
rect 14868 -851 14880 -842
rect 14932 -851 14944 -842
rect 14996 -851 15008 -842
rect 15060 -851 15072 -842
rect 15124 -851 15136 -799
rect 14805 -857 15136 -851
rect 15206 -799 15537 -793
rect 15206 -851 15217 -799
rect 15269 -808 15281 -799
rect 15333 -808 15345 -799
rect 15397 -808 15409 -799
rect 15461 -808 15473 -799
rect 15461 -842 15465 -808
rect 15269 -851 15281 -842
rect 15333 -851 15345 -842
rect 15397 -851 15409 -842
rect 15461 -851 15473 -842
rect 15525 -851 15537 -799
rect 15206 -857 15537 -851
rect 15565 -799 15617 -793
rect 15565 -857 15617 -851
rect 15645 -799 15816 -793
rect 15645 -851 15672 -799
rect 15724 -851 15736 -799
rect 15788 -851 15816 -799
rect 15645 -857 15816 -851
rect -94 -908 -36 -902
rect -94 -910 -82 -908
rect -106 -940 -82 -910
rect -94 -942 -82 -940
rect -48 -910 -36 -908
rect 706 -908 764 -902
rect 706 -910 718 -908
rect -48 -940 718 -910
rect -48 -942 -36 -940
rect -94 -948 -36 -942
rect 706 -942 718 -940
rect 752 -910 764 -908
rect 1506 -908 1564 -902
rect 1506 -910 1518 -908
rect 752 -940 1518 -910
rect 752 -942 764 -940
rect 706 -948 764 -942
rect 1506 -942 1518 -940
rect 1552 -910 1564 -908
rect 2306 -908 2364 -902
rect 2306 -910 2318 -908
rect 1552 -940 2318 -910
rect 1552 -942 1564 -940
rect 1506 -948 1564 -942
rect 2306 -942 2318 -940
rect 2352 -910 2364 -908
rect 3106 -908 3164 -902
rect 3106 -910 3118 -908
rect 2352 -940 3118 -910
rect 2352 -942 2364 -940
rect 2306 -948 2364 -942
rect 3106 -942 3118 -940
rect 3152 -910 3164 -908
rect 3906 -908 3964 -902
rect 3906 -910 3918 -908
rect 3152 -940 3918 -910
rect 3152 -942 3164 -940
rect 3106 -948 3164 -942
rect 3906 -942 3918 -940
rect 3952 -910 3964 -908
rect 4706 -908 4764 -902
rect 4706 -910 4718 -908
rect 3952 -940 4718 -910
rect 3952 -942 3964 -940
rect 3906 -948 3964 -942
rect 4706 -942 4718 -940
rect 4752 -910 4764 -908
rect 5506 -908 5564 -902
rect 5506 -910 5518 -908
rect 4752 -940 5518 -910
rect 4752 -942 4764 -940
rect 4706 -948 4764 -942
rect 5506 -942 5518 -940
rect 5552 -910 5564 -908
rect 6306 -908 6364 -902
rect 6306 -910 6318 -908
rect 5552 -940 6318 -910
rect 5552 -942 5564 -940
rect 5506 -948 5564 -942
rect 6306 -942 6318 -940
rect 6352 -910 6364 -908
rect 7106 -908 7164 -902
rect 7106 -910 7118 -908
rect 6352 -940 7118 -910
rect 6352 -942 6364 -940
rect 6306 -948 6364 -942
rect 7106 -942 7118 -940
rect 7152 -910 7164 -908
rect 7906 -908 7964 -902
rect 7906 -910 7918 -908
rect 7152 -940 7918 -910
rect 7152 -942 7164 -940
rect 7106 -948 7164 -942
rect 7906 -942 7918 -940
rect 7952 -910 7964 -908
rect 8706 -908 8764 -902
rect 8706 -910 8718 -908
rect 7952 -940 8718 -910
rect 7952 -942 7964 -940
rect 7906 -948 7964 -942
rect 8706 -942 8718 -940
rect 8752 -910 8764 -908
rect 9506 -908 9564 -902
rect 9506 -910 9518 -908
rect 8752 -940 9518 -910
rect 8752 -942 8764 -940
rect 8706 -948 8764 -942
rect 9506 -942 9518 -940
rect 9552 -910 9564 -908
rect 10306 -908 10364 -902
rect 10306 -910 10318 -908
rect 9552 -940 10318 -910
rect 9552 -942 9564 -940
rect 9506 -948 9564 -942
rect 10306 -942 10318 -940
rect 10352 -910 10364 -908
rect 11106 -908 11164 -902
rect 11106 -910 11118 -908
rect 10352 -940 11118 -910
rect 10352 -942 10364 -940
rect 10306 -948 10364 -942
rect 11106 -942 11118 -940
rect 11152 -910 11164 -908
rect 11906 -908 11964 -902
rect 11906 -910 11918 -908
rect 11152 -940 11918 -910
rect 11152 -942 11164 -940
rect 11106 -948 11164 -942
rect 11906 -942 11918 -940
rect 11952 -910 11964 -908
rect 12706 -908 12764 -902
rect 12706 -910 12718 -908
rect 11952 -940 12718 -910
rect 11952 -942 11964 -940
rect 11906 -948 11964 -942
rect 12706 -942 12718 -940
rect 12752 -910 12764 -908
rect 14520 -908 15136 -902
rect 14520 -910 14560 -908
rect 12752 -940 12776 -910
rect 14400 -940 14560 -910
rect 12752 -942 12764 -940
rect 12706 -948 12764 -942
rect 14520 -942 14560 -940
rect 14594 -942 14632 -908
rect 14666 -942 14841 -908
rect 14875 -942 14913 -908
rect 14947 -942 14985 -908
rect 15019 -942 15057 -908
rect 15091 -942 15136 -908
rect 14520 -948 15136 -942
rect 15206 -951 15212 -899
rect 15264 -902 15270 -899
rect 15264 -908 15822 -902
rect 15285 -942 15323 -908
rect 15357 -942 15395 -908
rect 15429 -942 15467 -908
rect 15501 -942 15676 -908
rect 15710 -942 15748 -908
rect 15782 -942 15822 -908
rect 15264 -948 15822 -942
rect 15264 -951 15270 -948
rect 14526 -999 14697 -993
rect -94 -1008 -36 -1002
rect -94 -1010 -82 -1008
rect -106 -1040 -82 -1010
rect -94 -1042 -82 -1040
rect -48 -1010 -36 -1008
rect 706 -1008 764 -1002
rect 706 -1010 718 -1008
rect -48 -1040 718 -1010
rect -48 -1042 -36 -1040
rect -94 -1048 -36 -1042
rect 706 -1042 718 -1040
rect 752 -1010 764 -1008
rect 1506 -1008 1564 -1002
rect 1506 -1010 1518 -1008
rect 752 -1040 1518 -1010
rect 752 -1042 764 -1040
rect 706 -1048 764 -1042
rect 1506 -1042 1518 -1040
rect 1552 -1010 1564 -1008
rect 2306 -1008 2364 -1002
rect 2306 -1010 2318 -1008
rect 1552 -1040 2318 -1010
rect 1552 -1042 1564 -1040
rect 1506 -1048 1564 -1042
rect 2306 -1042 2318 -1040
rect 2352 -1010 2364 -1008
rect 3106 -1008 3164 -1002
rect 3106 -1010 3118 -1008
rect 2352 -1040 3118 -1010
rect 2352 -1042 2364 -1040
rect 2306 -1048 2364 -1042
rect 3106 -1042 3118 -1040
rect 3152 -1010 3164 -1008
rect 3906 -1008 3964 -1002
rect 3906 -1010 3918 -1008
rect 3152 -1040 3918 -1010
rect 3152 -1042 3164 -1040
rect 3106 -1048 3164 -1042
rect 3906 -1042 3918 -1040
rect 3952 -1010 3964 -1008
rect 4706 -1008 4764 -1002
rect 4706 -1010 4718 -1008
rect 3952 -1040 4718 -1010
rect 3952 -1042 3964 -1040
rect 3906 -1048 3964 -1042
rect 4706 -1042 4718 -1040
rect 4752 -1010 4764 -1008
rect 5506 -1008 5564 -1002
rect 5506 -1010 5518 -1008
rect 4752 -1040 5518 -1010
rect 4752 -1042 4764 -1040
rect 4706 -1048 4764 -1042
rect 5506 -1042 5518 -1040
rect 5552 -1010 5564 -1008
rect 6306 -1008 6364 -1002
rect 6306 -1010 6318 -1008
rect 5552 -1040 6318 -1010
rect 5552 -1042 5564 -1040
rect 5506 -1048 5564 -1042
rect 6306 -1042 6318 -1040
rect 6352 -1010 6364 -1008
rect 7106 -1008 7164 -1002
rect 7106 -1010 7118 -1008
rect 6352 -1040 7118 -1010
rect 6352 -1042 6364 -1040
rect 6306 -1048 6364 -1042
rect 7106 -1042 7118 -1040
rect 7152 -1010 7164 -1008
rect 7906 -1008 7964 -1002
rect 7906 -1010 7918 -1008
rect 7152 -1040 7918 -1010
rect 7152 -1042 7164 -1040
rect 7106 -1048 7164 -1042
rect 7906 -1042 7918 -1040
rect 7952 -1010 7964 -1008
rect 8706 -1008 8764 -1002
rect 8706 -1010 8718 -1008
rect 7952 -1040 8718 -1010
rect 7952 -1042 7964 -1040
rect 7906 -1048 7964 -1042
rect 8706 -1042 8718 -1040
rect 8752 -1010 8764 -1008
rect 9506 -1008 9564 -1002
rect 9506 -1010 9518 -1008
rect 8752 -1040 9518 -1010
rect 8752 -1042 8764 -1040
rect 8706 -1048 8764 -1042
rect 9506 -1042 9518 -1040
rect 9552 -1010 9564 -1008
rect 10306 -1008 10364 -1002
rect 10306 -1010 10318 -1008
rect 9552 -1040 10318 -1010
rect 9552 -1042 9564 -1040
rect 9506 -1048 9564 -1042
rect 10306 -1042 10318 -1040
rect 10352 -1010 10364 -1008
rect 11106 -1008 11164 -1002
rect 11106 -1010 11118 -1008
rect 10352 -1040 11118 -1010
rect 10352 -1042 10364 -1040
rect 10306 -1048 10364 -1042
rect 11106 -1042 11118 -1040
rect 11152 -1010 11164 -1008
rect 11906 -1008 11964 -1002
rect 11906 -1010 11918 -1008
rect 11152 -1040 11918 -1010
rect 11152 -1042 11164 -1040
rect 11106 -1048 11164 -1042
rect 11906 -1042 11918 -1040
rect 11952 -1010 11964 -1008
rect 12706 -1008 12764 -1002
rect 12706 -1010 12718 -1008
rect 11952 -1040 12718 -1010
rect 11952 -1042 11964 -1040
rect 11906 -1048 11964 -1042
rect 12706 -1042 12718 -1040
rect 12752 -1010 12764 -1008
rect 14434 -1010 14440 -999
rect 12752 -1040 12776 -1010
rect 14400 -1040 14440 -1010
rect 12752 -1042 12764 -1040
rect 12706 -1048 12764 -1042
rect 14434 -1051 14440 -1040
rect 14492 -1051 14498 -999
rect 14526 -1051 14553 -999
rect 14605 -1051 14617 -999
rect 14669 -1051 14697 -999
rect 14526 -1057 14697 -1051
rect 14725 -999 14777 -993
rect 14725 -1057 14777 -1051
rect 14805 -999 15136 -993
rect 14805 -1051 14816 -999
rect 14868 -1008 14880 -999
rect 14932 -1008 14944 -999
rect 14996 -1008 15008 -999
rect 15060 -1008 15072 -999
rect 14876 -1042 14880 -1008
rect 14868 -1051 14880 -1042
rect 14932 -1051 14944 -1042
rect 14996 -1051 15008 -1042
rect 15060 -1051 15072 -1042
rect 15124 -1051 15136 -999
rect 14805 -1057 15136 -1051
rect 15206 -999 15537 -993
rect 15206 -1051 15217 -999
rect 15269 -1008 15281 -999
rect 15333 -1008 15345 -999
rect 15397 -1008 15409 -999
rect 15461 -1008 15473 -999
rect 15461 -1042 15465 -1008
rect 15269 -1051 15281 -1042
rect 15333 -1051 15345 -1042
rect 15397 -1051 15409 -1042
rect 15461 -1051 15473 -1042
rect 15525 -1051 15537 -999
rect 15206 -1057 15537 -1051
rect 15565 -999 15617 -993
rect 15565 -1057 15617 -1051
rect 15645 -999 15816 -993
rect 15645 -1051 15672 -999
rect 15724 -1051 15736 -999
rect 15788 -1051 15816 -999
rect 15645 -1057 15816 -1051
rect -94 -1108 -36 -1102
rect -94 -1110 -82 -1108
rect -106 -1140 -82 -1110
rect -94 -1142 -82 -1140
rect -48 -1110 -36 -1108
rect 706 -1108 764 -1102
rect 706 -1110 718 -1108
rect -48 -1140 718 -1110
rect -48 -1142 -36 -1140
rect -94 -1148 -36 -1142
rect 706 -1142 718 -1140
rect 752 -1110 764 -1108
rect 1506 -1108 1564 -1102
rect 1506 -1110 1518 -1108
rect 752 -1140 1518 -1110
rect 752 -1142 764 -1140
rect 706 -1148 764 -1142
rect 1506 -1142 1518 -1140
rect 1552 -1110 1564 -1108
rect 2306 -1108 2364 -1102
rect 2306 -1110 2318 -1108
rect 1552 -1140 2318 -1110
rect 1552 -1142 1564 -1140
rect 1506 -1148 1564 -1142
rect 2306 -1142 2318 -1140
rect 2352 -1110 2364 -1108
rect 3106 -1108 3164 -1102
rect 3106 -1110 3118 -1108
rect 2352 -1140 3118 -1110
rect 2352 -1142 2364 -1140
rect 2306 -1148 2364 -1142
rect 3106 -1142 3118 -1140
rect 3152 -1110 3164 -1108
rect 3906 -1108 3964 -1102
rect 3906 -1110 3918 -1108
rect 3152 -1140 3918 -1110
rect 3152 -1142 3164 -1140
rect 3106 -1148 3164 -1142
rect 3906 -1142 3918 -1140
rect 3952 -1110 3964 -1108
rect 4706 -1108 4764 -1102
rect 4706 -1110 4718 -1108
rect 3952 -1140 4718 -1110
rect 3952 -1142 3964 -1140
rect 3906 -1148 3964 -1142
rect 4706 -1142 4718 -1140
rect 4752 -1110 4764 -1108
rect 5506 -1108 5564 -1102
rect 5506 -1110 5518 -1108
rect 4752 -1140 5518 -1110
rect 4752 -1142 4764 -1140
rect 4706 -1148 4764 -1142
rect 5506 -1142 5518 -1140
rect 5552 -1110 5564 -1108
rect 6306 -1108 6364 -1102
rect 6306 -1110 6318 -1108
rect 5552 -1140 6318 -1110
rect 5552 -1142 5564 -1140
rect 5506 -1148 5564 -1142
rect 6306 -1142 6318 -1140
rect 6352 -1110 6364 -1108
rect 7106 -1108 7164 -1102
rect 7106 -1110 7118 -1108
rect 6352 -1140 7118 -1110
rect 6352 -1142 6364 -1140
rect 6306 -1148 6364 -1142
rect 7106 -1142 7118 -1140
rect 7152 -1110 7164 -1108
rect 7906 -1108 7964 -1102
rect 7906 -1110 7918 -1108
rect 7152 -1140 7918 -1110
rect 7152 -1142 7164 -1140
rect 7106 -1148 7164 -1142
rect 7906 -1142 7918 -1140
rect 7952 -1110 7964 -1108
rect 8706 -1108 8764 -1102
rect 8706 -1110 8718 -1108
rect 7952 -1140 8718 -1110
rect 7952 -1142 7964 -1140
rect 7906 -1148 7964 -1142
rect 8706 -1142 8718 -1140
rect 8752 -1110 8764 -1108
rect 9506 -1108 9564 -1102
rect 9506 -1110 9518 -1108
rect 8752 -1140 9518 -1110
rect 8752 -1142 8764 -1140
rect 8706 -1148 8764 -1142
rect 9506 -1142 9518 -1140
rect 9552 -1110 9564 -1108
rect 10306 -1108 10364 -1102
rect 10306 -1110 10318 -1108
rect 9552 -1140 10318 -1110
rect 9552 -1142 9564 -1140
rect 9506 -1148 9564 -1142
rect 10306 -1142 10318 -1140
rect 10352 -1110 10364 -1108
rect 11106 -1108 11164 -1102
rect 11106 -1110 11118 -1108
rect 10352 -1140 11118 -1110
rect 10352 -1142 10364 -1140
rect 10306 -1148 10364 -1142
rect 11106 -1142 11118 -1140
rect 11152 -1110 11164 -1108
rect 11906 -1108 11964 -1102
rect 11906 -1110 11918 -1108
rect 11152 -1140 11918 -1110
rect 11152 -1142 11164 -1140
rect 11106 -1148 11164 -1142
rect 11906 -1142 11918 -1140
rect 11952 -1110 11964 -1108
rect 12706 -1108 12764 -1102
rect 12706 -1110 12718 -1108
rect 11952 -1140 12718 -1110
rect 11952 -1142 11964 -1140
rect 11906 -1148 11964 -1142
rect 12706 -1142 12718 -1140
rect 12752 -1110 12764 -1108
rect 14520 -1108 15136 -1102
rect 14520 -1110 14560 -1108
rect 12752 -1140 12776 -1110
rect 14400 -1140 14560 -1110
rect 12752 -1142 12764 -1140
rect 12706 -1148 12764 -1142
rect 14520 -1142 14560 -1140
rect 14594 -1142 14632 -1108
rect 14666 -1142 14841 -1108
rect 14875 -1142 14913 -1108
rect 14947 -1142 14985 -1108
rect 15019 -1142 15057 -1108
rect 15091 -1142 15136 -1108
rect 14520 -1148 15136 -1142
rect 15206 -1151 15212 -1099
rect 15264 -1102 15270 -1099
rect 15264 -1108 15822 -1102
rect 15285 -1142 15323 -1108
rect 15357 -1142 15395 -1108
rect 15429 -1142 15467 -1108
rect 15501 -1142 15676 -1108
rect 15710 -1142 15748 -1108
rect 15782 -1142 15822 -1108
rect 15264 -1148 15822 -1142
rect 15264 -1151 15270 -1148
rect 14526 -1199 14697 -1193
rect -94 -1208 -36 -1202
rect -94 -1210 -82 -1208
rect -106 -1240 -82 -1210
rect -94 -1242 -82 -1240
rect -48 -1210 -36 -1208
rect 706 -1208 764 -1202
rect 706 -1210 718 -1208
rect -48 -1240 718 -1210
rect -48 -1242 -36 -1240
rect -94 -1248 -36 -1242
rect 706 -1242 718 -1240
rect 752 -1210 764 -1208
rect 1506 -1208 1564 -1202
rect 1506 -1210 1518 -1208
rect 752 -1240 1518 -1210
rect 752 -1242 764 -1240
rect 706 -1248 764 -1242
rect 1506 -1242 1518 -1240
rect 1552 -1210 1564 -1208
rect 2306 -1208 2364 -1202
rect 2306 -1210 2318 -1208
rect 1552 -1240 2318 -1210
rect 1552 -1242 1564 -1240
rect 1506 -1248 1564 -1242
rect 2306 -1242 2318 -1240
rect 2352 -1210 2364 -1208
rect 3106 -1208 3164 -1202
rect 3106 -1210 3118 -1208
rect 2352 -1240 3118 -1210
rect 2352 -1242 2364 -1240
rect 2306 -1248 2364 -1242
rect 3106 -1242 3118 -1240
rect 3152 -1210 3164 -1208
rect 3906 -1208 3964 -1202
rect 3906 -1210 3918 -1208
rect 3152 -1240 3918 -1210
rect 3152 -1242 3164 -1240
rect 3106 -1248 3164 -1242
rect 3906 -1242 3918 -1240
rect 3952 -1210 3964 -1208
rect 4706 -1208 4764 -1202
rect 4706 -1210 4718 -1208
rect 3952 -1240 4718 -1210
rect 3952 -1242 3964 -1240
rect 3906 -1248 3964 -1242
rect 4706 -1242 4718 -1240
rect 4752 -1210 4764 -1208
rect 5506 -1208 5564 -1202
rect 5506 -1210 5518 -1208
rect 4752 -1240 5518 -1210
rect 4752 -1242 4764 -1240
rect 4706 -1248 4764 -1242
rect 5506 -1242 5518 -1240
rect 5552 -1210 5564 -1208
rect 6306 -1208 6364 -1202
rect 6306 -1210 6318 -1208
rect 5552 -1240 6318 -1210
rect 5552 -1242 5564 -1240
rect 5506 -1248 5564 -1242
rect 6306 -1242 6318 -1240
rect 6352 -1210 6364 -1208
rect 7106 -1208 7164 -1202
rect 7106 -1210 7118 -1208
rect 6352 -1240 7118 -1210
rect 6352 -1242 6364 -1240
rect 6306 -1248 6364 -1242
rect 7106 -1242 7118 -1240
rect 7152 -1210 7164 -1208
rect 7906 -1208 7964 -1202
rect 7906 -1210 7918 -1208
rect 7152 -1240 7918 -1210
rect 7152 -1242 7164 -1240
rect 7106 -1248 7164 -1242
rect 7906 -1242 7918 -1240
rect 7952 -1210 7964 -1208
rect 8706 -1208 8764 -1202
rect 8706 -1210 8718 -1208
rect 7952 -1240 8718 -1210
rect 7952 -1242 7964 -1240
rect 7906 -1248 7964 -1242
rect 8706 -1242 8718 -1240
rect 8752 -1210 8764 -1208
rect 9506 -1208 9564 -1202
rect 9506 -1210 9518 -1208
rect 8752 -1240 9518 -1210
rect 8752 -1242 8764 -1240
rect 8706 -1248 8764 -1242
rect 9506 -1242 9518 -1240
rect 9552 -1210 9564 -1208
rect 10306 -1208 10364 -1202
rect 10306 -1210 10318 -1208
rect 9552 -1240 10318 -1210
rect 9552 -1242 9564 -1240
rect 9506 -1248 9564 -1242
rect 10306 -1242 10318 -1240
rect 10352 -1210 10364 -1208
rect 11106 -1208 11164 -1202
rect 11106 -1210 11118 -1208
rect 10352 -1240 11118 -1210
rect 10352 -1242 10364 -1240
rect 10306 -1248 10364 -1242
rect 11106 -1242 11118 -1240
rect 11152 -1210 11164 -1208
rect 11906 -1208 11964 -1202
rect 11906 -1210 11918 -1208
rect 11152 -1240 11918 -1210
rect 11152 -1242 11164 -1240
rect 11106 -1248 11164 -1242
rect 11906 -1242 11918 -1240
rect 11952 -1210 11964 -1208
rect 12706 -1208 12764 -1202
rect 12706 -1210 12718 -1208
rect 11952 -1240 12718 -1210
rect 11952 -1242 11964 -1240
rect 11906 -1248 11964 -1242
rect 12706 -1242 12718 -1240
rect 12752 -1210 12764 -1208
rect 14434 -1210 14440 -1199
rect 12752 -1240 12776 -1210
rect 14400 -1240 14440 -1210
rect 12752 -1242 12764 -1240
rect 12706 -1248 12764 -1242
rect 14434 -1251 14440 -1240
rect 14492 -1251 14498 -1199
rect 14526 -1251 14553 -1199
rect 14605 -1251 14617 -1199
rect 14669 -1251 14697 -1199
rect 14526 -1257 14697 -1251
rect 14725 -1199 14777 -1193
rect 14725 -1257 14777 -1251
rect 14805 -1199 15136 -1193
rect 14805 -1251 14816 -1199
rect 14868 -1208 14880 -1199
rect 14932 -1208 14944 -1199
rect 14996 -1208 15008 -1199
rect 15060 -1208 15072 -1199
rect 14876 -1242 14880 -1208
rect 14868 -1251 14880 -1242
rect 14932 -1251 14944 -1242
rect 14996 -1251 15008 -1242
rect 15060 -1251 15072 -1242
rect 15124 -1251 15136 -1199
rect 14805 -1257 15136 -1251
rect 15206 -1199 15537 -1193
rect 15206 -1251 15217 -1199
rect 15269 -1208 15281 -1199
rect 15333 -1208 15345 -1199
rect 15397 -1208 15409 -1199
rect 15461 -1208 15473 -1199
rect 15461 -1242 15465 -1208
rect 15269 -1251 15281 -1242
rect 15333 -1251 15345 -1242
rect 15397 -1251 15409 -1242
rect 15461 -1251 15473 -1242
rect 15525 -1251 15537 -1199
rect 15206 -1257 15537 -1251
rect 15565 -1199 15617 -1193
rect 15565 -1257 15617 -1251
rect 15645 -1199 15816 -1193
rect 15645 -1251 15672 -1199
rect 15724 -1251 15736 -1199
rect 15788 -1251 15816 -1199
rect 15645 -1257 15816 -1251
rect -94 -1308 -36 -1302
rect -94 -1310 -82 -1308
rect -106 -1340 -82 -1310
rect -94 -1342 -82 -1340
rect -48 -1310 -36 -1308
rect 706 -1308 764 -1302
rect 706 -1310 718 -1308
rect -48 -1340 718 -1310
rect -48 -1342 -36 -1340
rect -94 -1348 -36 -1342
rect 706 -1342 718 -1340
rect 752 -1310 764 -1308
rect 1506 -1308 1564 -1302
rect 1506 -1310 1518 -1308
rect 752 -1340 1518 -1310
rect 752 -1342 764 -1340
rect 706 -1348 764 -1342
rect 1506 -1342 1518 -1340
rect 1552 -1310 1564 -1308
rect 2306 -1308 2364 -1302
rect 2306 -1310 2318 -1308
rect 1552 -1340 2318 -1310
rect 1552 -1342 1564 -1340
rect 1506 -1348 1564 -1342
rect 2306 -1342 2318 -1340
rect 2352 -1310 2364 -1308
rect 3106 -1308 3164 -1302
rect 3106 -1310 3118 -1308
rect 2352 -1340 3118 -1310
rect 2352 -1342 2364 -1340
rect 2306 -1348 2364 -1342
rect 3106 -1342 3118 -1340
rect 3152 -1310 3164 -1308
rect 3906 -1308 3964 -1302
rect 3906 -1310 3918 -1308
rect 3152 -1340 3918 -1310
rect 3152 -1342 3164 -1340
rect 3106 -1348 3164 -1342
rect 3906 -1342 3918 -1340
rect 3952 -1310 3964 -1308
rect 4706 -1308 4764 -1302
rect 4706 -1310 4718 -1308
rect 3952 -1340 4718 -1310
rect 3952 -1342 3964 -1340
rect 3906 -1348 3964 -1342
rect 4706 -1342 4718 -1340
rect 4752 -1310 4764 -1308
rect 5506 -1308 5564 -1302
rect 5506 -1310 5518 -1308
rect 4752 -1340 5518 -1310
rect 4752 -1342 4764 -1340
rect 4706 -1348 4764 -1342
rect 5506 -1342 5518 -1340
rect 5552 -1310 5564 -1308
rect 6306 -1308 6364 -1302
rect 6306 -1310 6318 -1308
rect 5552 -1340 6318 -1310
rect 5552 -1342 5564 -1340
rect 5506 -1348 5564 -1342
rect 6306 -1342 6318 -1340
rect 6352 -1310 6364 -1308
rect 7106 -1308 7164 -1302
rect 7106 -1310 7118 -1308
rect 6352 -1340 7118 -1310
rect 6352 -1342 6364 -1340
rect 6306 -1348 6364 -1342
rect 7106 -1342 7118 -1340
rect 7152 -1310 7164 -1308
rect 7906 -1308 7964 -1302
rect 7906 -1310 7918 -1308
rect 7152 -1340 7918 -1310
rect 7152 -1342 7164 -1340
rect 7106 -1348 7164 -1342
rect 7906 -1342 7918 -1340
rect 7952 -1310 7964 -1308
rect 8706 -1308 8764 -1302
rect 8706 -1310 8718 -1308
rect 7952 -1340 8718 -1310
rect 7952 -1342 7964 -1340
rect 7906 -1348 7964 -1342
rect 8706 -1342 8718 -1340
rect 8752 -1310 8764 -1308
rect 9506 -1308 9564 -1302
rect 9506 -1310 9518 -1308
rect 8752 -1340 9518 -1310
rect 8752 -1342 8764 -1340
rect 8706 -1348 8764 -1342
rect 9506 -1342 9518 -1340
rect 9552 -1310 9564 -1308
rect 10306 -1308 10364 -1302
rect 10306 -1310 10318 -1308
rect 9552 -1340 10318 -1310
rect 9552 -1342 9564 -1340
rect 9506 -1348 9564 -1342
rect 10306 -1342 10318 -1340
rect 10352 -1310 10364 -1308
rect 11106 -1308 11164 -1302
rect 11106 -1310 11118 -1308
rect 10352 -1340 11118 -1310
rect 10352 -1342 10364 -1340
rect 10306 -1348 10364 -1342
rect 11106 -1342 11118 -1340
rect 11152 -1310 11164 -1308
rect 11906 -1308 11964 -1302
rect 11906 -1310 11918 -1308
rect 11152 -1340 11918 -1310
rect 11152 -1342 11164 -1340
rect 11106 -1348 11164 -1342
rect 11906 -1342 11918 -1340
rect 11952 -1310 11964 -1308
rect 12706 -1308 12764 -1302
rect 12706 -1310 12718 -1308
rect 11952 -1340 12718 -1310
rect 11952 -1342 11964 -1340
rect 11906 -1348 11964 -1342
rect 12706 -1342 12718 -1340
rect 12752 -1310 12764 -1308
rect 14520 -1308 15136 -1302
rect 14520 -1310 14560 -1308
rect 12752 -1340 12776 -1310
rect 14400 -1340 14560 -1310
rect 12752 -1342 12764 -1340
rect 12706 -1348 12764 -1342
rect 14520 -1342 14560 -1340
rect 14594 -1342 14632 -1308
rect 14666 -1342 14841 -1308
rect 14875 -1342 14913 -1308
rect 14947 -1342 14985 -1308
rect 15019 -1342 15057 -1308
rect 15091 -1342 15136 -1308
rect 14520 -1348 15136 -1342
rect 15206 -1351 15212 -1299
rect 15264 -1302 15270 -1299
rect 15264 -1308 15822 -1302
rect 15285 -1342 15323 -1308
rect 15357 -1342 15395 -1308
rect 15429 -1342 15467 -1308
rect 15501 -1342 15676 -1308
rect 15710 -1342 15748 -1308
rect 15782 -1342 15822 -1308
rect 15264 -1348 15822 -1342
rect 15264 -1351 15270 -1348
rect 14526 -1399 14697 -1393
rect -94 -1408 -36 -1402
rect -94 -1410 -82 -1408
rect -106 -1440 -82 -1410
rect -94 -1442 -82 -1440
rect -48 -1410 -36 -1408
rect 706 -1408 764 -1402
rect 706 -1410 718 -1408
rect -48 -1440 718 -1410
rect -48 -1442 -36 -1440
rect -94 -1448 -36 -1442
rect 706 -1442 718 -1440
rect 752 -1410 764 -1408
rect 1506 -1408 1564 -1402
rect 1506 -1410 1518 -1408
rect 752 -1440 1518 -1410
rect 752 -1442 764 -1440
rect 706 -1448 764 -1442
rect 1506 -1442 1518 -1440
rect 1552 -1410 1564 -1408
rect 2306 -1408 2364 -1402
rect 2306 -1410 2318 -1408
rect 1552 -1440 2318 -1410
rect 1552 -1442 1564 -1440
rect 1506 -1448 1564 -1442
rect 2306 -1442 2318 -1440
rect 2352 -1410 2364 -1408
rect 3106 -1408 3164 -1402
rect 3106 -1410 3118 -1408
rect 2352 -1440 3118 -1410
rect 2352 -1442 2364 -1440
rect 2306 -1448 2364 -1442
rect 3106 -1442 3118 -1440
rect 3152 -1410 3164 -1408
rect 3906 -1408 3964 -1402
rect 3906 -1410 3918 -1408
rect 3152 -1440 3918 -1410
rect 3152 -1442 3164 -1440
rect 3106 -1448 3164 -1442
rect 3906 -1442 3918 -1440
rect 3952 -1410 3964 -1408
rect 4706 -1408 4764 -1402
rect 4706 -1410 4718 -1408
rect 3952 -1440 4718 -1410
rect 3952 -1442 3964 -1440
rect 3906 -1448 3964 -1442
rect 4706 -1442 4718 -1440
rect 4752 -1410 4764 -1408
rect 5506 -1408 5564 -1402
rect 5506 -1410 5518 -1408
rect 4752 -1440 5518 -1410
rect 4752 -1442 4764 -1440
rect 4706 -1448 4764 -1442
rect 5506 -1442 5518 -1440
rect 5552 -1410 5564 -1408
rect 6306 -1408 6364 -1402
rect 6306 -1410 6318 -1408
rect 5552 -1440 6318 -1410
rect 5552 -1442 5564 -1440
rect 5506 -1448 5564 -1442
rect 6306 -1442 6318 -1440
rect 6352 -1410 6364 -1408
rect 7106 -1408 7164 -1402
rect 7106 -1410 7118 -1408
rect 6352 -1440 7118 -1410
rect 6352 -1442 6364 -1440
rect 6306 -1448 6364 -1442
rect 7106 -1442 7118 -1440
rect 7152 -1410 7164 -1408
rect 7906 -1408 7964 -1402
rect 7906 -1410 7918 -1408
rect 7152 -1440 7918 -1410
rect 7152 -1442 7164 -1440
rect 7106 -1448 7164 -1442
rect 7906 -1442 7918 -1440
rect 7952 -1410 7964 -1408
rect 8706 -1408 8764 -1402
rect 8706 -1410 8718 -1408
rect 7952 -1440 8718 -1410
rect 7952 -1442 7964 -1440
rect 7906 -1448 7964 -1442
rect 8706 -1442 8718 -1440
rect 8752 -1410 8764 -1408
rect 9506 -1408 9564 -1402
rect 9506 -1410 9518 -1408
rect 8752 -1440 9518 -1410
rect 8752 -1442 8764 -1440
rect 8706 -1448 8764 -1442
rect 9506 -1442 9518 -1440
rect 9552 -1410 9564 -1408
rect 10306 -1408 10364 -1402
rect 10306 -1410 10318 -1408
rect 9552 -1440 10318 -1410
rect 9552 -1442 9564 -1440
rect 9506 -1448 9564 -1442
rect 10306 -1442 10318 -1440
rect 10352 -1410 10364 -1408
rect 11106 -1408 11164 -1402
rect 11106 -1410 11118 -1408
rect 10352 -1440 11118 -1410
rect 10352 -1442 10364 -1440
rect 10306 -1448 10364 -1442
rect 11106 -1442 11118 -1440
rect 11152 -1410 11164 -1408
rect 11906 -1408 11964 -1402
rect 11906 -1410 11918 -1408
rect 11152 -1440 11918 -1410
rect 11152 -1442 11164 -1440
rect 11106 -1448 11164 -1442
rect 11906 -1442 11918 -1440
rect 11952 -1410 11964 -1408
rect 12706 -1408 12764 -1402
rect 12706 -1410 12718 -1408
rect 11952 -1440 12718 -1410
rect 11952 -1442 11964 -1440
rect 11906 -1448 11964 -1442
rect 12706 -1442 12718 -1440
rect 12752 -1410 12764 -1408
rect 14434 -1410 14440 -1399
rect 12752 -1440 12776 -1410
rect 14400 -1440 14440 -1410
rect 12752 -1442 12764 -1440
rect 12706 -1448 12764 -1442
rect 14434 -1451 14440 -1440
rect 14492 -1451 14498 -1399
rect 14526 -1451 14553 -1399
rect 14605 -1451 14617 -1399
rect 14669 -1451 14697 -1399
rect 14526 -1457 14697 -1451
rect 14725 -1399 14777 -1393
rect 14725 -1457 14777 -1451
rect 14805 -1399 15136 -1393
rect 14805 -1451 14816 -1399
rect 14868 -1408 14880 -1399
rect 14932 -1408 14944 -1399
rect 14996 -1408 15008 -1399
rect 15060 -1408 15072 -1399
rect 14876 -1442 14880 -1408
rect 14868 -1451 14880 -1442
rect 14932 -1451 14944 -1442
rect 14996 -1451 15008 -1442
rect 15060 -1451 15072 -1442
rect 15124 -1451 15136 -1399
rect 14805 -1457 15136 -1451
rect 15206 -1399 15537 -1393
rect 15206 -1451 15217 -1399
rect 15269 -1408 15281 -1399
rect 15333 -1408 15345 -1399
rect 15397 -1408 15409 -1399
rect 15461 -1408 15473 -1399
rect 15461 -1442 15465 -1408
rect 15269 -1451 15281 -1442
rect 15333 -1451 15345 -1442
rect 15397 -1451 15409 -1442
rect 15461 -1451 15473 -1442
rect 15525 -1451 15537 -1399
rect 15206 -1457 15537 -1451
rect 15565 -1399 15617 -1393
rect 15565 -1457 15617 -1451
rect 15645 -1399 15816 -1393
rect 15645 -1451 15672 -1399
rect 15724 -1451 15736 -1399
rect 15788 -1451 15816 -1399
rect 15645 -1457 15816 -1451
rect -94 -1508 -36 -1502
rect -94 -1510 -82 -1508
rect -106 -1540 -82 -1510
rect -94 -1542 -82 -1540
rect -48 -1510 -36 -1508
rect 706 -1508 764 -1502
rect 706 -1510 718 -1508
rect -48 -1540 718 -1510
rect -48 -1542 -36 -1540
rect -94 -1548 -36 -1542
rect 706 -1542 718 -1540
rect 752 -1510 764 -1508
rect 1506 -1508 1564 -1502
rect 1506 -1510 1518 -1508
rect 752 -1540 1518 -1510
rect 752 -1542 764 -1540
rect 706 -1548 764 -1542
rect 1506 -1542 1518 -1540
rect 1552 -1510 1564 -1508
rect 2306 -1508 2364 -1502
rect 2306 -1510 2318 -1508
rect 1552 -1540 2318 -1510
rect 1552 -1542 1564 -1540
rect 1506 -1548 1564 -1542
rect 2306 -1542 2318 -1540
rect 2352 -1510 2364 -1508
rect 3106 -1508 3164 -1502
rect 3106 -1510 3118 -1508
rect 2352 -1540 3118 -1510
rect 2352 -1542 2364 -1540
rect 2306 -1548 2364 -1542
rect 3106 -1542 3118 -1540
rect 3152 -1510 3164 -1508
rect 3906 -1508 3964 -1502
rect 3906 -1510 3918 -1508
rect 3152 -1540 3918 -1510
rect 3152 -1542 3164 -1540
rect 3106 -1548 3164 -1542
rect 3906 -1542 3918 -1540
rect 3952 -1510 3964 -1508
rect 4706 -1508 4764 -1502
rect 4706 -1510 4718 -1508
rect 3952 -1540 4718 -1510
rect 3952 -1542 3964 -1540
rect 3906 -1548 3964 -1542
rect 4706 -1542 4718 -1540
rect 4752 -1510 4764 -1508
rect 5506 -1508 5564 -1502
rect 5506 -1510 5518 -1508
rect 4752 -1540 5518 -1510
rect 4752 -1542 4764 -1540
rect 4706 -1548 4764 -1542
rect 5506 -1542 5518 -1540
rect 5552 -1510 5564 -1508
rect 6306 -1508 6364 -1502
rect 6306 -1510 6318 -1508
rect 5552 -1540 6318 -1510
rect 5552 -1542 5564 -1540
rect 5506 -1548 5564 -1542
rect 6306 -1542 6318 -1540
rect 6352 -1510 6364 -1508
rect 7106 -1508 7164 -1502
rect 7106 -1510 7118 -1508
rect 6352 -1540 7118 -1510
rect 6352 -1542 6364 -1540
rect 6306 -1548 6364 -1542
rect 7106 -1542 7118 -1540
rect 7152 -1510 7164 -1508
rect 7906 -1508 7964 -1502
rect 7906 -1510 7918 -1508
rect 7152 -1540 7918 -1510
rect 7152 -1542 7164 -1540
rect 7106 -1548 7164 -1542
rect 7906 -1542 7918 -1540
rect 7952 -1510 7964 -1508
rect 8706 -1508 8764 -1502
rect 8706 -1510 8718 -1508
rect 7952 -1540 8718 -1510
rect 7952 -1542 7964 -1540
rect 7906 -1548 7964 -1542
rect 8706 -1542 8718 -1540
rect 8752 -1510 8764 -1508
rect 9506 -1508 9564 -1502
rect 9506 -1510 9518 -1508
rect 8752 -1540 9518 -1510
rect 8752 -1542 8764 -1540
rect 8706 -1548 8764 -1542
rect 9506 -1542 9518 -1540
rect 9552 -1510 9564 -1508
rect 10306 -1508 10364 -1502
rect 10306 -1510 10318 -1508
rect 9552 -1540 10318 -1510
rect 9552 -1542 9564 -1540
rect 9506 -1548 9564 -1542
rect 10306 -1542 10318 -1540
rect 10352 -1510 10364 -1508
rect 11106 -1508 11164 -1502
rect 11106 -1510 11118 -1508
rect 10352 -1540 11118 -1510
rect 10352 -1542 10364 -1540
rect 10306 -1548 10364 -1542
rect 11106 -1542 11118 -1540
rect 11152 -1510 11164 -1508
rect 11906 -1508 11964 -1502
rect 11906 -1510 11918 -1508
rect 11152 -1540 11918 -1510
rect 11152 -1542 11164 -1540
rect 11106 -1548 11164 -1542
rect 11906 -1542 11918 -1540
rect 11952 -1510 11964 -1508
rect 12706 -1508 12764 -1502
rect 12706 -1510 12718 -1508
rect 11952 -1540 12718 -1510
rect 11952 -1542 11964 -1540
rect 11906 -1548 11964 -1542
rect 12706 -1542 12718 -1540
rect 12752 -1510 12764 -1508
rect 14520 -1508 15136 -1502
rect 14520 -1510 14560 -1508
rect 12752 -1540 12776 -1510
rect 14400 -1540 14560 -1510
rect 12752 -1542 12764 -1540
rect 12706 -1548 12764 -1542
rect 14520 -1542 14560 -1540
rect 14594 -1542 14632 -1508
rect 14666 -1542 14841 -1508
rect 14875 -1542 14913 -1508
rect 14947 -1542 14985 -1508
rect 15019 -1542 15057 -1508
rect 15091 -1542 15136 -1508
rect 14520 -1548 15136 -1542
rect 15206 -1551 15212 -1499
rect 15264 -1502 15270 -1499
rect 15264 -1508 15822 -1502
rect 15285 -1542 15323 -1508
rect 15357 -1542 15395 -1508
rect 15429 -1542 15467 -1508
rect 15501 -1542 15676 -1508
rect 15710 -1542 15748 -1508
rect 15782 -1542 15822 -1508
rect 15264 -1548 15822 -1542
rect 15264 -1551 15270 -1548
rect 14526 -1599 14697 -1593
rect -94 -1608 -36 -1602
rect -94 -1610 -82 -1608
rect -106 -1640 -82 -1610
rect -94 -1642 -82 -1640
rect -48 -1610 -36 -1608
rect 706 -1608 764 -1602
rect 706 -1610 718 -1608
rect -48 -1640 718 -1610
rect -48 -1642 -36 -1640
rect -94 -1648 -36 -1642
rect 706 -1642 718 -1640
rect 752 -1610 764 -1608
rect 1506 -1608 1564 -1602
rect 1506 -1610 1518 -1608
rect 752 -1640 1518 -1610
rect 752 -1642 764 -1640
rect 706 -1648 764 -1642
rect 1506 -1642 1518 -1640
rect 1552 -1610 1564 -1608
rect 2306 -1608 2364 -1602
rect 2306 -1610 2318 -1608
rect 1552 -1640 2318 -1610
rect 1552 -1642 1564 -1640
rect 1506 -1648 1564 -1642
rect 2306 -1642 2318 -1640
rect 2352 -1610 2364 -1608
rect 3106 -1608 3164 -1602
rect 3106 -1610 3118 -1608
rect 2352 -1640 3118 -1610
rect 2352 -1642 2364 -1640
rect 2306 -1648 2364 -1642
rect 3106 -1642 3118 -1640
rect 3152 -1610 3164 -1608
rect 3906 -1608 3964 -1602
rect 3906 -1610 3918 -1608
rect 3152 -1640 3918 -1610
rect 3152 -1642 3164 -1640
rect 3106 -1648 3164 -1642
rect 3906 -1642 3918 -1640
rect 3952 -1610 3964 -1608
rect 4706 -1608 4764 -1602
rect 4706 -1610 4718 -1608
rect 3952 -1640 4718 -1610
rect 3952 -1642 3964 -1640
rect 3906 -1648 3964 -1642
rect 4706 -1642 4718 -1640
rect 4752 -1610 4764 -1608
rect 5506 -1608 5564 -1602
rect 5506 -1610 5518 -1608
rect 4752 -1640 5518 -1610
rect 4752 -1642 4764 -1640
rect 4706 -1648 4764 -1642
rect 5506 -1642 5518 -1640
rect 5552 -1610 5564 -1608
rect 6306 -1608 6364 -1602
rect 6306 -1610 6318 -1608
rect 5552 -1640 6318 -1610
rect 5552 -1642 5564 -1640
rect 5506 -1648 5564 -1642
rect 6306 -1642 6318 -1640
rect 6352 -1610 6364 -1608
rect 7106 -1608 7164 -1602
rect 7106 -1610 7118 -1608
rect 6352 -1640 7118 -1610
rect 6352 -1642 6364 -1640
rect 6306 -1648 6364 -1642
rect 7106 -1642 7118 -1640
rect 7152 -1610 7164 -1608
rect 7906 -1608 7964 -1602
rect 7906 -1610 7918 -1608
rect 7152 -1640 7918 -1610
rect 7152 -1642 7164 -1640
rect 7106 -1648 7164 -1642
rect 7906 -1642 7918 -1640
rect 7952 -1610 7964 -1608
rect 8706 -1608 8764 -1602
rect 8706 -1610 8718 -1608
rect 7952 -1640 8718 -1610
rect 7952 -1642 7964 -1640
rect 7906 -1648 7964 -1642
rect 8706 -1642 8718 -1640
rect 8752 -1610 8764 -1608
rect 9506 -1608 9564 -1602
rect 9506 -1610 9518 -1608
rect 8752 -1640 9518 -1610
rect 8752 -1642 8764 -1640
rect 8706 -1648 8764 -1642
rect 9506 -1642 9518 -1640
rect 9552 -1610 9564 -1608
rect 10306 -1608 10364 -1602
rect 10306 -1610 10318 -1608
rect 9552 -1640 10318 -1610
rect 9552 -1642 9564 -1640
rect 9506 -1648 9564 -1642
rect 10306 -1642 10318 -1640
rect 10352 -1610 10364 -1608
rect 11106 -1608 11164 -1602
rect 11106 -1610 11118 -1608
rect 10352 -1640 11118 -1610
rect 10352 -1642 10364 -1640
rect 10306 -1648 10364 -1642
rect 11106 -1642 11118 -1640
rect 11152 -1610 11164 -1608
rect 11906 -1608 11964 -1602
rect 11906 -1610 11918 -1608
rect 11152 -1640 11918 -1610
rect 11152 -1642 11164 -1640
rect 11106 -1648 11164 -1642
rect 11906 -1642 11918 -1640
rect 11952 -1610 11964 -1608
rect 12706 -1608 12764 -1602
rect 12706 -1610 12718 -1608
rect 11952 -1640 12718 -1610
rect 11952 -1642 11964 -1640
rect 11906 -1648 11964 -1642
rect 12706 -1642 12718 -1640
rect 12752 -1610 12764 -1608
rect 14434 -1610 14440 -1599
rect 12752 -1640 12776 -1610
rect 14400 -1640 14440 -1610
rect 12752 -1642 12764 -1640
rect 12706 -1648 12764 -1642
rect 14434 -1651 14440 -1640
rect 14492 -1651 14498 -1599
rect 14526 -1651 14553 -1599
rect 14605 -1651 14617 -1599
rect 14669 -1651 14697 -1599
rect 14526 -1657 14697 -1651
rect 14725 -1599 14777 -1593
rect 14725 -1657 14777 -1651
rect 14805 -1599 15136 -1593
rect 14805 -1651 14816 -1599
rect 14868 -1608 14880 -1599
rect 14932 -1608 14944 -1599
rect 14996 -1608 15008 -1599
rect 15060 -1608 15072 -1599
rect 14876 -1642 14880 -1608
rect 14868 -1651 14880 -1642
rect 14932 -1651 14944 -1642
rect 14996 -1651 15008 -1642
rect 15060 -1651 15072 -1642
rect 15124 -1651 15136 -1599
rect 14805 -1657 15136 -1651
rect 15206 -1599 15537 -1593
rect 15206 -1651 15217 -1599
rect 15269 -1608 15281 -1599
rect 15333 -1608 15345 -1599
rect 15397 -1608 15409 -1599
rect 15461 -1608 15473 -1599
rect 15461 -1642 15465 -1608
rect 15269 -1651 15281 -1642
rect 15333 -1651 15345 -1642
rect 15397 -1651 15409 -1642
rect 15461 -1651 15473 -1642
rect 15525 -1651 15537 -1599
rect 15206 -1657 15537 -1651
rect 15565 -1599 15617 -1593
rect 15565 -1657 15617 -1651
rect 15645 -1599 15816 -1593
rect 15645 -1651 15672 -1599
rect 15724 -1651 15736 -1599
rect 15788 -1651 15816 -1599
rect 15645 -1657 15816 -1651
rect -94 -1708 -36 -1702
rect -94 -1710 -82 -1708
rect -106 -1740 -82 -1710
rect -94 -1742 -82 -1740
rect -48 -1710 -36 -1708
rect 706 -1708 764 -1702
rect 706 -1710 718 -1708
rect -48 -1740 718 -1710
rect -48 -1742 -36 -1740
rect -94 -1748 -36 -1742
rect 706 -1742 718 -1740
rect 752 -1710 764 -1708
rect 1506 -1708 1564 -1702
rect 1506 -1710 1518 -1708
rect 752 -1740 1518 -1710
rect 752 -1742 764 -1740
rect 706 -1748 764 -1742
rect 1506 -1742 1518 -1740
rect 1552 -1710 1564 -1708
rect 2306 -1708 2364 -1702
rect 2306 -1710 2318 -1708
rect 1552 -1740 2318 -1710
rect 1552 -1742 1564 -1740
rect 1506 -1748 1564 -1742
rect 2306 -1742 2318 -1740
rect 2352 -1710 2364 -1708
rect 3106 -1708 3164 -1702
rect 3106 -1710 3118 -1708
rect 2352 -1740 3118 -1710
rect 2352 -1742 2364 -1740
rect 2306 -1748 2364 -1742
rect 3106 -1742 3118 -1740
rect 3152 -1710 3164 -1708
rect 3906 -1708 3964 -1702
rect 3906 -1710 3918 -1708
rect 3152 -1740 3918 -1710
rect 3152 -1742 3164 -1740
rect 3106 -1748 3164 -1742
rect 3906 -1742 3918 -1740
rect 3952 -1710 3964 -1708
rect 4706 -1708 4764 -1702
rect 4706 -1710 4718 -1708
rect 3952 -1740 4718 -1710
rect 3952 -1742 3964 -1740
rect 3906 -1748 3964 -1742
rect 4706 -1742 4718 -1740
rect 4752 -1710 4764 -1708
rect 5506 -1708 5564 -1702
rect 5506 -1710 5518 -1708
rect 4752 -1740 5518 -1710
rect 4752 -1742 4764 -1740
rect 4706 -1748 4764 -1742
rect 5506 -1742 5518 -1740
rect 5552 -1710 5564 -1708
rect 6306 -1708 6364 -1702
rect 6306 -1710 6318 -1708
rect 5552 -1740 6318 -1710
rect 5552 -1742 5564 -1740
rect 5506 -1748 5564 -1742
rect 6306 -1742 6318 -1740
rect 6352 -1710 6364 -1708
rect 7106 -1708 7164 -1702
rect 7106 -1710 7118 -1708
rect 6352 -1740 7118 -1710
rect 6352 -1742 6364 -1740
rect 6306 -1748 6364 -1742
rect 7106 -1742 7118 -1740
rect 7152 -1710 7164 -1708
rect 7906 -1708 7964 -1702
rect 7906 -1710 7918 -1708
rect 7152 -1740 7918 -1710
rect 7152 -1742 7164 -1740
rect 7106 -1748 7164 -1742
rect 7906 -1742 7918 -1740
rect 7952 -1710 7964 -1708
rect 8706 -1708 8764 -1702
rect 8706 -1710 8718 -1708
rect 7952 -1740 8718 -1710
rect 7952 -1742 7964 -1740
rect 7906 -1748 7964 -1742
rect 8706 -1742 8718 -1740
rect 8752 -1710 8764 -1708
rect 9506 -1708 9564 -1702
rect 9506 -1710 9518 -1708
rect 8752 -1740 9518 -1710
rect 8752 -1742 8764 -1740
rect 8706 -1748 8764 -1742
rect 9506 -1742 9518 -1740
rect 9552 -1710 9564 -1708
rect 10306 -1708 10364 -1702
rect 10306 -1710 10318 -1708
rect 9552 -1740 10318 -1710
rect 9552 -1742 9564 -1740
rect 9506 -1748 9564 -1742
rect 10306 -1742 10318 -1740
rect 10352 -1710 10364 -1708
rect 11106 -1708 11164 -1702
rect 11106 -1710 11118 -1708
rect 10352 -1740 11118 -1710
rect 10352 -1742 10364 -1740
rect 10306 -1748 10364 -1742
rect 11106 -1742 11118 -1740
rect 11152 -1710 11164 -1708
rect 11906 -1708 11964 -1702
rect 11906 -1710 11918 -1708
rect 11152 -1740 11918 -1710
rect 11152 -1742 11164 -1740
rect 11106 -1748 11164 -1742
rect 11906 -1742 11918 -1740
rect 11952 -1710 11964 -1708
rect 12706 -1708 12764 -1702
rect 12706 -1710 12718 -1708
rect 11952 -1740 12718 -1710
rect 11952 -1742 11964 -1740
rect 11906 -1748 11964 -1742
rect 12706 -1742 12718 -1740
rect 12752 -1710 12764 -1708
rect 14520 -1708 15136 -1702
rect 14520 -1710 14560 -1708
rect 12752 -1740 12776 -1710
rect 14400 -1740 14560 -1710
rect 12752 -1742 12764 -1740
rect 12706 -1748 12764 -1742
rect 14520 -1742 14560 -1740
rect 14594 -1742 14632 -1708
rect 14666 -1742 14841 -1708
rect 14875 -1742 14913 -1708
rect 14947 -1742 14985 -1708
rect 15019 -1742 15057 -1708
rect 15091 -1742 15136 -1708
rect 14520 -1748 15136 -1742
rect 15206 -1751 15212 -1699
rect 15264 -1702 15270 -1699
rect 15264 -1708 15822 -1702
rect 15285 -1742 15323 -1708
rect 15357 -1742 15395 -1708
rect 15429 -1742 15467 -1708
rect 15501 -1742 15676 -1708
rect 15710 -1742 15748 -1708
rect 15782 -1742 15822 -1708
rect 15264 -1748 15822 -1742
rect 15264 -1751 15270 -1748
rect 14526 -1799 14697 -1793
rect -94 -1808 -36 -1802
rect -94 -1810 -82 -1808
rect -106 -1840 -82 -1810
rect -94 -1842 -82 -1840
rect -48 -1810 -36 -1808
rect 706 -1808 764 -1802
rect 706 -1810 718 -1808
rect -48 -1840 718 -1810
rect -48 -1842 -36 -1840
rect -94 -1848 -36 -1842
rect 706 -1842 718 -1840
rect 752 -1810 764 -1808
rect 1506 -1808 1564 -1802
rect 1506 -1810 1518 -1808
rect 752 -1840 1518 -1810
rect 752 -1842 764 -1840
rect 706 -1848 764 -1842
rect 1506 -1842 1518 -1840
rect 1552 -1810 1564 -1808
rect 2306 -1808 2364 -1802
rect 2306 -1810 2318 -1808
rect 1552 -1840 2318 -1810
rect 1552 -1842 1564 -1840
rect 1506 -1848 1564 -1842
rect 2306 -1842 2318 -1840
rect 2352 -1810 2364 -1808
rect 3106 -1808 3164 -1802
rect 3106 -1810 3118 -1808
rect 2352 -1840 3118 -1810
rect 2352 -1842 2364 -1840
rect 2306 -1848 2364 -1842
rect 3106 -1842 3118 -1840
rect 3152 -1810 3164 -1808
rect 3906 -1808 3964 -1802
rect 3906 -1810 3918 -1808
rect 3152 -1840 3918 -1810
rect 3152 -1842 3164 -1840
rect 3106 -1848 3164 -1842
rect 3906 -1842 3918 -1840
rect 3952 -1810 3964 -1808
rect 4706 -1808 4764 -1802
rect 4706 -1810 4718 -1808
rect 3952 -1840 4718 -1810
rect 3952 -1842 3964 -1840
rect 3906 -1848 3964 -1842
rect 4706 -1842 4718 -1840
rect 4752 -1810 4764 -1808
rect 5506 -1808 5564 -1802
rect 5506 -1810 5518 -1808
rect 4752 -1840 5518 -1810
rect 4752 -1842 4764 -1840
rect 4706 -1848 4764 -1842
rect 5506 -1842 5518 -1840
rect 5552 -1810 5564 -1808
rect 6306 -1808 6364 -1802
rect 6306 -1810 6318 -1808
rect 5552 -1840 6318 -1810
rect 5552 -1842 5564 -1840
rect 5506 -1848 5564 -1842
rect 6306 -1842 6318 -1840
rect 6352 -1810 6364 -1808
rect 7106 -1808 7164 -1802
rect 7106 -1810 7118 -1808
rect 6352 -1840 7118 -1810
rect 6352 -1842 6364 -1840
rect 6306 -1848 6364 -1842
rect 7106 -1842 7118 -1840
rect 7152 -1810 7164 -1808
rect 7906 -1808 7964 -1802
rect 7906 -1810 7918 -1808
rect 7152 -1840 7918 -1810
rect 7152 -1842 7164 -1840
rect 7106 -1848 7164 -1842
rect 7906 -1842 7918 -1840
rect 7952 -1810 7964 -1808
rect 8706 -1808 8764 -1802
rect 8706 -1810 8718 -1808
rect 7952 -1840 8718 -1810
rect 7952 -1842 7964 -1840
rect 7906 -1848 7964 -1842
rect 8706 -1842 8718 -1840
rect 8752 -1810 8764 -1808
rect 9506 -1808 9564 -1802
rect 9506 -1810 9518 -1808
rect 8752 -1840 9518 -1810
rect 8752 -1842 8764 -1840
rect 8706 -1848 8764 -1842
rect 9506 -1842 9518 -1840
rect 9552 -1810 9564 -1808
rect 10306 -1808 10364 -1802
rect 10306 -1810 10318 -1808
rect 9552 -1840 10318 -1810
rect 9552 -1842 9564 -1840
rect 9506 -1848 9564 -1842
rect 10306 -1842 10318 -1840
rect 10352 -1810 10364 -1808
rect 11106 -1808 11164 -1802
rect 11106 -1810 11118 -1808
rect 10352 -1840 11118 -1810
rect 10352 -1842 10364 -1840
rect 10306 -1848 10364 -1842
rect 11106 -1842 11118 -1840
rect 11152 -1810 11164 -1808
rect 11906 -1808 11964 -1802
rect 11906 -1810 11918 -1808
rect 11152 -1840 11918 -1810
rect 11152 -1842 11164 -1840
rect 11106 -1848 11164 -1842
rect 11906 -1842 11918 -1840
rect 11952 -1810 11964 -1808
rect 12706 -1808 12764 -1802
rect 12706 -1810 12718 -1808
rect 11952 -1840 12718 -1810
rect 11952 -1842 11964 -1840
rect 11906 -1848 11964 -1842
rect 12706 -1842 12718 -1840
rect 12752 -1810 12764 -1808
rect 14434 -1810 14440 -1799
rect 12752 -1840 12776 -1810
rect 14400 -1840 14440 -1810
rect 12752 -1842 12764 -1840
rect 12706 -1848 12764 -1842
rect 14434 -1851 14440 -1840
rect 14492 -1851 14498 -1799
rect 14526 -1851 14553 -1799
rect 14605 -1851 14617 -1799
rect 14669 -1851 14697 -1799
rect 14526 -1857 14697 -1851
rect 14725 -1799 14777 -1793
rect 14725 -1857 14777 -1851
rect 14805 -1799 15136 -1793
rect 14805 -1851 14816 -1799
rect 14868 -1808 14880 -1799
rect 14932 -1808 14944 -1799
rect 14996 -1808 15008 -1799
rect 15060 -1808 15072 -1799
rect 14876 -1842 14880 -1808
rect 14868 -1851 14880 -1842
rect 14932 -1851 14944 -1842
rect 14996 -1851 15008 -1842
rect 15060 -1851 15072 -1842
rect 15124 -1851 15136 -1799
rect 14805 -1857 15136 -1851
rect 15206 -1799 15537 -1793
rect 15206 -1851 15217 -1799
rect 15269 -1808 15281 -1799
rect 15333 -1808 15345 -1799
rect 15397 -1808 15409 -1799
rect 15461 -1808 15473 -1799
rect 15461 -1842 15465 -1808
rect 15269 -1851 15281 -1842
rect 15333 -1851 15345 -1842
rect 15397 -1851 15409 -1842
rect 15461 -1851 15473 -1842
rect 15525 -1851 15537 -1799
rect 15206 -1857 15537 -1851
rect 15565 -1799 15617 -1793
rect 15565 -1857 15617 -1851
rect 15645 -1799 15816 -1793
rect 15645 -1851 15672 -1799
rect 15724 -1851 15736 -1799
rect 15788 -1851 15816 -1799
rect 15645 -1857 15816 -1851
rect -94 -1908 -36 -1902
rect -94 -1910 -82 -1908
rect -106 -1940 -82 -1910
rect -94 -1942 -82 -1940
rect -48 -1910 -36 -1908
rect 706 -1908 764 -1902
rect 706 -1910 718 -1908
rect -48 -1940 718 -1910
rect -48 -1942 -36 -1940
rect -94 -1948 -36 -1942
rect 706 -1942 718 -1940
rect 752 -1910 764 -1908
rect 1506 -1908 1564 -1902
rect 1506 -1910 1518 -1908
rect 752 -1940 1518 -1910
rect 752 -1942 764 -1940
rect 706 -1948 764 -1942
rect 1506 -1942 1518 -1940
rect 1552 -1910 1564 -1908
rect 2306 -1908 2364 -1902
rect 2306 -1910 2318 -1908
rect 1552 -1940 2318 -1910
rect 1552 -1942 1564 -1940
rect 1506 -1948 1564 -1942
rect 2306 -1942 2318 -1940
rect 2352 -1910 2364 -1908
rect 3106 -1908 3164 -1902
rect 3106 -1910 3118 -1908
rect 2352 -1940 3118 -1910
rect 2352 -1942 2364 -1940
rect 2306 -1948 2364 -1942
rect 3106 -1942 3118 -1940
rect 3152 -1910 3164 -1908
rect 3906 -1908 3964 -1902
rect 3906 -1910 3918 -1908
rect 3152 -1940 3918 -1910
rect 3152 -1942 3164 -1940
rect 3106 -1948 3164 -1942
rect 3906 -1942 3918 -1940
rect 3952 -1910 3964 -1908
rect 4706 -1908 4764 -1902
rect 4706 -1910 4718 -1908
rect 3952 -1940 4718 -1910
rect 3952 -1942 3964 -1940
rect 3906 -1948 3964 -1942
rect 4706 -1942 4718 -1940
rect 4752 -1910 4764 -1908
rect 5506 -1908 5564 -1902
rect 5506 -1910 5518 -1908
rect 4752 -1940 5518 -1910
rect 4752 -1942 4764 -1940
rect 4706 -1948 4764 -1942
rect 5506 -1942 5518 -1940
rect 5552 -1910 5564 -1908
rect 6306 -1908 6364 -1902
rect 6306 -1910 6318 -1908
rect 5552 -1940 6318 -1910
rect 5552 -1942 5564 -1940
rect 5506 -1948 5564 -1942
rect 6306 -1942 6318 -1940
rect 6352 -1910 6364 -1908
rect 7106 -1908 7164 -1902
rect 7106 -1910 7118 -1908
rect 6352 -1940 7118 -1910
rect 6352 -1942 6364 -1940
rect 6306 -1948 6364 -1942
rect 7106 -1942 7118 -1940
rect 7152 -1910 7164 -1908
rect 7906 -1908 7964 -1902
rect 7906 -1910 7918 -1908
rect 7152 -1940 7918 -1910
rect 7152 -1942 7164 -1940
rect 7106 -1948 7164 -1942
rect 7906 -1942 7918 -1940
rect 7952 -1910 7964 -1908
rect 8706 -1908 8764 -1902
rect 8706 -1910 8718 -1908
rect 7952 -1940 8718 -1910
rect 7952 -1942 7964 -1940
rect 7906 -1948 7964 -1942
rect 8706 -1942 8718 -1940
rect 8752 -1910 8764 -1908
rect 9506 -1908 9564 -1902
rect 9506 -1910 9518 -1908
rect 8752 -1940 9518 -1910
rect 8752 -1942 8764 -1940
rect 8706 -1948 8764 -1942
rect 9506 -1942 9518 -1940
rect 9552 -1910 9564 -1908
rect 10306 -1908 10364 -1902
rect 10306 -1910 10318 -1908
rect 9552 -1940 10318 -1910
rect 9552 -1942 9564 -1940
rect 9506 -1948 9564 -1942
rect 10306 -1942 10318 -1940
rect 10352 -1910 10364 -1908
rect 11106 -1908 11164 -1902
rect 11106 -1910 11118 -1908
rect 10352 -1940 11118 -1910
rect 10352 -1942 10364 -1940
rect 10306 -1948 10364 -1942
rect 11106 -1942 11118 -1940
rect 11152 -1910 11164 -1908
rect 11906 -1908 11964 -1902
rect 11906 -1910 11918 -1908
rect 11152 -1940 11918 -1910
rect 11152 -1942 11164 -1940
rect 11106 -1948 11164 -1942
rect 11906 -1942 11918 -1940
rect 11952 -1910 11964 -1908
rect 12706 -1908 12764 -1902
rect 12706 -1910 12718 -1908
rect 11952 -1940 12718 -1910
rect 11952 -1942 11964 -1940
rect 11906 -1948 11964 -1942
rect 12706 -1942 12718 -1940
rect 12752 -1910 12764 -1908
rect 14520 -1908 15136 -1902
rect 14520 -1910 14560 -1908
rect 12752 -1940 12776 -1910
rect 14400 -1940 14560 -1910
rect 12752 -1942 12764 -1940
rect 12706 -1948 12764 -1942
rect 14520 -1942 14560 -1940
rect 14594 -1942 14632 -1908
rect 14666 -1942 14841 -1908
rect 14875 -1942 14913 -1908
rect 14947 -1942 14985 -1908
rect 15019 -1942 15057 -1908
rect 15091 -1942 15136 -1908
rect 14520 -1948 15136 -1942
rect 15206 -1951 15212 -1899
rect 15264 -1902 15270 -1899
rect 15264 -1908 15822 -1902
rect 15285 -1942 15323 -1908
rect 15357 -1942 15395 -1908
rect 15429 -1942 15467 -1908
rect 15501 -1942 15676 -1908
rect 15710 -1942 15748 -1908
rect 15782 -1942 15822 -1908
rect 15264 -1948 15822 -1942
rect 15264 -1951 15270 -1948
rect 14526 -1999 14697 -1993
rect -94 -2008 -36 -2002
rect -94 -2010 -82 -2008
rect -106 -2040 -82 -2010
rect -94 -2042 -82 -2040
rect -48 -2010 -36 -2008
rect 706 -2008 764 -2002
rect 706 -2010 718 -2008
rect -48 -2040 718 -2010
rect -48 -2042 -36 -2040
rect -94 -2048 -36 -2042
rect 706 -2042 718 -2040
rect 752 -2010 764 -2008
rect 1506 -2008 1564 -2002
rect 1506 -2010 1518 -2008
rect 752 -2040 1518 -2010
rect 752 -2042 764 -2040
rect 706 -2048 764 -2042
rect 1506 -2042 1518 -2040
rect 1552 -2010 1564 -2008
rect 2306 -2008 2364 -2002
rect 2306 -2010 2318 -2008
rect 1552 -2040 2318 -2010
rect 1552 -2042 1564 -2040
rect 1506 -2048 1564 -2042
rect 2306 -2042 2318 -2040
rect 2352 -2010 2364 -2008
rect 3106 -2008 3164 -2002
rect 3106 -2010 3118 -2008
rect 2352 -2040 3118 -2010
rect 2352 -2042 2364 -2040
rect 2306 -2048 2364 -2042
rect 3106 -2042 3118 -2040
rect 3152 -2010 3164 -2008
rect 3906 -2008 3964 -2002
rect 3906 -2010 3918 -2008
rect 3152 -2040 3918 -2010
rect 3152 -2042 3164 -2040
rect 3106 -2048 3164 -2042
rect 3906 -2042 3918 -2040
rect 3952 -2010 3964 -2008
rect 4706 -2008 4764 -2002
rect 4706 -2010 4718 -2008
rect 3952 -2040 4718 -2010
rect 3952 -2042 3964 -2040
rect 3906 -2048 3964 -2042
rect 4706 -2042 4718 -2040
rect 4752 -2010 4764 -2008
rect 5506 -2008 5564 -2002
rect 5506 -2010 5518 -2008
rect 4752 -2040 5518 -2010
rect 4752 -2042 4764 -2040
rect 4706 -2048 4764 -2042
rect 5506 -2042 5518 -2040
rect 5552 -2010 5564 -2008
rect 6306 -2008 6364 -2002
rect 6306 -2010 6318 -2008
rect 5552 -2040 6318 -2010
rect 5552 -2042 5564 -2040
rect 5506 -2048 5564 -2042
rect 6306 -2042 6318 -2040
rect 6352 -2010 6364 -2008
rect 7106 -2008 7164 -2002
rect 7106 -2010 7118 -2008
rect 6352 -2040 7118 -2010
rect 6352 -2042 6364 -2040
rect 6306 -2048 6364 -2042
rect 7106 -2042 7118 -2040
rect 7152 -2010 7164 -2008
rect 7906 -2008 7964 -2002
rect 7906 -2010 7918 -2008
rect 7152 -2040 7918 -2010
rect 7152 -2042 7164 -2040
rect 7106 -2048 7164 -2042
rect 7906 -2042 7918 -2040
rect 7952 -2010 7964 -2008
rect 8706 -2008 8764 -2002
rect 8706 -2010 8718 -2008
rect 7952 -2040 8718 -2010
rect 7952 -2042 7964 -2040
rect 7906 -2048 7964 -2042
rect 8706 -2042 8718 -2040
rect 8752 -2010 8764 -2008
rect 9506 -2008 9564 -2002
rect 9506 -2010 9518 -2008
rect 8752 -2040 9518 -2010
rect 8752 -2042 8764 -2040
rect 8706 -2048 8764 -2042
rect 9506 -2042 9518 -2040
rect 9552 -2010 9564 -2008
rect 10306 -2008 10364 -2002
rect 10306 -2010 10318 -2008
rect 9552 -2040 10318 -2010
rect 9552 -2042 9564 -2040
rect 9506 -2048 9564 -2042
rect 10306 -2042 10318 -2040
rect 10352 -2010 10364 -2008
rect 11106 -2008 11164 -2002
rect 11106 -2010 11118 -2008
rect 10352 -2040 11118 -2010
rect 10352 -2042 10364 -2040
rect 10306 -2048 10364 -2042
rect 11106 -2042 11118 -2040
rect 11152 -2010 11164 -2008
rect 11906 -2008 11964 -2002
rect 11906 -2010 11918 -2008
rect 11152 -2040 11918 -2010
rect 11152 -2042 11164 -2040
rect 11106 -2048 11164 -2042
rect 11906 -2042 11918 -2040
rect 11952 -2010 11964 -2008
rect 12706 -2008 12764 -2002
rect 12706 -2010 12718 -2008
rect 11952 -2040 12718 -2010
rect 11952 -2042 11964 -2040
rect 11906 -2048 11964 -2042
rect 12706 -2042 12718 -2040
rect 12752 -2010 12764 -2008
rect 14434 -2010 14440 -1999
rect 12752 -2040 12776 -2010
rect 14400 -2040 14440 -2010
rect 12752 -2042 12764 -2040
rect 12706 -2048 12764 -2042
rect 14434 -2051 14440 -2040
rect 14492 -2051 14498 -1999
rect 14526 -2051 14553 -1999
rect 14605 -2051 14617 -1999
rect 14669 -2051 14697 -1999
rect 14526 -2057 14697 -2051
rect 14725 -1999 14777 -1993
rect 14725 -2057 14777 -2051
rect 14805 -1999 15136 -1993
rect 14805 -2051 14816 -1999
rect 14868 -2008 14880 -1999
rect 14932 -2008 14944 -1999
rect 14996 -2008 15008 -1999
rect 15060 -2008 15072 -1999
rect 14876 -2042 14880 -2008
rect 14868 -2051 14880 -2042
rect 14932 -2051 14944 -2042
rect 14996 -2051 15008 -2042
rect 15060 -2051 15072 -2042
rect 15124 -2051 15136 -1999
rect 14805 -2057 15136 -2051
rect 15206 -1999 15537 -1993
rect 15206 -2051 15217 -1999
rect 15269 -2008 15281 -1999
rect 15333 -2008 15345 -1999
rect 15397 -2008 15409 -1999
rect 15461 -2008 15473 -1999
rect 15461 -2042 15465 -2008
rect 15269 -2051 15281 -2042
rect 15333 -2051 15345 -2042
rect 15397 -2051 15409 -2042
rect 15461 -2051 15473 -2042
rect 15525 -2051 15537 -1999
rect 15206 -2057 15537 -2051
rect 15565 -1999 15617 -1993
rect 15565 -2057 15617 -2051
rect 15645 -1999 15816 -1993
rect 15645 -2051 15672 -1999
rect 15724 -2051 15736 -1999
rect 15788 -2051 15816 -1999
rect 15645 -2057 15816 -2051
rect -65 -2135 12735 -2117
rect -65 -2169 -4 -2135
rect 30 -2169 68 -2135
rect 102 -2169 168 -2135
rect 202 -2169 240 -2135
rect 274 -2169 396 -2135
rect 430 -2169 468 -2135
rect 502 -2169 568 -2135
rect 602 -2169 640 -2135
rect 674 -2169 796 -2135
rect 830 -2169 868 -2135
rect 902 -2169 968 -2135
rect 1002 -2169 1040 -2135
rect 1074 -2169 1196 -2135
rect 1230 -2169 1268 -2135
rect 1302 -2169 1368 -2135
rect 1402 -2169 1440 -2135
rect 1474 -2169 1596 -2135
rect 1630 -2169 1668 -2135
rect 1702 -2169 1768 -2135
rect 1802 -2169 1840 -2135
rect 1874 -2169 1996 -2135
rect 2030 -2169 2068 -2135
rect 2102 -2169 2168 -2135
rect 2202 -2169 2240 -2135
rect 2274 -2169 2396 -2135
rect 2430 -2169 2468 -2135
rect 2502 -2169 2568 -2135
rect 2602 -2169 2640 -2135
rect 2674 -2169 2796 -2135
rect 2830 -2169 2868 -2135
rect 2902 -2169 2968 -2135
rect 3002 -2169 3040 -2135
rect 3074 -2169 3196 -2135
rect 3230 -2169 3268 -2135
rect 3302 -2169 3368 -2135
rect 3402 -2169 3440 -2135
rect 3474 -2169 3596 -2135
rect 3630 -2169 3668 -2135
rect 3702 -2169 3768 -2135
rect 3802 -2169 3840 -2135
rect 3874 -2169 3996 -2135
rect 4030 -2169 4068 -2135
rect 4102 -2169 4168 -2135
rect 4202 -2169 4240 -2135
rect 4274 -2169 4396 -2135
rect 4430 -2169 4468 -2135
rect 4502 -2169 4568 -2135
rect 4602 -2169 4640 -2135
rect 4674 -2169 4796 -2135
rect 4830 -2169 4868 -2135
rect 4902 -2169 4968 -2135
rect 5002 -2169 5040 -2135
rect 5074 -2169 5196 -2135
rect 5230 -2169 5268 -2135
rect 5302 -2169 5368 -2135
rect 5402 -2169 5440 -2135
rect 5474 -2169 5596 -2135
rect 5630 -2169 5668 -2135
rect 5702 -2169 5768 -2135
rect 5802 -2169 5840 -2135
rect 5874 -2169 5996 -2135
rect 6030 -2169 6068 -2135
rect 6102 -2169 6168 -2135
rect 6202 -2169 6240 -2135
rect 6274 -2169 6396 -2135
rect 6430 -2169 6468 -2135
rect 6502 -2169 6568 -2135
rect 6602 -2169 6640 -2135
rect 6674 -2169 6796 -2135
rect 6830 -2169 6868 -2135
rect 6902 -2169 6968 -2135
rect 7002 -2169 7040 -2135
rect 7074 -2169 7196 -2135
rect 7230 -2169 7268 -2135
rect 7302 -2169 7368 -2135
rect 7402 -2169 7440 -2135
rect 7474 -2169 7596 -2135
rect 7630 -2169 7668 -2135
rect 7702 -2169 7768 -2135
rect 7802 -2169 7840 -2135
rect 7874 -2169 7996 -2135
rect 8030 -2169 8068 -2135
rect 8102 -2169 8168 -2135
rect 8202 -2169 8240 -2135
rect 8274 -2169 8396 -2135
rect 8430 -2169 8468 -2135
rect 8502 -2169 8568 -2135
rect 8602 -2169 8640 -2135
rect 8674 -2169 8796 -2135
rect 8830 -2169 8868 -2135
rect 8902 -2169 8968 -2135
rect 9002 -2169 9040 -2135
rect 9074 -2169 9196 -2135
rect 9230 -2169 9268 -2135
rect 9302 -2169 9368 -2135
rect 9402 -2169 9440 -2135
rect 9474 -2169 9596 -2135
rect 9630 -2169 9668 -2135
rect 9702 -2169 9768 -2135
rect 9802 -2169 9840 -2135
rect 9874 -2169 9996 -2135
rect 10030 -2169 10068 -2135
rect 10102 -2169 10168 -2135
rect 10202 -2169 10240 -2135
rect 10274 -2169 10396 -2135
rect 10430 -2169 10468 -2135
rect 10502 -2169 10568 -2135
rect 10602 -2169 10640 -2135
rect 10674 -2169 10796 -2135
rect 10830 -2169 10868 -2135
rect 10902 -2169 10968 -2135
rect 11002 -2169 11040 -2135
rect 11074 -2169 11196 -2135
rect 11230 -2169 11268 -2135
rect 11302 -2169 11368 -2135
rect 11402 -2169 11440 -2135
rect 11474 -2169 11596 -2135
rect 11630 -2169 11668 -2135
rect 11702 -2169 11768 -2135
rect 11802 -2169 11840 -2135
rect 11874 -2169 11996 -2135
rect 12030 -2169 12068 -2135
rect 12102 -2169 12168 -2135
rect 12202 -2169 12240 -2135
rect 12274 -2169 12396 -2135
rect 12430 -2169 12468 -2135
rect 12502 -2169 12568 -2135
rect 12602 -2169 12640 -2135
rect 12674 -2169 12735 -2135
rect -65 -2187 12735 -2169
<< via1 >>
rect 9 4894 61 4903
rect 9 4860 18 4894
rect 18 4860 52 4894
rect 52 4860 61 4894
rect 9 4851 61 4860
rect 9 4753 18 4761
rect 18 4753 52 4761
rect 52 4753 61 4761
rect 9 4709 61 4753
rect 209 4910 261 4919
rect 209 4876 218 4910
rect 218 4876 252 4910
rect 252 4876 261 4910
rect 209 4867 261 4876
rect 9 4613 18 4621
rect 18 4613 52 4621
rect 52 4613 61 4621
rect 9 4569 61 4613
rect 209 4787 261 4831
rect 209 4779 218 4787
rect 218 4779 252 4787
rect 252 4779 261 4787
rect 409 4894 461 4903
rect 409 4860 418 4894
rect 418 4860 452 4894
rect 452 4860 461 4894
rect 409 4851 461 4860
rect 9 4473 18 4481
rect 18 4473 52 4481
rect 52 4473 61 4481
rect 9 4429 61 4473
rect 209 4647 261 4691
rect 209 4639 218 4647
rect 218 4639 252 4647
rect 252 4639 261 4647
rect 409 4753 418 4761
rect 418 4753 452 4761
rect 452 4753 461 4761
rect 409 4709 461 4753
rect 609 4910 661 4919
rect 609 4876 618 4910
rect 618 4876 652 4910
rect 652 4876 661 4910
rect 609 4867 661 4876
rect 9 4333 18 4341
rect 18 4333 52 4341
rect 52 4333 61 4341
rect 9 4289 61 4333
rect 209 4507 261 4551
rect 209 4499 218 4507
rect 218 4499 252 4507
rect 252 4499 261 4507
rect 409 4613 418 4621
rect 418 4613 452 4621
rect 452 4613 461 4621
rect 409 4569 461 4613
rect 609 4787 661 4831
rect 609 4779 618 4787
rect 618 4779 652 4787
rect 652 4779 661 4787
rect 809 4894 861 4903
rect 809 4860 818 4894
rect 818 4860 852 4894
rect 852 4860 861 4894
rect 809 4851 861 4860
rect 9 4193 18 4201
rect 18 4193 52 4201
rect 52 4193 61 4201
rect 9 4149 61 4193
rect 209 4367 261 4411
rect 209 4359 218 4367
rect 218 4359 252 4367
rect 252 4359 261 4367
rect 409 4473 418 4481
rect 418 4473 452 4481
rect 452 4473 461 4481
rect 409 4429 461 4473
rect 609 4647 661 4691
rect 609 4639 618 4647
rect 618 4639 652 4647
rect 652 4639 661 4647
rect 809 4753 818 4761
rect 818 4753 852 4761
rect 852 4753 861 4761
rect 809 4709 861 4753
rect 1009 4910 1061 4919
rect 1009 4876 1018 4910
rect 1018 4876 1052 4910
rect 1052 4876 1061 4910
rect 1009 4867 1061 4876
rect 9 4053 18 4061
rect 18 4053 52 4061
rect 52 4053 61 4061
rect 9 4009 61 4053
rect 209 4227 261 4271
rect 209 4219 218 4227
rect 218 4219 252 4227
rect 252 4219 261 4227
rect 409 4333 418 4341
rect 418 4333 452 4341
rect 452 4333 461 4341
rect 409 4289 461 4333
rect 609 4507 661 4551
rect 609 4499 618 4507
rect 618 4499 652 4507
rect 652 4499 661 4507
rect 809 4613 818 4621
rect 818 4613 852 4621
rect 852 4613 861 4621
rect 809 4569 861 4613
rect 1009 4787 1061 4831
rect 1009 4779 1018 4787
rect 1018 4779 1052 4787
rect 1052 4779 1061 4787
rect 1209 4894 1261 4903
rect 1209 4860 1218 4894
rect 1218 4860 1252 4894
rect 1252 4860 1261 4894
rect 1209 4851 1261 4860
rect 9 3913 18 3921
rect 18 3913 52 3921
rect 52 3913 61 3921
rect 9 3869 61 3913
rect 209 4087 261 4131
rect 209 4079 218 4087
rect 218 4079 252 4087
rect 252 4079 261 4087
rect 409 4193 418 4201
rect 418 4193 452 4201
rect 452 4193 461 4201
rect 409 4149 461 4193
rect 609 4367 661 4411
rect 609 4359 618 4367
rect 618 4359 652 4367
rect 652 4359 661 4367
rect 809 4473 818 4481
rect 818 4473 852 4481
rect 852 4473 861 4481
rect 809 4429 861 4473
rect 1009 4647 1061 4691
rect 1009 4639 1018 4647
rect 1018 4639 1052 4647
rect 1052 4639 1061 4647
rect 1209 4753 1218 4761
rect 1218 4753 1252 4761
rect 1252 4753 1261 4761
rect 1209 4709 1261 4753
rect 1409 4910 1461 4919
rect 1409 4876 1418 4910
rect 1418 4876 1452 4910
rect 1452 4876 1461 4910
rect 1409 4867 1461 4876
rect 9 3773 18 3781
rect 18 3773 52 3781
rect 52 3773 61 3781
rect 9 3729 61 3773
rect 209 3947 261 3991
rect 209 3939 218 3947
rect 218 3939 252 3947
rect 252 3939 261 3947
rect 409 4053 418 4061
rect 418 4053 452 4061
rect 452 4053 461 4061
rect 409 4009 461 4053
rect 609 4227 661 4271
rect 609 4219 618 4227
rect 618 4219 652 4227
rect 652 4219 661 4227
rect 809 4333 818 4341
rect 818 4333 852 4341
rect 852 4333 861 4341
rect 809 4289 861 4333
rect 1009 4507 1061 4551
rect 1009 4499 1018 4507
rect 1018 4499 1052 4507
rect 1052 4499 1061 4507
rect 1209 4613 1218 4621
rect 1218 4613 1252 4621
rect 1252 4613 1261 4621
rect 1209 4569 1261 4613
rect 1409 4787 1461 4831
rect 1409 4779 1418 4787
rect 1418 4779 1452 4787
rect 1452 4779 1461 4787
rect 1609 4894 1661 4903
rect 1609 4860 1618 4894
rect 1618 4860 1652 4894
rect 1652 4860 1661 4894
rect 1609 4851 1661 4860
rect 9 3684 61 3693
rect 9 3650 18 3684
rect 18 3650 52 3684
rect 52 3650 61 3684
rect 9 3641 61 3650
rect 9 3543 18 3551
rect 18 3543 52 3551
rect 52 3543 61 3551
rect 9 3499 61 3543
rect 209 3807 261 3851
rect 209 3799 218 3807
rect 218 3799 252 3807
rect 252 3799 261 3807
rect 409 3913 418 3921
rect 418 3913 452 3921
rect 452 3913 461 3921
rect 409 3869 461 3913
rect 609 4087 661 4131
rect 609 4079 618 4087
rect 618 4079 652 4087
rect 652 4079 661 4087
rect 809 4193 818 4201
rect 818 4193 852 4201
rect 852 4193 861 4201
rect 809 4149 861 4193
rect 1009 4367 1061 4411
rect 1009 4359 1018 4367
rect 1018 4359 1052 4367
rect 1052 4359 1061 4367
rect 1209 4473 1218 4481
rect 1218 4473 1252 4481
rect 1252 4473 1261 4481
rect 1209 4429 1261 4473
rect 1409 4647 1461 4691
rect 1409 4639 1418 4647
rect 1418 4639 1452 4647
rect 1452 4639 1461 4647
rect 1609 4753 1618 4761
rect 1618 4753 1652 4761
rect 1652 4753 1661 4761
rect 1609 4709 1661 4753
rect 1809 4910 1861 4919
rect 1809 4876 1818 4910
rect 1818 4876 1852 4910
rect 1852 4876 1861 4910
rect 1809 4867 1861 4876
rect 209 3700 261 3709
rect 209 3666 218 3700
rect 218 3666 252 3700
rect 252 3666 261 3700
rect 209 3657 261 3666
rect 9 3403 18 3411
rect 18 3403 52 3411
rect 52 3403 61 3411
rect 9 3359 61 3403
rect 209 3577 261 3621
rect 209 3569 218 3577
rect 218 3569 252 3577
rect 252 3569 261 3577
rect 409 3773 418 3781
rect 418 3773 452 3781
rect 452 3773 461 3781
rect 409 3729 461 3773
rect 609 3947 661 3991
rect 609 3939 618 3947
rect 618 3939 652 3947
rect 652 3939 661 3947
rect 809 4053 818 4061
rect 818 4053 852 4061
rect 852 4053 861 4061
rect 809 4009 861 4053
rect 1009 4227 1061 4271
rect 1009 4219 1018 4227
rect 1018 4219 1052 4227
rect 1052 4219 1061 4227
rect 1209 4333 1218 4341
rect 1218 4333 1252 4341
rect 1252 4333 1261 4341
rect 1209 4289 1261 4333
rect 1409 4507 1461 4551
rect 1409 4499 1418 4507
rect 1418 4499 1452 4507
rect 1452 4499 1461 4507
rect 1609 4613 1618 4621
rect 1618 4613 1652 4621
rect 1652 4613 1661 4621
rect 1609 4569 1661 4613
rect 1809 4787 1861 4831
rect 1809 4779 1818 4787
rect 1818 4779 1852 4787
rect 1852 4779 1861 4787
rect 2009 4894 2061 4903
rect 2009 4860 2018 4894
rect 2018 4860 2052 4894
rect 2052 4860 2061 4894
rect 2009 4851 2061 4860
rect 409 3684 461 3693
rect 409 3650 418 3684
rect 418 3650 452 3684
rect 452 3650 461 3684
rect 409 3641 461 3650
rect 9 3263 18 3271
rect 18 3263 52 3271
rect 52 3263 61 3271
rect 9 3219 61 3263
rect 209 3437 261 3481
rect 209 3429 218 3437
rect 218 3429 252 3437
rect 252 3429 261 3437
rect 409 3543 418 3551
rect 418 3543 452 3551
rect 452 3543 461 3551
rect 409 3499 461 3543
rect 609 3807 661 3851
rect 609 3799 618 3807
rect 618 3799 652 3807
rect 652 3799 661 3807
rect 809 3913 818 3921
rect 818 3913 852 3921
rect 852 3913 861 3921
rect 809 3869 861 3913
rect 1009 4087 1061 4131
rect 1009 4079 1018 4087
rect 1018 4079 1052 4087
rect 1052 4079 1061 4087
rect 1209 4193 1218 4201
rect 1218 4193 1252 4201
rect 1252 4193 1261 4201
rect 1209 4149 1261 4193
rect 1409 4367 1461 4411
rect 1409 4359 1418 4367
rect 1418 4359 1452 4367
rect 1452 4359 1461 4367
rect 1609 4473 1618 4481
rect 1618 4473 1652 4481
rect 1652 4473 1661 4481
rect 1609 4429 1661 4473
rect 1809 4647 1861 4691
rect 1809 4639 1818 4647
rect 1818 4639 1852 4647
rect 1852 4639 1861 4647
rect 2009 4753 2018 4761
rect 2018 4753 2052 4761
rect 2052 4753 2061 4761
rect 2009 4709 2061 4753
rect 2209 4910 2261 4919
rect 2209 4876 2218 4910
rect 2218 4876 2252 4910
rect 2252 4876 2261 4910
rect 2209 4867 2261 4876
rect 609 3700 661 3709
rect 609 3666 618 3700
rect 618 3666 652 3700
rect 652 3666 661 3700
rect 609 3657 661 3666
rect 9 3123 18 3131
rect 18 3123 52 3131
rect 52 3123 61 3131
rect 9 3079 61 3123
rect 209 3297 261 3341
rect 209 3289 218 3297
rect 218 3289 252 3297
rect 252 3289 261 3297
rect 409 3403 418 3411
rect 418 3403 452 3411
rect 452 3403 461 3411
rect 409 3359 461 3403
rect 609 3577 661 3621
rect 609 3569 618 3577
rect 618 3569 652 3577
rect 652 3569 661 3577
rect 809 3773 818 3781
rect 818 3773 852 3781
rect 852 3773 861 3781
rect 809 3729 861 3773
rect 1009 3947 1061 3991
rect 1009 3939 1018 3947
rect 1018 3939 1052 3947
rect 1052 3939 1061 3947
rect 1209 4053 1218 4061
rect 1218 4053 1252 4061
rect 1252 4053 1261 4061
rect 1209 4009 1261 4053
rect 1409 4227 1461 4271
rect 1409 4219 1418 4227
rect 1418 4219 1452 4227
rect 1452 4219 1461 4227
rect 1609 4333 1618 4341
rect 1618 4333 1652 4341
rect 1652 4333 1661 4341
rect 1609 4289 1661 4333
rect 1809 4507 1861 4551
rect 1809 4499 1818 4507
rect 1818 4499 1852 4507
rect 1852 4499 1861 4507
rect 2009 4613 2018 4621
rect 2018 4613 2052 4621
rect 2052 4613 2061 4621
rect 2009 4569 2061 4613
rect 2209 4787 2261 4831
rect 2209 4779 2218 4787
rect 2218 4779 2252 4787
rect 2252 4779 2261 4787
rect 2409 4894 2461 4903
rect 2409 4860 2418 4894
rect 2418 4860 2452 4894
rect 2452 4860 2461 4894
rect 2409 4851 2461 4860
rect 809 3684 861 3693
rect 809 3650 818 3684
rect 818 3650 852 3684
rect 852 3650 861 3684
rect 809 3641 861 3650
rect 9 2983 18 2991
rect 18 2983 52 2991
rect 52 2983 61 2991
rect 9 2939 61 2983
rect 209 3157 261 3201
rect 209 3149 218 3157
rect 218 3149 252 3157
rect 252 3149 261 3157
rect 409 3263 418 3271
rect 418 3263 452 3271
rect 452 3263 461 3271
rect 409 3219 461 3263
rect 609 3437 661 3481
rect 609 3429 618 3437
rect 618 3429 652 3437
rect 652 3429 661 3437
rect 809 3543 818 3551
rect 818 3543 852 3551
rect 852 3543 861 3551
rect 809 3499 861 3543
rect 1009 3807 1061 3851
rect 1009 3799 1018 3807
rect 1018 3799 1052 3807
rect 1052 3799 1061 3807
rect 1209 3913 1218 3921
rect 1218 3913 1252 3921
rect 1252 3913 1261 3921
rect 1209 3869 1261 3913
rect 1409 4087 1461 4131
rect 1409 4079 1418 4087
rect 1418 4079 1452 4087
rect 1452 4079 1461 4087
rect 1609 4193 1618 4201
rect 1618 4193 1652 4201
rect 1652 4193 1661 4201
rect 1609 4149 1661 4193
rect 1809 4367 1861 4411
rect 1809 4359 1818 4367
rect 1818 4359 1852 4367
rect 1852 4359 1861 4367
rect 2009 4473 2018 4481
rect 2018 4473 2052 4481
rect 2052 4473 2061 4481
rect 2009 4429 2061 4473
rect 2209 4647 2261 4691
rect 2209 4639 2218 4647
rect 2218 4639 2252 4647
rect 2252 4639 2261 4647
rect 2409 4753 2418 4761
rect 2418 4753 2452 4761
rect 2452 4753 2461 4761
rect 2409 4709 2461 4753
rect 2609 4910 2661 4919
rect 2609 4876 2618 4910
rect 2618 4876 2652 4910
rect 2652 4876 2661 4910
rect 2609 4867 2661 4876
rect 1009 3700 1061 3709
rect 1009 3666 1018 3700
rect 1018 3666 1052 3700
rect 1052 3666 1061 3700
rect 1009 3657 1061 3666
rect 9 2843 18 2851
rect 18 2843 52 2851
rect 52 2843 61 2851
rect 9 2799 61 2843
rect 209 3017 261 3061
rect 209 3009 218 3017
rect 218 3009 252 3017
rect 252 3009 261 3017
rect 409 3123 418 3131
rect 418 3123 452 3131
rect 452 3123 461 3131
rect 409 3079 461 3123
rect 609 3297 661 3341
rect 609 3289 618 3297
rect 618 3289 652 3297
rect 652 3289 661 3297
rect 809 3403 818 3411
rect 818 3403 852 3411
rect 852 3403 861 3411
rect 809 3359 861 3403
rect 1009 3577 1061 3621
rect 1009 3569 1018 3577
rect 1018 3569 1052 3577
rect 1052 3569 1061 3577
rect 1209 3773 1218 3781
rect 1218 3773 1252 3781
rect 1252 3773 1261 3781
rect 1209 3729 1261 3773
rect 1409 3947 1461 3991
rect 1409 3939 1418 3947
rect 1418 3939 1452 3947
rect 1452 3939 1461 3947
rect 1609 4053 1618 4061
rect 1618 4053 1652 4061
rect 1652 4053 1661 4061
rect 1609 4009 1661 4053
rect 1809 4227 1861 4271
rect 1809 4219 1818 4227
rect 1818 4219 1852 4227
rect 1852 4219 1861 4227
rect 2009 4333 2018 4341
rect 2018 4333 2052 4341
rect 2052 4333 2061 4341
rect 2009 4289 2061 4333
rect 2209 4507 2261 4551
rect 2209 4499 2218 4507
rect 2218 4499 2252 4507
rect 2252 4499 2261 4507
rect 2409 4613 2418 4621
rect 2418 4613 2452 4621
rect 2452 4613 2461 4621
rect 2409 4569 2461 4613
rect 2609 4787 2661 4831
rect 2609 4779 2618 4787
rect 2618 4779 2652 4787
rect 2652 4779 2661 4787
rect 2809 4894 2861 4903
rect 2809 4860 2818 4894
rect 2818 4860 2852 4894
rect 2852 4860 2861 4894
rect 2809 4851 2861 4860
rect 1209 3684 1261 3693
rect 1209 3650 1218 3684
rect 1218 3650 1252 3684
rect 1252 3650 1261 3684
rect 1209 3641 1261 3650
rect 9 2703 18 2711
rect 18 2703 52 2711
rect 52 2703 61 2711
rect 9 2659 61 2703
rect 209 2877 261 2921
rect 209 2869 218 2877
rect 218 2869 252 2877
rect 252 2869 261 2877
rect 409 2983 418 2991
rect 418 2983 452 2991
rect 452 2983 461 2991
rect 409 2939 461 2983
rect 609 3157 661 3201
rect 609 3149 618 3157
rect 618 3149 652 3157
rect 652 3149 661 3157
rect 809 3263 818 3271
rect 818 3263 852 3271
rect 852 3263 861 3271
rect 809 3219 861 3263
rect 1009 3437 1061 3481
rect 1009 3429 1018 3437
rect 1018 3429 1052 3437
rect 1052 3429 1061 3437
rect 1209 3543 1218 3551
rect 1218 3543 1252 3551
rect 1252 3543 1261 3551
rect 1209 3499 1261 3543
rect 1409 3807 1461 3851
rect 1409 3799 1418 3807
rect 1418 3799 1452 3807
rect 1452 3799 1461 3807
rect 1609 3913 1618 3921
rect 1618 3913 1652 3921
rect 1652 3913 1661 3921
rect 1609 3869 1661 3913
rect 1809 4087 1861 4131
rect 1809 4079 1818 4087
rect 1818 4079 1852 4087
rect 1852 4079 1861 4087
rect 2009 4193 2018 4201
rect 2018 4193 2052 4201
rect 2052 4193 2061 4201
rect 2009 4149 2061 4193
rect 2209 4367 2261 4411
rect 2209 4359 2218 4367
rect 2218 4359 2252 4367
rect 2252 4359 2261 4367
rect 2409 4473 2418 4481
rect 2418 4473 2452 4481
rect 2452 4473 2461 4481
rect 2409 4429 2461 4473
rect 2609 4647 2661 4691
rect 2609 4639 2618 4647
rect 2618 4639 2652 4647
rect 2652 4639 2661 4647
rect 2809 4753 2818 4761
rect 2818 4753 2852 4761
rect 2852 4753 2861 4761
rect 2809 4709 2861 4753
rect 3009 4910 3061 4919
rect 3009 4876 3018 4910
rect 3018 4876 3052 4910
rect 3052 4876 3061 4910
rect 3009 4867 3061 4876
rect 1409 3700 1461 3709
rect 1409 3666 1418 3700
rect 1418 3666 1452 3700
rect 1452 3666 1461 3700
rect 1409 3657 1461 3666
rect 9 2563 18 2571
rect 18 2563 52 2571
rect 52 2563 61 2571
rect 9 2519 61 2563
rect 209 2737 261 2781
rect 209 2729 218 2737
rect 218 2729 252 2737
rect 252 2729 261 2737
rect 409 2843 418 2851
rect 418 2843 452 2851
rect 452 2843 461 2851
rect 409 2799 461 2843
rect 609 3017 661 3061
rect 609 3009 618 3017
rect 618 3009 652 3017
rect 652 3009 661 3017
rect 809 3123 818 3131
rect 818 3123 852 3131
rect 852 3123 861 3131
rect 809 3079 861 3123
rect 1009 3297 1061 3341
rect 1009 3289 1018 3297
rect 1018 3289 1052 3297
rect 1052 3289 1061 3297
rect 1209 3403 1218 3411
rect 1218 3403 1252 3411
rect 1252 3403 1261 3411
rect 1209 3359 1261 3403
rect 1409 3577 1461 3621
rect 1409 3569 1418 3577
rect 1418 3569 1452 3577
rect 1452 3569 1461 3577
rect 1609 3773 1618 3781
rect 1618 3773 1652 3781
rect 1652 3773 1661 3781
rect 1609 3729 1661 3773
rect 1809 3947 1861 3991
rect 1809 3939 1818 3947
rect 1818 3939 1852 3947
rect 1852 3939 1861 3947
rect 2009 4053 2018 4061
rect 2018 4053 2052 4061
rect 2052 4053 2061 4061
rect 2009 4009 2061 4053
rect 2209 4227 2261 4271
rect 2209 4219 2218 4227
rect 2218 4219 2252 4227
rect 2252 4219 2261 4227
rect 2409 4333 2418 4341
rect 2418 4333 2452 4341
rect 2452 4333 2461 4341
rect 2409 4289 2461 4333
rect 2609 4507 2661 4551
rect 2609 4499 2618 4507
rect 2618 4499 2652 4507
rect 2652 4499 2661 4507
rect 2809 4613 2818 4621
rect 2818 4613 2852 4621
rect 2852 4613 2861 4621
rect 2809 4569 2861 4613
rect 3009 4787 3061 4831
rect 3009 4779 3018 4787
rect 3018 4779 3052 4787
rect 3052 4779 3061 4787
rect 3209 4894 3261 4903
rect 3209 4860 3218 4894
rect 3218 4860 3252 4894
rect 3252 4860 3261 4894
rect 3209 4851 3261 4860
rect 1609 3684 1661 3693
rect 1609 3650 1618 3684
rect 1618 3650 1652 3684
rect 1652 3650 1661 3684
rect 1609 3641 1661 3650
rect 9 2474 61 2483
rect 9 2440 18 2474
rect 18 2440 52 2474
rect 52 2440 61 2474
rect 9 2431 61 2440
rect 9 2333 18 2341
rect 18 2333 52 2341
rect 52 2333 61 2341
rect 9 2289 61 2333
rect 209 2597 261 2641
rect 209 2589 218 2597
rect 218 2589 252 2597
rect 252 2589 261 2597
rect 409 2703 418 2711
rect 418 2703 452 2711
rect 452 2703 461 2711
rect 409 2659 461 2703
rect 609 2877 661 2921
rect 609 2869 618 2877
rect 618 2869 652 2877
rect 652 2869 661 2877
rect 809 2983 818 2991
rect 818 2983 852 2991
rect 852 2983 861 2991
rect 809 2939 861 2983
rect 1009 3157 1061 3201
rect 1009 3149 1018 3157
rect 1018 3149 1052 3157
rect 1052 3149 1061 3157
rect 1209 3263 1218 3271
rect 1218 3263 1252 3271
rect 1252 3263 1261 3271
rect 1209 3219 1261 3263
rect 1409 3437 1461 3481
rect 1409 3429 1418 3437
rect 1418 3429 1452 3437
rect 1452 3429 1461 3437
rect 1609 3543 1618 3551
rect 1618 3543 1652 3551
rect 1652 3543 1661 3551
rect 1609 3499 1661 3543
rect 1809 3807 1861 3851
rect 1809 3799 1818 3807
rect 1818 3799 1852 3807
rect 1852 3799 1861 3807
rect 2009 3913 2018 3921
rect 2018 3913 2052 3921
rect 2052 3913 2061 3921
rect 2009 3869 2061 3913
rect 2209 4087 2261 4131
rect 2209 4079 2218 4087
rect 2218 4079 2252 4087
rect 2252 4079 2261 4087
rect 2409 4193 2418 4201
rect 2418 4193 2452 4201
rect 2452 4193 2461 4201
rect 2409 4149 2461 4193
rect 2609 4367 2661 4411
rect 2609 4359 2618 4367
rect 2618 4359 2652 4367
rect 2652 4359 2661 4367
rect 2809 4473 2818 4481
rect 2818 4473 2852 4481
rect 2852 4473 2861 4481
rect 2809 4429 2861 4473
rect 3009 4647 3061 4691
rect 3009 4639 3018 4647
rect 3018 4639 3052 4647
rect 3052 4639 3061 4647
rect 3209 4753 3218 4761
rect 3218 4753 3252 4761
rect 3252 4753 3261 4761
rect 3209 4709 3261 4753
rect 3409 4910 3461 4919
rect 3409 4876 3418 4910
rect 3418 4876 3452 4910
rect 3452 4876 3461 4910
rect 3409 4867 3461 4876
rect 1809 3700 1861 3709
rect 1809 3666 1818 3700
rect 1818 3666 1852 3700
rect 1852 3666 1861 3700
rect 1809 3657 1861 3666
rect 209 2490 261 2499
rect 209 2456 218 2490
rect 218 2456 252 2490
rect 252 2456 261 2490
rect 209 2447 261 2456
rect 9 2193 18 2201
rect 18 2193 52 2201
rect 52 2193 61 2201
rect 9 2149 61 2193
rect 209 2367 261 2411
rect 209 2359 218 2367
rect 218 2359 252 2367
rect 252 2359 261 2367
rect 409 2563 418 2571
rect 418 2563 452 2571
rect 452 2563 461 2571
rect 409 2519 461 2563
rect 609 2737 661 2781
rect 609 2729 618 2737
rect 618 2729 652 2737
rect 652 2729 661 2737
rect 809 2843 818 2851
rect 818 2843 852 2851
rect 852 2843 861 2851
rect 809 2799 861 2843
rect 1009 3017 1061 3061
rect 1009 3009 1018 3017
rect 1018 3009 1052 3017
rect 1052 3009 1061 3017
rect 1209 3123 1218 3131
rect 1218 3123 1252 3131
rect 1252 3123 1261 3131
rect 1209 3079 1261 3123
rect 1409 3297 1461 3341
rect 1409 3289 1418 3297
rect 1418 3289 1452 3297
rect 1452 3289 1461 3297
rect 1609 3403 1618 3411
rect 1618 3403 1652 3411
rect 1652 3403 1661 3411
rect 1609 3359 1661 3403
rect 1809 3577 1861 3621
rect 1809 3569 1818 3577
rect 1818 3569 1852 3577
rect 1852 3569 1861 3577
rect 2009 3773 2018 3781
rect 2018 3773 2052 3781
rect 2052 3773 2061 3781
rect 2009 3729 2061 3773
rect 2209 3947 2261 3991
rect 2209 3939 2218 3947
rect 2218 3939 2252 3947
rect 2252 3939 2261 3947
rect 2409 4053 2418 4061
rect 2418 4053 2452 4061
rect 2452 4053 2461 4061
rect 2409 4009 2461 4053
rect 2609 4227 2661 4271
rect 2609 4219 2618 4227
rect 2618 4219 2652 4227
rect 2652 4219 2661 4227
rect 2809 4333 2818 4341
rect 2818 4333 2852 4341
rect 2852 4333 2861 4341
rect 2809 4289 2861 4333
rect 3009 4507 3061 4551
rect 3009 4499 3018 4507
rect 3018 4499 3052 4507
rect 3052 4499 3061 4507
rect 3209 4613 3218 4621
rect 3218 4613 3252 4621
rect 3252 4613 3261 4621
rect 3209 4569 3261 4613
rect 3409 4787 3461 4831
rect 3409 4779 3418 4787
rect 3418 4779 3452 4787
rect 3452 4779 3461 4787
rect 3609 4894 3661 4903
rect 3609 4860 3618 4894
rect 3618 4860 3652 4894
rect 3652 4860 3661 4894
rect 3609 4851 3661 4860
rect 2009 3684 2061 3693
rect 2009 3650 2018 3684
rect 2018 3650 2052 3684
rect 2052 3650 2061 3684
rect 2009 3641 2061 3650
rect 409 2474 461 2483
rect 409 2440 418 2474
rect 418 2440 452 2474
rect 452 2440 461 2474
rect 409 2431 461 2440
rect 9 2053 18 2061
rect 18 2053 52 2061
rect 52 2053 61 2061
rect 9 2009 61 2053
rect 209 2227 261 2271
rect 209 2219 218 2227
rect 218 2219 252 2227
rect 252 2219 261 2227
rect 409 2333 418 2341
rect 418 2333 452 2341
rect 452 2333 461 2341
rect 409 2289 461 2333
rect 609 2597 661 2641
rect 609 2589 618 2597
rect 618 2589 652 2597
rect 652 2589 661 2597
rect 809 2703 818 2711
rect 818 2703 852 2711
rect 852 2703 861 2711
rect 809 2659 861 2703
rect 1009 2877 1061 2921
rect 1009 2869 1018 2877
rect 1018 2869 1052 2877
rect 1052 2869 1061 2877
rect 1209 2983 1218 2991
rect 1218 2983 1252 2991
rect 1252 2983 1261 2991
rect 1209 2939 1261 2983
rect 1409 3157 1461 3201
rect 1409 3149 1418 3157
rect 1418 3149 1452 3157
rect 1452 3149 1461 3157
rect 1609 3263 1618 3271
rect 1618 3263 1652 3271
rect 1652 3263 1661 3271
rect 1609 3219 1661 3263
rect 1809 3437 1861 3481
rect 1809 3429 1818 3437
rect 1818 3429 1852 3437
rect 1852 3429 1861 3437
rect 2009 3543 2018 3551
rect 2018 3543 2052 3551
rect 2052 3543 2061 3551
rect 2009 3499 2061 3543
rect 2209 3807 2261 3851
rect 2209 3799 2218 3807
rect 2218 3799 2252 3807
rect 2252 3799 2261 3807
rect 2409 3913 2418 3921
rect 2418 3913 2452 3921
rect 2452 3913 2461 3921
rect 2409 3869 2461 3913
rect 2609 4087 2661 4131
rect 2609 4079 2618 4087
rect 2618 4079 2652 4087
rect 2652 4079 2661 4087
rect 2809 4193 2818 4201
rect 2818 4193 2852 4201
rect 2852 4193 2861 4201
rect 2809 4149 2861 4193
rect 3009 4367 3061 4411
rect 3009 4359 3018 4367
rect 3018 4359 3052 4367
rect 3052 4359 3061 4367
rect 3209 4473 3218 4481
rect 3218 4473 3252 4481
rect 3252 4473 3261 4481
rect 3209 4429 3261 4473
rect 3409 4647 3461 4691
rect 3409 4639 3418 4647
rect 3418 4639 3452 4647
rect 3452 4639 3461 4647
rect 3609 4753 3618 4761
rect 3618 4753 3652 4761
rect 3652 4753 3661 4761
rect 3609 4709 3661 4753
rect 3809 4910 3861 4919
rect 3809 4876 3818 4910
rect 3818 4876 3852 4910
rect 3852 4876 3861 4910
rect 3809 4867 3861 4876
rect 2209 3700 2261 3709
rect 2209 3666 2218 3700
rect 2218 3666 2252 3700
rect 2252 3666 2261 3700
rect 2209 3657 2261 3666
rect 609 2490 661 2499
rect 609 2456 618 2490
rect 618 2456 652 2490
rect 652 2456 661 2490
rect 609 2447 661 2456
rect 9 1913 18 1921
rect 18 1913 52 1921
rect 52 1913 61 1921
rect 9 1869 61 1913
rect 209 2087 261 2131
rect 209 2079 218 2087
rect 218 2079 252 2087
rect 252 2079 261 2087
rect 409 2193 418 2201
rect 418 2193 452 2201
rect 452 2193 461 2201
rect 409 2149 461 2193
rect 609 2367 661 2411
rect 609 2359 618 2367
rect 618 2359 652 2367
rect 652 2359 661 2367
rect 809 2563 818 2571
rect 818 2563 852 2571
rect 852 2563 861 2571
rect 809 2519 861 2563
rect 1009 2737 1061 2781
rect 1009 2729 1018 2737
rect 1018 2729 1052 2737
rect 1052 2729 1061 2737
rect 1209 2843 1218 2851
rect 1218 2843 1252 2851
rect 1252 2843 1261 2851
rect 1209 2799 1261 2843
rect 1409 3017 1461 3061
rect 1409 3009 1418 3017
rect 1418 3009 1452 3017
rect 1452 3009 1461 3017
rect 1609 3123 1618 3131
rect 1618 3123 1652 3131
rect 1652 3123 1661 3131
rect 1609 3079 1661 3123
rect 1809 3297 1861 3341
rect 1809 3289 1818 3297
rect 1818 3289 1852 3297
rect 1852 3289 1861 3297
rect 2009 3403 2018 3411
rect 2018 3403 2052 3411
rect 2052 3403 2061 3411
rect 2009 3359 2061 3403
rect 2209 3577 2261 3621
rect 2209 3569 2218 3577
rect 2218 3569 2252 3577
rect 2252 3569 2261 3577
rect 2409 3773 2418 3781
rect 2418 3773 2452 3781
rect 2452 3773 2461 3781
rect 2409 3729 2461 3773
rect 2609 3947 2661 3991
rect 2609 3939 2618 3947
rect 2618 3939 2652 3947
rect 2652 3939 2661 3947
rect 2809 4053 2818 4061
rect 2818 4053 2852 4061
rect 2852 4053 2861 4061
rect 2809 4009 2861 4053
rect 3009 4227 3061 4271
rect 3009 4219 3018 4227
rect 3018 4219 3052 4227
rect 3052 4219 3061 4227
rect 3209 4333 3218 4341
rect 3218 4333 3252 4341
rect 3252 4333 3261 4341
rect 3209 4289 3261 4333
rect 3409 4507 3461 4551
rect 3409 4499 3418 4507
rect 3418 4499 3452 4507
rect 3452 4499 3461 4507
rect 3609 4613 3618 4621
rect 3618 4613 3652 4621
rect 3652 4613 3661 4621
rect 3609 4569 3661 4613
rect 3809 4787 3861 4831
rect 3809 4779 3818 4787
rect 3818 4779 3852 4787
rect 3852 4779 3861 4787
rect 4009 4894 4061 4903
rect 4009 4860 4018 4894
rect 4018 4860 4052 4894
rect 4052 4860 4061 4894
rect 4009 4851 4061 4860
rect 2409 3684 2461 3693
rect 2409 3650 2418 3684
rect 2418 3650 2452 3684
rect 2452 3650 2461 3684
rect 2409 3641 2461 3650
rect 809 2474 861 2483
rect 809 2440 818 2474
rect 818 2440 852 2474
rect 852 2440 861 2474
rect 809 2431 861 2440
rect 9 1773 18 1781
rect 18 1773 52 1781
rect 52 1773 61 1781
rect 9 1729 61 1773
rect 209 1947 261 1991
rect 209 1939 218 1947
rect 218 1939 252 1947
rect 252 1939 261 1947
rect 409 2053 418 2061
rect 418 2053 452 2061
rect 452 2053 461 2061
rect 409 2009 461 2053
rect 609 2227 661 2271
rect 609 2219 618 2227
rect 618 2219 652 2227
rect 652 2219 661 2227
rect 809 2333 818 2341
rect 818 2333 852 2341
rect 852 2333 861 2341
rect 809 2289 861 2333
rect 1009 2597 1061 2641
rect 1009 2589 1018 2597
rect 1018 2589 1052 2597
rect 1052 2589 1061 2597
rect 1209 2703 1218 2711
rect 1218 2703 1252 2711
rect 1252 2703 1261 2711
rect 1209 2659 1261 2703
rect 1409 2877 1461 2921
rect 1409 2869 1418 2877
rect 1418 2869 1452 2877
rect 1452 2869 1461 2877
rect 1609 2983 1618 2991
rect 1618 2983 1652 2991
rect 1652 2983 1661 2991
rect 1609 2939 1661 2983
rect 1809 3157 1861 3201
rect 1809 3149 1818 3157
rect 1818 3149 1852 3157
rect 1852 3149 1861 3157
rect 2009 3263 2018 3271
rect 2018 3263 2052 3271
rect 2052 3263 2061 3271
rect 2009 3219 2061 3263
rect 2209 3437 2261 3481
rect 2209 3429 2218 3437
rect 2218 3429 2252 3437
rect 2252 3429 2261 3437
rect 2409 3543 2418 3551
rect 2418 3543 2452 3551
rect 2452 3543 2461 3551
rect 2409 3499 2461 3543
rect 2609 3807 2661 3851
rect 2609 3799 2618 3807
rect 2618 3799 2652 3807
rect 2652 3799 2661 3807
rect 2809 3913 2818 3921
rect 2818 3913 2852 3921
rect 2852 3913 2861 3921
rect 2809 3869 2861 3913
rect 3009 4087 3061 4131
rect 3009 4079 3018 4087
rect 3018 4079 3052 4087
rect 3052 4079 3061 4087
rect 3209 4193 3218 4201
rect 3218 4193 3252 4201
rect 3252 4193 3261 4201
rect 3209 4149 3261 4193
rect 3409 4367 3461 4411
rect 3409 4359 3418 4367
rect 3418 4359 3452 4367
rect 3452 4359 3461 4367
rect 3609 4473 3618 4481
rect 3618 4473 3652 4481
rect 3652 4473 3661 4481
rect 3609 4429 3661 4473
rect 3809 4647 3861 4691
rect 3809 4639 3818 4647
rect 3818 4639 3852 4647
rect 3852 4639 3861 4647
rect 4009 4753 4018 4761
rect 4018 4753 4052 4761
rect 4052 4753 4061 4761
rect 4009 4709 4061 4753
rect 4209 4910 4261 4919
rect 4209 4876 4218 4910
rect 4218 4876 4252 4910
rect 4252 4876 4261 4910
rect 4209 4867 4261 4876
rect 2609 3700 2661 3709
rect 2609 3666 2618 3700
rect 2618 3666 2652 3700
rect 2652 3666 2661 3700
rect 2609 3657 2661 3666
rect 1009 2490 1061 2499
rect 1009 2456 1018 2490
rect 1018 2456 1052 2490
rect 1052 2456 1061 2490
rect 1009 2447 1061 2456
rect 9 1633 18 1641
rect 18 1633 52 1641
rect 52 1633 61 1641
rect 9 1589 61 1633
rect 209 1807 261 1851
rect 209 1799 218 1807
rect 218 1799 252 1807
rect 252 1799 261 1807
rect 409 1913 418 1921
rect 418 1913 452 1921
rect 452 1913 461 1921
rect 409 1869 461 1913
rect 609 2087 661 2131
rect 609 2079 618 2087
rect 618 2079 652 2087
rect 652 2079 661 2087
rect 809 2193 818 2201
rect 818 2193 852 2201
rect 852 2193 861 2201
rect 809 2149 861 2193
rect 1009 2367 1061 2411
rect 1009 2359 1018 2367
rect 1018 2359 1052 2367
rect 1052 2359 1061 2367
rect 1209 2563 1218 2571
rect 1218 2563 1252 2571
rect 1252 2563 1261 2571
rect 1209 2519 1261 2563
rect 1409 2737 1461 2781
rect 1409 2729 1418 2737
rect 1418 2729 1452 2737
rect 1452 2729 1461 2737
rect 1609 2843 1618 2851
rect 1618 2843 1652 2851
rect 1652 2843 1661 2851
rect 1609 2799 1661 2843
rect 1809 3017 1861 3061
rect 1809 3009 1818 3017
rect 1818 3009 1852 3017
rect 1852 3009 1861 3017
rect 2009 3123 2018 3131
rect 2018 3123 2052 3131
rect 2052 3123 2061 3131
rect 2009 3079 2061 3123
rect 2209 3297 2261 3341
rect 2209 3289 2218 3297
rect 2218 3289 2252 3297
rect 2252 3289 2261 3297
rect 2409 3403 2418 3411
rect 2418 3403 2452 3411
rect 2452 3403 2461 3411
rect 2409 3359 2461 3403
rect 2609 3577 2661 3621
rect 2609 3569 2618 3577
rect 2618 3569 2652 3577
rect 2652 3569 2661 3577
rect 2809 3773 2818 3781
rect 2818 3773 2852 3781
rect 2852 3773 2861 3781
rect 2809 3729 2861 3773
rect 3009 3947 3061 3991
rect 3009 3939 3018 3947
rect 3018 3939 3052 3947
rect 3052 3939 3061 3947
rect 3209 4053 3218 4061
rect 3218 4053 3252 4061
rect 3252 4053 3261 4061
rect 3209 4009 3261 4053
rect 3409 4227 3461 4271
rect 3409 4219 3418 4227
rect 3418 4219 3452 4227
rect 3452 4219 3461 4227
rect 3609 4333 3618 4341
rect 3618 4333 3652 4341
rect 3652 4333 3661 4341
rect 3609 4289 3661 4333
rect 3809 4507 3861 4551
rect 3809 4499 3818 4507
rect 3818 4499 3852 4507
rect 3852 4499 3861 4507
rect 4009 4613 4018 4621
rect 4018 4613 4052 4621
rect 4052 4613 4061 4621
rect 4009 4569 4061 4613
rect 4209 4787 4261 4831
rect 4209 4779 4218 4787
rect 4218 4779 4252 4787
rect 4252 4779 4261 4787
rect 4409 4894 4461 4903
rect 4409 4860 4418 4894
rect 4418 4860 4452 4894
rect 4452 4860 4461 4894
rect 4409 4851 4461 4860
rect 2809 3684 2861 3693
rect 2809 3650 2818 3684
rect 2818 3650 2852 3684
rect 2852 3650 2861 3684
rect 2809 3641 2861 3650
rect 1209 2474 1261 2483
rect 1209 2440 1218 2474
rect 1218 2440 1252 2474
rect 1252 2440 1261 2474
rect 1209 2431 1261 2440
rect 9 1493 18 1501
rect 18 1493 52 1501
rect 52 1493 61 1501
rect 9 1449 61 1493
rect 209 1667 261 1711
rect 209 1659 218 1667
rect 218 1659 252 1667
rect 252 1659 261 1667
rect 409 1773 418 1781
rect 418 1773 452 1781
rect 452 1773 461 1781
rect 409 1729 461 1773
rect 609 1947 661 1991
rect 609 1939 618 1947
rect 618 1939 652 1947
rect 652 1939 661 1947
rect 809 2053 818 2061
rect 818 2053 852 2061
rect 852 2053 861 2061
rect 809 2009 861 2053
rect 1009 2227 1061 2271
rect 1009 2219 1018 2227
rect 1018 2219 1052 2227
rect 1052 2219 1061 2227
rect 1209 2333 1218 2341
rect 1218 2333 1252 2341
rect 1252 2333 1261 2341
rect 1209 2289 1261 2333
rect 1409 2597 1461 2641
rect 1409 2589 1418 2597
rect 1418 2589 1452 2597
rect 1452 2589 1461 2597
rect 1609 2703 1618 2711
rect 1618 2703 1652 2711
rect 1652 2703 1661 2711
rect 1609 2659 1661 2703
rect 1809 2877 1861 2921
rect 1809 2869 1818 2877
rect 1818 2869 1852 2877
rect 1852 2869 1861 2877
rect 2009 2983 2018 2991
rect 2018 2983 2052 2991
rect 2052 2983 2061 2991
rect 2009 2939 2061 2983
rect 2209 3157 2261 3201
rect 2209 3149 2218 3157
rect 2218 3149 2252 3157
rect 2252 3149 2261 3157
rect 2409 3263 2418 3271
rect 2418 3263 2452 3271
rect 2452 3263 2461 3271
rect 2409 3219 2461 3263
rect 2609 3437 2661 3481
rect 2609 3429 2618 3437
rect 2618 3429 2652 3437
rect 2652 3429 2661 3437
rect 2809 3543 2818 3551
rect 2818 3543 2852 3551
rect 2852 3543 2861 3551
rect 2809 3499 2861 3543
rect 3009 3807 3061 3851
rect 3009 3799 3018 3807
rect 3018 3799 3052 3807
rect 3052 3799 3061 3807
rect 3209 3913 3218 3921
rect 3218 3913 3252 3921
rect 3252 3913 3261 3921
rect 3209 3869 3261 3913
rect 3409 4087 3461 4131
rect 3409 4079 3418 4087
rect 3418 4079 3452 4087
rect 3452 4079 3461 4087
rect 3609 4193 3618 4201
rect 3618 4193 3652 4201
rect 3652 4193 3661 4201
rect 3609 4149 3661 4193
rect 3809 4367 3861 4411
rect 3809 4359 3818 4367
rect 3818 4359 3852 4367
rect 3852 4359 3861 4367
rect 4009 4473 4018 4481
rect 4018 4473 4052 4481
rect 4052 4473 4061 4481
rect 4009 4429 4061 4473
rect 4209 4647 4261 4691
rect 4209 4639 4218 4647
rect 4218 4639 4252 4647
rect 4252 4639 4261 4647
rect 4409 4753 4418 4761
rect 4418 4753 4452 4761
rect 4452 4753 4461 4761
rect 4409 4709 4461 4753
rect 4609 4910 4661 4919
rect 4609 4876 4618 4910
rect 4618 4876 4652 4910
rect 4652 4876 4661 4910
rect 4609 4867 4661 4876
rect 3009 3700 3061 3709
rect 3009 3666 3018 3700
rect 3018 3666 3052 3700
rect 3052 3666 3061 3700
rect 3009 3657 3061 3666
rect 1409 2490 1461 2499
rect 1409 2456 1418 2490
rect 1418 2456 1452 2490
rect 1452 2456 1461 2490
rect 1409 2447 1461 2456
rect 9 1353 18 1361
rect 18 1353 52 1361
rect 52 1353 61 1361
rect 9 1309 61 1353
rect 209 1527 261 1571
rect 209 1519 218 1527
rect 218 1519 252 1527
rect 252 1519 261 1527
rect 409 1633 418 1641
rect 418 1633 452 1641
rect 452 1633 461 1641
rect 409 1589 461 1633
rect 609 1807 661 1851
rect 609 1799 618 1807
rect 618 1799 652 1807
rect 652 1799 661 1807
rect 809 1913 818 1921
rect 818 1913 852 1921
rect 852 1913 861 1921
rect 809 1869 861 1913
rect 1009 2087 1061 2131
rect 1009 2079 1018 2087
rect 1018 2079 1052 2087
rect 1052 2079 1061 2087
rect 1209 2193 1218 2201
rect 1218 2193 1252 2201
rect 1252 2193 1261 2201
rect 1209 2149 1261 2193
rect 1409 2367 1461 2411
rect 1409 2359 1418 2367
rect 1418 2359 1452 2367
rect 1452 2359 1461 2367
rect 1609 2563 1618 2571
rect 1618 2563 1652 2571
rect 1652 2563 1661 2571
rect 1609 2519 1661 2563
rect 1809 2737 1861 2781
rect 1809 2729 1818 2737
rect 1818 2729 1852 2737
rect 1852 2729 1861 2737
rect 2009 2843 2018 2851
rect 2018 2843 2052 2851
rect 2052 2843 2061 2851
rect 2009 2799 2061 2843
rect 2209 3017 2261 3061
rect 2209 3009 2218 3017
rect 2218 3009 2252 3017
rect 2252 3009 2261 3017
rect 2409 3123 2418 3131
rect 2418 3123 2452 3131
rect 2452 3123 2461 3131
rect 2409 3079 2461 3123
rect 2609 3297 2661 3341
rect 2609 3289 2618 3297
rect 2618 3289 2652 3297
rect 2652 3289 2661 3297
rect 2809 3403 2818 3411
rect 2818 3403 2852 3411
rect 2852 3403 2861 3411
rect 2809 3359 2861 3403
rect 3009 3577 3061 3621
rect 3009 3569 3018 3577
rect 3018 3569 3052 3577
rect 3052 3569 3061 3577
rect 3209 3773 3218 3781
rect 3218 3773 3252 3781
rect 3252 3773 3261 3781
rect 3209 3729 3261 3773
rect 3409 3947 3461 3991
rect 3409 3939 3418 3947
rect 3418 3939 3452 3947
rect 3452 3939 3461 3947
rect 3609 4053 3618 4061
rect 3618 4053 3652 4061
rect 3652 4053 3661 4061
rect 3609 4009 3661 4053
rect 3809 4227 3861 4271
rect 3809 4219 3818 4227
rect 3818 4219 3852 4227
rect 3852 4219 3861 4227
rect 4009 4333 4018 4341
rect 4018 4333 4052 4341
rect 4052 4333 4061 4341
rect 4009 4289 4061 4333
rect 4209 4507 4261 4551
rect 4209 4499 4218 4507
rect 4218 4499 4252 4507
rect 4252 4499 4261 4507
rect 4409 4613 4418 4621
rect 4418 4613 4452 4621
rect 4452 4613 4461 4621
rect 4409 4569 4461 4613
rect 4609 4787 4661 4831
rect 4609 4779 4618 4787
rect 4618 4779 4652 4787
rect 4652 4779 4661 4787
rect 4809 4894 4861 4903
rect 4809 4860 4818 4894
rect 4818 4860 4852 4894
rect 4852 4860 4861 4894
rect 4809 4851 4861 4860
rect 3209 3684 3261 3693
rect 3209 3650 3218 3684
rect 3218 3650 3252 3684
rect 3252 3650 3261 3684
rect 3209 3641 3261 3650
rect 1609 2474 1661 2483
rect 1609 2440 1618 2474
rect 1618 2440 1652 2474
rect 1652 2440 1661 2474
rect 1609 2431 1661 2440
rect 9 1264 61 1273
rect 9 1230 18 1264
rect 18 1230 52 1264
rect 52 1230 61 1264
rect 9 1221 61 1230
rect 9 1123 18 1131
rect 18 1123 52 1131
rect 52 1123 61 1131
rect 9 1079 61 1123
rect 209 1387 261 1431
rect 209 1379 218 1387
rect 218 1379 252 1387
rect 252 1379 261 1387
rect 409 1493 418 1501
rect 418 1493 452 1501
rect 452 1493 461 1501
rect 409 1449 461 1493
rect 609 1667 661 1711
rect 609 1659 618 1667
rect 618 1659 652 1667
rect 652 1659 661 1667
rect 809 1773 818 1781
rect 818 1773 852 1781
rect 852 1773 861 1781
rect 809 1729 861 1773
rect 1009 1947 1061 1991
rect 1009 1939 1018 1947
rect 1018 1939 1052 1947
rect 1052 1939 1061 1947
rect 1209 2053 1218 2061
rect 1218 2053 1252 2061
rect 1252 2053 1261 2061
rect 1209 2009 1261 2053
rect 1409 2227 1461 2271
rect 1409 2219 1418 2227
rect 1418 2219 1452 2227
rect 1452 2219 1461 2227
rect 1609 2333 1618 2341
rect 1618 2333 1652 2341
rect 1652 2333 1661 2341
rect 1609 2289 1661 2333
rect 1809 2597 1861 2641
rect 1809 2589 1818 2597
rect 1818 2589 1852 2597
rect 1852 2589 1861 2597
rect 2009 2703 2018 2711
rect 2018 2703 2052 2711
rect 2052 2703 2061 2711
rect 2009 2659 2061 2703
rect 2209 2877 2261 2921
rect 2209 2869 2218 2877
rect 2218 2869 2252 2877
rect 2252 2869 2261 2877
rect 2409 2983 2418 2991
rect 2418 2983 2452 2991
rect 2452 2983 2461 2991
rect 2409 2939 2461 2983
rect 2609 3157 2661 3201
rect 2609 3149 2618 3157
rect 2618 3149 2652 3157
rect 2652 3149 2661 3157
rect 2809 3263 2818 3271
rect 2818 3263 2852 3271
rect 2852 3263 2861 3271
rect 2809 3219 2861 3263
rect 3009 3437 3061 3481
rect 3009 3429 3018 3437
rect 3018 3429 3052 3437
rect 3052 3429 3061 3437
rect 3209 3543 3218 3551
rect 3218 3543 3252 3551
rect 3252 3543 3261 3551
rect 3209 3499 3261 3543
rect 3409 3807 3461 3851
rect 3409 3799 3418 3807
rect 3418 3799 3452 3807
rect 3452 3799 3461 3807
rect 3609 3913 3618 3921
rect 3618 3913 3652 3921
rect 3652 3913 3661 3921
rect 3609 3869 3661 3913
rect 3809 4087 3861 4131
rect 3809 4079 3818 4087
rect 3818 4079 3852 4087
rect 3852 4079 3861 4087
rect 4009 4193 4018 4201
rect 4018 4193 4052 4201
rect 4052 4193 4061 4201
rect 4009 4149 4061 4193
rect 4209 4367 4261 4411
rect 4209 4359 4218 4367
rect 4218 4359 4252 4367
rect 4252 4359 4261 4367
rect 4409 4473 4418 4481
rect 4418 4473 4452 4481
rect 4452 4473 4461 4481
rect 4409 4429 4461 4473
rect 4609 4647 4661 4691
rect 4609 4639 4618 4647
rect 4618 4639 4652 4647
rect 4652 4639 4661 4647
rect 4809 4753 4818 4761
rect 4818 4753 4852 4761
rect 4852 4753 4861 4761
rect 4809 4709 4861 4753
rect 5009 4910 5061 4919
rect 5009 4876 5018 4910
rect 5018 4876 5052 4910
rect 5052 4876 5061 4910
rect 5009 4867 5061 4876
rect 3409 3700 3461 3709
rect 3409 3666 3418 3700
rect 3418 3666 3452 3700
rect 3452 3666 3461 3700
rect 3409 3657 3461 3666
rect 1809 2490 1861 2499
rect 1809 2456 1818 2490
rect 1818 2456 1852 2490
rect 1852 2456 1861 2490
rect 1809 2447 1861 2456
rect 209 1280 261 1289
rect 209 1246 218 1280
rect 218 1246 252 1280
rect 252 1246 261 1280
rect 209 1237 261 1246
rect 9 983 18 991
rect 18 983 52 991
rect 52 983 61 991
rect 9 939 61 983
rect 209 1157 261 1201
rect 209 1149 218 1157
rect 218 1149 252 1157
rect 252 1149 261 1157
rect 409 1353 418 1361
rect 418 1353 452 1361
rect 452 1353 461 1361
rect 409 1309 461 1353
rect 609 1527 661 1571
rect 609 1519 618 1527
rect 618 1519 652 1527
rect 652 1519 661 1527
rect 809 1633 818 1641
rect 818 1633 852 1641
rect 852 1633 861 1641
rect 809 1589 861 1633
rect 1009 1807 1061 1851
rect 1009 1799 1018 1807
rect 1018 1799 1052 1807
rect 1052 1799 1061 1807
rect 1209 1913 1218 1921
rect 1218 1913 1252 1921
rect 1252 1913 1261 1921
rect 1209 1869 1261 1913
rect 1409 2087 1461 2131
rect 1409 2079 1418 2087
rect 1418 2079 1452 2087
rect 1452 2079 1461 2087
rect 1609 2193 1618 2201
rect 1618 2193 1652 2201
rect 1652 2193 1661 2201
rect 1609 2149 1661 2193
rect 1809 2367 1861 2411
rect 1809 2359 1818 2367
rect 1818 2359 1852 2367
rect 1852 2359 1861 2367
rect 2009 2563 2018 2571
rect 2018 2563 2052 2571
rect 2052 2563 2061 2571
rect 2009 2519 2061 2563
rect 2209 2737 2261 2781
rect 2209 2729 2218 2737
rect 2218 2729 2252 2737
rect 2252 2729 2261 2737
rect 2409 2843 2418 2851
rect 2418 2843 2452 2851
rect 2452 2843 2461 2851
rect 2409 2799 2461 2843
rect 2609 3017 2661 3061
rect 2609 3009 2618 3017
rect 2618 3009 2652 3017
rect 2652 3009 2661 3017
rect 2809 3123 2818 3131
rect 2818 3123 2852 3131
rect 2852 3123 2861 3131
rect 2809 3079 2861 3123
rect 3009 3297 3061 3341
rect 3009 3289 3018 3297
rect 3018 3289 3052 3297
rect 3052 3289 3061 3297
rect 3209 3403 3218 3411
rect 3218 3403 3252 3411
rect 3252 3403 3261 3411
rect 3209 3359 3261 3403
rect 3409 3577 3461 3621
rect 3409 3569 3418 3577
rect 3418 3569 3452 3577
rect 3452 3569 3461 3577
rect 3609 3773 3618 3781
rect 3618 3773 3652 3781
rect 3652 3773 3661 3781
rect 3609 3729 3661 3773
rect 3809 3947 3861 3991
rect 3809 3939 3818 3947
rect 3818 3939 3852 3947
rect 3852 3939 3861 3947
rect 4009 4053 4018 4061
rect 4018 4053 4052 4061
rect 4052 4053 4061 4061
rect 4009 4009 4061 4053
rect 4209 4227 4261 4271
rect 4209 4219 4218 4227
rect 4218 4219 4252 4227
rect 4252 4219 4261 4227
rect 4409 4333 4418 4341
rect 4418 4333 4452 4341
rect 4452 4333 4461 4341
rect 4409 4289 4461 4333
rect 4609 4507 4661 4551
rect 4609 4499 4618 4507
rect 4618 4499 4652 4507
rect 4652 4499 4661 4507
rect 4809 4613 4818 4621
rect 4818 4613 4852 4621
rect 4852 4613 4861 4621
rect 4809 4569 4861 4613
rect 5009 4787 5061 4831
rect 5009 4779 5018 4787
rect 5018 4779 5052 4787
rect 5052 4779 5061 4787
rect 5209 4894 5261 4903
rect 5209 4860 5218 4894
rect 5218 4860 5252 4894
rect 5252 4860 5261 4894
rect 5209 4851 5261 4860
rect 3609 3684 3661 3693
rect 3609 3650 3618 3684
rect 3618 3650 3652 3684
rect 3652 3650 3661 3684
rect 3609 3641 3661 3650
rect 2009 2474 2061 2483
rect 2009 2440 2018 2474
rect 2018 2440 2052 2474
rect 2052 2440 2061 2474
rect 2009 2431 2061 2440
rect 409 1264 461 1273
rect 409 1230 418 1264
rect 418 1230 452 1264
rect 452 1230 461 1264
rect 409 1221 461 1230
rect 9 843 18 851
rect 18 843 52 851
rect 52 843 61 851
rect 9 799 61 843
rect 209 1017 261 1061
rect 209 1009 218 1017
rect 218 1009 252 1017
rect 252 1009 261 1017
rect 409 1123 418 1131
rect 418 1123 452 1131
rect 452 1123 461 1131
rect 409 1079 461 1123
rect 609 1387 661 1431
rect 609 1379 618 1387
rect 618 1379 652 1387
rect 652 1379 661 1387
rect 809 1493 818 1501
rect 818 1493 852 1501
rect 852 1493 861 1501
rect 809 1449 861 1493
rect 1009 1667 1061 1711
rect 1009 1659 1018 1667
rect 1018 1659 1052 1667
rect 1052 1659 1061 1667
rect 1209 1773 1218 1781
rect 1218 1773 1252 1781
rect 1252 1773 1261 1781
rect 1209 1729 1261 1773
rect 1409 1947 1461 1991
rect 1409 1939 1418 1947
rect 1418 1939 1452 1947
rect 1452 1939 1461 1947
rect 1609 2053 1618 2061
rect 1618 2053 1652 2061
rect 1652 2053 1661 2061
rect 1609 2009 1661 2053
rect 1809 2227 1861 2271
rect 1809 2219 1818 2227
rect 1818 2219 1852 2227
rect 1852 2219 1861 2227
rect 2009 2333 2018 2341
rect 2018 2333 2052 2341
rect 2052 2333 2061 2341
rect 2009 2289 2061 2333
rect 2209 2597 2261 2641
rect 2209 2589 2218 2597
rect 2218 2589 2252 2597
rect 2252 2589 2261 2597
rect 2409 2703 2418 2711
rect 2418 2703 2452 2711
rect 2452 2703 2461 2711
rect 2409 2659 2461 2703
rect 2609 2877 2661 2921
rect 2609 2869 2618 2877
rect 2618 2869 2652 2877
rect 2652 2869 2661 2877
rect 2809 2983 2818 2991
rect 2818 2983 2852 2991
rect 2852 2983 2861 2991
rect 2809 2939 2861 2983
rect 3009 3157 3061 3201
rect 3009 3149 3018 3157
rect 3018 3149 3052 3157
rect 3052 3149 3061 3157
rect 3209 3263 3218 3271
rect 3218 3263 3252 3271
rect 3252 3263 3261 3271
rect 3209 3219 3261 3263
rect 3409 3437 3461 3481
rect 3409 3429 3418 3437
rect 3418 3429 3452 3437
rect 3452 3429 3461 3437
rect 3609 3543 3618 3551
rect 3618 3543 3652 3551
rect 3652 3543 3661 3551
rect 3609 3499 3661 3543
rect 3809 3807 3861 3851
rect 3809 3799 3818 3807
rect 3818 3799 3852 3807
rect 3852 3799 3861 3807
rect 4009 3913 4018 3921
rect 4018 3913 4052 3921
rect 4052 3913 4061 3921
rect 4009 3869 4061 3913
rect 4209 4087 4261 4131
rect 4209 4079 4218 4087
rect 4218 4079 4252 4087
rect 4252 4079 4261 4087
rect 4409 4193 4418 4201
rect 4418 4193 4452 4201
rect 4452 4193 4461 4201
rect 4409 4149 4461 4193
rect 4609 4367 4661 4411
rect 4609 4359 4618 4367
rect 4618 4359 4652 4367
rect 4652 4359 4661 4367
rect 4809 4473 4818 4481
rect 4818 4473 4852 4481
rect 4852 4473 4861 4481
rect 4809 4429 4861 4473
rect 5009 4647 5061 4691
rect 5009 4639 5018 4647
rect 5018 4639 5052 4647
rect 5052 4639 5061 4647
rect 5209 4753 5218 4761
rect 5218 4753 5252 4761
rect 5252 4753 5261 4761
rect 5209 4709 5261 4753
rect 5409 4910 5461 4919
rect 5409 4876 5418 4910
rect 5418 4876 5452 4910
rect 5452 4876 5461 4910
rect 5409 4867 5461 4876
rect 3809 3700 3861 3709
rect 3809 3666 3818 3700
rect 3818 3666 3852 3700
rect 3852 3666 3861 3700
rect 3809 3657 3861 3666
rect 2209 2490 2261 2499
rect 2209 2456 2218 2490
rect 2218 2456 2252 2490
rect 2252 2456 2261 2490
rect 2209 2447 2261 2456
rect 609 1280 661 1289
rect 609 1246 618 1280
rect 618 1246 652 1280
rect 652 1246 661 1280
rect 609 1237 661 1246
rect 9 703 18 711
rect 18 703 52 711
rect 52 703 61 711
rect 9 659 61 703
rect 209 877 261 921
rect 209 869 218 877
rect 218 869 252 877
rect 252 869 261 877
rect 409 983 418 991
rect 418 983 452 991
rect 452 983 461 991
rect 409 939 461 983
rect 609 1157 661 1201
rect 609 1149 618 1157
rect 618 1149 652 1157
rect 652 1149 661 1157
rect 809 1353 818 1361
rect 818 1353 852 1361
rect 852 1353 861 1361
rect 809 1309 861 1353
rect 1009 1527 1061 1571
rect 1009 1519 1018 1527
rect 1018 1519 1052 1527
rect 1052 1519 1061 1527
rect 1209 1633 1218 1641
rect 1218 1633 1252 1641
rect 1252 1633 1261 1641
rect 1209 1589 1261 1633
rect 1409 1807 1461 1851
rect 1409 1799 1418 1807
rect 1418 1799 1452 1807
rect 1452 1799 1461 1807
rect 1609 1913 1618 1921
rect 1618 1913 1652 1921
rect 1652 1913 1661 1921
rect 1609 1869 1661 1913
rect 1809 2087 1861 2131
rect 1809 2079 1818 2087
rect 1818 2079 1852 2087
rect 1852 2079 1861 2087
rect 2009 2193 2018 2201
rect 2018 2193 2052 2201
rect 2052 2193 2061 2201
rect 2009 2149 2061 2193
rect 2209 2367 2261 2411
rect 2209 2359 2218 2367
rect 2218 2359 2252 2367
rect 2252 2359 2261 2367
rect 2409 2563 2418 2571
rect 2418 2563 2452 2571
rect 2452 2563 2461 2571
rect 2409 2519 2461 2563
rect 2609 2737 2661 2781
rect 2609 2729 2618 2737
rect 2618 2729 2652 2737
rect 2652 2729 2661 2737
rect 2809 2843 2818 2851
rect 2818 2843 2852 2851
rect 2852 2843 2861 2851
rect 2809 2799 2861 2843
rect 3009 3017 3061 3061
rect 3009 3009 3018 3017
rect 3018 3009 3052 3017
rect 3052 3009 3061 3017
rect 3209 3123 3218 3131
rect 3218 3123 3252 3131
rect 3252 3123 3261 3131
rect 3209 3079 3261 3123
rect 3409 3297 3461 3341
rect 3409 3289 3418 3297
rect 3418 3289 3452 3297
rect 3452 3289 3461 3297
rect 3609 3403 3618 3411
rect 3618 3403 3652 3411
rect 3652 3403 3661 3411
rect 3609 3359 3661 3403
rect 3809 3577 3861 3621
rect 3809 3569 3818 3577
rect 3818 3569 3852 3577
rect 3852 3569 3861 3577
rect 4009 3773 4018 3781
rect 4018 3773 4052 3781
rect 4052 3773 4061 3781
rect 4009 3729 4061 3773
rect 4209 3947 4261 3991
rect 4209 3939 4218 3947
rect 4218 3939 4252 3947
rect 4252 3939 4261 3947
rect 4409 4053 4418 4061
rect 4418 4053 4452 4061
rect 4452 4053 4461 4061
rect 4409 4009 4461 4053
rect 4609 4227 4661 4271
rect 4609 4219 4618 4227
rect 4618 4219 4652 4227
rect 4652 4219 4661 4227
rect 4809 4333 4818 4341
rect 4818 4333 4852 4341
rect 4852 4333 4861 4341
rect 4809 4289 4861 4333
rect 5009 4507 5061 4551
rect 5009 4499 5018 4507
rect 5018 4499 5052 4507
rect 5052 4499 5061 4507
rect 5209 4613 5218 4621
rect 5218 4613 5252 4621
rect 5252 4613 5261 4621
rect 5209 4569 5261 4613
rect 5409 4787 5461 4831
rect 5409 4779 5418 4787
rect 5418 4779 5452 4787
rect 5452 4779 5461 4787
rect 5609 4894 5661 4903
rect 5609 4860 5618 4894
rect 5618 4860 5652 4894
rect 5652 4860 5661 4894
rect 5609 4851 5661 4860
rect 4009 3684 4061 3693
rect 4009 3650 4018 3684
rect 4018 3650 4052 3684
rect 4052 3650 4061 3684
rect 4009 3641 4061 3650
rect 2409 2474 2461 2483
rect 2409 2440 2418 2474
rect 2418 2440 2452 2474
rect 2452 2440 2461 2474
rect 2409 2431 2461 2440
rect 809 1264 861 1273
rect 809 1230 818 1264
rect 818 1230 852 1264
rect 852 1230 861 1264
rect 809 1221 861 1230
rect 9 563 18 571
rect 18 563 52 571
rect 52 563 61 571
rect 9 519 61 563
rect 209 737 261 781
rect 209 729 218 737
rect 218 729 252 737
rect 252 729 261 737
rect 409 843 418 851
rect 418 843 452 851
rect 452 843 461 851
rect 409 799 461 843
rect 609 1017 661 1061
rect 609 1009 618 1017
rect 618 1009 652 1017
rect 652 1009 661 1017
rect 809 1123 818 1131
rect 818 1123 852 1131
rect 852 1123 861 1131
rect 809 1079 861 1123
rect 1009 1387 1061 1431
rect 1009 1379 1018 1387
rect 1018 1379 1052 1387
rect 1052 1379 1061 1387
rect 1209 1493 1218 1501
rect 1218 1493 1252 1501
rect 1252 1493 1261 1501
rect 1209 1449 1261 1493
rect 1409 1667 1461 1711
rect 1409 1659 1418 1667
rect 1418 1659 1452 1667
rect 1452 1659 1461 1667
rect 1609 1773 1618 1781
rect 1618 1773 1652 1781
rect 1652 1773 1661 1781
rect 1609 1729 1661 1773
rect 1809 1947 1861 1991
rect 1809 1939 1818 1947
rect 1818 1939 1852 1947
rect 1852 1939 1861 1947
rect 2009 2053 2018 2061
rect 2018 2053 2052 2061
rect 2052 2053 2061 2061
rect 2009 2009 2061 2053
rect 2209 2227 2261 2271
rect 2209 2219 2218 2227
rect 2218 2219 2252 2227
rect 2252 2219 2261 2227
rect 2409 2333 2418 2341
rect 2418 2333 2452 2341
rect 2452 2333 2461 2341
rect 2409 2289 2461 2333
rect 2609 2597 2661 2641
rect 2609 2589 2618 2597
rect 2618 2589 2652 2597
rect 2652 2589 2661 2597
rect 2809 2703 2818 2711
rect 2818 2703 2852 2711
rect 2852 2703 2861 2711
rect 2809 2659 2861 2703
rect 3009 2877 3061 2921
rect 3009 2869 3018 2877
rect 3018 2869 3052 2877
rect 3052 2869 3061 2877
rect 3209 2983 3218 2991
rect 3218 2983 3252 2991
rect 3252 2983 3261 2991
rect 3209 2939 3261 2983
rect 3409 3157 3461 3201
rect 3409 3149 3418 3157
rect 3418 3149 3452 3157
rect 3452 3149 3461 3157
rect 3609 3263 3618 3271
rect 3618 3263 3652 3271
rect 3652 3263 3661 3271
rect 3609 3219 3661 3263
rect 3809 3437 3861 3481
rect 3809 3429 3818 3437
rect 3818 3429 3852 3437
rect 3852 3429 3861 3437
rect 4009 3543 4018 3551
rect 4018 3543 4052 3551
rect 4052 3543 4061 3551
rect 4009 3499 4061 3543
rect 4209 3807 4261 3851
rect 4209 3799 4218 3807
rect 4218 3799 4252 3807
rect 4252 3799 4261 3807
rect 4409 3913 4418 3921
rect 4418 3913 4452 3921
rect 4452 3913 4461 3921
rect 4409 3869 4461 3913
rect 4609 4087 4661 4131
rect 4609 4079 4618 4087
rect 4618 4079 4652 4087
rect 4652 4079 4661 4087
rect 4809 4193 4818 4201
rect 4818 4193 4852 4201
rect 4852 4193 4861 4201
rect 4809 4149 4861 4193
rect 5009 4367 5061 4411
rect 5009 4359 5018 4367
rect 5018 4359 5052 4367
rect 5052 4359 5061 4367
rect 5209 4473 5218 4481
rect 5218 4473 5252 4481
rect 5252 4473 5261 4481
rect 5209 4429 5261 4473
rect 5409 4647 5461 4691
rect 5409 4639 5418 4647
rect 5418 4639 5452 4647
rect 5452 4639 5461 4647
rect 5609 4753 5618 4761
rect 5618 4753 5652 4761
rect 5652 4753 5661 4761
rect 5609 4709 5661 4753
rect 5809 4910 5861 4919
rect 5809 4876 5818 4910
rect 5818 4876 5852 4910
rect 5852 4876 5861 4910
rect 5809 4867 5861 4876
rect 4209 3700 4261 3709
rect 4209 3666 4218 3700
rect 4218 3666 4252 3700
rect 4252 3666 4261 3700
rect 4209 3657 4261 3666
rect 2609 2490 2661 2499
rect 2609 2456 2618 2490
rect 2618 2456 2652 2490
rect 2652 2456 2661 2490
rect 2609 2447 2661 2456
rect 1009 1280 1061 1289
rect 1009 1246 1018 1280
rect 1018 1246 1052 1280
rect 1052 1246 1061 1280
rect 1009 1237 1061 1246
rect 9 423 18 431
rect 18 423 52 431
rect 52 423 61 431
rect 9 379 61 423
rect 209 597 261 641
rect 209 589 218 597
rect 218 589 252 597
rect 252 589 261 597
rect 409 703 418 711
rect 418 703 452 711
rect 452 703 461 711
rect 409 659 461 703
rect 609 877 661 921
rect 609 869 618 877
rect 618 869 652 877
rect 652 869 661 877
rect 809 983 818 991
rect 818 983 852 991
rect 852 983 861 991
rect 809 939 861 983
rect 1009 1157 1061 1201
rect 1009 1149 1018 1157
rect 1018 1149 1052 1157
rect 1052 1149 1061 1157
rect 1209 1353 1218 1361
rect 1218 1353 1252 1361
rect 1252 1353 1261 1361
rect 1209 1309 1261 1353
rect 1409 1527 1461 1571
rect 1409 1519 1418 1527
rect 1418 1519 1452 1527
rect 1452 1519 1461 1527
rect 1609 1633 1618 1641
rect 1618 1633 1652 1641
rect 1652 1633 1661 1641
rect 1609 1589 1661 1633
rect 1809 1807 1861 1851
rect 1809 1799 1818 1807
rect 1818 1799 1852 1807
rect 1852 1799 1861 1807
rect 2009 1913 2018 1921
rect 2018 1913 2052 1921
rect 2052 1913 2061 1921
rect 2009 1869 2061 1913
rect 2209 2087 2261 2131
rect 2209 2079 2218 2087
rect 2218 2079 2252 2087
rect 2252 2079 2261 2087
rect 2409 2193 2418 2201
rect 2418 2193 2452 2201
rect 2452 2193 2461 2201
rect 2409 2149 2461 2193
rect 2609 2367 2661 2411
rect 2609 2359 2618 2367
rect 2618 2359 2652 2367
rect 2652 2359 2661 2367
rect 2809 2563 2818 2571
rect 2818 2563 2852 2571
rect 2852 2563 2861 2571
rect 2809 2519 2861 2563
rect 3009 2737 3061 2781
rect 3009 2729 3018 2737
rect 3018 2729 3052 2737
rect 3052 2729 3061 2737
rect 3209 2843 3218 2851
rect 3218 2843 3252 2851
rect 3252 2843 3261 2851
rect 3209 2799 3261 2843
rect 3409 3017 3461 3061
rect 3409 3009 3418 3017
rect 3418 3009 3452 3017
rect 3452 3009 3461 3017
rect 3609 3123 3618 3131
rect 3618 3123 3652 3131
rect 3652 3123 3661 3131
rect 3609 3079 3661 3123
rect 3809 3297 3861 3341
rect 3809 3289 3818 3297
rect 3818 3289 3852 3297
rect 3852 3289 3861 3297
rect 4009 3403 4018 3411
rect 4018 3403 4052 3411
rect 4052 3403 4061 3411
rect 4009 3359 4061 3403
rect 4209 3577 4261 3621
rect 4209 3569 4218 3577
rect 4218 3569 4252 3577
rect 4252 3569 4261 3577
rect 4409 3773 4418 3781
rect 4418 3773 4452 3781
rect 4452 3773 4461 3781
rect 4409 3729 4461 3773
rect 4609 3947 4661 3991
rect 4609 3939 4618 3947
rect 4618 3939 4652 3947
rect 4652 3939 4661 3947
rect 4809 4053 4818 4061
rect 4818 4053 4852 4061
rect 4852 4053 4861 4061
rect 4809 4009 4861 4053
rect 5009 4227 5061 4271
rect 5009 4219 5018 4227
rect 5018 4219 5052 4227
rect 5052 4219 5061 4227
rect 5209 4333 5218 4341
rect 5218 4333 5252 4341
rect 5252 4333 5261 4341
rect 5209 4289 5261 4333
rect 5409 4507 5461 4551
rect 5409 4499 5418 4507
rect 5418 4499 5452 4507
rect 5452 4499 5461 4507
rect 5609 4613 5618 4621
rect 5618 4613 5652 4621
rect 5652 4613 5661 4621
rect 5609 4569 5661 4613
rect 5809 4787 5861 4831
rect 5809 4779 5818 4787
rect 5818 4779 5852 4787
rect 5852 4779 5861 4787
rect 6009 4894 6061 4903
rect 6009 4860 6018 4894
rect 6018 4860 6052 4894
rect 6052 4860 6061 4894
rect 6009 4851 6061 4860
rect 4409 3684 4461 3693
rect 4409 3650 4418 3684
rect 4418 3650 4452 3684
rect 4452 3650 4461 3684
rect 4409 3641 4461 3650
rect 2809 2474 2861 2483
rect 2809 2440 2818 2474
rect 2818 2440 2852 2474
rect 2852 2440 2861 2474
rect 2809 2431 2861 2440
rect 1209 1264 1261 1273
rect 1209 1230 1218 1264
rect 1218 1230 1252 1264
rect 1252 1230 1261 1264
rect 1209 1221 1261 1230
rect 9 283 18 291
rect 18 283 52 291
rect 52 283 61 291
rect 9 239 61 283
rect 209 457 261 501
rect 209 449 218 457
rect 218 449 252 457
rect 252 449 261 457
rect 409 563 418 571
rect 418 563 452 571
rect 452 563 461 571
rect 409 519 461 563
rect 609 737 661 781
rect 609 729 618 737
rect 618 729 652 737
rect 652 729 661 737
rect 809 843 818 851
rect 818 843 852 851
rect 852 843 861 851
rect 809 799 861 843
rect 1009 1017 1061 1061
rect 1009 1009 1018 1017
rect 1018 1009 1052 1017
rect 1052 1009 1061 1017
rect 1209 1123 1218 1131
rect 1218 1123 1252 1131
rect 1252 1123 1261 1131
rect 1209 1079 1261 1123
rect 1409 1387 1461 1431
rect 1409 1379 1418 1387
rect 1418 1379 1452 1387
rect 1452 1379 1461 1387
rect 1609 1493 1618 1501
rect 1618 1493 1652 1501
rect 1652 1493 1661 1501
rect 1609 1449 1661 1493
rect 1809 1667 1861 1711
rect 1809 1659 1818 1667
rect 1818 1659 1852 1667
rect 1852 1659 1861 1667
rect 2009 1773 2018 1781
rect 2018 1773 2052 1781
rect 2052 1773 2061 1781
rect 2009 1729 2061 1773
rect 2209 1947 2261 1991
rect 2209 1939 2218 1947
rect 2218 1939 2252 1947
rect 2252 1939 2261 1947
rect 2409 2053 2418 2061
rect 2418 2053 2452 2061
rect 2452 2053 2461 2061
rect 2409 2009 2461 2053
rect 2609 2227 2661 2271
rect 2609 2219 2618 2227
rect 2618 2219 2652 2227
rect 2652 2219 2661 2227
rect 2809 2333 2818 2341
rect 2818 2333 2852 2341
rect 2852 2333 2861 2341
rect 2809 2289 2861 2333
rect 3009 2597 3061 2641
rect 3009 2589 3018 2597
rect 3018 2589 3052 2597
rect 3052 2589 3061 2597
rect 3209 2703 3218 2711
rect 3218 2703 3252 2711
rect 3252 2703 3261 2711
rect 3209 2659 3261 2703
rect 3409 2877 3461 2921
rect 3409 2869 3418 2877
rect 3418 2869 3452 2877
rect 3452 2869 3461 2877
rect 3609 2983 3618 2991
rect 3618 2983 3652 2991
rect 3652 2983 3661 2991
rect 3609 2939 3661 2983
rect 3809 3157 3861 3201
rect 3809 3149 3818 3157
rect 3818 3149 3852 3157
rect 3852 3149 3861 3157
rect 4009 3263 4018 3271
rect 4018 3263 4052 3271
rect 4052 3263 4061 3271
rect 4009 3219 4061 3263
rect 4209 3437 4261 3481
rect 4209 3429 4218 3437
rect 4218 3429 4252 3437
rect 4252 3429 4261 3437
rect 4409 3543 4418 3551
rect 4418 3543 4452 3551
rect 4452 3543 4461 3551
rect 4409 3499 4461 3543
rect 4609 3807 4661 3851
rect 4609 3799 4618 3807
rect 4618 3799 4652 3807
rect 4652 3799 4661 3807
rect 4809 3913 4818 3921
rect 4818 3913 4852 3921
rect 4852 3913 4861 3921
rect 4809 3869 4861 3913
rect 5009 4087 5061 4131
rect 5009 4079 5018 4087
rect 5018 4079 5052 4087
rect 5052 4079 5061 4087
rect 5209 4193 5218 4201
rect 5218 4193 5252 4201
rect 5252 4193 5261 4201
rect 5209 4149 5261 4193
rect 5409 4367 5461 4411
rect 5409 4359 5418 4367
rect 5418 4359 5452 4367
rect 5452 4359 5461 4367
rect 5609 4473 5618 4481
rect 5618 4473 5652 4481
rect 5652 4473 5661 4481
rect 5609 4429 5661 4473
rect 5809 4647 5861 4691
rect 5809 4639 5818 4647
rect 5818 4639 5852 4647
rect 5852 4639 5861 4647
rect 6009 4753 6018 4761
rect 6018 4753 6052 4761
rect 6052 4753 6061 4761
rect 6009 4709 6061 4753
rect 6209 4910 6261 4919
rect 6209 4876 6218 4910
rect 6218 4876 6252 4910
rect 6252 4876 6261 4910
rect 6209 4867 6261 4876
rect 4609 3700 4661 3709
rect 4609 3666 4618 3700
rect 4618 3666 4652 3700
rect 4652 3666 4661 3700
rect 4609 3657 4661 3666
rect 3009 2490 3061 2499
rect 3009 2456 3018 2490
rect 3018 2456 3052 2490
rect 3052 2456 3061 2490
rect 3009 2447 3061 2456
rect 1409 1280 1461 1289
rect 1409 1246 1418 1280
rect 1418 1246 1452 1280
rect 1452 1246 1461 1280
rect 1409 1237 1461 1246
rect 9 143 18 151
rect 18 143 52 151
rect 52 143 61 151
rect 9 99 61 143
rect 209 317 261 361
rect 209 309 218 317
rect 218 309 252 317
rect 252 309 261 317
rect 409 423 418 431
rect 418 423 452 431
rect 452 423 461 431
rect 409 379 461 423
rect 609 597 661 641
rect 609 589 618 597
rect 618 589 652 597
rect 652 589 661 597
rect 809 703 818 711
rect 818 703 852 711
rect 852 703 861 711
rect 809 659 861 703
rect 1009 877 1061 921
rect 1009 869 1018 877
rect 1018 869 1052 877
rect 1052 869 1061 877
rect 1209 983 1218 991
rect 1218 983 1252 991
rect 1252 983 1261 991
rect 1209 939 1261 983
rect 1409 1157 1461 1201
rect 1409 1149 1418 1157
rect 1418 1149 1452 1157
rect 1452 1149 1461 1157
rect 1609 1353 1618 1361
rect 1618 1353 1652 1361
rect 1652 1353 1661 1361
rect 1609 1309 1661 1353
rect 1809 1527 1861 1571
rect 1809 1519 1818 1527
rect 1818 1519 1852 1527
rect 1852 1519 1861 1527
rect 2009 1633 2018 1641
rect 2018 1633 2052 1641
rect 2052 1633 2061 1641
rect 2009 1589 2061 1633
rect 2209 1807 2261 1851
rect 2209 1799 2218 1807
rect 2218 1799 2252 1807
rect 2252 1799 2261 1807
rect 2409 1913 2418 1921
rect 2418 1913 2452 1921
rect 2452 1913 2461 1921
rect 2409 1869 2461 1913
rect 2609 2087 2661 2131
rect 2609 2079 2618 2087
rect 2618 2079 2652 2087
rect 2652 2079 2661 2087
rect 2809 2193 2818 2201
rect 2818 2193 2852 2201
rect 2852 2193 2861 2201
rect 2809 2149 2861 2193
rect 3009 2367 3061 2411
rect 3009 2359 3018 2367
rect 3018 2359 3052 2367
rect 3052 2359 3061 2367
rect 3209 2563 3218 2571
rect 3218 2563 3252 2571
rect 3252 2563 3261 2571
rect 3209 2519 3261 2563
rect 3409 2737 3461 2781
rect 3409 2729 3418 2737
rect 3418 2729 3452 2737
rect 3452 2729 3461 2737
rect 3609 2843 3618 2851
rect 3618 2843 3652 2851
rect 3652 2843 3661 2851
rect 3609 2799 3661 2843
rect 3809 3017 3861 3061
rect 3809 3009 3818 3017
rect 3818 3009 3852 3017
rect 3852 3009 3861 3017
rect 4009 3123 4018 3131
rect 4018 3123 4052 3131
rect 4052 3123 4061 3131
rect 4009 3079 4061 3123
rect 4209 3297 4261 3341
rect 4209 3289 4218 3297
rect 4218 3289 4252 3297
rect 4252 3289 4261 3297
rect 4409 3403 4418 3411
rect 4418 3403 4452 3411
rect 4452 3403 4461 3411
rect 4409 3359 4461 3403
rect 4609 3577 4661 3621
rect 4609 3569 4618 3577
rect 4618 3569 4652 3577
rect 4652 3569 4661 3577
rect 4809 3773 4818 3781
rect 4818 3773 4852 3781
rect 4852 3773 4861 3781
rect 4809 3729 4861 3773
rect 5009 3947 5061 3991
rect 5009 3939 5018 3947
rect 5018 3939 5052 3947
rect 5052 3939 5061 3947
rect 5209 4053 5218 4061
rect 5218 4053 5252 4061
rect 5252 4053 5261 4061
rect 5209 4009 5261 4053
rect 5409 4227 5461 4271
rect 5409 4219 5418 4227
rect 5418 4219 5452 4227
rect 5452 4219 5461 4227
rect 5609 4333 5618 4341
rect 5618 4333 5652 4341
rect 5652 4333 5661 4341
rect 5609 4289 5661 4333
rect 5809 4507 5861 4551
rect 5809 4499 5818 4507
rect 5818 4499 5852 4507
rect 5852 4499 5861 4507
rect 6009 4613 6018 4621
rect 6018 4613 6052 4621
rect 6052 4613 6061 4621
rect 6009 4569 6061 4613
rect 6209 4787 6261 4831
rect 6209 4779 6218 4787
rect 6218 4779 6252 4787
rect 6252 4779 6261 4787
rect 6409 4894 6461 4903
rect 6409 4860 6418 4894
rect 6418 4860 6452 4894
rect 6452 4860 6461 4894
rect 6409 4851 6461 4860
rect 4809 3684 4861 3693
rect 4809 3650 4818 3684
rect 4818 3650 4852 3684
rect 4852 3650 4861 3684
rect 4809 3641 4861 3650
rect 3209 2474 3261 2483
rect 3209 2440 3218 2474
rect 3218 2440 3252 2474
rect 3252 2440 3261 2474
rect 3209 2431 3261 2440
rect 1609 1264 1661 1273
rect 1609 1230 1618 1264
rect 1618 1230 1652 1264
rect 1652 1230 1661 1264
rect 1609 1221 1661 1230
rect 9 54 61 63
rect 9 20 18 54
rect 18 20 52 54
rect 52 20 61 54
rect 9 11 61 20
rect -91 -60 -39 -15
rect -91 -67 -82 -60
rect -82 -67 -48 -60
rect -48 -67 -39 -60
rect -91 -94 -82 -79
rect -82 -94 -48 -79
rect -48 -94 -39 -79
rect -91 -131 -39 -94
rect 9 -74 61 -22
rect 209 177 261 221
rect 209 169 218 177
rect 218 169 252 177
rect 252 169 261 177
rect 409 283 418 291
rect 418 283 452 291
rect 452 283 461 291
rect 409 239 461 283
rect 609 457 661 501
rect 609 449 618 457
rect 618 449 652 457
rect 652 449 661 457
rect 809 563 818 571
rect 818 563 852 571
rect 852 563 861 571
rect 809 519 861 563
rect 1009 737 1061 781
rect 1009 729 1018 737
rect 1018 729 1052 737
rect 1052 729 1061 737
rect 1209 843 1218 851
rect 1218 843 1252 851
rect 1252 843 1261 851
rect 1209 799 1261 843
rect 1409 1017 1461 1061
rect 1409 1009 1418 1017
rect 1418 1009 1452 1017
rect 1452 1009 1461 1017
rect 1609 1123 1618 1131
rect 1618 1123 1652 1131
rect 1652 1123 1661 1131
rect 1609 1079 1661 1123
rect 1809 1387 1861 1431
rect 1809 1379 1818 1387
rect 1818 1379 1852 1387
rect 1852 1379 1861 1387
rect 2009 1493 2018 1501
rect 2018 1493 2052 1501
rect 2052 1493 2061 1501
rect 2009 1449 2061 1493
rect 2209 1667 2261 1711
rect 2209 1659 2218 1667
rect 2218 1659 2252 1667
rect 2252 1659 2261 1667
rect 2409 1773 2418 1781
rect 2418 1773 2452 1781
rect 2452 1773 2461 1781
rect 2409 1729 2461 1773
rect 2609 1947 2661 1991
rect 2609 1939 2618 1947
rect 2618 1939 2652 1947
rect 2652 1939 2661 1947
rect 2809 2053 2818 2061
rect 2818 2053 2852 2061
rect 2852 2053 2861 2061
rect 2809 2009 2861 2053
rect 3009 2227 3061 2271
rect 3009 2219 3018 2227
rect 3018 2219 3052 2227
rect 3052 2219 3061 2227
rect 3209 2333 3218 2341
rect 3218 2333 3252 2341
rect 3252 2333 3261 2341
rect 3209 2289 3261 2333
rect 3409 2597 3461 2641
rect 3409 2589 3418 2597
rect 3418 2589 3452 2597
rect 3452 2589 3461 2597
rect 3609 2703 3618 2711
rect 3618 2703 3652 2711
rect 3652 2703 3661 2711
rect 3609 2659 3661 2703
rect 3809 2877 3861 2921
rect 3809 2869 3818 2877
rect 3818 2869 3852 2877
rect 3852 2869 3861 2877
rect 4009 2983 4018 2991
rect 4018 2983 4052 2991
rect 4052 2983 4061 2991
rect 4009 2939 4061 2983
rect 4209 3157 4261 3201
rect 4209 3149 4218 3157
rect 4218 3149 4252 3157
rect 4252 3149 4261 3157
rect 4409 3263 4418 3271
rect 4418 3263 4452 3271
rect 4452 3263 4461 3271
rect 4409 3219 4461 3263
rect 4609 3437 4661 3481
rect 4609 3429 4618 3437
rect 4618 3429 4652 3437
rect 4652 3429 4661 3437
rect 4809 3543 4818 3551
rect 4818 3543 4852 3551
rect 4852 3543 4861 3551
rect 4809 3499 4861 3543
rect 5009 3807 5061 3851
rect 5009 3799 5018 3807
rect 5018 3799 5052 3807
rect 5052 3799 5061 3807
rect 5209 3913 5218 3921
rect 5218 3913 5252 3921
rect 5252 3913 5261 3921
rect 5209 3869 5261 3913
rect 5409 4087 5461 4131
rect 5409 4079 5418 4087
rect 5418 4079 5452 4087
rect 5452 4079 5461 4087
rect 5609 4193 5618 4201
rect 5618 4193 5652 4201
rect 5652 4193 5661 4201
rect 5609 4149 5661 4193
rect 5809 4367 5861 4411
rect 5809 4359 5818 4367
rect 5818 4359 5852 4367
rect 5852 4359 5861 4367
rect 6009 4473 6018 4481
rect 6018 4473 6052 4481
rect 6052 4473 6061 4481
rect 6009 4429 6061 4473
rect 6209 4647 6261 4691
rect 6209 4639 6218 4647
rect 6218 4639 6252 4647
rect 6252 4639 6261 4647
rect 6409 4753 6418 4761
rect 6418 4753 6452 4761
rect 6452 4753 6461 4761
rect 6409 4709 6461 4753
rect 6609 4910 6661 4919
rect 6609 4876 6618 4910
rect 6618 4876 6652 4910
rect 6652 4876 6661 4910
rect 6609 4867 6661 4876
rect 5009 3700 5061 3709
rect 5009 3666 5018 3700
rect 5018 3666 5052 3700
rect 5052 3666 5061 3700
rect 5009 3657 5061 3666
rect 3409 2490 3461 2499
rect 3409 2456 3418 2490
rect 3418 2456 3452 2490
rect 3452 2456 3461 2490
rect 3409 2447 3461 2456
rect 1809 1280 1861 1289
rect 1809 1246 1818 1280
rect 1818 1246 1852 1280
rect 1852 1246 1861 1280
rect 1809 1237 1861 1246
rect 209 70 261 79
rect 209 36 218 70
rect 218 36 252 70
rect 252 36 261 70
rect 209 27 261 36
rect 109 -60 161 -15
rect 109 -67 118 -60
rect 118 -67 152 -60
rect 152 -67 161 -60
rect -91 -166 -82 -143
rect -82 -166 -48 -143
rect -48 -166 -39 -143
rect -91 -195 -39 -166
rect -75 -248 -23 -239
rect -75 -282 -66 -248
rect -66 -282 -32 -248
rect -32 -282 -23 -248
rect -75 -291 -23 -282
rect -91 -363 -39 -326
rect -91 -378 -82 -363
rect -82 -378 -48 -363
rect -48 -378 -39 -363
rect -91 -397 -82 -390
rect -82 -397 -48 -390
rect -48 -397 -39 -390
rect -91 -435 -39 -397
rect -91 -442 -82 -435
rect -82 -442 -48 -435
rect -48 -442 -39 -435
rect -91 -469 -82 -454
rect -82 -469 -48 -454
rect -48 -469 -39 -454
rect -91 -506 -39 -469
rect 109 -94 118 -79
rect 118 -94 152 -79
rect 152 -94 161 -79
rect 109 -131 161 -94
rect 209 -74 261 -22
rect 409 143 418 151
rect 418 143 452 151
rect 452 143 461 151
rect 409 99 461 143
rect 609 317 661 361
rect 609 309 618 317
rect 618 309 652 317
rect 652 309 661 317
rect 809 423 818 431
rect 818 423 852 431
rect 852 423 861 431
rect 809 379 861 423
rect 1009 597 1061 641
rect 1009 589 1018 597
rect 1018 589 1052 597
rect 1052 589 1061 597
rect 1209 703 1218 711
rect 1218 703 1252 711
rect 1252 703 1261 711
rect 1209 659 1261 703
rect 1409 877 1461 921
rect 1409 869 1418 877
rect 1418 869 1452 877
rect 1452 869 1461 877
rect 1609 983 1618 991
rect 1618 983 1652 991
rect 1652 983 1661 991
rect 1609 939 1661 983
rect 1809 1157 1861 1201
rect 1809 1149 1818 1157
rect 1818 1149 1852 1157
rect 1852 1149 1861 1157
rect 2009 1353 2018 1361
rect 2018 1353 2052 1361
rect 2052 1353 2061 1361
rect 2009 1309 2061 1353
rect 2209 1527 2261 1571
rect 2209 1519 2218 1527
rect 2218 1519 2252 1527
rect 2252 1519 2261 1527
rect 2409 1633 2418 1641
rect 2418 1633 2452 1641
rect 2452 1633 2461 1641
rect 2409 1589 2461 1633
rect 2609 1807 2661 1851
rect 2609 1799 2618 1807
rect 2618 1799 2652 1807
rect 2652 1799 2661 1807
rect 2809 1913 2818 1921
rect 2818 1913 2852 1921
rect 2852 1913 2861 1921
rect 2809 1869 2861 1913
rect 3009 2087 3061 2131
rect 3009 2079 3018 2087
rect 3018 2079 3052 2087
rect 3052 2079 3061 2087
rect 3209 2193 3218 2201
rect 3218 2193 3252 2201
rect 3252 2193 3261 2201
rect 3209 2149 3261 2193
rect 3409 2367 3461 2411
rect 3409 2359 3418 2367
rect 3418 2359 3452 2367
rect 3452 2359 3461 2367
rect 3609 2563 3618 2571
rect 3618 2563 3652 2571
rect 3652 2563 3661 2571
rect 3609 2519 3661 2563
rect 3809 2737 3861 2781
rect 3809 2729 3818 2737
rect 3818 2729 3852 2737
rect 3852 2729 3861 2737
rect 4009 2843 4018 2851
rect 4018 2843 4052 2851
rect 4052 2843 4061 2851
rect 4009 2799 4061 2843
rect 4209 3017 4261 3061
rect 4209 3009 4218 3017
rect 4218 3009 4252 3017
rect 4252 3009 4261 3017
rect 4409 3123 4418 3131
rect 4418 3123 4452 3131
rect 4452 3123 4461 3131
rect 4409 3079 4461 3123
rect 4609 3297 4661 3341
rect 4609 3289 4618 3297
rect 4618 3289 4652 3297
rect 4652 3289 4661 3297
rect 4809 3403 4818 3411
rect 4818 3403 4852 3411
rect 4852 3403 4861 3411
rect 4809 3359 4861 3403
rect 5009 3577 5061 3621
rect 5009 3569 5018 3577
rect 5018 3569 5052 3577
rect 5052 3569 5061 3577
rect 5209 3773 5218 3781
rect 5218 3773 5252 3781
rect 5252 3773 5261 3781
rect 5209 3729 5261 3773
rect 5409 3947 5461 3991
rect 5409 3939 5418 3947
rect 5418 3939 5452 3947
rect 5452 3939 5461 3947
rect 5609 4053 5618 4061
rect 5618 4053 5652 4061
rect 5652 4053 5661 4061
rect 5609 4009 5661 4053
rect 5809 4227 5861 4271
rect 5809 4219 5818 4227
rect 5818 4219 5852 4227
rect 5852 4219 5861 4227
rect 6009 4333 6018 4341
rect 6018 4333 6052 4341
rect 6052 4333 6061 4341
rect 6009 4289 6061 4333
rect 6209 4507 6261 4551
rect 6209 4499 6218 4507
rect 6218 4499 6252 4507
rect 6252 4499 6261 4507
rect 6409 4613 6418 4621
rect 6418 4613 6452 4621
rect 6452 4613 6461 4621
rect 6409 4569 6461 4613
rect 6609 4787 6661 4831
rect 6609 4779 6618 4787
rect 6618 4779 6652 4787
rect 6652 4779 6661 4787
rect 6809 4894 6861 4903
rect 6809 4860 6818 4894
rect 6818 4860 6852 4894
rect 6852 4860 6861 4894
rect 6809 4851 6861 4860
rect 5209 3684 5261 3693
rect 5209 3650 5218 3684
rect 5218 3650 5252 3684
rect 5252 3650 5261 3684
rect 5209 3641 5261 3650
rect 3609 2474 3661 2483
rect 3609 2440 3618 2474
rect 3618 2440 3652 2474
rect 3652 2440 3661 2474
rect 3609 2431 3661 2440
rect 2009 1264 2061 1273
rect 2009 1230 2018 1264
rect 2018 1230 2052 1264
rect 2052 1230 2061 1264
rect 2009 1221 2061 1230
rect 409 54 461 63
rect 409 20 418 54
rect 418 20 452 54
rect 452 20 461 54
rect 409 11 461 20
rect 309 -60 361 -15
rect 309 -67 318 -60
rect 318 -67 352 -60
rect 352 -67 361 -60
rect 109 -166 118 -143
rect 118 -166 152 -143
rect 152 -166 161 -143
rect 109 -195 161 -166
rect 125 -248 177 -239
rect 125 -282 134 -248
rect 134 -282 168 -248
rect 168 -282 177 -248
rect 125 -291 177 -282
rect 109 -363 161 -326
rect 109 -378 118 -363
rect 118 -378 152 -363
rect 152 -378 161 -363
rect 109 -397 118 -390
rect 118 -397 152 -390
rect 152 -397 161 -390
rect 109 -435 161 -397
rect 109 -442 118 -435
rect 118 -442 152 -435
rect 152 -442 161 -435
rect 109 -469 118 -454
rect 118 -469 152 -454
rect 152 -469 161 -454
rect 109 -506 161 -469
rect 309 -94 318 -79
rect 318 -94 352 -79
rect 352 -94 361 -79
rect 309 -131 361 -94
rect 409 -74 461 -22
rect 609 177 661 221
rect 609 169 618 177
rect 618 169 652 177
rect 652 169 661 177
rect 809 283 818 291
rect 818 283 852 291
rect 852 283 861 291
rect 809 239 861 283
rect 1009 457 1061 501
rect 1009 449 1018 457
rect 1018 449 1052 457
rect 1052 449 1061 457
rect 1209 563 1218 571
rect 1218 563 1252 571
rect 1252 563 1261 571
rect 1209 519 1261 563
rect 1409 737 1461 781
rect 1409 729 1418 737
rect 1418 729 1452 737
rect 1452 729 1461 737
rect 1609 843 1618 851
rect 1618 843 1652 851
rect 1652 843 1661 851
rect 1609 799 1661 843
rect 1809 1017 1861 1061
rect 1809 1009 1818 1017
rect 1818 1009 1852 1017
rect 1852 1009 1861 1017
rect 2009 1123 2018 1131
rect 2018 1123 2052 1131
rect 2052 1123 2061 1131
rect 2009 1079 2061 1123
rect 2209 1387 2261 1431
rect 2209 1379 2218 1387
rect 2218 1379 2252 1387
rect 2252 1379 2261 1387
rect 2409 1493 2418 1501
rect 2418 1493 2452 1501
rect 2452 1493 2461 1501
rect 2409 1449 2461 1493
rect 2609 1667 2661 1711
rect 2609 1659 2618 1667
rect 2618 1659 2652 1667
rect 2652 1659 2661 1667
rect 2809 1773 2818 1781
rect 2818 1773 2852 1781
rect 2852 1773 2861 1781
rect 2809 1729 2861 1773
rect 3009 1947 3061 1991
rect 3009 1939 3018 1947
rect 3018 1939 3052 1947
rect 3052 1939 3061 1947
rect 3209 2053 3218 2061
rect 3218 2053 3252 2061
rect 3252 2053 3261 2061
rect 3209 2009 3261 2053
rect 3409 2227 3461 2271
rect 3409 2219 3418 2227
rect 3418 2219 3452 2227
rect 3452 2219 3461 2227
rect 3609 2333 3618 2341
rect 3618 2333 3652 2341
rect 3652 2333 3661 2341
rect 3609 2289 3661 2333
rect 3809 2597 3861 2641
rect 3809 2589 3818 2597
rect 3818 2589 3852 2597
rect 3852 2589 3861 2597
rect 4009 2703 4018 2711
rect 4018 2703 4052 2711
rect 4052 2703 4061 2711
rect 4009 2659 4061 2703
rect 4209 2877 4261 2921
rect 4209 2869 4218 2877
rect 4218 2869 4252 2877
rect 4252 2869 4261 2877
rect 4409 2983 4418 2991
rect 4418 2983 4452 2991
rect 4452 2983 4461 2991
rect 4409 2939 4461 2983
rect 4609 3157 4661 3201
rect 4609 3149 4618 3157
rect 4618 3149 4652 3157
rect 4652 3149 4661 3157
rect 4809 3263 4818 3271
rect 4818 3263 4852 3271
rect 4852 3263 4861 3271
rect 4809 3219 4861 3263
rect 5009 3437 5061 3481
rect 5009 3429 5018 3437
rect 5018 3429 5052 3437
rect 5052 3429 5061 3437
rect 5209 3543 5218 3551
rect 5218 3543 5252 3551
rect 5252 3543 5261 3551
rect 5209 3499 5261 3543
rect 5409 3807 5461 3851
rect 5409 3799 5418 3807
rect 5418 3799 5452 3807
rect 5452 3799 5461 3807
rect 5609 3913 5618 3921
rect 5618 3913 5652 3921
rect 5652 3913 5661 3921
rect 5609 3869 5661 3913
rect 5809 4087 5861 4131
rect 5809 4079 5818 4087
rect 5818 4079 5852 4087
rect 5852 4079 5861 4087
rect 6009 4193 6018 4201
rect 6018 4193 6052 4201
rect 6052 4193 6061 4201
rect 6009 4149 6061 4193
rect 6209 4367 6261 4411
rect 6209 4359 6218 4367
rect 6218 4359 6252 4367
rect 6252 4359 6261 4367
rect 6409 4473 6418 4481
rect 6418 4473 6452 4481
rect 6452 4473 6461 4481
rect 6409 4429 6461 4473
rect 6609 4647 6661 4691
rect 6609 4639 6618 4647
rect 6618 4639 6652 4647
rect 6652 4639 6661 4647
rect 6809 4753 6818 4761
rect 6818 4753 6852 4761
rect 6852 4753 6861 4761
rect 6809 4709 6861 4753
rect 7009 4910 7061 4919
rect 7009 4876 7018 4910
rect 7018 4876 7052 4910
rect 7052 4876 7061 4910
rect 7009 4867 7061 4876
rect 5409 3700 5461 3709
rect 5409 3666 5418 3700
rect 5418 3666 5452 3700
rect 5452 3666 5461 3700
rect 5409 3657 5461 3666
rect 3809 2490 3861 2499
rect 3809 2456 3818 2490
rect 3818 2456 3852 2490
rect 3852 2456 3861 2490
rect 3809 2447 3861 2456
rect 2209 1280 2261 1289
rect 2209 1246 2218 1280
rect 2218 1246 2252 1280
rect 2252 1246 2261 1280
rect 2209 1237 2261 1246
rect 609 70 661 79
rect 609 36 618 70
rect 618 36 652 70
rect 652 36 661 70
rect 609 27 661 36
rect 509 -60 561 -15
rect 509 -67 518 -60
rect 518 -67 552 -60
rect 552 -67 561 -60
rect 309 -166 318 -143
rect 318 -166 352 -143
rect 352 -166 361 -143
rect 309 -195 361 -166
rect 325 -248 377 -239
rect 325 -282 334 -248
rect 334 -282 368 -248
rect 368 -282 377 -248
rect 325 -291 377 -282
rect 309 -363 361 -326
rect 309 -378 318 -363
rect 318 -378 352 -363
rect 352 -378 361 -363
rect 309 -397 318 -390
rect 318 -397 352 -390
rect 352 -397 361 -390
rect 309 -435 361 -397
rect 309 -442 318 -435
rect 318 -442 352 -435
rect 352 -442 361 -435
rect 309 -469 318 -454
rect 318 -469 352 -454
rect 352 -469 361 -454
rect 309 -506 361 -469
rect 509 -94 518 -79
rect 518 -94 552 -79
rect 552 -94 561 -79
rect 509 -131 561 -94
rect 609 -74 661 -22
rect 809 143 818 151
rect 818 143 852 151
rect 852 143 861 151
rect 809 99 861 143
rect 1009 317 1061 361
rect 1009 309 1018 317
rect 1018 309 1052 317
rect 1052 309 1061 317
rect 1209 423 1218 431
rect 1218 423 1252 431
rect 1252 423 1261 431
rect 1209 379 1261 423
rect 1409 597 1461 641
rect 1409 589 1418 597
rect 1418 589 1452 597
rect 1452 589 1461 597
rect 1609 703 1618 711
rect 1618 703 1652 711
rect 1652 703 1661 711
rect 1609 659 1661 703
rect 1809 877 1861 921
rect 1809 869 1818 877
rect 1818 869 1852 877
rect 1852 869 1861 877
rect 2009 983 2018 991
rect 2018 983 2052 991
rect 2052 983 2061 991
rect 2009 939 2061 983
rect 2209 1157 2261 1201
rect 2209 1149 2218 1157
rect 2218 1149 2252 1157
rect 2252 1149 2261 1157
rect 2409 1353 2418 1361
rect 2418 1353 2452 1361
rect 2452 1353 2461 1361
rect 2409 1309 2461 1353
rect 2609 1527 2661 1571
rect 2609 1519 2618 1527
rect 2618 1519 2652 1527
rect 2652 1519 2661 1527
rect 2809 1633 2818 1641
rect 2818 1633 2852 1641
rect 2852 1633 2861 1641
rect 2809 1589 2861 1633
rect 3009 1807 3061 1851
rect 3009 1799 3018 1807
rect 3018 1799 3052 1807
rect 3052 1799 3061 1807
rect 3209 1913 3218 1921
rect 3218 1913 3252 1921
rect 3252 1913 3261 1921
rect 3209 1869 3261 1913
rect 3409 2087 3461 2131
rect 3409 2079 3418 2087
rect 3418 2079 3452 2087
rect 3452 2079 3461 2087
rect 3609 2193 3618 2201
rect 3618 2193 3652 2201
rect 3652 2193 3661 2201
rect 3609 2149 3661 2193
rect 3809 2367 3861 2411
rect 3809 2359 3818 2367
rect 3818 2359 3852 2367
rect 3852 2359 3861 2367
rect 4009 2563 4018 2571
rect 4018 2563 4052 2571
rect 4052 2563 4061 2571
rect 4009 2519 4061 2563
rect 4209 2737 4261 2781
rect 4209 2729 4218 2737
rect 4218 2729 4252 2737
rect 4252 2729 4261 2737
rect 4409 2843 4418 2851
rect 4418 2843 4452 2851
rect 4452 2843 4461 2851
rect 4409 2799 4461 2843
rect 4609 3017 4661 3061
rect 4609 3009 4618 3017
rect 4618 3009 4652 3017
rect 4652 3009 4661 3017
rect 4809 3123 4818 3131
rect 4818 3123 4852 3131
rect 4852 3123 4861 3131
rect 4809 3079 4861 3123
rect 5009 3297 5061 3341
rect 5009 3289 5018 3297
rect 5018 3289 5052 3297
rect 5052 3289 5061 3297
rect 5209 3403 5218 3411
rect 5218 3403 5252 3411
rect 5252 3403 5261 3411
rect 5209 3359 5261 3403
rect 5409 3577 5461 3621
rect 5409 3569 5418 3577
rect 5418 3569 5452 3577
rect 5452 3569 5461 3577
rect 5609 3773 5618 3781
rect 5618 3773 5652 3781
rect 5652 3773 5661 3781
rect 5609 3729 5661 3773
rect 5809 3947 5861 3991
rect 5809 3939 5818 3947
rect 5818 3939 5852 3947
rect 5852 3939 5861 3947
rect 6009 4053 6018 4061
rect 6018 4053 6052 4061
rect 6052 4053 6061 4061
rect 6009 4009 6061 4053
rect 6209 4227 6261 4271
rect 6209 4219 6218 4227
rect 6218 4219 6252 4227
rect 6252 4219 6261 4227
rect 6409 4333 6418 4341
rect 6418 4333 6452 4341
rect 6452 4333 6461 4341
rect 6409 4289 6461 4333
rect 6609 4507 6661 4551
rect 6609 4499 6618 4507
rect 6618 4499 6652 4507
rect 6652 4499 6661 4507
rect 6809 4613 6818 4621
rect 6818 4613 6852 4621
rect 6852 4613 6861 4621
rect 6809 4569 6861 4613
rect 7009 4787 7061 4831
rect 7009 4779 7018 4787
rect 7018 4779 7052 4787
rect 7052 4779 7061 4787
rect 7209 4894 7261 4903
rect 7209 4860 7218 4894
rect 7218 4860 7252 4894
rect 7252 4860 7261 4894
rect 7209 4851 7261 4860
rect 5609 3684 5661 3693
rect 5609 3650 5618 3684
rect 5618 3650 5652 3684
rect 5652 3650 5661 3684
rect 5609 3641 5661 3650
rect 4009 2474 4061 2483
rect 4009 2440 4018 2474
rect 4018 2440 4052 2474
rect 4052 2440 4061 2474
rect 4009 2431 4061 2440
rect 2409 1264 2461 1273
rect 2409 1230 2418 1264
rect 2418 1230 2452 1264
rect 2452 1230 2461 1264
rect 2409 1221 2461 1230
rect 809 54 861 63
rect 809 20 818 54
rect 818 20 852 54
rect 852 20 861 54
rect 809 11 861 20
rect 709 -60 761 -15
rect 709 -67 718 -60
rect 718 -67 752 -60
rect 752 -67 761 -60
rect 509 -166 518 -143
rect 518 -166 552 -143
rect 552 -166 561 -143
rect 509 -195 561 -166
rect 525 -248 577 -239
rect 525 -282 534 -248
rect 534 -282 568 -248
rect 568 -282 577 -248
rect 525 -291 577 -282
rect 509 -363 561 -326
rect 509 -378 518 -363
rect 518 -378 552 -363
rect 552 -378 561 -363
rect 509 -397 518 -390
rect 518 -397 552 -390
rect 552 -397 561 -390
rect 509 -435 561 -397
rect 509 -442 518 -435
rect 518 -442 552 -435
rect 552 -442 561 -435
rect 509 -469 518 -454
rect 518 -469 552 -454
rect 552 -469 561 -454
rect 509 -506 561 -469
rect 709 -94 718 -79
rect 718 -94 752 -79
rect 752 -94 761 -79
rect 709 -131 761 -94
rect 809 -74 861 -22
rect 1009 177 1061 221
rect 1009 169 1018 177
rect 1018 169 1052 177
rect 1052 169 1061 177
rect 1209 283 1218 291
rect 1218 283 1252 291
rect 1252 283 1261 291
rect 1209 239 1261 283
rect 1409 457 1461 501
rect 1409 449 1418 457
rect 1418 449 1452 457
rect 1452 449 1461 457
rect 1609 563 1618 571
rect 1618 563 1652 571
rect 1652 563 1661 571
rect 1609 519 1661 563
rect 1809 737 1861 781
rect 1809 729 1818 737
rect 1818 729 1852 737
rect 1852 729 1861 737
rect 2009 843 2018 851
rect 2018 843 2052 851
rect 2052 843 2061 851
rect 2009 799 2061 843
rect 2209 1017 2261 1061
rect 2209 1009 2218 1017
rect 2218 1009 2252 1017
rect 2252 1009 2261 1017
rect 2409 1123 2418 1131
rect 2418 1123 2452 1131
rect 2452 1123 2461 1131
rect 2409 1079 2461 1123
rect 2609 1387 2661 1431
rect 2609 1379 2618 1387
rect 2618 1379 2652 1387
rect 2652 1379 2661 1387
rect 2809 1493 2818 1501
rect 2818 1493 2852 1501
rect 2852 1493 2861 1501
rect 2809 1449 2861 1493
rect 3009 1667 3061 1711
rect 3009 1659 3018 1667
rect 3018 1659 3052 1667
rect 3052 1659 3061 1667
rect 3209 1773 3218 1781
rect 3218 1773 3252 1781
rect 3252 1773 3261 1781
rect 3209 1729 3261 1773
rect 3409 1947 3461 1991
rect 3409 1939 3418 1947
rect 3418 1939 3452 1947
rect 3452 1939 3461 1947
rect 3609 2053 3618 2061
rect 3618 2053 3652 2061
rect 3652 2053 3661 2061
rect 3609 2009 3661 2053
rect 3809 2227 3861 2271
rect 3809 2219 3818 2227
rect 3818 2219 3852 2227
rect 3852 2219 3861 2227
rect 4009 2333 4018 2341
rect 4018 2333 4052 2341
rect 4052 2333 4061 2341
rect 4009 2289 4061 2333
rect 4209 2597 4261 2641
rect 4209 2589 4218 2597
rect 4218 2589 4252 2597
rect 4252 2589 4261 2597
rect 4409 2703 4418 2711
rect 4418 2703 4452 2711
rect 4452 2703 4461 2711
rect 4409 2659 4461 2703
rect 4609 2877 4661 2921
rect 4609 2869 4618 2877
rect 4618 2869 4652 2877
rect 4652 2869 4661 2877
rect 4809 2983 4818 2991
rect 4818 2983 4852 2991
rect 4852 2983 4861 2991
rect 4809 2939 4861 2983
rect 5009 3157 5061 3201
rect 5009 3149 5018 3157
rect 5018 3149 5052 3157
rect 5052 3149 5061 3157
rect 5209 3263 5218 3271
rect 5218 3263 5252 3271
rect 5252 3263 5261 3271
rect 5209 3219 5261 3263
rect 5409 3437 5461 3481
rect 5409 3429 5418 3437
rect 5418 3429 5452 3437
rect 5452 3429 5461 3437
rect 5609 3543 5618 3551
rect 5618 3543 5652 3551
rect 5652 3543 5661 3551
rect 5609 3499 5661 3543
rect 5809 3807 5861 3851
rect 5809 3799 5818 3807
rect 5818 3799 5852 3807
rect 5852 3799 5861 3807
rect 6009 3913 6018 3921
rect 6018 3913 6052 3921
rect 6052 3913 6061 3921
rect 6009 3869 6061 3913
rect 6209 4087 6261 4131
rect 6209 4079 6218 4087
rect 6218 4079 6252 4087
rect 6252 4079 6261 4087
rect 6409 4193 6418 4201
rect 6418 4193 6452 4201
rect 6452 4193 6461 4201
rect 6409 4149 6461 4193
rect 6609 4367 6661 4411
rect 6609 4359 6618 4367
rect 6618 4359 6652 4367
rect 6652 4359 6661 4367
rect 6809 4473 6818 4481
rect 6818 4473 6852 4481
rect 6852 4473 6861 4481
rect 6809 4429 6861 4473
rect 7009 4647 7061 4691
rect 7009 4639 7018 4647
rect 7018 4639 7052 4647
rect 7052 4639 7061 4647
rect 7209 4753 7218 4761
rect 7218 4753 7252 4761
rect 7252 4753 7261 4761
rect 7209 4709 7261 4753
rect 7409 4910 7461 4919
rect 7409 4876 7418 4910
rect 7418 4876 7452 4910
rect 7452 4876 7461 4910
rect 7409 4867 7461 4876
rect 5809 3700 5861 3709
rect 5809 3666 5818 3700
rect 5818 3666 5852 3700
rect 5852 3666 5861 3700
rect 5809 3657 5861 3666
rect 4209 2490 4261 2499
rect 4209 2456 4218 2490
rect 4218 2456 4252 2490
rect 4252 2456 4261 2490
rect 4209 2447 4261 2456
rect 2609 1280 2661 1289
rect 2609 1246 2618 1280
rect 2618 1246 2652 1280
rect 2652 1246 2661 1280
rect 2609 1237 2661 1246
rect 1009 70 1061 79
rect 1009 36 1018 70
rect 1018 36 1052 70
rect 1052 36 1061 70
rect 1009 27 1061 36
rect 909 -60 961 -15
rect 909 -67 918 -60
rect 918 -67 952 -60
rect 952 -67 961 -60
rect 709 -166 718 -143
rect 718 -166 752 -143
rect 752 -166 761 -143
rect 709 -195 761 -166
rect 725 -248 777 -239
rect 725 -282 734 -248
rect 734 -282 768 -248
rect 768 -282 777 -248
rect 725 -291 777 -282
rect 709 -363 761 -326
rect 709 -378 718 -363
rect 718 -378 752 -363
rect 752 -378 761 -363
rect 709 -397 718 -390
rect 718 -397 752 -390
rect 752 -397 761 -390
rect 709 -435 761 -397
rect 709 -442 718 -435
rect 718 -442 752 -435
rect 752 -442 761 -435
rect 709 -469 718 -454
rect 718 -469 752 -454
rect 752 -469 761 -454
rect 709 -506 761 -469
rect 909 -94 918 -79
rect 918 -94 952 -79
rect 952 -94 961 -79
rect 909 -131 961 -94
rect 1009 -74 1061 -22
rect 1209 143 1218 151
rect 1218 143 1252 151
rect 1252 143 1261 151
rect 1209 99 1261 143
rect 1409 317 1461 361
rect 1409 309 1418 317
rect 1418 309 1452 317
rect 1452 309 1461 317
rect 1609 423 1618 431
rect 1618 423 1652 431
rect 1652 423 1661 431
rect 1609 379 1661 423
rect 1809 597 1861 641
rect 1809 589 1818 597
rect 1818 589 1852 597
rect 1852 589 1861 597
rect 2009 703 2018 711
rect 2018 703 2052 711
rect 2052 703 2061 711
rect 2009 659 2061 703
rect 2209 877 2261 921
rect 2209 869 2218 877
rect 2218 869 2252 877
rect 2252 869 2261 877
rect 2409 983 2418 991
rect 2418 983 2452 991
rect 2452 983 2461 991
rect 2409 939 2461 983
rect 2609 1157 2661 1201
rect 2609 1149 2618 1157
rect 2618 1149 2652 1157
rect 2652 1149 2661 1157
rect 2809 1353 2818 1361
rect 2818 1353 2852 1361
rect 2852 1353 2861 1361
rect 2809 1309 2861 1353
rect 3009 1527 3061 1571
rect 3009 1519 3018 1527
rect 3018 1519 3052 1527
rect 3052 1519 3061 1527
rect 3209 1633 3218 1641
rect 3218 1633 3252 1641
rect 3252 1633 3261 1641
rect 3209 1589 3261 1633
rect 3409 1807 3461 1851
rect 3409 1799 3418 1807
rect 3418 1799 3452 1807
rect 3452 1799 3461 1807
rect 3609 1913 3618 1921
rect 3618 1913 3652 1921
rect 3652 1913 3661 1921
rect 3609 1869 3661 1913
rect 3809 2087 3861 2131
rect 3809 2079 3818 2087
rect 3818 2079 3852 2087
rect 3852 2079 3861 2087
rect 4009 2193 4018 2201
rect 4018 2193 4052 2201
rect 4052 2193 4061 2201
rect 4009 2149 4061 2193
rect 4209 2367 4261 2411
rect 4209 2359 4218 2367
rect 4218 2359 4252 2367
rect 4252 2359 4261 2367
rect 4409 2563 4418 2571
rect 4418 2563 4452 2571
rect 4452 2563 4461 2571
rect 4409 2519 4461 2563
rect 4609 2737 4661 2781
rect 4609 2729 4618 2737
rect 4618 2729 4652 2737
rect 4652 2729 4661 2737
rect 4809 2843 4818 2851
rect 4818 2843 4852 2851
rect 4852 2843 4861 2851
rect 4809 2799 4861 2843
rect 5009 3017 5061 3061
rect 5009 3009 5018 3017
rect 5018 3009 5052 3017
rect 5052 3009 5061 3017
rect 5209 3123 5218 3131
rect 5218 3123 5252 3131
rect 5252 3123 5261 3131
rect 5209 3079 5261 3123
rect 5409 3297 5461 3341
rect 5409 3289 5418 3297
rect 5418 3289 5452 3297
rect 5452 3289 5461 3297
rect 5609 3403 5618 3411
rect 5618 3403 5652 3411
rect 5652 3403 5661 3411
rect 5609 3359 5661 3403
rect 5809 3577 5861 3621
rect 5809 3569 5818 3577
rect 5818 3569 5852 3577
rect 5852 3569 5861 3577
rect 6009 3773 6018 3781
rect 6018 3773 6052 3781
rect 6052 3773 6061 3781
rect 6009 3729 6061 3773
rect 6209 3947 6261 3991
rect 6209 3939 6218 3947
rect 6218 3939 6252 3947
rect 6252 3939 6261 3947
rect 6409 4053 6418 4061
rect 6418 4053 6452 4061
rect 6452 4053 6461 4061
rect 6409 4009 6461 4053
rect 6609 4227 6661 4271
rect 6609 4219 6618 4227
rect 6618 4219 6652 4227
rect 6652 4219 6661 4227
rect 6809 4333 6818 4341
rect 6818 4333 6852 4341
rect 6852 4333 6861 4341
rect 6809 4289 6861 4333
rect 7009 4507 7061 4551
rect 7009 4499 7018 4507
rect 7018 4499 7052 4507
rect 7052 4499 7061 4507
rect 7209 4613 7218 4621
rect 7218 4613 7252 4621
rect 7252 4613 7261 4621
rect 7209 4569 7261 4613
rect 7409 4787 7461 4831
rect 7409 4779 7418 4787
rect 7418 4779 7452 4787
rect 7452 4779 7461 4787
rect 7609 4894 7661 4903
rect 7609 4860 7618 4894
rect 7618 4860 7652 4894
rect 7652 4860 7661 4894
rect 7609 4851 7661 4860
rect 6009 3684 6061 3693
rect 6009 3650 6018 3684
rect 6018 3650 6052 3684
rect 6052 3650 6061 3684
rect 6009 3641 6061 3650
rect 4409 2474 4461 2483
rect 4409 2440 4418 2474
rect 4418 2440 4452 2474
rect 4452 2440 4461 2474
rect 4409 2431 4461 2440
rect 2809 1264 2861 1273
rect 2809 1230 2818 1264
rect 2818 1230 2852 1264
rect 2852 1230 2861 1264
rect 2809 1221 2861 1230
rect 1209 54 1261 63
rect 1209 20 1218 54
rect 1218 20 1252 54
rect 1252 20 1261 54
rect 1209 11 1261 20
rect 1109 -60 1161 -15
rect 1109 -67 1118 -60
rect 1118 -67 1152 -60
rect 1152 -67 1161 -60
rect 909 -166 918 -143
rect 918 -166 952 -143
rect 952 -166 961 -143
rect 909 -195 961 -166
rect 925 -248 977 -239
rect 925 -282 934 -248
rect 934 -282 968 -248
rect 968 -282 977 -248
rect 925 -291 977 -282
rect 909 -363 961 -326
rect 909 -378 918 -363
rect 918 -378 952 -363
rect 952 -378 961 -363
rect 909 -397 918 -390
rect 918 -397 952 -390
rect 952 -397 961 -390
rect 909 -435 961 -397
rect 909 -442 918 -435
rect 918 -442 952 -435
rect 952 -442 961 -435
rect 909 -469 918 -454
rect 918 -469 952 -454
rect 952 -469 961 -454
rect 909 -506 961 -469
rect 1109 -94 1118 -79
rect 1118 -94 1152 -79
rect 1152 -94 1161 -79
rect 1109 -131 1161 -94
rect 1209 -74 1261 -22
rect 1409 177 1461 221
rect 1409 169 1418 177
rect 1418 169 1452 177
rect 1452 169 1461 177
rect 1609 283 1618 291
rect 1618 283 1652 291
rect 1652 283 1661 291
rect 1609 239 1661 283
rect 1809 457 1861 501
rect 1809 449 1818 457
rect 1818 449 1852 457
rect 1852 449 1861 457
rect 2009 563 2018 571
rect 2018 563 2052 571
rect 2052 563 2061 571
rect 2009 519 2061 563
rect 2209 737 2261 781
rect 2209 729 2218 737
rect 2218 729 2252 737
rect 2252 729 2261 737
rect 2409 843 2418 851
rect 2418 843 2452 851
rect 2452 843 2461 851
rect 2409 799 2461 843
rect 2609 1017 2661 1061
rect 2609 1009 2618 1017
rect 2618 1009 2652 1017
rect 2652 1009 2661 1017
rect 2809 1123 2818 1131
rect 2818 1123 2852 1131
rect 2852 1123 2861 1131
rect 2809 1079 2861 1123
rect 3009 1387 3061 1431
rect 3009 1379 3018 1387
rect 3018 1379 3052 1387
rect 3052 1379 3061 1387
rect 3209 1493 3218 1501
rect 3218 1493 3252 1501
rect 3252 1493 3261 1501
rect 3209 1449 3261 1493
rect 3409 1667 3461 1711
rect 3409 1659 3418 1667
rect 3418 1659 3452 1667
rect 3452 1659 3461 1667
rect 3609 1773 3618 1781
rect 3618 1773 3652 1781
rect 3652 1773 3661 1781
rect 3609 1729 3661 1773
rect 3809 1947 3861 1991
rect 3809 1939 3818 1947
rect 3818 1939 3852 1947
rect 3852 1939 3861 1947
rect 4009 2053 4018 2061
rect 4018 2053 4052 2061
rect 4052 2053 4061 2061
rect 4009 2009 4061 2053
rect 4209 2227 4261 2271
rect 4209 2219 4218 2227
rect 4218 2219 4252 2227
rect 4252 2219 4261 2227
rect 4409 2333 4418 2341
rect 4418 2333 4452 2341
rect 4452 2333 4461 2341
rect 4409 2289 4461 2333
rect 4609 2597 4661 2641
rect 4609 2589 4618 2597
rect 4618 2589 4652 2597
rect 4652 2589 4661 2597
rect 4809 2703 4818 2711
rect 4818 2703 4852 2711
rect 4852 2703 4861 2711
rect 4809 2659 4861 2703
rect 5009 2877 5061 2921
rect 5009 2869 5018 2877
rect 5018 2869 5052 2877
rect 5052 2869 5061 2877
rect 5209 2983 5218 2991
rect 5218 2983 5252 2991
rect 5252 2983 5261 2991
rect 5209 2939 5261 2983
rect 5409 3157 5461 3201
rect 5409 3149 5418 3157
rect 5418 3149 5452 3157
rect 5452 3149 5461 3157
rect 5609 3263 5618 3271
rect 5618 3263 5652 3271
rect 5652 3263 5661 3271
rect 5609 3219 5661 3263
rect 5809 3437 5861 3481
rect 5809 3429 5818 3437
rect 5818 3429 5852 3437
rect 5852 3429 5861 3437
rect 6009 3543 6018 3551
rect 6018 3543 6052 3551
rect 6052 3543 6061 3551
rect 6009 3499 6061 3543
rect 6209 3807 6261 3851
rect 6209 3799 6218 3807
rect 6218 3799 6252 3807
rect 6252 3799 6261 3807
rect 6409 3913 6418 3921
rect 6418 3913 6452 3921
rect 6452 3913 6461 3921
rect 6409 3869 6461 3913
rect 6609 4087 6661 4131
rect 6609 4079 6618 4087
rect 6618 4079 6652 4087
rect 6652 4079 6661 4087
rect 6809 4193 6818 4201
rect 6818 4193 6852 4201
rect 6852 4193 6861 4201
rect 6809 4149 6861 4193
rect 7009 4367 7061 4411
rect 7009 4359 7018 4367
rect 7018 4359 7052 4367
rect 7052 4359 7061 4367
rect 7209 4473 7218 4481
rect 7218 4473 7252 4481
rect 7252 4473 7261 4481
rect 7209 4429 7261 4473
rect 7409 4647 7461 4691
rect 7409 4639 7418 4647
rect 7418 4639 7452 4647
rect 7452 4639 7461 4647
rect 7609 4753 7618 4761
rect 7618 4753 7652 4761
rect 7652 4753 7661 4761
rect 7609 4709 7661 4753
rect 7809 4910 7861 4919
rect 7809 4876 7818 4910
rect 7818 4876 7852 4910
rect 7852 4876 7861 4910
rect 7809 4867 7861 4876
rect 6209 3700 6261 3709
rect 6209 3666 6218 3700
rect 6218 3666 6252 3700
rect 6252 3666 6261 3700
rect 6209 3657 6261 3666
rect 4609 2490 4661 2499
rect 4609 2456 4618 2490
rect 4618 2456 4652 2490
rect 4652 2456 4661 2490
rect 4609 2447 4661 2456
rect 3009 1280 3061 1289
rect 3009 1246 3018 1280
rect 3018 1246 3052 1280
rect 3052 1246 3061 1280
rect 3009 1237 3061 1246
rect 1409 70 1461 79
rect 1409 36 1418 70
rect 1418 36 1452 70
rect 1452 36 1461 70
rect 1409 27 1461 36
rect 1309 -60 1361 -15
rect 1309 -67 1318 -60
rect 1318 -67 1352 -60
rect 1352 -67 1361 -60
rect 1109 -166 1118 -143
rect 1118 -166 1152 -143
rect 1152 -166 1161 -143
rect 1109 -195 1161 -166
rect 1125 -248 1177 -239
rect 1125 -282 1134 -248
rect 1134 -282 1168 -248
rect 1168 -282 1177 -248
rect 1125 -291 1177 -282
rect 1109 -363 1161 -326
rect 1109 -378 1118 -363
rect 1118 -378 1152 -363
rect 1152 -378 1161 -363
rect 1109 -397 1118 -390
rect 1118 -397 1152 -390
rect 1152 -397 1161 -390
rect 1109 -435 1161 -397
rect 1109 -442 1118 -435
rect 1118 -442 1152 -435
rect 1152 -442 1161 -435
rect 1109 -469 1118 -454
rect 1118 -469 1152 -454
rect 1152 -469 1161 -454
rect 1109 -506 1161 -469
rect 1309 -94 1318 -79
rect 1318 -94 1352 -79
rect 1352 -94 1361 -79
rect 1309 -131 1361 -94
rect 1409 -74 1461 -22
rect 1609 143 1618 151
rect 1618 143 1652 151
rect 1652 143 1661 151
rect 1609 99 1661 143
rect 1809 317 1861 361
rect 1809 309 1818 317
rect 1818 309 1852 317
rect 1852 309 1861 317
rect 2009 423 2018 431
rect 2018 423 2052 431
rect 2052 423 2061 431
rect 2009 379 2061 423
rect 2209 597 2261 641
rect 2209 589 2218 597
rect 2218 589 2252 597
rect 2252 589 2261 597
rect 2409 703 2418 711
rect 2418 703 2452 711
rect 2452 703 2461 711
rect 2409 659 2461 703
rect 2609 877 2661 921
rect 2609 869 2618 877
rect 2618 869 2652 877
rect 2652 869 2661 877
rect 2809 983 2818 991
rect 2818 983 2852 991
rect 2852 983 2861 991
rect 2809 939 2861 983
rect 3009 1157 3061 1201
rect 3009 1149 3018 1157
rect 3018 1149 3052 1157
rect 3052 1149 3061 1157
rect 3209 1353 3218 1361
rect 3218 1353 3252 1361
rect 3252 1353 3261 1361
rect 3209 1309 3261 1353
rect 3409 1527 3461 1571
rect 3409 1519 3418 1527
rect 3418 1519 3452 1527
rect 3452 1519 3461 1527
rect 3609 1633 3618 1641
rect 3618 1633 3652 1641
rect 3652 1633 3661 1641
rect 3609 1589 3661 1633
rect 3809 1807 3861 1851
rect 3809 1799 3818 1807
rect 3818 1799 3852 1807
rect 3852 1799 3861 1807
rect 4009 1913 4018 1921
rect 4018 1913 4052 1921
rect 4052 1913 4061 1921
rect 4009 1869 4061 1913
rect 4209 2087 4261 2131
rect 4209 2079 4218 2087
rect 4218 2079 4252 2087
rect 4252 2079 4261 2087
rect 4409 2193 4418 2201
rect 4418 2193 4452 2201
rect 4452 2193 4461 2201
rect 4409 2149 4461 2193
rect 4609 2367 4661 2411
rect 4609 2359 4618 2367
rect 4618 2359 4652 2367
rect 4652 2359 4661 2367
rect 4809 2563 4818 2571
rect 4818 2563 4852 2571
rect 4852 2563 4861 2571
rect 4809 2519 4861 2563
rect 5009 2737 5061 2781
rect 5009 2729 5018 2737
rect 5018 2729 5052 2737
rect 5052 2729 5061 2737
rect 5209 2843 5218 2851
rect 5218 2843 5252 2851
rect 5252 2843 5261 2851
rect 5209 2799 5261 2843
rect 5409 3017 5461 3061
rect 5409 3009 5418 3017
rect 5418 3009 5452 3017
rect 5452 3009 5461 3017
rect 5609 3123 5618 3131
rect 5618 3123 5652 3131
rect 5652 3123 5661 3131
rect 5609 3079 5661 3123
rect 5809 3297 5861 3341
rect 5809 3289 5818 3297
rect 5818 3289 5852 3297
rect 5852 3289 5861 3297
rect 6009 3403 6018 3411
rect 6018 3403 6052 3411
rect 6052 3403 6061 3411
rect 6009 3359 6061 3403
rect 6209 3577 6261 3621
rect 6209 3569 6218 3577
rect 6218 3569 6252 3577
rect 6252 3569 6261 3577
rect 6409 3773 6418 3781
rect 6418 3773 6452 3781
rect 6452 3773 6461 3781
rect 6409 3729 6461 3773
rect 6609 3947 6661 3991
rect 6609 3939 6618 3947
rect 6618 3939 6652 3947
rect 6652 3939 6661 3947
rect 6809 4053 6818 4061
rect 6818 4053 6852 4061
rect 6852 4053 6861 4061
rect 6809 4009 6861 4053
rect 7009 4227 7061 4271
rect 7009 4219 7018 4227
rect 7018 4219 7052 4227
rect 7052 4219 7061 4227
rect 7209 4333 7218 4341
rect 7218 4333 7252 4341
rect 7252 4333 7261 4341
rect 7209 4289 7261 4333
rect 7409 4507 7461 4551
rect 7409 4499 7418 4507
rect 7418 4499 7452 4507
rect 7452 4499 7461 4507
rect 7609 4613 7618 4621
rect 7618 4613 7652 4621
rect 7652 4613 7661 4621
rect 7609 4569 7661 4613
rect 7809 4787 7861 4831
rect 7809 4779 7818 4787
rect 7818 4779 7852 4787
rect 7852 4779 7861 4787
rect 8009 4894 8061 4903
rect 8009 4860 8018 4894
rect 8018 4860 8052 4894
rect 8052 4860 8061 4894
rect 8009 4851 8061 4860
rect 6409 3684 6461 3693
rect 6409 3650 6418 3684
rect 6418 3650 6452 3684
rect 6452 3650 6461 3684
rect 6409 3641 6461 3650
rect 4809 2474 4861 2483
rect 4809 2440 4818 2474
rect 4818 2440 4852 2474
rect 4852 2440 4861 2474
rect 4809 2431 4861 2440
rect 3209 1264 3261 1273
rect 3209 1230 3218 1264
rect 3218 1230 3252 1264
rect 3252 1230 3261 1264
rect 3209 1221 3261 1230
rect 1609 54 1661 63
rect 1609 20 1618 54
rect 1618 20 1652 54
rect 1652 20 1661 54
rect 1609 11 1661 20
rect 1509 -60 1561 -15
rect 1509 -67 1518 -60
rect 1518 -67 1552 -60
rect 1552 -67 1561 -60
rect 1309 -166 1318 -143
rect 1318 -166 1352 -143
rect 1352 -166 1361 -143
rect 1309 -195 1361 -166
rect 1325 -248 1377 -239
rect 1325 -282 1334 -248
rect 1334 -282 1368 -248
rect 1368 -282 1377 -248
rect 1325 -291 1377 -282
rect 1309 -363 1361 -326
rect 1309 -378 1318 -363
rect 1318 -378 1352 -363
rect 1352 -378 1361 -363
rect 1309 -397 1318 -390
rect 1318 -397 1352 -390
rect 1352 -397 1361 -390
rect 1309 -435 1361 -397
rect 1309 -442 1318 -435
rect 1318 -442 1352 -435
rect 1352 -442 1361 -435
rect 1309 -469 1318 -454
rect 1318 -469 1352 -454
rect 1352 -469 1361 -454
rect 1309 -506 1361 -469
rect 1509 -94 1518 -79
rect 1518 -94 1552 -79
rect 1552 -94 1561 -79
rect 1509 -131 1561 -94
rect 1609 -74 1661 -22
rect 1809 177 1861 221
rect 1809 169 1818 177
rect 1818 169 1852 177
rect 1852 169 1861 177
rect 2009 283 2018 291
rect 2018 283 2052 291
rect 2052 283 2061 291
rect 2009 239 2061 283
rect 2209 457 2261 501
rect 2209 449 2218 457
rect 2218 449 2252 457
rect 2252 449 2261 457
rect 2409 563 2418 571
rect 2418 563 2452 571
rect 2452 563 2461 571
rect 2409 519 2461 563
rect 2609 737 2661 781
rect 2609 729 2618 737
rect 2618 729 2652 737
rect 2652 729 2661 737
rect 2809 843 2818 851
rect 2818 843 2852 851
rect 2852 843 2861 851
rect 2809 799 2861 843
rect 3009 1017 3061 1061
rect 3009 1009 3018 1017
rect 3018 1009 3052 1017
rect 3052 1009 3061 1017
rect 3209 1123 3218 1131
rect 3218 1123 3252 1131
rect 3252 1123 3261 1131
rect 3209 1079 3261 1123
rect 3409 1387 3461 1431
rect 3409 1379 3418 1387
rect 3418 1379 3452 1387
rect 3452 1379 3461 1387
rect 3609 1493 3618 1501
rect 3618 1493 3652 1501
rect 3652 1493 3661 1501
rect 3609 1449 3661 1493
rect 3809 1667 3861 1711
rect 3809 1659 3818 1667
rect 3818 1659 3852 1667
rect 3852 1659 3861 1667
rect 4009 1773 4018 1781
rect 4018 1773 4052 1781
rect 4052 1773 4061 1781
rect 4009 1729 4061 1773
rect 4209 1947 4261 1991
rect 4209 1939 4218 1947
rect 4218 1939 4252 1947
rect 4252 1939 4261 1947
rect 4409 2053 4418 2061
rect 4418 2053 4452 2061
rect 4452 2053 4461 2061
rect 4409 2009 4461 2053
rect 4609 2227 4661 2271
rect 4609 2219 4618 2227
rect 4618 2219 4652 2227
rect 4652 2219 4661 2227
rect 4809 2333 4818 2341
rect 4818 2333 4852 2341
rect 4852 2333 4861 2341
rect 4809 2289 4861 2333
rect 5009 2597 5061 2641
rect 5009 2589 5018 2597
rect 5018 2589 5052 2597
rect 5052 2589 5061 2597
rect 5209 2703 5218 2711
rect 5218 2703 5252 2711
rect 5252 2703 5261 2711
rect 5209 2659 5261 2703
rect 5409 2877 5461 2921
rect 5409 2869 5418 2877
rect 5418 2869 5452 2877
rect 5452 2869 5461 2877
rect 5609 2983 5618 2991
rect 5618 2983 5652 2991
rect 5652 2983 5661 2991
rect 5609 2939 5661 2983
rect 5809 3157 5861 3201
rect 5809 3149 5818 3157
rect 5818 3149 5852 3157
rect 5852 3149 5861 3157
rect 6009 3263 6018 3271
rect 6018 3263 6052 3271
rect 6052 3263 6061 3271
rect 6009 3219 6061 3263
rect 6209 3437 6261 3481
rect 6209 3429 6218 3437
rect 6218 3429 6252 3437
rect 6252 3429 6261 3437
rect 6409 3543 6418 3551
rect 6418 3543 6452 3551
rect 6452 3543 6461 3551
rect 6409 3499 6461 3543
rect 6609 3807 6661 3851
rect 6609 3799 6618 3807
rect 6618 3799 6652 3807
rect 6652 3799 6661 3807
rect 6809 3913 6818 3921
rect 6818 3913 6852 3921
rect 6852 3913 6861 3921
rect 6809 3869 6861 3913
rect 7009 4087 7061 4131
rect 7009 4079 7018 4087
rect 7018 4079 7052 4087
rect 7052 4079 7061 4087
rect 7209 4193 7218 4201
rect 7218 4193 7252 4201
rect 7252 4193 7261 4201
rect 7209 4149 7261 4193
rect 7409 4367 7461 4411
rect 7409 4359 7418 4367
rect 7418 4359 7452 4367
rect 7452 4359 7461 4367
rect 7609 4473 7618 4481
rect 7618 4473 7652 4481
rect 7652 4473 7661 4481
rect 7609 4429 7661 4473
rect 7809 4647 7861 4691
rect 7809 4639 7818 4647
rect 7818 4639 7852 4647
rect 7852 4639 7861 4647
rect 8009 4753 8018 4761
rect 8018 4753 8052 4761
rect 8052 4753 8061 4761
rect 8009 4709 8061 4753
rect 8209 4910 8261 4919
rect 8209 4876 8218 4910
rect 8218 4876 8252 4910
rect 8252 4876 8261 4910
rect 8209 4867 8261 4876
rect 6609 3700 6661 3709
rect 6609 3666 6618 3700
rect 6618 3666 6652 3700
rect 6652 3666 6661 3700
rect 6609 3657 6661 3666
rect 5009 2490 5061 2499
rect 5009 2456 5018 2490
rect 5018 2456 5052 2490
rect 5052 2456 5061 2490
rect 5009 2447 5061 2456
rect 3409 1280 3461 1289
rect 3409 1246 3418 1280
rect 3418 1246 3452 1280
rect 3452 1246 3461 1280
rect 3409 1237 3461 1246
rect 1809 70 1861 79
rect 1809 36 1818 70
rect 1818 36 1852 70
rect 1852 36 1861 70
rect 1809 27 1861 36
rect 1709 -60 1761 -15
rect 1709 -67 1718 -60
rect 1718 -67 1752 -60
rect 1752 -67 1761 -60
rect 1509 -166 1518 -143
rect 1518 -166 1552 -143
rect 1552 -166 1561 -143
rect 1509 -195 1561 -166
rect 1525 -248 1577 -239
rect 1525 -282 1534 -248
rect 1534 -282 1568 -248
rect 1568 -282 1577 -248
rect 1525 -291 1577 -282
rect 1509 -363 1561 -326
rect 1509 -378 1518 -363
rect 1518 -378 1552 -363
rect 1552 -378 1561 -363
rect 1509 -397 1518 -390
rect 1518 -397 1552 -390
rect 1552 -397 1561 -390
rect 1509 -435 1561 -397
rect 1509 -442 1518 -435
rect 1518 -442 1552 -435
rect 1552 -442 1561 -435
rect 1509 -469 1518 -454
rect 1518 -469 1552 -454
rect 1552 -469 1561 -454
rect 1509 -506 1561 -469
rect 1709 -94 1718 -79
rect 1718 -94 1752 -79
rect 1752 -94 1761 -79
rect 1709 -131 1761 -94
rect 1809 -74 1861 -22
rect 2009 143 2018 151
rect 2018 143 2052 151
rect 2052 143 2061 151
rect 2009 99 2061 143
rect 2209 317 2261 361
rect 2209 309 2218 317
rect 2218 309 2252 317
rect 2252 309 2261 317
rect 2409 423 2418 431
rect 2418 423 2452 431
rect 2452 423 2461 431
rect 2409 379 2461 423
rect 2609 597 2661 641
rect 2609 589 2618 597
rect 2618 589 2652 597
rect 2652 589 2661 597
rect 2809 703 2818 711
rect 2818 703 2852 711
rect 2852 703 2861 711
rect 2809 659 2861 703
rect 3009 877 3061 921
rect 3009 869 3018 877
rect 3018 869 3052 877
rect 3052 869 3061 877
rect 3209 983 3218 991
rect 3218 983 3252 991
rect 3252 983 3261 991
rect 3209 939 3261 983
rect 3409 1157 3461 1201
rect 3409 1149 3418 1157
rect 3418 1149 3452 1157
rect 3452 1149 3461 1157
rect 3609 1353 3618 1361
rect 3618 1353 3652 1361
rect 3652 1353 3661 1361
rect 3609 1309 3661 1353
rect 3809 1527 3861 1571
rect 3809 1519 3818 1527
rect 3818 1519 3852 1527
rect 3852 1519 3861 1527
rect 4009 1633 4018 1641
rect 4018 1633 4052 1641
rect 4052 1633 4061 1641
rect 4009 1589 4061 1633
rect 4209 1807 4261 1851
rect 4209 1799 4218 1807
rect 4218 1799 4252 1807
rect 4252 1799 4261 1807
rect 4409 1913 4418 1921
rect 4418 1913 4452 1921
rect 4452 1913 4461 1921
rect 4409 1869 4461 1913
rect 4609 2087 4661 2131
rect 4609 2079 4618 2087
rect 4618 2079 4652 2087
rect 4652 2079 4661 2087
rect 4809 2193 4818 2201
rect 4818 2193 4852 2201
rect 4852 2193 4861 2201
rect 4809 2149 4861 2193
rect 5009 2367 5061 2411
rect 5009 2359 5018 2367
rect 5018 2359 5052 2367
rect 5052 2359 5061 2367
rect 5209 2563 5218 2571
rect 5218 2563 5252 2571
rect 5252 2563 5261 2571
rect 5209 2519 5261 2563
rect 5409 2737 5461 2781
rect 5409 2729 5418 2737
rect 5418 2729 5452 2737
rect 5452 2729 5461 2737
rect 5609 2843 5618 2851
rect 5618 2843 5652 2851
rect 5652 2843 5661 2851
rect 5609 2799 5661 2843
rect 5809 3017 5861 3061
rect 5809 3009 5818 3017
rect 5818 3009 5852 3017
rect 5852 3009 5861 3017
rect 6009 3123 6018 3131
rect 6018 3123 6052 3131
rect 6052 3123 6061 3131
rect 6009 3079 6061 3123
rect 6209 3297 6261 3341
rect 6209 3289 6218 3297
rect 6218 3289 6252 3297
rect 6252 3289 6261 3297
rect 6409 3403 6418 3411
rect 6418 3403 6452 3411
rect 6452 3403 6461 3411
rect 6409 3359 6461 3403
rect 6609 3577 6661 3621
rect 6609 3569 6618 3577
rect 6618 3569 6652 3577
rect 6652 3569 6661 3577
rect 6809 3773 6818 3781
rect 6818 3773 6852 3781
rect 6852 3773 6861 3781
rect 6809 3729 6861 3773
rect 7009 3947 7061 3991
rect 7009 3939 7018 3947
rect 7018 3939 7052 3947
rect 7052 3939 7061 3947
rect 7209 4053 7218 4061
rect 7218 4053 7252 4061
rect 7252 4053 7261 4061
rect 7209 4009 7261 4053
rect 7409 4227 7461 4271
rect 7409 4219 7418 4227
rect 7418 4219 7452 4227
rect 7452 4219 7461 4227
rect 7609 4333 7618 4341
rect 7618 4333 7652 4341
rect 7652 4333 7661 4341
rect 7609 4289 7661 4333
rect 7809 4507 7861 4551
rect 7809 4499 7818 4507
rect 7818 4499 7852 4507
rect 7852 4499 7861 4507
rect 8009 4613 8018 4621
rect 8018 4613 8052 4621
rect 8052 4613 8061 4621
rect 8009 4569 8061 4613
rect 8209 4787 8261 4831
rect 8209 4779 8218 4787
rect 8218 4779 8252 4787
rect 8252 4779 8261 4787
rect 8409 4894 8461 4903
rect 8409 4860 8418 4894
rect 8418 4860 8452 4894
rect 8452 4860 8461 4894
rect 8409 4851 8461 4860
rect 6809 3684 6861 3693
rect 6809 3650 6818 3684
rect 6818 3650 6852 3684
rect 6852 3650 6861 3684
rect 6809 3641 6861 3650
rect 5209 2474 5261 2483
rect 5209 2440 5218 2474
rect 5218 2440 5252 2474
rect 5252 2440 5261 2474
rect 5209 2431 5261 2440
rect 3609 1264 3661 1273
rect 3609 1230 3618 1264
rect 3618 1230 3652 1264
rect 3652 1230 3661 1264
rect 3609 1221 3661 1230
rect 2009 54 2061 63
rect 2009 20 2018 54
rect 2018 20 2052 54
rect 2052 20 2061 54
rect 2009 11 2061 20
rect 1909 -60 1961 -15
rect 1909 -67 1918 -60
rect 1918 -67 1952 -60
rect 1952 -67 1961 -60
rect 1709 -166 1718 -143
rect 1718 -166 1752 -143
rect 1752 -166 1761 -143
rect 1709 -195 1761 -166
rect 1725 -248 1777 -239
rect 1725 -282 1734 -248
rect 1734 -282 1768 -248
rect 1768 -282 1777 -248
rect 1725 -291 1777 -282
rect 1709 -363 1761 -326
rect 1709 -378 1718 -363
rect 1718 -378 1752 -363
rect 1752 -378 1761 -363
rect 1709 -397 1718 -390
rect 1718 -397 1752 -390
rect 1752 -397 1761 -390
rect 1709 -435 1761 -397
rect 1709 -442 1718 -435
rect 1718 -442 1752 -435
rect 1752 -442 1761 -435
rect 1709 -469 1718 -454
rect 1718 -469 1752 -454
rect 1752 -469 1761 -454
rect 1709 -506 1761 -469
rect 1909 -94 1918 -79
rect 1918 -94 1952 -79
rect 1952 -94 1961 -79
rect 1909 -131 1961 -94
rect 2009 -74 2061 -22
rect 2209 177 2261 221
rect 2209 169 2218 177
rect 2218 169 2252 177
rect 2252 169 2261 177
rect 2409 283 2418 291
rect 2418 283 2452 291
rect 2452 283 2461 291
rect 2409 239 2461 283
rect 2609 457 2661 501
rect 2609 449 2618 457
rect 2618 449 2652 457
rect 2652 449 2661 457
rect 2809 563 2818 571
rect 2818 563 2852 571
rect 2852 563 2861 571
rect 2809 519 2861 563
rect 3009 737 3061 781
rect 3009 729 3018 737
rect 3018 729 3052 737
rect 3052 729 3061 737
rect 3209 843 3218 851
rect 3218 843 3252 851
rect 3252 843 3261 851
rect 3209 799 3261 843
rect 3409 1017 3461 1061
rect 3409 1009 3418 1017
rect 3418 1009 3452 1017
rect 3452 1009 3461 1017
rect 3609 1123 3618 1131
rect 3618 1123 3652 1131
rect 3652 1123 3661 1131
rect 3609 1079 3661 1123
rect 3809 1387 3861 1431
rect 3809 1379 3818 1387
rect 3818 1379 3852 1387
rect 3852 1379 3861 1387
rect 4009 1493 4018 1501
rect 4018 1493 4052 1501
rect 4052 1493 4061 1501
rect 4009 1449 4061 1493
rect 4209 1667 4261 1711
rect 4209 1659 4218 1667
rect 4218 1659 4252 1667
rect 4252 1659 4261 1667
rect 4409 1773 4418 1781
rect 4418 1773 4452 1781
rect 4452 1773 4461 1781
rect 4409 1729 4461 1773
rect 4609 1947 4661 1991
rect 4609 1939 4618 1947
rect 4618 1939 4652 1947
rect 4652 1939 4661 1947
rect 4809 2053 4818 2061
rect 4818 2053 4852 2061
rect 4852 2053 4861 2061
rect 4809 2009 4861 2053
rect 5009 2227 5061 2271
rect 5009 2219 5018 2227
rect 5018 2219 5052 2227
rect 5052 2219 5061 2227
rect 5209 2333 5218 2341
rect 5218 2333 5252 2341
rect 5252 2333 5261 2341
rect 5209 2289 5261 2333
rect 5409 2597 5461 2641
rect 5409 2589 5418 2597
rect 5418 2589 5452 2597
rect 5452 2589 5461 2597
rect 5609 2703 5618 2711
rect 5618 2703 5652 2711
rect 5652 2703 5661 2711
rect 5609 2659 5661 2703
rect 5809 2877 5861 2921
rect 5809 2869 5818 2877
rect 5818 2869 5852 2877
rect 5852 2869 5861 2877
rect 6009 2983 6018 2991
rect 6018 2983 6052 2991
rect 6052 2983 6061 2991
rect 6009 2939 6061 2983
rect 6209 3157 6261 3201
rect 6209 3149 6218 3157
rect 6218 3149 6252 3157
rect 6252 3149 6261 3157
rect 6409 3263 6418 3271
rect 6418 3263 6452 3271
rect 6452 3263 6461 3271
rect 6409 3219 6461 3263
rect 6609 3437 6661 3481
rect 6609 3429 6618 3437
rect 6618 3429 6652 3437
rect 6652 3429 6661 3437
rect 6809 3543 6818 3551
rect 6818 3543 6852 3551
rect 6852 3543 6861 3551
rect 6809 3499 6861 3543
rect 7009 3807 7061 3851
rect 7009 3799 7018 3807
rect 7018 3799 7052 3807
rect 7052 3799 7061 3807
rect 7209 3913 7218 3921
rect 7218 3913 7252 3921
rect 7252 3913 7261 3921
rect 7209 3869 7261 3913
rect 7409 4087 7461 4131
rect 7409 4079 7418 4087
rect 7418 4079 7452 4087
rect 7452 4079 7461 4087
rect 7609 4193 7618 4201
rect 7618 4193 7652 4201
rect 7652 4193 7661 4201
rect 7609 4149 7661 4193
rect 7809 4367 7861 4411
rect 7809 4359 7818 4367
rect 7818 4359 7852 4367
rect 7852 4359 7861 4367
rect 8009 4473 8018 4481
rect 8018 4473 8052 4481
rect 8052 4473 8061 4481
rect 8009 4429 8061 4473
rect 8209 4647 8261 4691
rect 8209 4639 8218 4647
rect 8218 4639 8252 4647
rect 8252 4639 8261 4647
rect 8409 4753 8418 4761
rect 8418 4753 8452 4761
rect 8452 4753 8461 4761
rect 8409 4709 8461 4753
rect 8609 4910 8661 4919
rect 8609 4876 8618 4910
rect 8618 4876 8652 4910
rect 8652 4876 8661 4910
rect 8609 4867 8661 4876
rect 7009 3700 7061 3709
rect 7009 3666 7018 3700
rect 7018 3666 7052 3700
rect 7052 3666 7061 3700
rect 7009 3657 7061 3666
rect 5409 2490 5461 2499
rect 5409 2456 5418 2490
rect 5418 2456 5452 2490
rect 5452 2456 5461 2490
rect 5409 2447 5461 2456
rect 3809 1280 3861 1289
rect 3809 1246 3818 1280
rect 3818 1246 3852 1280
rect 3852 1246 3861 1280
rect 3809 1237 3861 1246
rect 2209 70 2261 79
rect 2209 36 2218 70
rect 2218 36 2252 70
rect 2252 36 2261 70
rect 2209 27 2261 36
rect 2109 -60 2161 -15
rect 2109 -67 2118 -60
rect 2118 -67 2152 -60
rect 2152 -67 2161 -60
rect 1909 -166 1918 -143
rect 1918 -166 1952 -143
rect 1952 -166 1961 -143
rect 1909 -195 1961 -166
rect 1925 -248 1977 -239
rect 1925 -282 1934 -248
rect 1934 -282 1968 -248
rect 1968 -282 1977 -248
rect 1925 -291 1977 -282
rect 1909 -363 1961 -326
rect 1909 -378 1918 -363
rect 1918 -378 1952 -363
rect 1952 -378 1961 -363
rect 1909 -397 1918 -390
rect 1918 -397 1952 -390
rect 1952 -397 1961 -390
rect 1909 -435 1961 -397
rect 1909 -442 1918 -435
rect 1918 -442 1952 -435
rect 1952 -442 1961 -435
rect 1909 -469 1918 -454
rect 1918 -469 1952 -454
rect 1952 -469 1961 -454
rect 1909 -506 1961 -469
rect 2109 -94 2118 -79
rect 2118 -94 2152 -79
rect 2152 -94 2161 -79
rect 2109 -131 2161 -94
rect 2209 -74 2261 -22
rect 2409 143 2418 151
rect 2418 143 2452 151
rect 2452 143 2461 151
rect 2409 99 2461 143
rect 2609 317 2661 361
rect 2609 309 2618 317
rect 2618 309 2652 317
rect 2652 309 2661 317
rect 2809 423 2818 431
rect 2818 423 2852 431
rect 2852 423 2861 431
rect 2809 379 2861 423
rect 3009 597 3061 641
rect 3009 589 3018 597
rect 3018 589 3052 597
rect 3052 589 3061 597
rect 3209 703 3218 711
rect 3218 703 3252 711
rect 3252 703 3261 711
rect 3209 659 3261 703
rect 3409 877 3461 921
rect 3409 869 3418 877
rect 3418 869 3452 877
rect 3452 869 3461 877
rect 3609 983 3618 991
rect 3618 983 3652 991
rect 3652 983 3661 991
rect 3609 939 3661 983
rect 3809 1157 3861 1201
rect 3809 1149 3818 1157
rect 3818 1149 3852 1157
rect 3852 1149 3861 1157
rect 4009 1353 4018 1361
rect 4018 1353 4052 1361
rect 4052 1353 4061 1361
rect 4009 1309 4061 1353
rect 4209 1527 4261 1571
rect 4209 1519 4218 1527
rect 4218 1519 4252 1527
rect 4252 1519 4261 1527
rect 4409 1633 4418 1641
rect 4418 1633 4452 1641
rect 4452 1633 4461 1641
rect 4409 1589 4461 1633
rect 4609 1807 4661 1851
rect 4609 1799 4618 1807
rect 4618 1799 4652 1807
rect 4652 1799 4661 1807
rect 4809 1913 4818 1921
rect 4818 1913 4852 1921
rect 4852 1913 4861 1921
rect 4809 1869 4861 1913
rect 5009 2087 5061 2131
rect 5009 2079 5018 2087
rect 5018 2079 5052 2087
rect 5052 2079 5061 2087
rect 5209 2193 5218 2201
rect 5218 2193 5252 2201
rect 5252 2193 5261 2201
rect 5209 2149 5261 2193
rect 5409 2367 5461 2411
rect 5409 2359 5418 2367
rect 5418 2359 5452 2367
rect 5452 2359 5461 2367
rect 5609 2563 5618 2571
rect 5618 2563 5652 2571
rect 5652 2563 5661 2571
rect 5609 2519 5661 2563
rect 5809 2737 5861 2781
rect 5809 2729 5818 2737
rect 5818 2729 5852 2737
rect 5852 2729 5861 2737
rect 6009 2843 6018 2851
rect 6018 2843 6052 2851
rect 6052 2843 6061 2851
rect 6009 2799 6061 2843
rect 6209 3017 6261 3061
rect 6209 3009 6218 3017
rect 6218 3009 6252 3017
rect 6252 3009 6261 3017
rect 6409 3123 6418 3131
rect 6418 3123 6452 3131
rect 6452 3123 6461 3131
rect 6409 3079 6461 3123
rect 6609 3297 6661 3341
rect 6609 3289 6618 3297
rect 6618 3289 6652 3297
rect 6652 3289 6661 3297
rect 6809 3403 6818 3411
rect 6818 3403 6852 3411
rect 6852 3403 6861 3411
rect 6809 3359 6861 3403
rect 7009 3577 7061 3621
rect 7009 3569 7018 3577
rect 7018 3569 7052 3577
rect 7052 3569 7061 3577
rect 7209 3773 7218 3781
rect 7218 3773 7252 3781
rect 7252 3773 7261 3781
rect 7209 3729 7261 3773
rect 7409 3947 7461 3991
rect 7409 3939 7418 3947
rect 7418 3939 7452 3947
rect 7452 3939 7461 3947
rect 7609 4053 7618 4061
rect 7618 4053 7652 4061
rect 7652 4053 7661 4061
rect 7609 4009 7661 4053
rect 7809 4227 7861 4271
rect 7809 4219 7818 4227
rect 7818 4219 7852 4227
rect 7852 4219 7861 4227
rect 8009 4333 8018 4341
rect 8018 4333 8052 4341
rect 8052 4333 8061 4341
rect 8009 4289 8061 4333
rect 8209 4507 8261 4551
rect 8209 4499 8218 4507
rect 8218 4499 8252 4507
rect 8252 4499 8261 4507
rect 8409 4613 8418 4621
rect 8418 4613 8452 4621
rect 8452 4613 8461 4621
rect 8409 4569 8461 4613
rect 8609 4787 8661 4831
rect 8609 4779 8618 4787
rect 8618 4779 8652 4787
rect 8652 4779 8661 4787
rect 8809 4894 8861 4903
rect 8809 4860 8818 4894
rect 8818 4860 8852 4894
rect 8852 4860 8861 4894
rect 8809 4851 8861 4860
rect 7209 3684 7261 3693
rect 7209 3650 7218 3684
rect 7218 3650 7252 3684
rect 7252 3650 7261 3684
rect 7209 3641 7261 3650
rect 5609 2474 5661 2483
rect 5609 2440 5618 2474
rect 5618 2440 5652 2474
rect 5652 2440 5661 2474
rect 5609 2431 5661 2440
rect 4009 1264 4061 1273
rect 4009 1230 4018 1264
rect 4018 1230 4052 1264
rect 4052 1230 4061 1264
rect 4009 1221 4061 1230
rect 2409 54 2461 63
rect 2409 20 2418 54
rect 2418 20 2452 54
rect 2452 20 2461 54
rect 2409 11 2461 20
rect 2309 -60 2361 -15
rect 2309 -67 2318 -60
rect 2318 -67 2352 -60
rect 2352 -67 2361 -60
rect 2109 -166 2118 -143
rect 2118 -166 2152 -143
rect 2152 -166 2161 -143
rect 2109 -195 2161 -166
rect 2125 -248 2177 -239
rect 2125 -282 2134 -248
rect 2134 -282 2168 -248
rect 2168 -282 2177 -248
rect 2125 -291 2177 -282
rect 2109 -363 2161 -326
rect 2109 -378 2118 -363
rect 2118 -378 2152 -363
rect 2152 -378 2161 -363
rect 2109 -397 2118 -390
rect 2118 -397 2152 -390
rect 2152 -397 2161 -390
rect 2109 -435 2161 -397
rect 2109 -442 2118 -435
rect 2118 -442 2152 -435
rect 2152 -442 2161 -435
rect 2109 -469 2118 -454
rect 2118 -469 2152 -454
rect 2152 -469 2161 -454
rect 2109 -506 2161 -469
rect 2309 -94 2318 -79
rect 2318 -94 2352 -79
rect 2352 -94 2361 -79
rect 2309 -131 2361 -94
rect 2409 -74 2461 -22
rect 2609 177 2661 221
rect 2609 169 2618 177
rect 2618 169 2652 177
rect 2652 169 2661 177
rect 2809 283 2818 291
rect 2818 283 2852 291
rect 2852 283 2861 291
rect 2809 239 2861 283
rect 3009 457 3061 501
rect 3009 449 3018 457
rect 3018 449 3052 457
rect 3052 449 3061 457
rect 3209 563 3218 571
rect 3218 563 3252 571
rect 3252 563 3261 571
rect 3209 519 3261 563
rect 3409 737 3461 781
rect 3409 729 3418 737
rect 3418 729 3452 737
rect 3452 729 3461 737
rect 3609 843 3618 851
rect 3618 843 3652 851
rect 3652 843 3661 851
rect 3609 799 3661 843
rect 3809 1017 3861 1061
rect 3809 1009 3818 1017
rect 3818 1009 3852 1017
rect 3852 1009 3861 1017
rect 4009 1123 4018 1131
rect 4018 1123 4052 1131
rect 4052 1123 4061 1131
rect 4009 1079 4061 1123
rect 4209 1387 4261 1431
rect 4209 1379 4218 1387
rect 4218 1379 4252 1387
rect 4252 1379 4261 1387
rect 4409 1493 4418 1501
rect 4418 1493 4452 1501
rect 4452 1493 4461 1501
rect 4409 1449 4461 1493
rect 4609 1667 4661 1711
rect 4609 1659 4618 1667
rect 4618 1659 4652 1667
rect 4652 1659 4661 1667
rect 4809 1773 4818 1781
rect 4818 1773 4852 1781
rect 4852 1773 4861 1781
rect 4809 1729 4861 1773
rect 5009 1947 5061 1991
rect 5009 1939 5018 1947
rect 5018 1939 5052 1947
rect 5052 1939 5061 1947
rect 5209 2053 5218 2061
rect 5218 2053 5252 2061
rect 5252 2053 5261 2061
rect 5209 2009 5261 2053
rect 5409 2227 5461 2271
rect 5409 2219 5418 2227
rect 5418 2219 5452 2227
rect 5452 2219 5461 2227
rect 5609 2333 5618 2341
rect 5618 2333 5652 2341
rect 5652 2333 5661 2341
rect 5609 2289 5661 2333
rect 5809 2597 5861 2641
rect 5809 2589 5818 2597
rect 5818 2589 5852 2597
rect 5852 2589 5861 2597
rect 6009 2703 6018 2711
rect 6018 2703 6052 2711
rect 6052 2703 6061 2711
rect 6009 2659 6061 2703
rect 6209 2877 6261 2921
rect 6209 2869 6218 2877
rect 6218 2869 6252 2877
rect 6252 2869 6261 2877
rect 6409 2983 6418 2991
rect 6418 2983 6452 2991
rect 6452 2983 6461 2991
rect 6409 2939 6461 2983
rect 6609 3157 6661 3201
rect 6609 3149 6618 3157
rect 6618 3149 6652 3157
rect 6652 3149 6661 3157
rect 6809 3263 6818 3271
rect 6818 3263 6852 3271
rect 6852 3263 6861 3271
rect 6809 3219 6861 3263
rect 7009 3437 7061 3481
rect 7009 3429 7018 3437
rect 7018 3429 7052 3437
rect 7052 3429 7061 3437
rect 7209 3543 7218 3551
rect 7218 3543 7252 3551
rect 7252 3543 7261 3551
rect 7209 3499 7261 3543
rect 7409 3807 7461 3851
rect 7409 3799 7418 3807
rect 7418 3799 7452 3807
rect 7452 3799 7461 3807
rect 7609 3913 7618 3921
rect 7618 3913 7652 3921
rect 7652 3913 7661 3921
rect 7609 3869 7661 3913
rect 7809 4087 7861 4131
rect 7809 4079 7818 4087
rect 7818 4079 7852 4087
rect 7852 4079 7861 4087
rect 8009 4193 8018 4201
rect 8018 4193 8052 4201
rect 8052 4193 8061 4201
rect 8009 4149 8061 4193
rect 8209 4367 8261 4411
rect 8209 4359 8218 4367
rect 8218 4359 8252 4367
rect 8252 4359 8261 4367
rect 8409 4473 8418 4481
rect 8418 4473 8452 4481
rect 8452 4473 8461 4481
rect 8409 4429 8461 4473
rect 8609 4647 8661 4691
rect 8609 4639 8618 4647
rect 8618 4639 8652 4647
rect 8652 4639 8661 4647
rect 8809 4753 8818 4761
rect 8818 4753 8852 4761
rect 8852 4753 8861 4761
rect 8809 4709 8861 4753
rect 9009 4910 9061 4919
rect 9009 4876 9018 4910
rect 9018 4876 9052 4910
rect 9052 4876 9061 4910
rect 9009 4867 9061 4876
rect 7409 3700 7461 3709
rect 7409 3666 7418 3700
rect 7418 3666 7452 3700
rect 7452 3666 7461 3700
rect 7409 3657 7461 3666
rect 5809 2490 5861 2499
rect 5809 2456 5818 2490
rect 5818 2456 5852 2490
rect 5852 2456 5861 2490
rect 5809 2447 5861 2456
rect 4209 1280 4261 1289
rect 4209 1246 4218 1280
rect 4218 1246 4252 1280
rect 4252 1246 4261 1280
rect 4209 1237 4261 1246
rect 2609 70 2661 79
rect 2609 36 2618 70
rect 2618 36 2652 70
rect 2652 36 2661 70
rect 2609 27 2661 36
rect 2509 -60 2561 -15
rect 2509 -67 2518 -60
rect 2518 -67 2552 -60
rect 2552 -67 2561 -60
rect 2309 -166 2318 -143
rect 2318 -166 2352 -143
rect 2352 -166 2361 -143
rect 2309 -195 2361 -166
rect 2325 -248 2377 -239
rect 2325 -282 2334 -248
rect 2334 -282 2368 -248
rect 2368 -282 2377 -248
rect 2325 -291 2377 -282
rect 2309 -363 2361 -326
rect 2309 -378 2318 -363
rect 2318 -378 2352 -363
rect 2352 -378 2361 -363
rect 2309 -397 2318 -390
rect 2318 -397 2352 -390
rect 2352 -397 2361 -390
rect 2309 -435 2361 -397
rect 2309 -442 2318 -435
rect 2318 -442 2352 -435
rect 2352 -442 2361 -435
rect 2309 -469 2318 -454
rect 2318 -469 2352 -454
rect 2352 -469 2361 -454
rect 2309 -506 2361 -469
rect 2509 -94 2518 -79
rect 2518 -94 2552 -79
rect 2552 -94 2561 -79
rect 2509 -131 2561 -94
rect 2609 -74 2661 -22
rect 2809 143 2818 151
rect 2818 143 2852 151
rect 2852 143 2861 151
rect 2809 99 2861 143
rect 3009 317 3061 361
rect 3009 309 3018 317
rect 3018 309 3052 317
rect 3052 309 3061 317
rect 3209 423 3218 431
rect 3218 423 3252 431
rect 3252 423 3261 431
rect 3209 379 3261 423
rect 3409 597 3461 641
rect 3409 589 3418 597
rect 3418 589 3452 597
rect 3452 589 3461 597
rect 3609 703 3618 711
rect 3618 703 3652 711
rect 3652 703 3661 711
rect 3609 659 3661 703
rect 3809 877 3861 921
rect 3809 869 3818 877
rect 3818 869 3852 877
rect 3852 869 3861 877
rect 4009 983 4018 991
rect 4018 983 4052 991
rect 4052 983 4061 991
rect 4009 939 4061 983
rect 4209 1157 4261 1201
rect 4209 1149 4218 1157
rect 4218 1149 4252 1157
rect 4252 1149 4261 1157
rect 4409 1353 4418 1361
rect 4418 1353 4452 1361
rect 4452 1353 4461 1361
rect 4409 1309 4461 1353
rect 4609 1527 4661 1571
rect 4609 1519 4618 1527
rect 4618 1519 4652 1527
rect 4652 1519 4661 1527
rect 4809 1633 4818 1641
rect 4818 1633 4852 1641
rect 4852 1633 4861 1641
rect 4809 1589 4861 1633
rect 5009 1807 5061 1851
rect 5009 1799 5018 1807
rect 5018 1799 5052 1807
rect 5052 1799 5061 1807
rect 5209 1913 5218 1921
rect 5218 1913 5252 1921
rect 5252 1913 5261 1921
rect 5209 1869 5261 1913
rect 5409 2087 5461 2131
rect 5409 2079 5418 2087
rect 5418 2079 5452 2087
rect 5452 2079 5461 2087
rect 5609 2193 5618 2201
rect 5618 2193 5652 2201
rect 5652 2193 5661 2201
rect 5609 2149 5661 2193
rect 5809 2367 5861 2411
rect 5809 2359 5818 2367
rect 5818 2359 5852 2367
rect 5852 2359 5861 2367
rect 6009 2563 6018 2571
rect 6018 2563 6052 2571
rect 6052 2563 6061 2571
rect 6009 2519 6061 2563
rect 6209 2737 6261 2781
rect 6209 2729 6218 2737
rect 6218 2729 6252 2737
rect 6252 2729 6261 2737
rect 6409 2843 6418 2851
rect 6418 2843 6452 2851
rect 6452 2843 6461 2851
rect 6409 2799 6461 2843
rect 6609 3017 6661 3061
rect 6609 3009 6618 3017
rect 6618 3009 6652 3017
rect 6652 3009 6661 3017
rect 6809 3123 6818 3131
rect 6818 3123 6852 3131
rect 6852 3123 6861 3131
rect 6809 3079 6861 3123
rect 7009 3297 7061 3341
rect 7009 3289 7018 3297
rect 7018 3289 7052 3297
rect 7052 3289 7061 3297
rect 7209 3403 7218 3411
rect 7218 3403 7252 3411
rect 7252 3403 7261 3411
rect 7209 3359 7261 3403
rect 7409 3577 7461 3621
rect 7409 3569 7418 3577
rect 7418 3569 7452 3577
rect 7452 3569 7461 3577
rect 7609 3773 7618 3781
rect 7618 3773 7652 3781
rect 7652 3773 7661 3781
rect 7609 3729 7661 3773
rect 7809 3947 7861 3991
rect 7809 3939 7818 3947
rect 7818 3939 7852 3947
rect 7852 3939 7861 3947
rect 8009 4053 8018 4061
rect 8018 4053 8052 4061
rect 8052 4053 8061 4061
rect 8009 4009 8061 4053
rect 8209 4227 8261 4271
rect 8209 4219 8218 4227
rect 8218 4219 8252 4227
rect 8252 4219 8261 4227
rect 8409 4333 8418 4341
rect 8418 4333 8452 4341
rect 8452 4333 8461 4341
rect 8409 4289 8461 4333
rect 8609 4507 8661 4551
rect 8609 4499 8618 4507
rect 8618 4499 8652 4507
rect 8652 4499 8661 4507
rect 8809 4613 8818 4621
rect 8818 4613 8852 4621
rect 8852 4613 8861 4621
rect 8809 4569 8861 4613
rect 9009 4787 9061 4831
rect 9009 4779 9018 4787
rect 9018 4779 9052 4787
rect 9052 4779 9061 4787
rect 9209 4894 9261 4903
rect 9209 4860 9218 4894
rect 9218 4860 9252 4894
rect 9252 4860 9261 4894
rect 9209 4851 9261 4860
rect 7609 3684 7661 3693
rect 7609 3650 7618 3684
rect 7618 3650 7652 3684
rect 7652 3650 7661 3684
rect 7609 3641 7661 3650
rect 6009 2474 6061 2483
rect 6009 2440 6018 2474
rect 6018 2440 6052 2474
rect 6052 2440 6061 2474
rect 6009 2431 6061 2440
rect 4409 1264 4461 1273
rect 4409 1230 4418 1264
rect 4418 1230 4452 1264
rect 4452 1230 4461 1264
rect 4409 1221 4461 1230
rect 2809 54 2861 63
rect 2809 20 2818 54
rect 2818 20 2852 54
rect 2852 20 2861 54
rect 2809 11 2861 20
rect 2709 -60 2761 -15
rect 2709 -67 2718 -60
rect 2718 -67 2752 -60
rect 2752 -67 2761 -60
rect 2509 -166 2518 -143
rect 2518 -166 2552 -143
rect 2552 -166 2561 -143
rect 2509 -195 2561 -166
rect 2525 -248 2577 -239
rect 2525 -282 2534 -248
rect 2534 -282 2568 -248
rect 2568 -282 2577 -248
rect 2525 -291 2577 -282
rect 2509 -363 2561 -326
rect 2509 -378 2518 -363
rect 2518 -378 2552 -363
rect 2552 -378 2561 -363
rect 2509 -397 2518 -390
rect 2518 -397 2552 -390
rect 2552 -397 2561 -390
rect 2509 -435 2561 -397
rect 2509 -442 2518 -435
rect 2518 -442 2552 -435
rect 2552 -442 2561 -435
rect 2509 -469 2518 -454
rect 2518 -469 2552 -454
rect 2552 -469 2561 -454
rect 2509 -506 2561 -469
rect 2709 -94 2718 -79
rect 2718 -94 2752 -79
rect 2752 -94 2761 -79
rect 2709 -131 2761 -94
rect 2809 -74 2861 -22
rect 3009 177 3061 221
rect 3009 169 3018 177
rect 3018 169 3052 177
rect 3052 169 3061 177
rect 3209 283 3218 291
rect 3218 283 3252 291
rect 3252 283 3261 291
rect 3209 239 3261 283
rect 3409 457 3461 501
rect 3409 449 3418 457
rect 3418 449 3452 457
rect 3452 449 3461 457
rect 3609 563 3618 571
rect 3618 563 3652 571
rect 3652 563 3661 571
rect 3609 519 3661 563
rect 3809 737 3861 781
rect 3809 729 3818 737
rect 3818 729 3852 737
rect 3852 729 3861 737
rect 4009 843 4018 851
rect 4018 843 4052 851
rect 4052 843 4061 851
rect 4009 799 4061 843
rect 4209 1017 4261 1061
rect 4209 1009 4218 1017
rect 4218 1009 4252 1017
rect 4252 1009 4261 1017
rect 4409 1123 4418 1131
rect 4418 1123 4452 1131
rect 4452 1123 4461 1131
rect 4409 1079 4461 1123
rect 4609 1387 4661 1431
rect 4609 1379 4618 1387
rect 4618 1379 4652 1387
rect 4652 1379 4661 1387
rect 4809 1493 4818 1501
rect 4818 1493 4852 1501
rect 4852 1493 4861 1501
rect 4809 1449 4861 1493
rect 5009 1667 5061 1711
rect 5009 1659 5018 1667
rect 5018 1659 5052 1667
rect 5052 1659 5061 1667
rect 5209 1773 5218 1781
rect 5218 1773 5252 1781
rect 5252 1773 5261 1781
rect 5209 1729 5261 1773
rect 5409 1947 5461 1991
rect 5409 1939 5418 1947
rect 5418 1939 5452 1947
rect 5452 1939 5461 1947
rect 5609 2053 5618 2061
rect 5618 2053 5652 2061
rect 5652 2053 5661 2061
rect 5609 2009 5661 2053
rect 5809 2227 5861 2271
rect 5809 2219 5818 2227
rect 5818 2219 5852 2227
rect 5852 2219 5861 2227
rect 6009 2333 6018 2341
rect 6018 2333 6052 2341
rect 6052 2333 6061 2341
rect 6009 2289 6061 2333
rect 6209 2597 6261 2641
rect 6209 2589 6218 2597
rect 6218 2589 6252 2597
rect 6252 2589 6261 2597
rect 6409 2703 6418 2711
rect 6418 2703 6452 2711
rect 6452 2703 6461 2711
rect 6409 2659 6461 2703
rect 6609 2877 6661 2921
rect 6609 2869 6618 2877
rect 6618 2869 6652 2877
rect 6652 2869 6661 2877
rect 6809 2983 6818 2991
rect 6818 2983 6852 2991
rect 6852 2983 6861 2991
rect 6809 2939 6861 2983
rect 7009 3157 7061 3201
rect 7009 3149 7018 3157
rect 7018 3149 7052 3157
rect 7052 3149 7061 3157
rect 7209 3263 7218 3271
rect 7218 3263 7252 3271
rect 7252 3263 7261 3271
rect 7209 3219 7261 3263
rect 7409 3437 7461 3481
rect 7409 3429 7418 3437
rect 7418 3429 7452 3437
rect 7452 3429 7461 3437
rect 7609 3543 7618 3551
rect 7618 3543 7652 3551
rect 7652 3543 7661 3551
rect 7609 3499 7661 3543
rect 7809 3807 7861 3851
rect 7809 3799 7818 3807
rect 7818 3799 7852 3807
rect 7852 3799 7861 3807
rect 8009 3913 8018 3921
rect 8018 3913 8052 3921
rect 8052 3913 8061 3921
rect 8009 3869 8061 3913
rect 8209 4087 8261 4131
rect 8209 4079 8218 4087
rect 8218 4079 8252 4087
rect 8252 4079 8261 4087
rect 8409 4193 8418 4201
rect 8418 4193 8452 4201
rect 8452 4193 8461 4201
rect 8409 4149 8461 4193
rect 8609 4367 8661 4411
rect 8609 4359 8618 4367
rect 8618 4359 8652 4367
rect 8652 4359 8661 4367
rect 8809 4473 8818 4481
rect 8818 4473 8852 4481
rect 8852 4473 8861 4481
rect 8809 4429 8861 4473
rect 9009 4647 9061 4691
rect 9009 4639 9018 4647
rect 9018 4639 9052 4647
rect 9052 4639 9061 4647
rect 9209 4753 9218 4761
rect 9218 4753 9252 4761
rect 9252 4753 9261 4761
rect 9209 4709 9261 4753
rect 9409 4910 9461 4919
rect 9409 4876 9418 4910
rect 9418 4876 9452 4910
rect 9452 4876 9461 4910
rect 9409 4867 9461 4876
rect 7809 3700 7861 3709
rect 7809 3666 7818 3700
rect 7818 3666 7852 3700
rect 7852 3666 7861 3700
rect 7809 3657 7861 3666
rect 6209 2490 6261 2499
rect 6209 2456 6218 2490
rect 6218 2456 6252 2490
rect 6252 2456 6261 2490
rect 6209 2447 6261 2456
rect 4609 1280 4661 1289
rect 4609 1246 4618 1280
rect 4618 1246 4652 1280
rect 4652 1246 4661 1280
rect 4609 1237 4661 1246
rect 3009 70 3061 79
rect 3009 36 3018 70
rect 3018 36 3052 70
rect 3052 36 3061 70
rect 3009 27 3061 36
rect 2909 -60 2961 -15
rect 2909 -67 2918 -60
rect 2918 -67 2952 -60
rect 2952 -67 2961 -60
rect 2709 -166 2718 -143
rect 2718 -166 2752 -143
rect 2752 -166 2761 -143
rect 2709 -195 2761 -166
rect 2725 -248 2777 -239
rect 2725 -282 2734 -248
rect 2734 -282 2768 -248
rect 2768 -282 2777 -248
rect 2725 -291 2777 -282
rect 2709 -363 2761 -326
rect 2709 -378 2718 -363
rect 2718 -378 2752 -363
rect 2752 -378 2761 -363
rect 2709 -397 2718 -390
rect 2718 -397 2752 -390
rect 2752 -397 2761 -390
rect 2709 -435 2761 -397
rect 2709 -442 2718 -435
rect 2718 -442 2752 -435
rect 2752 -442 2761 -435
rect 2709 -469 2718 -454
rect 2718 -469 2752 -454
rect 2752 -469 2761 -454
rect 2709 -506 2761 -469
rect 2909 -94 2918 -79
rect 2918 -94 2952 -79
rect 2952 -94 2961 -79
rect 2909 -131 2961 -94
rect 3009 -74 3061 -22
rect 3209 143 3218 151
rect 3218 143 3252 151
rect 3252 143 3261 151
rect 3209 99 3261 143
rect 3409 317 3461 361
rect 3409 309 3418 317
rect 3418 309 3452 317
rect 3452 309 3461 317
rect 3609 423 3618 431
rect 3618 423 3652 431
rect 3652 423 3661 431
rect 3609 379 3661 423
rect 3809 597 3861 641
rect 3809 589 3818 597
rect 3818 589 3852 597
rect 3852 589 3861 597
rect 4009 703 4018 711
rect 4018 703 4052 711
rect 4052 703 4061 711
rect 4009 659 4061 703
rect 4209 877 4261 921
rect 4209 869 4218 877
rect 4218 869 4252 877
rect 4252 869 4261 877
rect 4409 983 4418 991
rect 4418 983 4452 991
rect 4452 983 4461 991
rect 4409 939 4461 983
rect 4609 1157 4661 1201
rect 4609 1149 4618 1157
rect 4618 1149 4652 1157
rect 4652 1149 4661 1157
rect 4809 1353 4818 1361
rect 4818 1353 4852 1361
rect 4852 1353 4861 1361
rect 4809 1309 4861 1353
rect 5009 1527 5061 1571
rect 5009 1519 5018 1527
rect 5018 1519 5052 1527
rect 5052 1519 5061 1527
rect 5209 1633 5218 1641
rect 5218 1633 5252 1641
rect 5252 1633 5261 1641
rect 5209 1589 5261 1633
rect 5409 1807 5461 1851
rect 5409 1799 5418 1807
rect 5418 1799 5452 1807
rect 5452 1799 5461 1807
rect 5609 1913 5618 1921
rect 5618 1913 5652 1921
rect 5652 1913 5661 1921
rect 5609 1869 5661 1913
rect 5809 2087 5861 2131
rect 5809 2079 5818 2087
rect 5818 2079 5852 2087
rect 5852 2079 5861 2087
rect 6009 2193 6018 2201
rect 6018 2193 6052 2201
rect 6052 2193 6061 2201
rect 6009 2149 6061 2193
rect 6209 2367 6261 2411
rect 6209 2359 6218 2367
rect 6218 2359 6252 2367
rect 6252 2359 6261 2367
rect 6409 2563 6418 2571
rect 6418 2563 6452 2571
rect 6452 2563 6461 2571
rect 6409 2519 6461 2563
rect 6609 2737 6661 2781
rect 6609 2729 6618 2737
rect 6618 2729 6652 2737
rect 6652 2729 6661 2737
rect 6809 2843 6818 2851
rect 6818 2843 6852 2851
rect 6852 2843 6861 2851
rect 6809 2799 6861 2843
rect 7009 3017 7061 3061
rect 7009 3009 7018 3017
rect 7018 3009 7052 3017
rect 7052 3009 7061 3017
rect 7209 3123 7218 3131
rect 7218 3123 7252 3131
rect 7252 3123 7261 3131
rect 7209 3079 7261 3123
rect 7409 3297 7461 3341
rect 7409 3289 7418 3297
rect 7418 3289 7452 3297
rect 7452 3289 7461 3297
rect 7609 3403 7618 3411
rect 7618 3403 7652 3411
rect 7652 3403 7661 3411
rect 7609 3359 7661 3403
rect 7809 3577 7861 3621
rect 7809 3569 7818 3577
rect 7818 3569 7852 3577
rect 7852 3569 7861 3577
rect 8009 3773 8018 3781
rect 8018 3773 8052 3781
rect 8052 3773 8061 3781
rect 8009 3729 8061 3773
rect 8209 3947 8261 3991
rect 8209 3939 8218 3947
rect 8218 3939 8252 3947
rect 8252 3939 8261 3947
rect 8409 4053 8418 4061
rect 8418 4053 8452 4061
rect 8452 4053 8461 4061
rect 8409 4009 8461 4053
rect 8609 4227 8661 4271
rect 8609 4219 8618 4227
rect 8618 4219 8652 4227
rect 8652 4219 8661 4227
rect 8809 4333 8818 4341
rect 8818 4333 8852 4341
rect 8852 4333 8861 4341
rect 8809 4289 8861 4333
rect 9009 4507 9061 4551
rect 9009 4499 9018 4507
rect 9018 4499 9052 4507
rect 9052 4499 9061 4507
rect 9209 4613 9218 4621
rect 9218 4613 9252 4621
rect 9252 4613 9261 4621
rect 9209 4569 9261 4613
rect 9409 4787 9461 4831
rect 9409 4779 9418 4787
rect 9418 4779 9452 4787
rect 9452 4779 9461 4787
rect 9609 4894 9661 4903
rect 9609 4860 9618 4894
rect 9618 4860 9652 4894
rect 9652 4860 9661 4894
rect 9609 4851 9661 4860
rect 8009 3684 8061 3693
rect 8009 3650 8018 3684
rect 8018 3650 8052 3684
rect 8052 3650 8061 3684
rect 8009 3641 8061 3650
rect 6409 2474 6461 2483
rect 6409 2440 6418 2474
rect 6418 2440 6452 2474
rect 6452 2440 6461 2474
rect 6409 2431 6461 2440
rect 4809 1264 4861 1273
rect 4809 1230 4818 1264
rect 4818 1230 4852 1264
rect 4852 1230 4861 1264
rect 4809 1221 4861 1230
rect 3209 54 3261 63
rect 3209 20 3218 54
rect 3218 20 3252 54
rect 3252 20 3261 54
rect 3209 11 3261 20
rect 3109 -60 3161 -15
rect 3109 -67 3118 -60
rect 3118 -67 3152 -60
rect 3152 -67 3161 -60
rect 2909 -166 2918 -143
rect 2918 -166 2952 -143
rect 2952 -166 2961 -143
rect 2909 -195 2961 -166
rect 2925 -248 2977 -239
rect 2925 -282 2934 -248
rect 2934 -282 2968 -248
rect 2968 -282 2977 -248
rect 2925 -291 2977 -282
rect 2909 -363 2961 -326
rect 2909 -378 2918 -363
rect 2918 -378 2952 -363
rect 2952 -378 2961 -363
rect 2909 -397 2918 -390
rect 2918 -397 2952 -390
rect 2952 -397 2961 -390
rect 2909 -435 2961 -397
rect 2909 -442 2918 -435
rect 2918 -442 2952 -435
rect 2952 -442 2961 -435
rect 2909 -469 2918 -454
rect 2918 -469 2952 -454
rect 2952 -469 2961 -454
rect 2909 -506 2961 -469
rect 3109 -94 3118 -79
rect 3118 -94 3152 -79
rect 3152 -94 3161 -79
rect 3109 -131 3161 -94
rect 3209 -74 3261 -22
rect 3409 177 3461 221
rect 3409 169 3418 177
rect 3418 169 3452 177
rect 3452 169 3461 177
rect 3609 283 3618 291
rect 3618 283 3652 291
rect 3652 283 3661 291
rect 3609 239 3661 283
rect 3809 457 3861 501
rect 3809 449 3818 457
rect 3818 449 3852 457
rect 3852 449 3861 457
rect 4009 563 4018 571
rect 4018 563 4052 571
rect 4052 563 4061 571
rect 4009 519 4061 563
rect 4209 737 4261 781
rect 4209 729 4218 737
rect 4218 729 4252 737
rect 4252 729 4261 737
rect 4409 843 4418 851
rect 4418 843 4452 851
rect 4452 843 4461 851
rect 4409 799 4461 843
rect 4609 1017 4661 1061
rect 4609 1009 4618 1017
rect 4618 1009 4652 1017
rect 4652 1009 4661 1017
rect 4809 1123 4818 1131
rect 4818 1123 4852 1131
rect 4852 1123 4861 1131
rect 4809 1079 4861 1123
rect 5009 1387 5061 1431
rect 5009 1379 5018 1387
rect 5018 1379 5052 1387
rect 5052 1379 5061 1387
rect 5209 1493 5218 1501
rect 5218 1493 5252 1501
rect 5252 1493 5261 1501
rect 5209 1449 5261 1493
rect 5409 1667 5461 1711
rect 5409 1659 5418 1667
rect 5418 1659 5452 1667
rect 5452 1659 5461 1667
rect 5609 1773 5618 1781
rect 5618 1773 5652 1781
rect 5652 1773 5661 1781
rect 5609 1729 5661 1773
rect 5809 1947 5861 1991
rect 5809 1939 5818 1947
rect 5818 1939 5852 1947
rect 5852 1939 5861 1947
rect 6009 2053 6018 2061
rect 6018 2053 6052 2061
rect 6052 2053 6061 2061
rect 6009 2009 6061 2053
rect 6209 2227 6261 2271
rect 6209 2219 6218 2227
rect 6218 2219 6252 2227
rect 6252 2219 6261 2227
rect 6409 2333 6418 2341
rect 6418 2333 6452 2341
rect 6452 2333 6461 2341
rect 6409 2289 6461 2333
rect 6609 2597 6661 2641
rect 6609 2589 6618 2597
rect 6618 2589 6652 2597
rect 6652 2589 6661 2597
rect 6809 2703 6818 2711
rect 6818 2703 6852 2711
rect 6852 2703 6861 2711
rect 6809 2659 6861 2703
rect 7009 2877 7061 2921
rect 7009 2869 7018 2877
rect 7018 2869 7052 2877
rect 7052 2869 7061 2877
rect 7209 2983 7218 2991
rect 7218 2983 7252 2991
rect 7252 2983 7261 2991
rect 7209 2939 7261 2983
rect 7409 3157 7461 3201
rect 7409 3149 7418 3157
rect 7418 3149 7452 3157
rect 7452 3149 7461 3157
rect 7609 3263 7618 3271
rect 7618 3263 7652 3271
rect 7652 3263 7661 3271
rect 7609 3219 7661 3263
rect 7809 3437 7861 3481
rect 7809 3429 7818 3437
rect 7818 3429 7852 3437
rect 7852 3429 7861 3437
rect 8009 3543 8018 3551
rect 8018 3543 8052 3551
rect 8052 3543 8061 3551
rect 8009 3499 8061 3543
rect 8209 3807 8261 3851
rect 8209 3799 8218 3807
rect 8218 3799 8252 3807
rect 8252 3799 8261 3807
rect 8409 3913 8418 3921
rect 8418 3913 8452 3921
rect 8452 3913 8461 3921
rect 8409 3869 8461 3913
rect 8609 4087 8661 4131
rect 8609 4079 8618 4087
rect 8618 4079 8652 4087
rect 8652 4079 8661 4087
rect 8809 4193 8818 4201
rect 8818 4193 8852 4201
rect 8852 4193 8861 4201
rect 8809 4149 8861 4193
rect 9009 4367 9061 4411
rect 9009 4359 9018 4367
rect 9018 4359 9052 4367
rect 9052 4359 9061 4367
rect 9209 4473 9218 4481
rect 9218 4473 9252 4481
rect 9252 4473 9261 4481
rect 9209 4429 9261 4473
rect 9409 4647 9461 4691
rect 9409 4639 9418 4647
rect 9418 4639 9452 4647
rect 9452 4639 9461 4647
rect 9609 4753 9618 4761
rect 9618 4753 9652 4761
rect 9652 4753 9661 4761
rect 9609 4709 9661 4753
rect 9809 4910 9861 4919
rect 9809 4876 9818 4910
rect 9818 4876 9852 4910
rect 9852 4876 9861 4910
rect 9809 4867 9861 4876
rect 8209 3700 8261 3709
rect 8209 3666 8218 3700
rect 8218 3666 8252 3700
rect 8252 3666 8261 3700
rect 8209 3657 8261 3666
rect 6609 2490 6661 2499
rect 6609 2456 6618 2490
rect 6618 2456 6652 2490
rect 6652 2456 6661 2490
rect 6609 2447 6661 2456
rect 5009 1280 5061 1289
rect 5009 1246 5018 1280
rect 5018 1246 5052 1280
rect 5052 1246 5061 1280
rect 5009 1237 5061 1246
rect 3409 70 3461 79
rect 3409 36 3418 70
rect 3418 36 3452 70
rect 3452 36 3461 70
rect 3409 27 3461 36
rect 3309 -60 3361 -15
rect 3309 -67 3318 -60
rect 3318 -67 3352 -60
rect 3352 -67 3361 -60
rect 3109 -166 3118 -143
rect 3118 -166 3152 -143
rect 3152 -166 3161 -143
rect 3109 -195 3161 -166
rect 3125 -248 3177 -239
rect 3125 -282 3134 -248
rect 3134 -282 3168 -248
rect 3168 -282 3177 -248
rect 3125 -291 3177 -282
rect 3109 -363 3161 -326
rect 3109 -378 3118 -363
rect 3118 -378 3152 -363
rect 3152 -378 3161 -363
rect 3109 -397 3118 -390
rect 3118 -397 3152 -390
rect 3152 -397 3161 -390
rect 3109 -435 3161 -397
rect 3109 -442 3118 -435
rect 3118 -442 3152 -435
rect 3152 -442 3161 -435
rect 3109 -469 3118 -454
rect 3118 -469 3152 -454
rect 3152 -469 3161 -454
rect 3109 -506 3161 -469
rect 3309 -94 3318 -79
rect 3318 -94 3352 -79
rect 3352 -94 3361 -79
rect 3309 -131 3361 -94
rect 3409 -74 3461 -22
rect 3609 143 3618 151
rect 3618 143 3652 151
rect 3652 143 3661 151
rect 3609 99 3661 143
rect 3809 317 3861 361
rect 3809 309 3818 317
rect 3818 309 3852 317
rect 3852 309 3861 317
rect 4009 423 4018 431
rect 4018 423 4052 431
rect 4052 423 4061 431
rect 4009 379 4061 423
rect 4209 597 4261 641
rect 4209 589 4218 597
rect 4218 589 4252 597
rect 4252 589 4261 597
rect 4409 703 4418 711
rect 4418 703 4452 711
rect 4452 703 4461 711
rect 4409 659 4461 703
rect 4609 877 4661 921
rect 4609 869 4618 877
rect 4618 869 4652 877
rect 4652 869 4661 877
rect 4809 983 4818 991
rect 4818 983 4852 991
rect 4852 983 4861 991
rect 4809 939 4861 983
rect 5009 1157 5061 1201
rect 5009 1149 5018 1157
rect 5018 1149 5052 1157
rect 5052 1149 5061 1157
rect 5209 1353 5218 1361
rect 5218 1353 5252 1361
rect 5252 1353 5261 1361
rect 5209 1309 5261 1353
rect 5409 1527 5461 1571
rect 5409 1519 5418 1527
rect 5418 1519 5452 1527
rect 5452 1519 5461 1527
rect 5609 1633 5618 1641
rect 5618 1633 5652 1641
rect 5652 1633 5661 1641
rect 5609 1589 5661 1633
rect 5809 1807 5861 1851
rect 5809 1799 5818 1807
rect 5818 1799 5852 1807
rect 5852 1799 5861 1807
rect 6009 1913 6018 1921
rect 6018 1913 6052 1921
rect 6052 1913 6061 1921
rect 6009 1869 6061 1913
rect 6209 2087 6261 2131
rect 6209 2079 6218 2087
rect 6218 2079 6252 2087
rect 6252 2079 6261 2087
rect 6409 2193 6418 2201
rect 6418 2193 6452 2201
rect 6452 2193 6461 2201
rect 6409 2149 6461 2193
rect 6609 2367 6661 2411
rect 6609 2359 6618 2367
rect 6618 2359 6652 2367
rect 6652 2359 6661 2367
rect 6809 2563 6818 2571
rect 6818 2563 6852 2571
rect 6852 2563 6861 2571
rect 6809 2519 6861 2563
rect 7009 2737 7061 2781
rect 7009 2729 7018 2737
rect 7018 2729 7052 2737
rect 7052 2729 7061 2737
rect 7209 2843 7218 2851
rect 7218 2843 7252 2851
rect 7252 2843 7261 2851
rect 7209 2799 7261 2843
rect 7409 3017 7461 3061
rect 7409 3009 7418 3017
rect 7418 3009 7452 3017
rect 7452 3009 7461 3017
rect 7609 3123 7618 3131
rect 7618 3123 7652 3131
rect 7652 3123 7661 3131
rect 7609 3079 7661 3123
rect 7809 3297 7861 3341
rect 7809 3289 7818 3297
rect 7818 3289 7852 3297
rect 7852 3289 7861 3297
rect 8009 3403 8018 3411
rect 8018 3403 8052 3411
rect 8052 3403 8061 3411
rect 8009 3359 8061 3403
rect 8209 3577 8261 3621
rect 8209 3569 8218 3577
rect 8218 3569 8252 3577
rect 8252 3569 8261 3577
rect 8409 3773 8418 3781
rect 8418 3773 8452 3781
rect 8452 3773 8461 3781
rect 8409 3729 8461 3773
rect 8609 3947 8661 3991
rect 8609 3939 8618 3947
rect 8618 3939 8652 3947
rect 8652 3939 8661 3947
rect 8809 4053 8818 4061
rect 8818 4053 8852 4061
rect 8852 4053 8861 4061
rect 8809 4009 8861 4053
rect 9009 4227 9061 4271
rect 9009 4219 9018 4227
rect 9018 4219 9052 4227
rect 9052 4219 9061 4227
rect 9209 4333 9218 4341
rect 9218 4333 9252 4341
rect 9252 4333 9261 4341
rect 9209 4289 9261 4333
rect 9409 4507 9461 4551
rect 9409 4499 9418 4507
rect 9418 4499 9452 4507
rect 9452 4499 9461 4507
rect 9609 4613 9618 4621
rect 9618 4613 9652 4621
rect 9652 4613 9661 4621
rect 9609 4569 9661 4613
rect 9809 4787 9861 4831
rect 9809 4779 9818 4787
rect 9818 4779 9852 4787
rect 9852 4779 9861 4787
rect 10009 4894 10061 4903
rect 10009 4860 10018 4894
rect 10018 4860 10052 4894
rect 10052 4860 10061 4894
rect 10009 4851 10061 4860
rect 8409 3684 8461 3693
rect 8409 3650 8418 3684
rect 8418 3650 8452 3684
rect 8452 3650 8461 3684
rect 8409 3641 8461 3650
rect 6809 2474 6861 2483
rect 6809 2440 6818 2474
rect 6818 2440 6852 2474
rect 6852 2440 6861 2474
rect 6809 2431 6861 2440
rect 5209 1264 5261 1273
rect 5209 1230 5218 1264
rect 5218 1230 5252 1264
rect 5252 1230 5261 1264
rect 5209 1221 5261 1230
rect 3609 54 3661 63
rect 3609 20 3618 54
rect 3618 20 3652 54
rect 3652 20 3661 54
rect 3609 11 3661 20
rect 3509 -60 3561 -15
rect 3509 -67 3518 -60
rect 3518 -67 3552 -60
rect 3552 -67 3561 -60
rect 3309 -166 3318 -143
rect 3318 -166 3352 -143
rect 3352 -166 3361 -143
rect 3309 -195 3361 -166
rect 3325 -248 3377 -239
rect 3325 -282 3334 -248
rect 3334 -282 3368 -248
rect 3368 -282 3377 -248
rect 3325 -291 3377 -282
rect 3309 -363 3361 -326
rect 3309 -378 3318 -363
rect 3318 -378 3352 -363
rect 3352 -378 3361 -363
rect 3309 -397 3318 -390
rect 3318 -397 3352 -390
rect 3352 -397 3361 -390
rect 3309 -435 3361 -397
rect 3309 -442 3318 -435
rect 3318 -442 3352 -435
rect 3352 -442 3361 -435
rect 3309 -469 3318 -454
rect 3318 -469 3352 -454
rect 3352 -469 3361 -454
rect 3309 -506 3361 -469
rect 3509 -94 3518 -79
rect 3518 -94 3552 -79
rect 3552 -94 3561 -79
rect 3509 -131 3561 -94
rect 3609 -74 3661 -22
rect 3809 177 3861 221
rect 3809 169 3818 177
rect 3818 169 3852 177
rect 3852 169 3861 177
rect 4009 283 4018 291
rect 4018 283 4052 291
rect 4052 283 4061 291
rect 4009 239 4061 283
rect 4209 457 4261 501
rect 4209 449 4218 457
rect 4218 449 4252 457
rect 4252 449 4261 457
rect 4409 563 4418 571
rect 4418 563 4452 571
rect 4452 563 4461 571
rect 4409 519 4461 563
rect 4609 737 4661 781
rect 4609 729 4618 737
rect 4618 729 4652 737
rect 4652 729 4661 737
rect 4809 843 4818 851
rect 4818 843 4852 851
rect 4852 843 4861 851
rect 4809 799 4861 843
rect 5009 1017 5061 1061
rect 5009 1009 5018 1017
rect 5018 1009 5052 1017
rect 5052 1009 5061 1017
rect 5209 1123 5218 1131
rect 5218 1123 5252 1131
rect 5252 1123 5261 1131
rect 5209 1079 5261 1123
rect 5409 1387 5461 1431
rect 5409 1379 5418 1387
rect 5418 1379 5452 1387
rect 5452 1379 5461 1387
rect 5609 1493 5618 1501
rect 5618 1493 5652 1501
rect 5652 1493 5661 1501
rect 5609 1449 5661 1493
rect 5809 1667 5861 1711
rect 5809 1659 5818 1667
rect 5818 1659 5852 1667
rect 5852 1659 5861 1667
rect 6009 1773 6018 1781
rect 6018 1773 6052 1781
rect 6052 1773 6061 1781
rect 6009 1729 6061 1773
rect 6209 1947 6261 1991
rect 6209 1939 6218 1947
rect 6218 1939 6252 1947
rect 6252 1939 6261 1947
rect 6409 2053 6418 2061
rect 6418 2053 6452 2061
rect 6452 2053 6461 2061
rect 6409 2009 6461 2053
rect 6609 2227 6661 2271
rect 6609 2219 6618 2227
rect 6618 2219 6652 2227
rect 6652 2219 6661 2227
rect 6809 2333 6818 2341
rect 6818 2333 6852 2341
rect 6852 2333 6861 2341
rect 6809 2289 6861 2333
rect 7009 2597 7061 2641
rect 7009 2589 7018 2597
rect 7018 2589 7052 2597
rect 7052 2589 7061 2597
rect 7209 2703 7218 2711
rect 7218 2703 7252 2711
rect 7252 2703 7261 2711
rect 7209 2659 7261 2703
rect 7409 2877 7461 2921
rect 7409 2869 7418 2877
rect 7418 2869 7452 2877
rect 7452 2869 7461 2877
rect 7609 2983 7618 2991
rect 7618 2983 7652 2991
rect 7652 2983 7661 2991
rect 7609 2939 7661 2983
rect 7809 3157 7861 3201
rect 7809 3149 7818 3157
rect 7818 3149 7852 3157
rect 7852 3149 7861 3157
rect 8009 3263 8018 3271
rect 8018 3263 8052 3271
rect 8052 3263 8061 3271
rect 8009 3219 8061 3263
rect 8209 3437 8261 3481
rect 8209 3429 8218 3437
rect 8218 3429 8252 3437
rect 8252 3429 8261 3437
rect 8409 3543 8418 3551
rect 8418 3543 8452 3551
rect 8452 3543 8461 3551
rect 8409 3499 8461 3543
rect 8609 3807 8661 3851
rect 8609 3799 8618 3807
rect 8618 3799 8652 3807
rect 8652 3799 8661 3807
rect 8809 3913 8818 3921
rect 8818 3913 8852 3921
rect 8852 3913 8861 3921
rect 8809 3869 8861 3913
rect 9009 4087 9061 4131
rect 9009 4079 9018 4087
rect 9018 4079 9052 4087
rect 9052 4079 9061 4087
rect 9209 4193 9218 4201
rect 9218 4193 9252 4201
rect 9252 4193 9261 4201
rect 9209 4149 9261 4193
rect 9409 4367 9461 4411
rect 9409 4359 9418 4367
rect 9418 4359 9452 4367
rect 9452 4359 9461 4367
rect 9609 4473 9618 4481
rect 9618 4473 9652 4481
rect 9652 4473 9661 4481
rect 9609 4429 9661 4473
rect 9809 4647 9861 4691
rect 9809 4639 9818 4647
rect 9818 4639 9852 4647
rect 9852 4639 9861 4647
rect 10009 4753 10018 4761
rect 10018 4753 10052 4761
rect 10052 4753 10061 4761
rect 10009 4709 10061 4753
rect 10209 4910 10261 4919
rect 10209 4876 10218 4910
rect 10218 4876 10252 4910
rect 10252 4876 10261 4910
rect 10209 4867 10261 4876
rect 8609 3700 8661 3709
rect 8609 3666 8618 3700
rect 8618 3666 8652 3700
rect 8652 3666 8661 3700
rect 8609 3657 8661 3666
rect 7009 2490 7061 2499
rect 7009 2456 7018 2490
rect 7018 2456 7052 2490
rect 7052 2456 7061 2490
rect 7009 2447 7061 2456
rect 5409 1280 5461 1289
rect 5409 1246 5418 1280
rect 5418 1246 5452 1280
rect 5452 1246 5461 1280
rect 5409 1237 5461 1246
rect 3809 70 3861 79
rect 3809 36 3818 70
rect 3818 36 3852 70
rect 3852 36 3861 70
rect 3809 27 3861 36
rect 3709 -60 3761 -15
rect 3709 -67 3718 -60
rect 3718 -67 3752 -60
rect 3752 -67 3761 -60
rect 3509 -166 3518 -143
rect 3518 -166 3552 -143
rect 3552 -166 3561 -143
rect 3509 -195 3561 -166
rect 3525 -248 3577 -239
rect 3525 -282 3534 -248
rect 3534 -282 3568 -248
rect 3568 -282 3577 -248
rect 3525 -291 3577 -282
rect 3509 -363 3561 -326
rect 3509 -378 3518 -363
rect 3518 -378 3552 -363
rect 3552 -378 3561 -363
rect 3509 -397 3518 -390
rect 3518 -397 3552 -390
rect 3552 -397 3561 -390
rect 3509 -435 3561 -397
rect 3509 -442 3518 -435
rect 3518 -442 3552 -435
rect 3552 -442 3561 -435
rect 3509 -469 3518 -454
rect 3518 -469 3552 -454
rect 3552 -469 3561 -454
rect 3509 -506 3561 -469
rect 3709 -94 3718 -79
rect 3718 -94 3752 -79
rect 3752 -94 3761 -79
rect 3709 -131 3761 -94
rect 3809 -74 3861 -22
rect 4009 143 4018 151
rect 4018 143 4052 151
rect 4052 143 4061 151
rect 4009 99 4061 143
rect 4209 317 4261 361
rect 4209 309 4218 317
rect 4218 309 4252 317
rect 4252 309 4261 317
rect 4409 423 4418 431
rect 4418 423 4452 431
rect 4452 423 4461 431
rect 4409 379 4461 423
rect 4609 597 4661 641
rect 4609 589 4618 597
rect 4618 589 4652 597
rect 4652 589 4661 597
rect 4809 703 4818 711
rect 4818 703 4852 711
rect 4852 703 4861 711
rect 4809 659 4861 703
rect 5009 877 5061 921
rect 5009 869 5018 877
rect 5018 869 5052 877
rect 5052 869 5061 877
rect 5209 983 5218 991
rect 5218 983 5252 991
rect 5252 983 5261 991
rect 5209 939 5261 983
rect 5409 1157 5461 1201
rect 5409 1149 5418 1157
rect 5418 1149 5452 1157
rect 5452 1149 5461 1157
rect 5609 1353 5618 1361
rect 5618 1353 5652 1361
rect 5652 1353 5661 1361
rect 5609 1309 5661 1353
rect 5809 1527 5861 1571
rect 5809 1519 5818 1527
rect 5818 1519 5852 1527
rect 5852 1519 5861 1527
rect 6009 1633 6018 1641
rect 6018 1633 6052 1641
rect 6052 1633 6061 1641
rect 6009 1589 6061 1633
rect 6209 1807 6261 1851
rect 6209 1799 6218 1807
rect 6218 1799 6252 1807
rect 6252 1799 6261 1807
rect 6409 1913 6418 1921
rect 6418 1913 6452 1921
rect 6452 1913 6461 1921
rect 6409 1869 6461 1913
rect 6609 2087 6661 2131
rect 6609 2079 6618 2087
rect 6618 2079 6652 2087
rect 6652 2079 6661 2087
rect 6809 2193 6818 2201
rect 6818 2193 6852 2201
rect 6852 2193 6861 2201
rect 6809 2149 6861 2193
rect 7009 2367 7061 2411
rect 7009 2359 7018 2367
rect 7018 2359 7052 2367
rect 7052 2359 7061 2367
rect 7209 2563 7218 2571
rect 7218 2563 7252 2571
rect 7252 2563 7261 2571
rect 7209 2519 7261 2563
rect 7409 2737 7461 2781
rect 7409 2729 7418 2737
rect 7418 2729 7452 2737
rect 7452 2729 7461 2737
rect 7609 2843 7618 2851
rect 7618 2843 7652 2851
rect 7652 2843 7661 2851
rect 7609 2799 7661 2843
rect 7809 3017 7861 3061
rect 7809 3009 7818 3017
rect 7818 3009 7852 3017
rect 7852 3009 7861 3017
rect 8009 3123 8018 3131
rect 8018 3123 8052 3131
rect 8052 3123 8061 3131
rect 8009 3079 8061 3123
rect 8209 3297 8261 3341
rect 8209 3289 8218 3297
rect 8218 3289 8252 3297
rect 8252 3289 8261 3297
rect 8409 3403 8418 3411
rect 8418 3403 8452 3411
rect 8452 3403 8461 3411
rect 8409 3359 8461 3403
rect 8609 3577 8661 3621
rect 8609 3569 8618 3577
rect 8618 3569 8652 3577
rect 8652 3569 8661 3577
rect 8809 3773 8818 3781
rect 8818 3773 8852 3781
rect 8852 3773 8861 3781
rect 8809 3729 8861 3773
rect 9009 3947 9061 3991
rect 9009 3939 9018 3947
rect 9018 3939 9052 3947
rect 9052 3939 9061 3947
rect 9209 4053 9218 4061
rect 9218 4053 9252 4061
rect 9252 4053 9261 4061
rect 9209 4009 9261 4053
rect 9409 4227 9461 4271
rect 9409 4219 9418 4227
rect 9418 4219 9452 4227
rect 9452 4219 9461 4227
rect 9609 4333 9618 4341
rect 9618 4333 9652 4341
rect 9652 4333 9661 4341
rect 9609 4289 9661 4333
rect 9809 4507 9861 4551
rect 9809 4499 9818 4507
rect 9818 4499 9852 4507
rect 9852 4499 9861 4507
rect 10009 4613 10018 4621
rect 10018 4613 10052 4621
rect 10052 4613 10061 4621
rect 10009 4569 10061 4613
rect 10209 4787 10261 4831
rect 10209 4779 10218 4787
rect 10218 4779 10252 4787
rect 10252 4779 10261 4787
rect 10409 4894 10461 4903
rect 10409 4860 10418 4894
rect 10418 4860 10452 4894
rect 10452 4860 10461 4894
rect 10409 4851 10461 4860
rect 8809 3684 8861 3693
rect 8809 3650 8818 3684
rect 8818 3650 8852 3684
rect 8852 3650 8861 3684
rect 8809 3641 8861 3650
rect 7209 2474 7261 2483
rect 7209 2440 7218 2474
rect 7218 2440 7252 2474
rect 7252 2440 7261 2474
rect 7209 2431 7261 2440
rect 5609 1264 5661 1273
rect 5609 1230 5618 1264
rect 5618 1230 5652 1264
rect 5652 1230 5661 1264
rect 5609 1221 5661 1230
rect 4009 54 4061 63
rect 4009 20 4018 54
rect 4018 20 4052 54
rect 4052 20 4061 54
rect 4009 11 4061 20
rect 3909 -60 3961 -15
rect 3909 -67 3918 -60
rect 3918 -67 3952 -60
rect 3952 -67 3961 -60
rect 3709 -166 3718 -143
rect 3718 -166 3752 -143
rect 3752 -166 3761 -143
rect 3709 -195 3761 -166
rect 3725 -248 3777 -239
rect 3725 -282 3734 -248
rect 3734 -282 3768 -248
rect 3768 -282 3777 -248
rect 3725 -291 3777 -282
rect 3709 -363 3761 -326
rect 3709 -378 3718 -363
rect 3718 -378 3752 -363
rect 3752 -378 3761 -363
rect 3709 -397 3718 -390
rect 3718 -397 3752 -390
rect 3752 -397 3761 -390
rect 3709 -435 3761 -397
rect 3709 -442 3718 -435
rect 3718 -442 3752 -435
rect 3752 -442 3761 -435
rect 3709 -469 3718 -454
rect 3718 -469 3752 -454
rect 3752 -469 3761 -454
rect 3709 -506 3761 -469
rect 3909 -94 3918 -79
rect 3918 -94 3952 -79
rect 3952 -94 3961 -79
rect 3909 -131 3961 -94
rect 4009 -74 4061 -22
rect 4209 177 4261 221
rect 4209 169 4218 177
rect 4218 169 4252 177
rect 4252 169 4261 177
rect 4409 283 4418 291
rect 4418 283 4452 291
rect 4452 283 4461 291
rect 4409 239 4461 283
rect 4609 457 4661 501
rect 4609 449 4618 457
rect 4618 449 4652 457
rect 4652 449 4661 457
rect 4809 563 4818 571
rect 4818 563 4852 571
rect 4852 563 4861 571
rect 4809 519 4861 563
rect 5009 737 5061 781
rect 5009 729 5018 737
rect 5018 729 5052 737
rect 5052 729 5061 737
rect 5209 843 5218 851
rect 5218 843 5252 851
rect 5252 843 5261 851
rect 5209 799 5261 843
rect 5409 1017 5461 1061
rect 5409 1009 5418 1017
rect 5418 1009 5452 1017
rect 5452 1009 5461 1017
rect 5609 1123 5618 1131
rect 5618 1123 5652 1131
rect 5652 1123 5661 1131
rect 5609 1079 5661 1123
rect 5809 1387 5861 1431
rect 5809 1379 5818 1387
rect 5818 1379 5852 1387
rect 5852 1379 5861 1387
rect 6009 1493 6018 1501
rect 6018 1493 6052 1501
rect 6052 1493 6061 1501
rect 6009 1449 6061 1493
rect 6209 1667 6261 1711
rect 6209 1659 6218 1667
rect 6218 1659 6252 1667
rect 6252 1659 6261 1667
rect 6409 1773 6418 1781
rect 6418 1773 6452 1781
rect 6452 1773 6461 1781
rect 6409 1729 6461 1773
rect 6609 1947 6661 1991
rect 6609 1939 6618 1947
rect 6618 1939 6652 1947
rect 6652 1939 6661 1947
rect 6809 2053 6818 2061
rect 6818 2053 6852 2061
rect 6852 2053 6861 2061
rect 6809 2009 6861 2053
rect 7009 2227 7061 2271
rect 7009 2219 7018 2227
rect 7018 2219 7052 2227
rect 7052 2219 7061 2227
rect 7209 2333 7218 2341
rect 7218 2333 7252 2341
rect 7252 2333 7261 2341
rect 7209 2289 7261 2333
rect 7409 2597 7461 2641
rect 7409 2589 7418 2597
rect 7418 2589 7452 2597
rect 7452 2589 7461 2597
rect 7609 2703 7618 2711
rect 7618 2703 7652 2711
rect 7652 2703 7661 2711
rect 7609 2659 7661 2703
rect 7809 2877 7861 2921
rect 7809 2869 7818 2877
rect 7818 2869 7852 2877
rect 7852 2869 7861 2877
rect 8009 2983 8018 2991
rect 8018 2983 8052 2991
rect 8052 2983 8061 2991
rect 8009 2939 8061 2983
rect 8209 3157 8261 3201
rect 8209 3149 8218 3157
rect 8218 3149 8252 3157
rect 8252 3149 8261 3157
rect 8409 3263 8418 3271
rect 8418 3263 8452 3271
rect 8452 3263 8461 3271
rect 8409 3219 8461 3263
rect 8609 3437 8661 3481
rect 8609 3429 8618 3437
rect 8618 3429 8652 3437
rect 8652 3429 8661 3437
rect 8809 3543 8818 3551
rect 8818 3543 8852 3551
rect 8852 3543 8861 3551
rect 8809 3499 8861 3543
rect 9009 3807 9061 3851
rect 9009 3799 9018 3807
rect 9018 3799 9052 3807
rect 9052 3799 9061 3807
rect 9209 3913 9218 3921
rect 9218 3913 9252 3921
rect 9252 3913 9261 3921
rect 9209 3869 9261 3913
rect 9409 4087 9461 4131
rect 9409 4079 9418 4087
rect 9418 4079 9452 4087
rect 9452 4079 9461 4087
rect 9609 4193 9618 4201
rect 9618 4193 9652 4201
rect 9652 4193 9661 4201
rect 9609 4149 9661 4193
rect 9809 4367 9861 4411
rect 9809 4359 9818 4367
rect 9818 4359 9852 4367
rect 9852 4359 9861 4367
rect 10009 4473 10018 4481
rect 10018 4473 10052 4481
rect 10052 4473 10061 4481
rect 10009 4429 10061 4473
rect 10209 4647 10261 4691
rect 10209 4639 10218 4647
rect 10218 4639 10252 4647
rect 10252 4639 10261 4647
rect 10409 4753 10418 4761
rect 10418 4753 10452 4761
rect 10452 4753 10461 4761
rect 10409 4709 10461 4753
rect 10609 4910 10661 4919
rect 10609 4876 10618 4910
rect 10618 4876 10652 4910
rect 10652 4876 10661 4910
rect 10609 4867 10661 4876
rect 9009 3700 9061 3709
rect 9009 3666 9018 3700
rect 9018 3666 9052 3700
rect 9052 3666 9061 3700
rect 9009 3657 9061 3666
rect 7409 2490 7461 2499
rect 7409 2456 7418 2490
rect 7418 2456 7452 2490
rect 7452 2456 7461 2490
rect 7409 2447 7461 2456
rect 5809 1280 5861 1289
rect 5809 1246 5818 1280
rect 5818 1246 5852 1280
rect 5852 1246 5861 1280
rect 5809 1237 5861 1246
rect 4209 70 4261 79
rect 4209 36 4218 70
rect 4218 36 4252 70
rect 4252 36 4261 70
rect 4209 27 4261 36
rect 4109 -60 4161 -15
rect 4109 -67 4118 -60
rect 4118 -67 4152 -60
rect 4152 -67 4161 -60
rect 3909 -166 3918 -143
rect 3918 -166 3952 -143
rect 3952 -166 3961 -143
rect 3909 -195 3961 -166
rect 3925 -248 3977 -239
rect 3925 -282 3934 -248
rect 3934 -282 3968 -248
rect 3968 -282 3977 -248
rect 3925 -291 3977 -282
rect 3909 -363 3961 -326
rect 3909 -378 3918 -363
rect 3918 -378 3952 -363
rect 3952 -378 3961 -363
rect 3909 -397 3918 -390
rect 3918 -397 3952 -390
rect 3952 -397 3961 -390
rect 3909 -435 3961 -397
rect 3909 -442 3918 -435
rect 3918 -442 3952 -435
rect 3952 -442 3961 -435
rect 3909 -469 3918 -454
rect 3918 -469 3952 -454
rect 3952 -469 3961 -454
rect 3909 -506 3961 -469
rect 4109 -94 4118 -79
rect 4118 -94 4152 -79
rect 4152 -94 4161 -79
rect 4109 -131 4161 -94
rect 4209 -74 4261 -22
rect 4409 143 4418 151
rect 4418 143 4452 151
rect 4452 143 4461 151
rect 4409 99 4461 143
rect 4609 317 4661 361
rect 4609 309 4618 317
rect 4618 309 4652 317
rect 4652 309 4661 317
rect 4809 423 4818 431
rect 4818 423 4852 431
rect 4852 423 4861 431
rect 4809 379 4861 423
rect 5009 597 5061 641
rect 5009 589 5018 597
rect 5018 589 5052 597
rect 5052 589 5061 597
rect 5209 703 5218 711
rect 5218 703 5252 711
rect 5252 703 5261 711
rect 5209 659 5261 703
rect 5409 877 5461 921
rect 5409 869 5418 877
rect 5418 869 5452 877
rect 5452 869 5461 877
rect 5609 983 5618 991
rect 5618 983 5652 991
rect 5652 983 5661 991
rect 5609 939 5661 983
rect 5809 1157 5861 1201
rect 5809 1149 5818 1157
rect 5818 1149 5852 1157
rect 5852 1149 5861 1157
rect 6009 1353 6018 1361
rect 6018 1353 6052 1361
rect 6052 1353 6061 1361
rect 6009 1309 6061 1353
rect 6209 1527 6261 1571
rect 6209 1519 6218 1527
rect 6218 1519 6252 1527
rect 6252 1519 6261 1527
rect 6409 1633 6418 1641
rect 6418 1633 6452 1641
rect 6452 1633 6461 1641
rect 6409 1589 6461 1633
rect 6609 1807 6661 1851
rect 6609 1799 6618 1807
rect 6618 1799 6652 1807
rect 6652 1799 6661 1807
rect 6809 1913 6818 1921
rect 6818 1913 6852 1921
rect 6852 1913 6861 1921
rect 6809 1869 6861 1913
rect 7009 2087 7061 2131
rect 7009 2079 7018 2087
rect 7018 2079 7052 2087
rect 7052 2079 7061 2087
rect 7209 2193 7218 2201
rect 7218 2193 7252 2201
rect 7252 2193 7261 2201
rect 7209 2149 7261 2193
rect 7409 2367 7461 2411
rect 7409 2359 7418 2367
rect 7418 2359 7452 2367
rect 7452 2359 7461 2367
rect 7609 2563 7618 2571
rect 7618 2563 7652 2571
rect 7652 2563 7661 2571
rect 7609 2519 7661 2563
rect 7809 2737 7861 2781
rect 7809 2729 7818 2737
rect 7818 2729 7852 2737
rect 7852 2729 7861 2737
rect 8009 2843 8018 2851
rect 8018 2843 8052 2851
rect 8052 2843 8061 2851
rect 8009 2799 8061 2843
rect 8209 3017 8261 3061
rect 8209 3009 8218 3017
rect 8218 3009 8252 3017
rect 8252 3009 8261 3017
rect 8409 3123 8418 3131
rect 8418 3123 8452 3131
rect 8452 3123 8461 3131
rect 8409 3079 8461 3123
rect 8609 3297 8661 3341
rect 8609 3289 8618 3297
rect 8618 3289 8652 3297
rect 8652 3289 8661 3297
rect 8809 3403 8818 3411
rect 8818 3403 8852 3411
rect 8852 3403 8861 3411
rect 8809 3359 8861 3403
rect 9009 3577 9061 3621
rect 9009 3569 9018 3577
rect 9018 3569 9052 3577
rect 9052 3569 9061 3577
rect 9209 3773 9218 3781
rect 9218 3773 9252 3781
rect 9252 3773 9261 3781
rect 9209 3729 9261 3773
rect 9409 3947 9461 3991
rect 9409 3939 9418 3947
rect 9418 3939 9452 3947
rect 9452 3939 9461 3947
rect 9609 4053 9618 4061
rect 9618 4053 9652 4061
rect 9652 4053 9661 4061
rect 9609 4009 9661 4053
rect 9809 4227 9861 4271
rect 9809 4219 9818 4227
rect 9818 4219 9852 4227
rect 9852 4219 9861 4227
rect 10009 4333 10018 4341
rect 10018 4333 10052 4341
rect 10052 4333 10061 4341
rect 10009 4289 10061 4333
rect 10209 4507 10261 4551
rect 10209 4499 10218 4507
rect 10218 4499 10252 4507
rect 10252 4499 10261 4507
rect 10409 4613 10418 4621
rect 10418 4613 10452 4621
rect 10452 4613 10461 4621
rect 10409 4569 10461 4613
rect 10609 4787 10661 4831
rect 10609 4779 10618 4787
rect 10618 4779 10652 4787
rect 10652 4779 10661 4787
rect 10809 4894 10861 4903
rect 10809 4860 10818 4894
rect 10818 4860 10852 4894
rect 10852 4860 10861 4894
rect 10809 4851 10861 4860
rect 9209 3684 9261 3693
rect 9209 3650 9218 3684
rect 9218 3650 9252 3684
rect 9252 3650 9261 3684
rect 9209 3641 9261 3650
rect 7609 2474 7661 2483
rect 7609 2440 7618 2474
rect 7618 2440 7652 2474
rect 7652 2440 7661 2474
rect 7609 2431 7661 2440
rect 6009 1264 6061 1273
rect 6009 1230 6018 1264
rect 6018 1230 6052 1264
rect 6052 1230 6061 1264
rect 6009 1221 6061 1230
rect 4409 54 4461 63
rect 4409 20 4418 54
rect 4418 20 4452 54
rect 4452 20 4461 54
rect 4409 11 4461 20
rect 4309 -60 4361 -15
rect 4309 -67 4318 -60
rect 4318 -67 4352 -60
rect 4352 -67 4361 -60
rect 4109 -166 4118 -143
rect 4118 -166 4152 -143
rect 4152 -166 4161 -143
rect 4109 -195 4161 -166
rect 4125 -248 4177 -239
rect 4125 -282 4134 -248
rect 4134 -282 4168 -248
rect 4168 -282 4177 -248
rect 4125 -291 4177 -282
rect 4109 -363 4161 -326
rect 4109 -378 4118 -363
rect 4118 -378 4152 -363
rect 4152 -378 4161 -363
rect 4109 -397 4118 -390
rect 4118 -397 4152 -390
rect 4152 -397 4161 -390
rect 4109 -435 4161 -397
rect 4109 -442 4118 -435
rect 4118 -442 4152 -435
rect 4152 -442 4161 -435
rect 4109 -469 4118 -454
rect 4118 -469 4152 -454
rect 4152 -469 4161 -454
rect 4109 -506 4161 -469
rect 4309 -94 4318 -79
rect 4318 -94 4352 -79
rect 4352 -94 4361 -79
rect 4309 -131 4361 -94
rect 4409 -74 4461 -22
rect 4609 177 4661 221
rect 4609 169 4618 177
rect 4618 169 4652 177
rect 4652 169 4661 177
rect 4809 283 4818 291
rect 4818 283 4852 291
rect 4852 283 4861 291
rect 4809 239 4861 283
rect 5009 457 5061 501
rect 5009 449 5018 457
rect 5018 449 5052 457
rect 5052 449 5061 457
rect 5209 563 5218 571
rect 5218 563 5252 571
rect 5252 563 5261 571
rect 5209 519 5261 563
rect 5409 737 5461 781
rect 5409 729 5418 737
rect 5418 729 5452 737
rect 5452 729 5461 737
rect 5609 843 5618 851
rect 5618 843 5652 851
rect 5652 843 5661 851
rect 5609 799 5661 843
rect 5809 1017 5861 1061
rect 5809 1009 5818 1017
rect 5818 1009 5852 1017
rect 5852 1009 5861 1017
rect 6009 1123 6018 1131
rect 6018 1123 6052 1131
rect 6052 1123 6061 1131
rect 6009 1079 6061 1123
rect 6209 1387 6261 1431
rect 6209 1379 6218 1387
rect 6218 1379 6252 1387
rect 6252 1379 6261 1387
rect 6409 1493 6418 1501
rect 6418 1493 6452 1501
rect 6452 1493 6461 1501
rect 6409 1449 6461 1493
rect 6609 1667 6661 1711
rect 6609 1659 6618 1667
rect 6618 1659 6652 1667
rect 6652 1659 6661 1667
rect 6809 1773 6818 1781
rect 6818 1773 6852 1781
rect 6852 1773 6861 1781
rect 6809 1729 6861 1773
rect 7009 1947 7061 1991
rect 7009 1939 7018 1947
rect 7018 1939 7052 1947
rect 7052 1939 7061 1947
rect 7209 2053 7218 2061
rect 7218 2053 7252 2061
rect 7252 2053 7261 2061
rect 7209 2009 7261 2053
rect 7409 2227 7461 2271
rect 7409 2219 7418 2227
rect 7418 2219 7452 2227
rect 7452 2219 7461 2227
rect 7609 2333 7618 2341
rect 7618 2333 7652 2341
rect 7652 2333 7661 2341
rect 7609 2289 7661 2333
rect 7809 2597 7861 2641
rect 7809 2589 7818 2597
rect 7818 2589 7852 2597
rect 7852 2589 7861 2597
rect 8009 2703 8018 2711
rect 8018 2703 8052 2711
rect 8052 2703 8061 2711
rect 8009 2659 8061 2703
rect 8209 2877 8261 2921
rect 8209 2869 8218 2877
rect 8218 2869 8252 2877
rect 8252 2869 8261 2877
rect 8409 2983 8418 2991
rect 8418 2983 8452 2991
rect 8452 2983 8461 2991
rect 8409 2939 8461 2983
rect 8609 3157 8661 3201
rect 8609 3149 8618 3157
rect 8618 3149 8652 3157
rect 8652 3149 8661 3157
rect 8809 3263 8818 3271
rect 8818 3263 8852 3271
rect 8852 3263 8861 3271
rect 8809 3219 8861 3263
rect 9009 3437 9061 3481
rect 9009 3429 9018 3437
rect 9018 3429 9052 3437
rect 9052 3429 9061 3437
rect 9209 3543 9218 3551
rect 9218 3543 9252 3551
rect 9252 3543 9261 3551
rect 9209 3499 9261 3543
rect 9409 3807 9461 3851
rect 9409 3799 9418 3807
rect 9418 3799 9452 3807
rect 9452 3799 9461 3807
rect 9609 3913 9618 3921
rect 9618 3913 9652 3921
rect 9652 3913 9661 3921
rect 9609 3869 9661 3913
rect 9809 4087 9861 4131
rect 9809 4079 9818 4087
rect 9818 4079 9852 4087
rect 9852 4079 9861 4087
rect 10009 4193 10018 4201
rect 10018 4193 10052 4201
rect 10052 4193 10061 4201
rect 10009 4149 10061 4193
rect 10209 4367 10261 4411
rect 10209 4359 10218 4367
rect 10218 4359 10252 4367
rect 10252 4359 10261 4367
rect 10409 4473 10418 4481
rect 10418 4473 10452 4481
rect 10452 4473 10461 4481
rect 10409 4429 10461 4473
rect 10609 4647 10661 4691
rect 10609 4639 10618 4647
rect 10618 4639 10652 4647
rect 10652 4639 10661 4647
rect 10809 4753 10818 4761
rect 10818 4753 10852 4761
rect 10852 4753 10861 4761
rect 10809 4709 10861 4753
rect 11009 4910 11061 4919
rect 11009 4876 11018 4910
rect 11018 4876 11052 4910
rect 11052 4876 11061 4910
rect 11009 4867 11061 4876
rect 9409 3700 9461 3709
rect 9409 3666 9418 3700
rect 9418 3666 9452 3700
rect 9452 3666 9461 3700
rect 9409 3657 9461 3666
rect 7809 2490 7861 2499
rect 7809 2456 7818 2490
rect 7818 2456 7852 2490
rect 7852 2456 7861 2490
rect 7809 2447 7861 2456
rect 6209 1280 6261 1289
rect 6209 1246 6218 1280
rect 6218 1246 6252 1280
rect 6252 1246 6261 1280
rect 6209 1237 6261 1246
rect 4609 70 4661 79
rect 4609 36 4618 70
rect 4618 36 4652 70
rect 4652 36 4661 70
rect 4609 27 4661 36
rect 4509 -60 4561 -15
rect 4509 -67 4518 -60
rect 4518 -67 4552 -60
rect 4552 -67 4561 -60
rect 4309 -166 4318 -143
rect 4318 -166 4352 -143
rect 4352 -166 4361 -143
rect 4309 -195 4361 -166
rect 4325 -248 4377 -239
rect 4325 -282 4334 -248
rect 4334 -282 4368 -248
rect 4368 -282 4377 -248
rect 4325 -291 4377 -282
rect 4309 -363 4361 -326
rect 4309 -378 4318 -363
rect 4318 -378 4352 -363
rect 4352 -378 4361 -363
rect 4309 -397 4318 -390
rect 4318 -397 4352 -390
rect 4352 -397 4361 -390
rect 4309 -435 4361 -397
rect 4309 -442 4318 -435
rect 4318 -442 4352 -435
rect 4352 -442 4361 -435
rect 4309 -469 4318 -454
rect 4318 -469 4352 -454
rect 4352 -469 4361 -454
rect 4309 -506 4361 -469
rect 4509 -94 4518 -79
rect 4518 -94 4552 -79
rect 4552 -94 4561 -79
rect 4509 -131 4561 -94
rect 4609 -74 4661 -22
rect 4809 143 4818 151
rect 4818 143 4852 151
rect 4852 143 4861 151
rect 4809 99 4861 143
rect 5009 317 5061 361
rect 5009 309 5018 317
rect 5018 309 5052 317
rect 5052 309 5061 317
rect 5209 423 5218 431
rect 5218 423 5252 431
rect 5252 423 5261 431
rect 5209 379 5261 423
rect 5409 597 5461 641
rect 5409 589 5418 597
rect 5418 589 5452 597
rect 5452 589 5461 597
rect 5609 703 5618 711
rect 5618 703 5652 711
rect 5652 703 5661 711
rect 5609 659 5661 703
rect 5809 877 5861 921
rect 5809 869 5818 877
rect 5818 869 5852 877
rect 5852 869 5861 877
rect 6009 983 6018 991
rect 6018 983 6052 991
rect 6052 983 6061 991
rect 6009 939 6061 983
rect 6209 1157 6261 1201
rect 6209 1149 6218 1157
rect 6218 1149 6252 1157
rect 6252 1149 6261 1157
rect 6409 1353 6418 1361
rect 6418 1353 6452 1361
rect 6452 1353 6461 1361
rect 6409 1309 6461 1353
rect 6609 1527 6661 1571
rect 6609 1519 6618 1527
rect 6618 1519 6652 1527
rect 6652 1519 6661 1527
rect 6809 1633 6818 1641
rect 6818 1633 6852 1641
rect 6852 1633 6861 1641
rect 6809 1589 6861 1633
rect 7009 1807 7061 1851
rect 7009 1799 7018 1807
rect 7018 1799 7052 1807
rect 7052 1799 7061 1807
rect 7209 1913 7218 1921
rect 7218 1913 7252 1921
rect 7252 1913 7261 1921
rect 7209 1869 7261 1913
rect 7409 2087 7461 2131
rect 7409 2079 7418 2087
rect 7418 2079 7452 2087
rect 7452 2079 7461 2087
rect 7609 2193 7618 2201
rect 7618 2193 7652 2201
rect 7652 2193 7661 2201
rect 7609 2149 7661 2193
rect 7809 2367 7861 2411
rect 7809 2359 7818 2367
rect 7818 2359 7852 2367
rect 7852 2359 7861 2367
rect 8009 2563 8018 2571
rect 8018 2563 8052 2571
rect 8052 2563 8061 2571
rect 8009 2519 8061 2563
rect 8209 2737 8261 2781
rect 8209 2729 8218 2737
rect 8218 2729 8252 2737
rect 8252 2729 8261 2737
rect 8409 2843 8418 2851
rect 8418 2843 8452 2851
rect 8452 2843 8461 2851
rect 8409 2799 8461 2843
rect 8609 3017 8661 3061
rect 8609 3009 8618 3017
rect 8618 3009 8652 3017
rect 8652 3009 8661 3017
rect 8809 3123 8818 3131
rect 8818 3123 8852 3131
rect 8852 3123 8861 3131
rect 8809 3079 8861 3123
rect 9009 3297 9061 3341
rect 9009 3289 9018 3297
rect 9018 3289 9052 3297
rect 9052 3289 9061 3297
rect 9209 3403 9218 3411
rect 9218 3403 9252 3411
rect 9252 3403 9261 3411
rect 9209 3359 9261 3403
rect 9409 3577 9461 3621
rect 9409 3569 9418 3577
rect 9418 3569 9452 3577
rect 9452 3569 9461 3577
rect 9609 3773 9618 3781
rect 9618 3773 9652 3781
rect 9652 3773 9661 3781
rect 9609 3729 9661 3773
rect 9809 3947 9861 3991
rect 9809 3939 9818 3947
rect 9818 3939 9852 3947
rect 9852 3939 9861 3947
rect 10009 4053 10018 4061
rect 10018 4053 10052 4061
rect 10052 4053 10061 4061
rect 10009 4009 10061 4053
rect 10209 4227 10261 4271
rect 10209 4219 10218 4227
rect 10218 4219 10252 4227
rect 10252 4219 10261 4227
rect 10409 4333 10418 4341
rect 10418 4333 10452 4341
rect 10452 4333 10461 4341
rect 10409 4289 10461 4333
rect 10609 4507 10661 4551
rect 10609 4499 10618 4507
rect 10618 4499 10652 4507
rect 10652 4499 10661 4507
rect 10809 4613 10818 4621
rect 10818 4613 10852 4621
rect 10852 4613 10861 4621
rect 10809 4569 10861 4613
rect 11009 4787 11061 4831
rect 11009 4779 11018 4787
rect 11018 4779 11052 4787
rect 11052 4779 11061 4787
rect 11209 4894 11261 4903
rect 11209 4860 11218 4894
rect 11218 4860 11252 4894
rect 11252 4860 11261 4894
rect 11209 4851 11261 4860
rect 9609 3684 9661 3693
rect 9609 3650 9618 3684
rect 9618 3650 9652 3684
rect 9652 3650 9661 3684
rect 9609 3641 9661 3650
rect 8009 2474 8061 2483
rect 8009 2440 8018 2474
rect 8018 2440 8052 2474
rect 8052 2440 8061 2474
rect 8009 2431 8061 2440
rect 6409 1264 6461 1273
rect 6409 1230 6418 1264
rect 6418 1230 6452 1264
rect 6452 1230 6461 1264
rect 6409 1221 6461 1230
rect 4809 54 4861 63
rect 4809 20 4818 54
rect 4818 20 4852 54
rect 4852 20 4861 54
rect 4809 11 4861 20
rect 4709 -60 4761 -15
rect 4709 -67 4718 -60
rect 4718 -67 4752 -60
rect 4752 -67 4761 -60
rect 4509 -166 4518 -143
rect 4518 -166 4552 -143
rect 4552 -166 4561 -143
rect 4509 -195 4561 -166
rect 4525 -248 4577 -239
rect 4525 -282 4534 -248
rect 4534 -282 4568 -248
rect 4568 -282 4577 -248
rect 4525 -291 4577 -282
rect 4509 -363 4561 -326
rect 4509 -378 4518 -363
rect 4518 -378 4552 -363
rect 4552 -378 4561 -363
rect 4509 -397 4518 -390
rect 4518 -397 4552 -390
rect 4552 -397 4561 -390
rect 4509 -435 4561 -397
rect 4509 -442 4518 -435
rect 4518 -442 4552 -435
rect 4552 -442 4561 -435
rect 4509 -469 4518 -454
rect 4518 -469 4552 -454
rect 4552 -469 4561 -454
rect 4509 -506 4561 -469
rect 4709 -94 4718 -79
rect 4718 -94 4752 -79
rect 4752 -94 4761 -79
rect 4709 -131 4761 -94
rect 4809 -74 4861 -22
rect 5009 177 5061 221
rect 5009 169 5018 177
rect 5018 169 5052 177
rect 5052 169 5061 177
rect 5209 283 5218 291
rect 5218 283 5252 291
rect 5252 283 5261 291
rect 5209 239 5261 283
rect 5409 457 5461 501
rect 5409 449 5418 457
rect 5418 449 5452 457
rect 5452 449 5461 457
rect 5609 563 5618 571
rect 5618 563 5652 571
rect 5652 563 5661 571
rect 5609 519 5661 563
rect 5809 737 5861 781
rect 5809 729 5818 737
rect 5818 729 5852 737
rect 5852 729 5861 737
rect 6009 843 6018 851
rect 6018 843 6052 851
rect 6052 843 6061 851
rect 6009 799 6061 843
rect 6209 1017 6261 1061
rect 6209 1009 6218 1017
rect 6218 1009 6252 1017
rect 6252 1009 6261 1017
rect 6409 1123 6418 1131
rect 6418 1123 6452 1131
rect 6452 1123 6461 1131
rect 6409 1079 6461 1123
rect 6609 1387 6661 1431
rect 6609 1379 6618 1387
rect 6618 1379 6652 1387
rect 6652 1379 6661 1387
rect 6809 1493 6818 1501
rect 6818 1493 6852 1501
rect 6852 1493 6861 1501
rect 6809 1449 6861 1493
rect 7009 1667 7061 1711
rect 7009 1659 7018 1667
rect 7018 1659 7052 1667
rect 7052 1659 7061 1667
rect 7209 1773 7218 1781
rect 7218 1773 7252 1781
rect 7252 1773 7261 1781
rect 7209 1729 7261 1773
rect 7409 1947 7461 1991
rect 7409 1939 7418 1947
rect 7418 1939 7452 1947
rect 7452 1939 7461 1947
rect 7609 2053 7618 2061
rect 7618 2053 7652 2061
rect 7652 2053 7661 2061
rect 7609 2009 7661 2053
rect 7809 2227 7861 2271
rect 7809 2219 7818 2227
rect 7818 2219 7852 2227
rect 7852 2219 7861 2227
rect 8009 2333 8018 2341
rect 8018 2333 8052 2341
rect 8052 2333 8061 2341
rect 8009 2289 8061 2333
rect 8209 2597 8261 2641
rect 8209 2589 8218 2597
rect 8218 2589 8252 2597
rect 8252 2589 8261 2597
rect 8409 2703 8418 2711
rect 8418 2703 8452 2711
rect 8452 2703 8461 2711
rect 8409 2659 8461 2703
rect 8609 2877 8661 2921
rect 8609 2869 8618 2877
rect 8618 2869 8652 2877
rect 8652 2869 8661 2877
rect 8809 2983 8818 2991
rect 8818 2983 8852 2991
rect 8852 2983 8861 2991
rect 8809 2939 8861 2983
rect 9009 3157 9061 3201
rect 9009 3149 9018 3157
rect 9018 3149 9052 3157
rect 9052 3149 9061 3157
rect 9209 3263 9218 3271
rect 9218 3263 9252 3271
rect 9252 3263 9261 3271
rect 9209 3219 9261 3263
rect 9409 3437 9461 3481
rect 9409 3429 9418 3437
rect 9418 3429 9452 3437
rect 9452 3429 9461 3437
rect 9609 3543 9618 3551
rect 9618 3543 9652 3551
rect 9652 3543 9661 3551
rect 9609 3499 9661 3543
rect 9809 3807 9861 3851
rect 9809 3799 9818 3807
rect 9818 3799 9852 3807
rect 9852 3799 9861 3807
rect 10009 3913 10018 3921
rect 10018 3913 10052 3921
rect 10052 3913 10061 3921
rect 10009 3869 10061 3913
rect 10209 4087 10261 4131
rect 10209 4079 10218 4087
rect 10218 4079 10252 4087
rect 10252 4079 10261 4087
rect 10409 4193 10418 4201
rect 10418 4193 10452 4201
rect 10452 4193 10461 4201
rect 10409 4149 10461 4193
rect 10609 4367 10661 4411
rect 10609 4359 10618 4367
rect 10618 4359 10652 4367
rect 10652 4359 10661 4367
rect 10809 4473 10818 4481
rect 10818 4473 10852 4481
rect 10852 4473 10861 4481
rect 10809 4429 10861 4473
rect 11009 4647 11061 4691
rect 11009 4639 11018 4647
rect 11018 4639 11052 4647
rect 11052 4639 11061 4647
rect 11209 4753 11218 4761
rect 11218 4753 11252 4761
rect 11252 4753 11261 4761
rect 11209 4709 11261 4753
rect 11409 4910 11461 4919
rect 11409 4876 11418 4910
rect 11418 4876 11452 4910
rect 11452 4876 11461 4910
rect 11409 4867 11461 4876
rect 9809 3700 9861 3709
rect 9809 3666 9818 3700
rect 9818 3666 9852 3700
rect 9852 3666 9861 3700
rect 9809 3657 9861 3666
rect 8209 2490 8261 2499
rect 8209 2456 8218 2490
rect 8218 2456 8252 2490
rect 8252 2456 8261 2490
rect 8209 2447 8261 2456
rect 6609 1280 6661 1289
rect 6609 1246 6618 1280
rect 6618 1246 6652 1280
rect 6652 1246 6661 1280
rect 6609 1237 6661 1246
rect 5009 70 5061 79
rect 5009 36 5018 70
rect 5018 36 5052 70
rect 5052 36 5061 70
rect 5009 27 5061 36
rect 4909 -60 4961 -15
rect 4909 -67 4918 -60
rect 4918 -67 4952 -60
rect 4952 -67 4961 -60
rect 4709 -166 4718 -143
rect 4718 -166 4752 -143
rect 4752 -166 4761 -143
rect 4709 -195 4761 -166
rect 4725 -248 4777 -239
rect 4725 -282 4734 -248
rect 4734 -282 4768 -248
rect 4768 -282 4777 -248
rect 4725 -291 4777 -282
rect 4709 -363 4761 -326
rect 4709 -378 4718 -363
rect 4718 -378 4752 -363
rect 4752 -378 4761 -363
rect 4709 -397 4718 -390
rect 4718 -397 4752 -390
rect 4752 -397 4761 -390
rect 4709 -435 4761 -397
rect 4709 -442 4718 -435
rect 4718 -442 4752 -435
rect 4752 -442 4761 -435
rect 4709 -469 4718 -454
rect 4718 -469 4752 -454
rect 4752 -469 4761 -454
rect 4709 -506 4761 -469
rect 4909 -94 4918 -79
rect 4918 -94 4952 -79
rect 4952 -94 4961 -79
rect 4909 -131 4961 -94
rect 5009 -74 5061 -22
rect 5209 143 5218 151
rect 5218 143 5252 151
rect 5252 143 5261 151
rect 5209 99 5261 143
rect 5409 317 5461 361
rect 5409 309 5418 317
rect 5418 309 5452 317
rect 5452 309 5461 317
rect 5609 423 5618 431
rect 5618 423 5652 431
rect 5652 423 5661 431
rect 5609 379 5661 423
rect 5809 597 5861 641
rect 5809 589 5818 597
rect 5818 589 5852 597
rect 5852 589 5861 597
rect 6009 703 6018 711
rect 6018 703 6052 711
rect 6052 703 6061 711
rect 6009 659 6061 703
rect 6209 877 6261 921
rect 6209 869 6218 877
rect 6218 869 6252 877
rect 6252 869 6261 877
rect 6409 983 6418 991
rect 6418 983 6452 991
rect 6452 983 6461 991
rect 6409 939 6461 983
rect 6609 1157 6661 1201
rect 6609 1149 6618 1157
rect 6618 1149 6652 1157
rect 6652 1149 6661 1157
rect 6809 1353 6818 1361
rect 6818 1353 6852 1361
rect 6852 1353 6861 1361
rect 6809 1309 6861 1353
rect 7009 1527 7061 1571
rect 7009 1519 7018 1527
rect 7018 1519 7052 1527
rect 7052 1519 7061 1527
rect 7209 1633 7218 1641
rect 7218 1633 7252 1641
rect 7252 1633 7261 1641
rect 7209 1589 7261 1633
rect 7409 1807 7461 1851
rect 7409 1799 7418 1807
rect 7418 1799 7452 1807
rect 7452 1799 7461 1807
rect 7609 1913 7618 1921
rect 7618 1913 7652 1921
rect 7652 1913 7661 1921
rect 7609 1869 7661 1913
rect 7809 2087 7861 2131
rect 7809 2079 7818 2087
rect 7818 2079 7852 2087
rect 7852 2079 7861 2087
rect 8009 2193 8018 2201
rect 8018 2193 8052 2201
rect 8052 2193 8061 2201
rect 8009 2149 8061 2193
rect 8209 2367 8261 2411
rect 8209 2359 8218 2367
rect 8218 2359 8252 2367
rect 8252 2359 8261 2367
rect 8409 2563 8418 2571
rect 8418 2563 8452 2571
rect 8452 2563 8461 2571
rect 8409 2519 8461 2563
rect 8609 2737 8661 2781
rect 8609 2729 8618 2737
rect 8618 2729 8652 2737
rect 8652 2729 8661 2737
rect 8809 2843 8818 2851
rect 8818 2843 8852 2851
rect 8852 2843 8861 2851
rect 8809 2799 8861 2843
rect 9009 3017 9061 3061
rect 9009 3009 9018 3017
rect 9018 3009 9052 3017
rect 9052 3009 9061 3017
rect 9209 3123 9218 3131
rect 9218 3123 9252 3131
rect 9252 3123 9261 3131
rect 9209 3079 9261 3123
rect 9409 3297 9461 3341
rect 9409 3289 9418 3297
rect 9418 3289 9452 3297
rect 9452 3289 9461 3297
rect 9609 3403 9618 3411
rect 9618 3403 9652 3411
rect 9652 3403 9661 3411
rect 9609 3359 9661 3403
rect 9809 3577 9861 3621
rect 9809 3569 9818 3577
rect 9818 3569 9852 3577
rect 9852 3569 9861 3577
rect 10009 3773 10018 3781
rect 10018 3773 10052 3781
rect 10052 3773 10061 3781
rect 10009 3729 10061 3773
rect 10209 3947 10261 3991
rect 10209 3939 10218 3947
rect 10218 3939 10252 3947
rect 10252 3939 10261 3947
rect 10409 4053 10418 4061
rect 10418 4053 10452 4061
rect 10452 4053 10461 4061
rect 10409 4009 10461 4053
rect 10609 4227 10661 4271
rect 10609 4219 10618 4227
rect 10618 4219 10652 4227
rect 10652 4219 10661 4227
rect 10809 4333 10818 4341
rect 10818 4333 10852 4341
rect 10852 4333 10861 4341
rect 10809 4289 10861 4333
rect 11009 4507 11061 4551
rect 11009 4499 11018 4507
rect 11018 4499 11052 4507
rect 11052 4499 11061 4507
rect 11209 4613 11218 4621
rect 11218 4613 11252 4621
rect 11252 4613 11261 4621
rect 11209 4569 11261 4613
rect 11409 4787 11461 4831
rect 11409 4779 11418 4787
rect 11418 4779 11452 4787
rect 11452 4779 11461 4787
rect 11609 4894 11661 4903
rect 11609 4860 11618 4894
rect 11618 4860 11652 4894
rect 11652 4860 11661 4894
rect 11609 4851 11661 4860
rect 10009 3684 10061 3693
rect 10009 3650 10018 3684
rect 10018 3650 10052 3684
rect 10052 3650 10061 3684
rect 10009 3641 10061 3650
rect 8409 2474 8461 2483
rect 8409 2440 8418 2474
rect 8418 2440 8452 2474
rect 8452 2440 8461 2474
rect 8409 2431 8461 2440
rect 6809 1264 6861 1273
rect 6809 1230 6818 1264
rect 6818 1230 6852 1264
rect 6852 1230 6861 1264
rect 6809 1221 6861 1230
rect 5209 54 5261 63
rect 5209 20 5218 54
rect 5218 20 5252 54
rect 5252 20 5261 54
rect 5209 11 5261 20
rect 5109 -60 5161 -15
rect 5109 -67 5118 -60
rect 5118 -67 5152 -60
rect 5152 -67 5161 -60
rect 4909 -166 4918 -143
rect 4918 -166 4952 -143
rect 4952 -166 4961 -143
rect 4909 -195 4961 -166
rect 4925 -248 4977 -239
rect 4925 -282 4934 -248
rect 4934 -282 4968 -248
rect 4968 -282 4977 -248
rect 4925 -291 4977 -282
rect 4909 -363 4961 -326
rect 4909 -378 4918 -363
rect 4918 -378 4952 -363
rect 4952 -378 4961 -363
rect 4909 -397 4918 -390
rect 4918 -397 4952 -390
rect 4952 -397 4961 -390
rect 4909 -435 4961 -397
rect 4909 -442 4918 -435
rect 4918 -442 4952 -435
rect 4952 -442 4961 -435
rect 4909 -469 4918 -454
rect 4918 -469 4952 -454
rect 4952 -469 4961 -454
rect 4909 -506 4961 -469
rect 5109 -94 5118 -79
rect 5118 -94 5152 -79
rect 5152 -94 5161 -79
rect 5109 -131 5161 -94
rect 5209 -74 5261 -22
rect 5409 177 5461 221
rect 5409 169 5418 177
rect 5418 169 5452 177
rect 5452 169 5461 177
rect 5609 283 5618 291
rect 5618 283 5652 291
rect 5652 283 5661 291
rect 5609 239 5661 283
rect 5809 457 5861 501
rect 5809 449 5818 457
rect 5818 449 5852 457
rect 5852 449 5861 457
rect 6009 563 6018 571
rect 6018 563 6052 571
rect 6052 563 6061 571
rect 6009 519 6061 563
rect 6209 737 6261 781
rect 6209 729 6218 737
rect 6218 729 6252 737
rect 6252 729 6261 737
rect 6409 843 6418 851
rect 6418 843 6452 851
rect 6452 843 6461 851
rect 6409 799 6461 843
rect 6609 1017 6661 1061
rect 6609 1009 6618 1017
rect 6618 1009 6652 1017
rect 6652 1009 6661 1017
rect 6809 1123 6818 1131
rect 6818 1123 6852 1131
rect 6852 1123 6861 1131
rect 6809 1079 6861 1123
rect 7009 1387 7061 1431
rect 7009 1379 7018 1387
rect 7018 1379 7052 1387
rect 7052 1379 7061 1387
rect 7209 1493 7218 1501
rect 7218 1493 7252 1501
rect 7252 1493 7261 1501
rect 7209 1449 7261 1493
rect 7409 1667 7461 1711
rect 7409 1659 7418 1667
rect 7418 1659 7452 1667
rect 7452 1659 7461 1667
rect 7609 1773 7618 1781
rect 7618 1773 7652 1781
rect 7652 1773 7661 1781
rect 7609 1729 7661 1773
rect 7809 1947 7861 1991
rect 7809 1939 7818 1947
rect 7818 1939 7852 1947
rect 7852 1939 7861 1947
rect 8009 2053 8018 2061
rect 8018 2053 8052 2061
rect 8052 2053 8061 2061
rect 8009 2009 8061 2053
rect 8209 2227 8261 2271
rect 8209 2219 8218 2227
rect 8218 2219 8252 2227
rect 8252 2219 8261 2227
rect 8409 2333 8418 2341
rect 8418 2333 8452 2341
rect 8452 2333 8461 2341
rect 8409 2289 8461 2333
rect 8609 2597 8661 2641
rect 8609 2589 8618 2597
rect 8618 2589 8652 2597
rect 8652 2589 8661 2597
rect 8809 2703 8818 2711
rect 8818 2703 8852 2711
rect 8852 2703 8861 2711
rect 8809 2659 8861 2703
rect 9009 2877 9061 2921
rect 9009 2869 9018 2877
rect 9018 2869 9052 2877
rect 9052 2869 9061 2877
rect 9209 2983 9218 2991
rect 9218 2983 9252 2991
rect 9252 2983 9261 2991
rect 9209 2939 9261 2983
rect 9409 3157 9461 3201
rect 9409 3149 9418 3157
rect 9418 3149 9452 3157
rect 9452 3149 9461 3157
rect 9609 3263 9618 3271
rect 9618 3263 9652 3271
rect 9652 3263 9661 3271
rect 9609 3219 9661 3263
rect 9809 3437 9861 3481
rect 9809 3429 9818 3437
rect 9818 3429 9852 3437
rect 9852 3429 9861 3437
rect 10009 3543 10018 3551
rect 10018 3543 10052 3551
rect 10052 3543 10061 3551
rect 10009 3499 10061 3543
rect 10209 3807 10261 3851
rect 10209 3799 10218 3807
rect 10218 3799 10252 3807
rect 10252 3799 10261 3807
rect 10409 3913 10418 3921
rect 10418 3913 10452 3921
rect 10452 3913 10461 3921
rect 10409 3869 10461 3913
rect 10609 4087 10661 4131
rect 10609 4079 10618 4087
rect 10618 4079 10652 4087
rect 10652 4079 10661 4087
rect 10809 4193 10818 4201
rect 10818 4193 10852 4201
rect 10852 4193 10861 4201
rect 10809 4149 10861 4193
rect 11009 4367 11061 4411
rect 11009 4359 11018 4367
rect 11018 4359 11052 4367
rect 11052 4359 11061 4367
rect 11209 4473 11218 4481
rect 11218 4473 11252 4481
rect 11252 4473 11261 4481
rect 11209 4429 11261 4473
rect 11409 4647 11461 4691
rect 11409 4639 11418 4647
rect 11418 4639 11452 4647
rect 11452 4639 11461 4647
rect 11609 4753 11618 4761
rect 11618 4753 11652 4761
rect 11652 4753 11661 4761
rect 11609 4709 11661 4753
rect 11809 4910 11861 4919
rect 11809 4876 11818 4910
rect 11818 4876 11852 4910
rect 11852 4876 11861 4910
rect 11809 4867 11861 4876
rect 10209 3700 10261 3709
rect 10209 3666 10218 3700
rect 10218 3666 10252 3700
rect 10252 3666 10261 3700
rect 10209 3657 10261 3666
rect 8609 2490 8661 2499
rect 8609 2456 8618 2490
rect 8618 2456 8652 2490
rect 8652 2456 8661 2490
rect 8609 2447 8661 2456
rect 7009 1280 7061 1289
rect 7009 1246 7018 1280
rect 7018 1246 7052 1280
rect 7052 1246 7061 1280
rect 7009 1237 7061 1246
rect 5409 70 5461 79
rect 5409 36 5418 70
rect 5418 36 5452 70
rect 5452 36 5461 70
rect 5409 27 5461 36
rect 5309 -60 5361 -15
rect 5309 -67 5318 -60
rect 5318 -67 5352 -60
rect 5352 -67 5361 -60
rect 5109 -166 5118 -143
rect 5118 -166 5152 -143
rect 5152 -166 5161 -143
rect 5109 -195 5161 -166
rect 5125 -248 5177 -239
rect 5125 -282 5134 -248
rect 5134 -282 5168 -248
rect 5168 -282 5177 -248
rect 5125 -291 5177 -282
rect 5109 -363 5161 -326
rect 5109 -378 5118 -363
rect 5118 -378 5152 -363
rect 5152 -378 5161 -363
rect 5109 -397 5118 -390
rect 5118 -397 5152 -390
rect 5152 -397 5161 -390
rect 5109 -435 5161 -397
rect 5109 -442 5118 -435
rect 5118 -442 5152 -435
rect 5152 -442 5161 -435
rect 5109 -469 5118 -454
rect 5118 -469 5152 -454
rect 5152 -469 5161 -454
rect 5109 -506 5161 -469
rect 5309 -94 5318 -79
rect 5318 -94 5352 -79
rect 5352 -94 5361 -79
rect 5309 -131 5361 -94
rect 5409 -74 5461 -22
rect 5609 143 5618 151
rect 5618 143 5652 151
rect 5652 143 5661 151
rect 5609 99 5661 143
rect 5809 317 5861 361
rect 5809 309 5818 317
rect 5818 309 5852 317
rect 5852 309 5861 317
rect 6009 423 6018 431
rect 6018 423 6052 431
rect 6052 423 6061 431
rect 6009 379 6061 423
rect 6209 597 6261 641
rect 6209 589 6218 597
rect 6218 589 6252 597
rect 6252 589 6261 597
rect 6409 703 6418 711
rect 6418 703 6452 711
rect 6452 703 6461 711
rect 6409 659 6461 703
rect 6609 877 6661 921
rect 6609 869 6618 877
rect 6618 869 6652 877
rect 6652 869 6661 877
rect 6809 983 6818 991
rect 6818 983 6852 991
rect 6852 983 6861 991
rect 6809 939 6861 983
rect 7009 1157 7061 1201
rect 7009 1149 7018 1157
rect 7018 1149 7052 1157
rect 7052 1149 7061 1157
rect 7209 1353 7218 1361
rect 7218 1353 7252 1361
rect 7252 1353 7261 1361
rect 7209 1309 7261 1353
rect 7409 1527 7461 1571
rect 7409 1519 7418 1527
rect 7418 1519 7452 1527
rect 7452 1519 7461 1527
rect 7609 1633 7618 1641
rect 7618 1633 7652 1641
rect 7652 1633 7661 1641
rect 7609 1589 7661 1633
rect 7809 1807 7861 1851
rect 7809 1799 7818 1807
rect 7818 1799 7852 1807
rect 7852 1799 7861 1807
rect 8009 1913 8018 1921
rect 8018 1913 8052 1921
rect 8052 1913 8061 1921
rect 8009 1869 8061 1913
rect 8209 2087 8261 2131
rect 8209 2079 8218 2087
rect 8218 2079 8252 2087
rect 8252 2079 8261 2087
rect 8409 2193 8418 2201
rect 8418 2193 8452 2201
rect 8452 2193 8461 2201
rect 8409 2149 8461 2193
rect 8609 2367 8661 2411
rect 8609 2359 8618 2367
rect 8618 2359 8652 2367
rect 8652 2359 8661 2367
rect 8809 2563 8818 2571
rect 8818 2563 8852 2571
rect 8852 2563 8861 2571
rect 8809 2519 8861 2563
rect 9009 2737 9061 2781
rect 9009 2729 9018 2737
rect 9018 2729 9052 2737
rect 9052 2729 9061 2737
rect 9209 2843 9218 2851
rect 9218 2843 9252 2851
rect 9252 2843 9261 2851
rect 9209 2799 9261 2843
rect 9409 3017 9461 3061
rect 9409 3009 9418 3017
rect 9418 3009 9452 3017
rect 9452 3009 9461 3017
rect 9609 3123 9618 3131
rect 9618 3123 9652 3131
rect 9652 3123 9661 3131
rect 9609 3079 9661 3123
rect 9809 3297 9861 3341
rect 9809 3289 9818 3297
rect 9818 3289 9852 3297
rect 9852 3289 9861 3297
rect 10009 3403 10018 3411
rect 10018 3403 10052 3411
rect 10052 3403 10061 3411
rect 10009 3359 10061 3403
rect 10209 3577 10261 3621
rect 10209 3569 10218 3577
rect 10218 3569 10252 3577
rect 10252 3569 10261 3577
rect 10409 3773 10418 3781
rect 10418 3773 10452 3781
rect 10452 3773 10461 3781
rect 10409 3729 10461 3773
rect 10609 3947 10661 3991
rect 10609 3939 10618 3947
rect 10618 3939 10652 3947
rect 10652 3939 10661 3947
rect 10809 4053 10818 4061
rect 10818 4053 10852 4061
rect 10852 4053 10861 4061
rect 10809 4009 10861 4053
rect 11009 4227 11061 4271
rect 11009 4219 11018 4227
rect 11018 4219 11052 4227
rect 11052 4219 11061 4227
rect 11209 4333 11218 4341
rect 11218 4333 11252 4341
rect 11252 4333 11261 4341
rect 11209 4289 11261 4333
rect 11409 4507 11461 4551
rect 11409 4499 11418 4507
rect 11418 4499 11452 4507
rect 11452 4499 11461 4507
rect 11609 4613 11618 4621
rect 11618 4613 11652 4621
rect 11652 4613 11661 4621
rect 11609 4569 11661 4613
rect 11809 4787 11861 4831
rect 11809 4779 11818 4787
rect 11818 4779 11852 4787
rect 11852 4779 11861 4787
rect 12009 4894 12061 4903
rect 12009 4860 12018 4894
rect 12018 4860 12052 4894
rect 12052 4860 12061 4894
rect 12009 4851 12061 4860
rect 10409 3684 10461 3693
rect 10409 3650 10418 3684
rect 10418 3650 10452 3684
rect 10452 3650 10461 3684
rect 10409 3641 10461 3650
rect 8809 2474 8861 2483
rect 8809 2440 8818 2474
rect 8818 2440 8852 2474
rect 8852 2440 8861 2474
rect 8809 2431 8861 2440
rect 7209 1264 7261 1273
rect 7209 1230 7218 1264
rect 7218 1230 7252 1264
rect 7252 1230 7261 1264
rect 7209 1221 7261 1230
rect 5609 54 5661 63
rect 5609 20 5618 54
rect 5618 20 5652 54
rect 5652 20 5661 54
rect 5609 11 5661 20
rect 5509 -60 5561 -15
rect 5509 -67 5518 -60
rect 5518 -67 5552 -60
rect 5552 -67 5561 -60
rect 5309 -166 5318 -143
rect 5318 -166 5352 -143
rect 5352 -166 5361 -143
rect 5309 -195 5361 -166
rect 5325 -248 5377 -239
rect 5325 -282 5334 -248
rect 5334 -282 5368 -248
rect 5368 -282 5377 -248
rect 5325 -291 5377 -282
rect 5309 -363 5361 -326
rect 5309 -378 5318 -363
rect 5318 -378 5352 -363
rect 5352 -378 5361 -363
rect 5309 -397 5318 -390
rect 5318 -397 5352 -390
rect 5352 -397 5361 -390
rect 5309 -435 5361 -397
rect 5309 -442 5318 -435
rect 5318 -442 5352 -435
rect 5352 -442 5361 -435
rect 5309 -469 5318 -454
rect 5318 -469 5352 -454
rect 5352 -469 5361 -454
rect 5309 -506 5361 -469
rect 5509 -94 5518 -79
rect 5518 -94 5552 -79
rect 5552 -94 5561 -79
rect 5509 -131 5561 -94
rect 5609 -74 5661 -22
rect 5809 177 5861 221
rect 5809 169 5818 177
rect 5818 169 5852 177
rect 5852 169 5861 177
rect 6009 283 6018 291
rect 6018 283 6052 291
rect 6052 283 6061 291
rect 6009 239 6061 283
rect 6209 457 6261 501
rect 6209 449 6218 457
rect 6218 449 6252 457
rect 6252 449 6261 457
rect 6409 563 6418 571
rect 6418 563 6452 571
rect 6452 563 6461 571
rect 6409 519 6461 563
rect 6609 737 6661 781
rect 6609 729 6618 737
rect 6618 729 6652 737
rect 6652 729 6661 737
rect 6809 843 6818 851
rect 6818 843 6852 851
rect 6852 843 6861 851
rect 6809 799 6861 843
rect 7009 1017 7061 1061
rect 7009 1009 7018 1017
rect 7018 1009 7052 1017
rect 7052 1009 7061 1017
rect 7209 1123 7218 1131
rect 7218 1123 7252 1131
rect 7252 1123 7261 1131
rect 7209 1079 7261 1123
rect 7409 1387 7461 1431
rect 7409 1379 7418 1387
rect 7418 1379 7452 1387
rect 7452 1379 7461 1387
rect 7609 1493 7618 1501
rect 7618 1493 7652 1501
rect 7652 1493 7661 1501
rect 7609 1449 7661 1493
rect 7809 1667 7861 1711
rect 7809 1659 7818 1667
rect 7818 1659 7852 1667
rect 7852 1659 7861 1667
rect 8009 1773 8018 1781
rect 8018 1773 8052 1781
rect 8052 1773 8061 1781
rect 8009 1729 8061 1773
rect 8209 1947 8261 1991
rect 8209 1939 8218 1947
rect 8218 1939 8252 1947
rect 8252 1939 8261 1947
rect 8409 2053 8418 2061
rect 8418 2053 8452 2061
rect 8452 2053 8461 2061
rect 8409 2009 8461 2053
rect 8609 2227 8661 2271
rect 8609 2219 8618 2227
rect 8618 2219 8652 2227
rect 8652 2219 8661 2227
rect 8809 2333 8818 2341
rect 8818 2333 8852 2341
rect 8852 2333 8861 2341
rect 8809 2289 8861 2333
rect 9009 2597 9061 2641
rect 9009 2589 9018 2597
rect 9018 2589 9052 2597
rect 9052 2589 9061 2597
rect 9209 2703 9218 2711
rect 9218 2703 9252 2711
rect 9252 2703 9261 2711
rect 9209 2659 9261 2703
rect 9409 2877 9461 2921
rect 9409 2869 9418 2877
rect 9418 2869 9452 2877
rect 9452 2869 9461 2877
rect 9609 2983 9618 2991
rect 9618 2983 9652 2991
rect 9652 2983 9661 2991
rect 9609 2939 9661 2983
rect 9809 3157 9861 3201
rect 9809 3149 9818 3157
rect 9818 3149 9852 3157
rect 9852 3149 9861 3157
rect 10009 3263 10018 3271
rect 10018 3263 10052 3271
rect 10052 3263 10061 3271
rect 10009 3219 10061 3263
rect 10209 3437 10261 3481
rect 10209 3429 10218 3437
rect 10218 3429 10252 3437
rect 10252 3429 10261 3437
rect 10409 3543 10418 3551
rect 10418 3543 10452 3551
rect 10452 3543 10461 3551
rect 10409 3499 10461 3543
rect 10609 3807 10661 3851
rect 10609 3799 10618 3807
rect 10618 3799 10652 3807
rect 10652 3799 10661 3807
rect 10809 3913 10818 3921
rect 10818 3913 10852 3921
rect 10852 3913 10861 3921
rect 10809 3869 10861 3913
rect 11009 4087 11061 4131
rect 11009 4079 11018 4087
rect 11018 4079 11052 4087
rect 11052 4079 11061 4087
rect 11209 4193 11218 4201
rect 11218 4193 11252 4201
rect 11252 4193 11261 4201
rect 11209 4149 11261 4193
rect 11409 4367 11461 4411
rect 11409 4359 11418 4367
rect 11418 4359 11452 4367
rect 11452 4359 11461 4367
rect 11609 4473 11618 4481
rect 11618 4473 11652 4481
rect 11652 4473 11661 4481
rect 11609 4429 11661 4473
rect 11809 4647 11861 4691
rect 11809 4639 11818 4647
rect 11818 4639 11852 4647
rect 11852 4639 11861 4647
rect 12009 4753 12018 4761
rect 12018 4753 12052 4761
rect 12052 4753 12061 4761
rect 12009 4709 12061 4753
rect 12209 4910 12261 4919
rect 12209 4876 12218 4910
rect 12218 4876 12252 4910
rect 12252 4876 12261 4910
rect 12209 4867 12261 4876
rect 10609 3700 10661 3709
rect 10609 3666 10618 3700
rect 10618 3666 10652 3700
rect 10652 3666 10661 3700
rect 10609 3657 10661 3666
rect 9009 2490 9061 2499
rect 9009 2456 9018 2490
rect 9018 2456 9052 2490
rect 9052 2456 9061 2490
rect 9009 2447 9061 2456
rect 7409 1280 7461 1289
rect 7409 1246 7418 1280
rect 7418 1246 7452 1280
rect 7452 1246 7461 1280
rect 7409 1237 7461 1246
rect 5809 70 5861 79
rect 5809 36 5818 70
rect 5818 36 5852 70
rect 5852 36 5861 70
rect 5809 27 5861 36
rect 5709 -60 5761 -15
rect 5709 -67 5718 -60
rect 5718 -67 5752 -60
rect 5752 -67 5761 -60
rect 5509 -166 5518 -143
rect 5518 -166 5552 -143
rect 5552 -166 5561 -143
rect 5509 -195 5561 -166
rect 5525 -248 5577 -239
rect 5525 -282 5534 -248
rect 5534 -282 5568 -248
rect 5568 -282 5577 -248
rect 5525 -291 5577 -282
rect 5509 -363 5561 -326
rect 5509 -378 5518 -363
rect 5518 -378 5552 -363
rect 5552 -378 5561 -363
rect 5509 -397 5518 -390
rect 5518 -397 5552 -390
rect 5552 -397 5561 -390
rect 5509 -435 5561 -397
rect 5509 -442 5518 -435
rect 5518 -442 5552 -435
rect 5552 -442 5561 -435
rect 5509 -469 5518 -454
rect 5518 -469 5552 -454
rect 5552 -469 5561 -454
rect 5509 -506 5561 -469
rect 5709 -94 5718 -79
rect 5718 -94 5752 -79
rect 5752 -94 5761 -79
rect 5709 -131 5761 -94
rect 5809 -74 5861 -22
rect 6009 143 6018 151
rect 6018 143 6052 151
rect 6052 143 6061 151
rect 6009 99 6061 143
rect 6209 317 6261 361
rect 6209 309 6218 317
rect 6218 309 6252 317
rect 6252 309 6261 317
rect 6409 423 6418 431
rect 6418 423 6452 431
rect 6452 423 6461 431
rect 6409 379 6461 423
rect 6609 597 6661 641
rect 6609 589 6618 597
rect 6618 589 6652 597
rect 6652 589 6661 597
rect 6809 703 6818 711
rect 6818 703 6852 711
rect 6852 703 6861 711
rect 6809 659 6861 703
rect 7009 877 7061 921
rect 7009 869 7018 877
rect 7018 869 7052 877
rect 7052 869 7061 877
rect 7209 983 7218 991
rect 7218 983 7252 991
rect 7252 983 7261 991
rect 7209 939 7261 983
rect 7409 1157 7461 1201
rect 7409 1149 7418 1157
rect 7418 1149 7452 1157
rect 7452 1149 7461 1157
rect 7609 1353 7618 1361
rect 7618 1353 7652 1361
rect 7652 1353 7661 1361
rect 7609 1309 7661 1353
rect 7809 1527 7861 1571
rect 7809 1519 7818 1527
rect 7818 1519 7852 1527
rect 7852 1519 7861 1527
rect 8009 1633 8018 1641
rect 8018 1633 8052 1641
rect 8052 1633 8061 1641
rect 8009 1589 8061 1633
rect 8209 1807 8261 1851
rect 8209 1799 8218 1807
rect 8218 1799 8252 1807
rect 8252 1799 8261 1807
rect 8409 1913 8418 1921
rect 8418 1913 8452 1921
rect 8452 1913 8461 1921
rect 8409 1869 8461 1913
rect 8609 2087 8661 2131
rect 8609 2079 8618 2087
rect 8618 2079 8652 2087
rect 8652 2079 8661 2087
rect 8809 2193 8818 2201
rect 8818 2193 8852 2201
rect 8852 2193 8861 2201
rect 8809 2149 8861 2193
rect 9009 2367 9061 2411
rect 9009 2359 9018 2367
rect 9018 2359 9052 2367
rect 9052 2359 9061 2367
rect 9209 2563 9218 2571
rect 9218 2563 9252 2571
rect 9252 2563 9261 2571
rect 9209 2519 9261 2563
rect 9409 2737 9461 2781
rect 9409 2729 9418 2737
rect 9418 2729 9452 2737
rect 9452 2729 9461 2737
rect 9609 2843 9618 2851
rect 9618 2843 9652 2851
rect 9652 2843 9661 2851
rect 9609 2799 9661 2843
rect 9809 3017 9861 3061
rect 9809 3009 9818 3017
rect 9818 3009 9852 3017
rect 9852 3009 9861 3017
rect 10009 3123 10018 3131
rect 10018 3123 10052 3131
rect 10052 3123 10061 3131
rect 10009 3079 10061 3123
rect 10209 3297 10261 3341
rect 10209 3289 10218 3297
rect 10218 3289 10252 3297
rect 10252 3289 10261 3297
rect 10409 3403 10418 3411
rect 10418 3403 10452 3411
rect 10452 3403 10461 3411
rect 10409 3359 10461 3403
rect 10609 3577 10661 3621
rect 10609 3569 10618 3577
rect 10618 3569 10652 3577
rect 10652 3569 10661 3577
rect 10809 3773 10818 3781
rect 10818 3773 10852 3781
rect 10852 3773 10861 3781
rect 10809 3729 10861 3773
rect 11009 3947 11061 3991
rect 11009 3939 11018 3947
rect 11018 3939 11052 3947
rect 11052 3939 11061 3947
rect 11209 4053 11218 4061
rect 11218 4053 11252 4061
rect 11252 4053 11261 4061
rect 11209 4009 11261 4053
rect 11409 4227 11461 4271
rect 11409 4219 11418 4227
rect 11418 4219 11452 4227
rect 11452 4219 11461 4227
rect 11609 4333 11618 4341
rect 11618 4333 11652 4341
rect 11652 4333 11661 4341
rect 11609 4289 11661 4333
rect 11809 4507 11861 4551
rect 11809 4499 11818 4507
rect 11818 4499 11852 4507
rect 11852 4499 11861 4507
rect 12009 4613 12018 4621
rect 12018 4613 12052 4621
rect 12052 4613 12061 4621
rect 12009 4569 12061 4613
rect 12209 4787 12261 4831
rect 12209 4779 12218 4787
rect 12218 4779 12252 4787
rect 12252 4779 12261 4787
rect 12409 4894 12461 4903
rect 12409 4860 12418 4894
rect 12418 4860 12452 4894
rect 12452 4860 12461 4894
rect 12409 4851 12461 4860
rect 10809 3684 10861 3693
rect 10809 3650 10818 3684
rect 10818 3650 10852 3684
rect 10852 3650 10861 3684
rect 10809 3641 10861 3650
rect 9209 2474 9261 2483
rect 9209 2440 9218 2474
rect 9218 2440 9252 2474
rect 9252 2440 9261 2474
rect 9209 2431 9261 2440
rect 7609 1264 7661 1273
rect 7609 1230 7618 1264
rect 7618 1230 7652 1264
rect 7652 1230 7661 1264
rect 7609 1221 7661 1230
rect 6009 54 6061 63
rect 6009 20 6018 54
rect 6018 20 6052 54
rect 6052 20 6061 54
rect 6009 11 6061 20
rect 5909 -60 5961 -15
rect 5909 -67 5918 -60
rect 5918 -67 5952 -60
rect 5952 -67 5961 -60
rect 5709 -166 5718 -143
rect 5718 -166 5752 -143
rect 5752 -166 5761 -143
rect 5709 -195 5761 -166
rect 5725 -248 5777 -239
rect 5725 -282 5734 -248
rect 5734 -282 5768 -248
rect 5768 -282 5777 -248
rect 5725 -291 5777 -282
rect 5709 -363 5761 -326
rect 5709 -378 5718 -363
rect 5718 -378 5752 -363
rect 5752 -378 5761 -363
rect 5709 -397 5718 -390
rect 5718 -397 5752 -390
rect 5752 -397 5761 -390
rect 5709 -435 5761 -397
rect 5709 -442 5718 -435
rect 5718 -442 5752 -435
rect 5752 -442 5761 -435
rect 5709 -469 5718 -454
rect 5718 -469 5752 -454
rect 5752 -469 5761 -454
rect 5709 -506 5761 -469
rect 5909 -94 5918 -79
rect 5918 -94 5952 -79
rect 5952 -94 5961 -79
rect 5909 -131 5961 -94
rect 6009 -74 6061 -22
rect 6209 177 6261 221
rect 6209 169 6218 177
rect 6218 169 6252 177
rect 6252 169 6261 177
rect 6409 283 6418 291
rect 6418 283 6452 291
rect 6452 283 6461 291
rect 6409 239 6461 283
rect 6609 457 6661 501
rect 6609 449 6618 457
rect 6618 449 6652 457
rect 6652 449 6661 457
rect 6809 563 6818 571
rect 6818 563 6852 571
rect 6852 563 6861 571
rect 6809 519 6861 563
rect 7009 737 7061 781
rect 7009 729 7018 737
rect 7018 729 7052 737
rect 7052 729 7061 737
rect 7209 843 7218 851
rect 7218 843 7252 851
rect 7252 843 7261 851
rect 7209 799 7261 843
rect 7409 1017 7461 1061
rect 7409 1009 7418 1017
rect 7418 1009 7452 1017
rect 7452 1009 7461 1017
rect 7609 1123 7618 1131
rect 7618 1123 7652 1131
rect 7652 1123 7661 1131
rect 7609 1079 7661 1123
rect 7809 1387 7861 1431
rect 7809 1379 7818 1387
rect 7818 1379 7852 1387
rect 7852 1379 7861 1387
rect 8009 1493 8018 1501
rect 8018 1493 8052 1501
rect 8052 1493 8061 1501
rect 8009 1449 8061 1493
rect 8209 1667 8261 1711
rect 8209 1659 8218 1667
rect 8218 1659 8252 1667
rect 8252 1659 8261 1667
rect 8409 1773 8418 1781
rect 8418 1773 8452 1781
rect 8452 1773 8461 1781
rect 8409 1729 8461 1773
rect 8609 1947 8661 1991
rect 8609 1939 8618 1947
rect 8618 1939 8652 1947
rect 8652 1939 8661 1947
rect 8809 2053 8818 2061
rect 8818 2053 8852 2061
rect 8852 2053 8861 2061
rect 8809 2009 8861 2053
rect 9009 2227 9061 2271
rect 9009 2219 9018 2227
rect 9018 2219 9052 2227
rect 9052 2219 9061 2227
rect 9209 2333 9218 2341
rect 9218 2333 9252 2341
rect 9252 2333 9261 2341
rect 9209 2289 9261 2333
rect 9409 2597 9461 2641
rect 9409 2589 9418 2597
rect 9418 2589 9452 2597
rect 9452 2589 9461 2597
rect 9609 2703 9618 2711
rect 9618 2703 9652 2711
rect 9652 2703 9661 2711
rect 9609 2659 9661 2703
rect 9809 2877 9861 2921
rect 9809 2869 9818 2877
rect 9818 2869 9852 2877
rect 9852 2869 9861 2877
rect 10009 2983 10018 2991
rect 10018 2983 10052 2991
rect 10052 2983 10061 2991
rect 10009 2939 10061 2983
rect 10209 3157 10261 3201
rect 10209 3149 10218 3157
rect 10218 3149 10252 3157
rect 10252 3149 10261 3157
rect 10409 3263 10418 3271
rect 10418 3263 10452 3271
rect 10452 3263 10461 3271
rect 10409 3219 10461 3263
rect 10609 3437 10661 3481
rect 10609 3429 10618 3437
rect 10618 3429 10652 3437
rect 10652 3429 10661 3437
rect 10809 3543 10818 3551
rect 10818 3543 10852 3551
rect 10852 3543 10861 3551
rect 10809 3499 10861 3543
rect 11009 3807 11061 3851
rect 11009 3799 11018 3807
rect 11018 3799 11052 3807
rect 11052 3799 11061 3807
rect 11209 3913 11218 3921
rect 11218 3913 11252 3921
rect 11252 3913 11261 3921
rect 11209 3869 11261 3913
rect 11409 4087 11461 4131
rect 11409 4079 11418 4087
rect 11418 4079 11452 4087
rect 11452 4079 11461 4087
rect 11609 4193 11618 4201
rect 11618 4193 11652 4201
rect 11652 4193 11661 4201
rect 11609 4149 11661 4193
rect 11809 4367 11861 4411
rect 11809 4359 11818 4367
rect 11818 4359 11852 4367
rect 11852 4359 11861 4367
rect 12009 4473 12018 4481
rect 12018 4473 12052 4481
rect 12052 4473 12061 4481
rect 12009 4429 12061 4473
rect 12209 4647 12261 4691
rect 12209 4639 12218 4647
rect 12218 4639 12252 4647
rect 12252 4639 12261 4647
rect 12409 4753 12418 4761
rect 12418 4753 12452 4761
rect 12452 4753 12461 4761
rect 12409 4709 12461 4753
rect 12609 4910 12661 4919
rect 12609 4876 12618 4910
rect 12618 4876 12652 4910
rect 12652 4876 12661 4910
rect 12609 4867 12661 4876
rect 11009 3700 11061 3709
rect 11009 3666 11018 3700
rect 11018 3666 11052 3700
rect 11052 3666 11061 3700
rect 11009 3657 11061 3666
rect 9409 2490 9461 2499
rect 9409 2456 9418 2490
rect 9418 2456 9452 2490
rect 9452 2456 9461 2490
rect 9409 2447 9461 2456
rect 7809 1280 7861 1289
rect 7809 1246 7818 1280
rect 7818 1246 7852 1280
rect 7852 1246 7861 1280
rect 7809 1237 7861 1246
rect 6209 70 6261 79
rect 6209 36 6218 70
rect 6218 36 6252 70
rect 6252 36 6261 70
rect 6209 27 6261 36
rect 6109 -60 6161 -15
rect 6109 -67 6118 -60
rect 6118 -67 6152 -60
rect 6152 -67 6161 -60
rect 5909 -166 5918 -143
rect 5918 -166 5952 -143
rect 5952 -166 5961 -143
rect 5909 -195 5961 -166
rect 5925 -248 5977 -239
rect 5925 -282 5934 -248
rect 5934 -282 5968 -248
rect 5968 -282 5977 -248
rect 5925 -291 5977 -282
rect 5909 -363 5961 -326
rect 5909 -378 5918 -363
rect 5918 -378 5952 -363
rect 5952 -378 5961 -363
rect 5909 -397 5918 -390
rect 5918 -397 5952 -390
rect 5952 -397 5961 -390
rect 5909 -435 5961 -397
rect 5909 -442 5918 -435
rect 5918 -442 5952 -435
rect 5952 -442 5961 -435
rect 5909 -469 5918 -454
rect 5918 -469 5952 -454
rect 5952 -469 5961 -454
rect 5909 -506 5961 -469
rect 6109 -94 6118 -79
rect 6118 -94 6152 -79
rect 6152 -94 6161 -79
rect 6109 -131 6161 -94
rect 6209 -74 6261 -22
rect 6409 143 6418 151
rect 6418 143 6452 151
rect 6452 143 6461 151
rect 6409 99 6461 143
rect 6609 317 6661 361
rect 6609 309 6618 317
rect 6618 309 6652 317
rect 6652 309 6661 317
rect 6809 423 6818 431
rect 6818 423 6852 431
rect 6852 423 6861 431
rect 6809 379 6861 423
rect 7009 597 7061 641
rect 7009 589 7018 597
rect 7018 589 7052 597
rect 7052 589 7061 597
rect 7209 703 7218 711
rect 7218 703 7252 711
rect 7252 703 7261 711
rect 7209 659 7261 703
rect 7409 877 7461 921
rect 7409 869 7418 877
rect 7418 869 7452 877
rect 7452 869 7461 877
rect 7609 983 7618 991
rect 7618 983 7652 991
rect 7652 983 7661 991
rect 7609 939 7661 983
rect 7809 1157 7861 1201
rect 7809 1149 7818 1157
rect 7818 1149 7852 1157
rect 7852 1149 7861 1157
rect 8009 1353 8018 1361
rect 8018 1353 8052 1361
rect 8052 1353 8061 1361
rect 8009 1309 8061 1353
rect 8209 1527 8261 1571
rect 8209 1519 8218 1527
rect 8218 1519 8252 1527
rect 8252 1519 8261 1527
rect 8409 1633 8418 1641
rect 8418 1633 8452 1641
rect 8452 1633 8461 1641
rect 8409 1589 8461 1633
rect 8609 1807 8661 1851
rect 8609 1799 8618 1807
rect 8618 1799 8652 1807
rect 8652 1799 8661 1807
rect 8809 1913 8818 1921
rect 8818 1913 8852 1921
rect 8852 1913 8861 1921
rect 8809 1869 8861 1913
rect 9009 2087 9061 2131
rect 9009 2079 9018 2087
rect 9018 2079 9052 2087
rect 9052 2079 9061 2087
rect 9209 2193 9218 2201
rect 9218 2193 9252 2201
rect 9252 2193 9261 2201
rect 9209 2149 9261 2193
rect 9409 2367 9461 2411
rect 9409 2359 9418 2367
rect 9418 2359 9452 2367
rect 9452 2359 9461 2367
rect 9609 2563 9618 2571
rect 9618 2563 9652 2571
rect 9652 2563 9661 2571
rect 9609 2519 9661 2563
rect 9809 2737 9861 2781
rect 9809 2729 9818 2737
rect 9818 2729 9852 2737
rect 9852 2729 9861 2737
rect 10009 2843 10018 2851
rect 10018 2843 10052 2851
rect 10052 2843 10061 2851
rect 10009 2799 10061 2843
rect 10209 3017 10261 3061
rect 10209 3009 10218 3017
rect 10218 3009 10252 3017
rect 10252 3009 10261 3017
rect 10409 3123 10418 3131
rect 10418 3123 10452 3131
rect 10452 3123 10461 3131
rect 10409 3079 10461 3123
rect 10609 3297 10661 3341
rect 10609 3289 10618 3297
rect 10618 3289 10652 3297
rect 10652 3289 10661 3297
rect 10809 3403 10818 3411
rect 10818 3403 10852 3411
rect 10852 3403 10861 3411
rect 10809 3359 10861 3403
rect 11009 3577 11061 3621
rect 11009 3569 11018 3577
rect 11018 3569 11052 3577
rect 11052 3569 11061 3577
rect 11209 3773 11218 3781
rect 11218 3773 11252 3781
rect 11252 3773 11261 3781
rect 11209 3729 11261 3773
rect 11409 3947 11461 3991
rect 11409 3939 11418 3947
rect 11418 3939 11452 3947
rect 11452 3939 11461 3947
rect 11609 4053 11618 4061
rect 11618 4053 11652 4061
rect 11652 4053 11661 4061
rect 11609 4009 11661 4053
rect 11809 4227 11861 4271
rect 11809 4219 11818 4227
rect 11818 4219 11852 4227
rect 11852 4219 11861 4227
rect 12009 4333 12018 4341
rect 12018 4333 12052 4341
rect 12052 4333 12061 4341
rect 12009 4289 12061 4333
rect 12209 4507 12261 4551
rect 12209 4499 12218 4507
rect 12218 4499 12252 4507
rect 12252 4499 12261 4507
rect 12409 4613 12418 4621
rect 12418 4613 12452 4621
rect 12452 4613 12461 4621
rect 12409 4569 12461 4613
rect 12609 4787 12661 4831
rect 12609 4779 12618 4787
rect 12618 4779 12652 4787
rect 12652 4779 12661 4787
rect 11209 3684 11261 3693
rect 11209 3650 11218 3684
rect 11218 3650 11252 3684
rect 11252 3650 11261 3684
rect 11209 3641 11261 3650
rect 9609 2474 9661 2483
rect 9609 2440 9618 2474
rect 9618 2440 9652 2474
rect 9652 2440 9661 2474
rect 9609 2431 9661 2440
rect 8009 1264 8061 1273
rect 8009 1230 8018 1264
rect 8018 1230 8052 1264
rect 8052 1230 8061 1264
rect 8009 1221 8061 1230
rect 6409 54 6461 63
rect 6409 20 6418 54
rect 6418 20 6452 54
rect 6452 20 6461 54
rect 6409 11 6461 20
rect 6309 -60 6361 -15
rect 6309 -67 6318 -60
rect 6318 -67 6352 -60
rect 6352 -67 6361 -60
rect 6109 -166 6118 -143
rect 6118 -166 6152 -143
rect 6152 -166 6161 -143
rect 6109 -195 6161 -166
rect 6125 -248 6177 -239
rect 6125 -282 6134 -248
rect 6134 -282 6168 -248
rect 6168 -282 6177 -248
rect 6125 -291 6177 -282
rect 6109 -363 6161 -326
rect 6109 -378 6118 -363
rect 6118 -378 6152 -363
rect 6152 -378 6161 -363
rect 6109 -397 6118 -390
rect 6118 -397 6152 -390
rect 6152 -397 6161 -390
rect 6109 -435 6161 -397
rect 6109 -442 6118 -435
rect 6118 -442 6152 -435
rect 6152 -442 6161 -435
rect 6109 -469 6118 -454
rect 6118 -469 6152 -454
rect 6152 -469 6161 -454
rect 6109 -506 6161 -469
rect 6309 -94 6318 -79
rect 6318 -94 6352 -79
rect 6352 -94 6361 -79
rect 6309 -131 6361 -94
rect 6409 -74 6461 -22
rect 6609 177 6661 221
rect 6609 169 6618 177
rect 6618 169 6652 177
rect 6652 169 6661 177
rect 6809 283 6818 291
rect 6818 283 6852 291
rect 6852 283 6861 291
rect 6809 239 6861 283
rect 7009 457 7061 501
rect 7009 449 7018 457
rect 7018 449 7052 457
rect 7052 449 7061 457
rect 7209 563 7218 571
rect 7218 563 7252 571
rect 7252 563 7261 571
rect 7209 519 7261 563
rect 7409 737 7461 781
rect 7409 729 7418 737
rect 7418 729 7452 737
rect 7452 729 7461 737
rect 7609 843 7618 851
rect 7618 843 7652 851
rect 7652 843 7661 851
rect 7609 799 7661 843
rect 7809 1017 7861 1061
rect 7809 1009 7818 1017
rect 7818 1009 7852 1017
rect 7852 1009 7861 1017
rect 8009 1123 8018 1131
rect 8018 1123 8052 1131
rect 8052 1123 8061 1131
rect 8009 1079 8061 1123
rect 8209 1387 8261 1431
rect 8209 1379 8218 1387
rect 8218 1379 8252 1387
rect 8252 1379 8261 1387
rect 8409 1493 8418 1501
rect 8418 1493 8452 1501
rect 8452 1493 8461 1501
rect 8409 1449 8461 1493
rect 8609 1667 8661 1711
rect 8609 1659 8618 1667
rect 8618 1659 8652 1667
rect 8652 1659 8661 1667
rect 8809 1773 8818 1781
rect 8818 1773 8852 1781
rect 8852 1773 8861 1781
rect 8809 1729 8861 1773
rect 9009 1947 9061 1991
rect 9009 1939 9018 1947
rect 9018 1939 9052 1947
rect 9052 1939 9061 1947
rect 9209 2053 9218 2061
rect 9218 2053 9252 2061
rect 9252 2053 9261 2061
rect 9209 2009 9261 2053
rect 9409 2227 9461 2271
rect 9409 2219 9418 2227
rect 9418 2219 9452 2227
rect 9452 2219 9461 2227
rect 9609 2333 9618 2341
rect 9618 2333 9652 2341
rect 9652 2333 9661 2341
rect 9609 2289 9661 2333
rect 9809 2597 9861 2641
rect 9809 2589 9818 2597
rect 9818 2589 9852 2597
rect 9852 2589 9861 2597
rect 10009 2703 10018 2711
rect 10018 2703 10052 2711
rect 10052 2703 10061 2711
rect 10009 2659 10061 2703
rect 10209 2877 10261 2921
rect 10209 2869 10218 2877
rect 10218 2869 10252 2877
rect 10252 2869 10261 2877
rect 10409 2983 10418 2991
rect 10418 2983 10452 2991
rect 10452 2983 10461 2991
rect 10409 2939 10461 2983
rect 10609 3157 10661 3201
rect 10609 3149 10618 3157
rect 10618 3149 10652 3157
rect 10652 3149 10661 3157
rect 10809 3263 10818 3271
rect 10818 3263 10852 3271
rect 10852 3263 10861 3271
rect 10809 3219 10861 3263
rect 11009 3437 11061 3481
rect 11009 3429 11018 3437
rect 11018 3429 11052 3437
rect 11052 3429 11061 3437
rect 11209 3543 11218 3551
rect 11218 3543 11252 3551
rect 11252 3543 11261 3551
rect 11209 3499 11261 3543
rect 11409 3807 11461 3851
rect 11409 3799 11418 3807
rect 11418 3799 11452 3807
rect 11452 3799 11461 3807
rect 11609 3913 11618 3921
rect 11618 3913 11652 3921
rect 11652 3913 11661 3921
rect 11609 3869 11661 3913
rect 11809 4087 11861 4131
rect 11809 4079 11818 4087
rect 11818 4079 11852 4087
rect 11852 4079 11861 4087
rect 12009 4193 12018 4201
rect 12018 4193 12052 4201
rect 12052 4193 12061 4201
rect 12009 4149 12061 4193
rect 12209 4367 12261 4411
rect 12209 4359 12218 4367
rect 12218 4359 12252 4367
rect 12252 4359 12261 4367
rect 12409 4473 12418 4481
rect 12418 4473 12452 4481
rect 12452 4473 12461 4481
rect 12409 4429 12461 4473
rect 12609 4647 12661 4691
rect 12609 4639 12618 4647
rect 12618 4639 12652 4647
rect 12652 4639 12661 4647
rect 12809 4753 12818 4761
rect 12818 4753 12852 4761
rect 12852 4753 12861 4761
rect 12809 4709 12861 4753
rect 12907 4709 12959 4761
rect 11409 3700 11461 3709
rect 11409 3666 11418 3700
rect 11418 3666 11452 3700
rect 11452 3666 11461 3700
rect 11409 3657 11461 3666
rect 9809 2490 9861 2499
rect 9809 2456 9818 2490
rect 9818 2456 9852 2490
rect 9852 2456 9861 2490
rect 9809 2447 9861 2456
rect 8209 1280 8261 1289
rect 8209 1246 8218 1280
rect 8218 1246 8252 1280
rect 8252 1246 8261 1280
rect 8209 1237 8261 1246
rect 6609 70 6661 79
rect 6609 36 6618 70
rect 6618 36 6652 70
rect 6652 36 6661 70
rect 6609 27 6661 36
rect 6509 -60 6561 -15
rect 6509 -67 6518 -60
rect 6518 -67 6552 -60
rect 6552 -67 6561 -60
rect 6309 -166 6318 -143
rect 6318 -166 6352 -143
rect 6352 -166 6361 -143
rect 6309 -195 6361 -166
rect 6325 -248 6377 -239
rect 6325 -282 6334 -248
rect 6334 -282 6368 -248
rect 6368 -282 6377 -248
rect 6325 -291 6377 -282
rect 6309 -363 6361 -326
rect 6309 -378 6318 -363
rect 6318 -378 6352 -363
rect 6352 -378 6361 -363
rect 6309 -397 6318 -390
rect 6318 -397 6352 -390
rect 6352 -397 6361 -390
rect 6309 -435 6361 -397
rect 6309 -442 6318 -435
rect 6318 -442 6352 -435
rect 6352 -442 6361 -435
rect 6309 -469 6318 -454
rect 6318 -469 6352 -454
rect 6352 -469 6361 -454
rect 6309 -506 6361 -469
rect 6509 -94 6518 -79
rect 6518 -94 6552 -79
rect 6552 -94 6561 -79
rect 6509 -131 6561 -94
rect 6609 -74 6661 -22
rect 6809 143 6818 151
rect 6818 143 6852 151
rect 6852 143 6861 151
rect 6809 99 6861 143
rect 7009 317 7061 361
rect 7009 309 7018 317
rect 7018 309 7052 317
rect 7052 309 7061 317
rect 7209 423 7218 431
rect 7218 423 7252 431
rect 7252 423 7261 431
rect 7209 379 7261 423
rect 7409 597 7461 641
rect 7409 589 7418 597
rect 7418 589 7452 597
rect 7452 589 7461 597
rect 7609 703 7618 711
rect 7618 703 7652 711
rect 7652 703 7661 711
rect 7609 659 7661 703
rect 7809 877 7861 921
rect 7809 869 7818 877
rect 7818 869 7852 877
rect 7852 869 7861 877
rect 8009 983 8018 991
rect 8018 983 8052 991
rect 8052 983 8061 991
rect 8009 939 8061 983
rect 8209 1157 8261 1201
rect 8209 1149 8218 1157
rect 8218 1149 8252 1157
rect 8252 1149 8261 1157
rect 8409 1353 8418 1361
rect 8418 1353 8452 1361
rect 8452 1353 8461 1361
rect 8409 1309 8461 1353
rect 8609 1527 8661 1571
rect 8609 1519 8618 1527
rect 8618 1519 8652 1527
rect 8652 1519 8661 1527
rect 8809 1633 8818 1641
rect 8818 1633 8852 1641
rect 8852 1633 8861 1641
rect 8809 1589 8861 1633
rect 9009 1807 9061 1851
rect 9009 1799 9018 1807
rect 9018 1799 9052 1807
rect 9052 1799 9061 1807
rect 9209 1913 9218 1921
rect 9218 1913 9252 1921
rect 9252 1913 9261 1921
rect 9209 1869 9261 1913
rect 9409 2087 9461 2131
rect 9409 2079 9418 2087
rect 9418 2079 9452 2087
rect 9452 2079 9461 2087
rect 9609 2193 9618 2201
rect 9618 2193 9652 2201
rect 9652 2193 9661 2201
rect 9609 2149 9661 2193
rect 9809 2367 9861 2411
rect 9809 2359 9818 2367
rect 9818 2359 9852 2367
rect 9852 2359 9861 2367
rect 10009 2563 10018 2571
rect 10018 2563 10052 2571
rect 10052 2563 10061 2571
rect 10009 2519 10061 2563
rect 10209 2737 10261 2781
rect 10209 2729 10218 2737
rect 10218 2729 10252 2737
rect 10252 2729 10261 2737
rect 10409 2843 10418 2851
rect 10418 2843 10452 2851
rect 10452 2843 10461 2851
rect 10409 2799 10461 2843
rect 10609 3017 10661 3061
rect 10609 3009 10618 3017
rect 10618 3009 10652 3017
rect 10652 3009 10661 3017
rect 10809 3123 10818 3131
rect 10818 3123 10852 3131
rect 10852 3123 10861 3131
rect 10809 3079 10861 3123
rect 11009 3297 11061 3341
rect 11009 3289 11018 3297
rect 11018 3289 11052 3297
rect 11052 3289 11061 3297
rect 11209 3403 11218 3411
rect 11218 3403 11252 3411
rect 11252 3403 11261 3411
rect 11209 3359 11261 3403
rect 11409 3577 11461 3621
rect 11409 3569 11418 3577
rect 11418 3569 11452 3577
rect 11452 3569 11461 3577
rect 11609 3773 11618 3781
rect 11618 3773 11652 3781
rect 11652 3773 11661 3781
rect 11609 3729 11661 3773
rect 11809 3947 11861 3991
rect 11809 3939 11818 3947
rect 11818 3939 11852 3947
rect 11852 3939 11861 3947
rect 12009 4053 12018 4061
rect 12018 4053 12052 4061
rect 12052 4053 12061 4061
rect 12009 4009 12061 4053
rect 12209 4227 12261 4271
rect 12209 4219 12218 4227
rect 12218 4219 12252 4227
rect 12252 4219 12261 4227
rect 12409 4333 12418 4341
rect 12418 4333 12452 4341
rect 12452 4333 12461 4341
rect 12409 4289 12461 4333
rect 12609 4507 12661 4551
rect 12609 4499 12618 4507
rect 12618 4499 12652 4507
rect 12652 4499 12661 4507
rect 12809 4613 12818 4621
rect 12818 4613 12852 4621
rect 12852 4613 12861 4621
rect 12809 4569 12861 4613
rect 12907 4569 12959 4621
rect 11609 3684 11661 3693
rect 11609 3650 11618 3684
rect 11618 3650 11652 3684
rect 11652 3650 11661 3684
rect 11609 3641 11661 3650
rect 10009 2474 10061 2483
rect 10009 2440 10018 2474
rect 10018 2440 10052 2474
rect 10052 2440 10061 2474
rect 10009 2431 10061 2440
rect 8409 1264 8461 1273
rect 8409 1230 8418 1264
rect 8418 1230 8452 1264
rect 8452 1230 8461 1264
rect 8409 1221 8461 1230
rect 6809 54 6861 63
rect 6809 20 6818 54
rect 6818 20 6852 54
rect 6852 20 6861 54
rect 6809 11 6861 20
rect 6709 -60 6761 -15
rect 6709 -67 6718 -60
rect 6718 -67 6752 -60
rect 6752 -67 6761 -60
rect 6509 -166 6518 -143
rect 6518 -166 6552 -143
rect 6552 -166 6561 -143
rect 6509 -195 6561 -166
rect 6525 -248 6577 -239
rect 6525 -282 6534 -248
rect 6534 -282 6568 -248
rect 6568 -282 6577 -248
rect 6525 -291 6577 -282
rect 6509 -363 6561 -326
rect 6509 -378 6518 -363
rect 6518 -378 6552 -363
rect 6552 -378 6561 -363
rect 6509 -397 6518 -390
rect 6518 -397 6552 -390
rect 6552 -397 6561 -390
rect 6509 -435 6561 -397
rect 6509 -442 6518 -435
rect 6518 -442 6552 -435
rect 6552 -442 6561 -435
rect 6509 -469 6518 -454
rect 6518 -469 6552 -454
rect 6552 -469 6561 -454
rect 6509 -506 6561 -469
rect 6709 -94 6718 -79
rect 6718 -94 6752 -79
rect 6752 -94 6761 -79
rect 6709 -131 6761 -94
rect 6809 -74 6861 -22
rect 7009 177 7061 221
rect 7009 169 7018 177
rect 7018 169 7052 177
rect 7052 169 7061 177
rect 7209 283 7218 291
rect 7218 283 7252 291
rect 7252 283 7261 291
rect 7209 239 7261 283
rect 7409 457 7461 501
rect 7409 449 7418 457
rect 7418 449 7452 457
rect 7452 449 7461 457
rect 7609 563 7618 571
rect 7618 563 7652 571
rect 7652 563 7661 571
rect 7609 519 7661 563
rect 7809 737 7861 781
rect 7809 729 7818 737
rect 7818 729 7852 737
rect 7852 729 7861 737
rect 8009 843 8018 851
rect 8018 843 8052 851
rect 8052 843 8061 851
rect 8009 799 8061 843
rect 8209 1017 8261 1061
rect 8209 1009 8218 1017
rect 8218 1009 8252 1017
rect 8252 1009 8261 1017
rect 8409 1123 8418 1131
rect 8418 1123 8452 1131
rect 8452 1123 8461 1131
rect 8409 1079 8461 1123
rect 8609 1387 8661 1431
rect 8609 1379 8618 1387
rect 8618 1379 8652 1387
rect 8652 1379 8661 1387
rect 8809 1493 8818 1501
rect 8818 1493 8852 1501
rect 8852 1493 8861 1501
rect 8809 1449 8861 1493
rect 9009 1667 9061 1711
rect 9009 1659 9018 1667
rect 9018 1659 9052 1667
rect 9052 1659 9061 1667
rect 9209 1773 9218 1781
rect 9218 1773 9252 1781
rect 9252 1773 9261 1781
rect 9209 1729 9261 1773
rect 9409 1947 9461 1991
rect 9409 1939 9418 1947
rect 9418 1939 9452 1947
rect 9452 1939 9461 1947
rect 9609 2053 9618 2061
rect 9618 2053 9652 2061
rect 9652 2053 9661 2061
rect 9609 2009 9661 2053
rect 9809 2227 9861 2271
rect 9809 2219 9818 2227
rect 9818 2219 9852 2227
rect 9852 2219 9861 2227
rect 10009 2333 10018 2341
rect 10018 2333 10052 2341
rect 10052 2333 10061 2341
rect 10009 2289 10061 2333
rect 10209 2597 10261 2641
rect 10209 2589 10218 2597
rect 10218 2589 10252 2597
rect 10252 2589 10261 2597
rect 10409 2703 10418 2711
rect 10418 2703 10452 2711
rect 10452 2703 10461 2711
rect 10409 2659 10461 2703
rect 10609 2877 10661 2921
rect 10609 2869 10618 2877
rect 10618 2869 10652 2877
rect 10652 2869 10661 2877
rect 10809 2983 10818 2991
rect 10818 2983 10852 2991
rect 10852 2983 10861 2991
rect 10809 2939 10861 2983
rect 11009 3157 11061 3201
rect 11009 3149 11018 3157
rect 11018 3149 11052 3157
rect 11052 3149 11061 3157
rect 11209 3263 11218 3271
rect 11218 3263 11252 3271
rect 11252 3263 11261 3271
rect 11209 3219 11261 3263
rect 11409 3437 11461 3481
rect 11409 3429 11418 3437
rect 11418 3429 11452 3437
rect 11452 3429 11461 3437
rect 11609 3543 11618 3551
rect 11618 3543 11652 3551
rect 11652 3543 11661 3551
rect 11609 3499 11661 3543
rect 11809 3807 11861 3851
rect 11809 3799 11818 3807
rect 11818 3799 11852 3807
rect 11852 3799 11861 3807
rect 12009 3913 12018 3921
rect 12018 3913 12052 3921
rect 12052 3913 12061 3921
rect 12009 3869 12061 3913
rect 12209 4087 12261 4131
rect 12209 4079 12218 4087
rect 12218 4079 12252 4087
rect 12252 4079 12261 4087
rect 12409 4193 12418 4201
rect 12418 4193 12452 4201
rect 12452 4193 12461 4201
rect 12409 4149 12461 4193
rect 12609 4367 12661 4411
rect 12609 4359 12618 4367
rect 12618 4359 12652 4367
rect 12652 4359 12661 4367
rect 12809 4473 12818 4481
rect 12818 4473 12852 4481
rect 12852 4473 12861 4481
rect 12809 4429 12861 4473
rect 12907 4429 12959 4481
rect 11809 3700 11861 3709
rect 11809 3666 11818 3700
rect 11818 3666 11852 3700
rect 11852 3666 11861 3700
rect 11809 3657 11861 3666
rect 10209 2490 10261 2499
rect 10209 2456 10218 2490
rect 10218 2456 10252 2490
rect 10252 2456 10261 2490
rect 10209 2447 10261 2456
rect 8609 1280 8661 1289
rect 8609 1246 8618 1280
rect 8618 1246 8652 1280
rect 8652 1246 8661 1280
rect 8609 1237 8661 1246
rect 7009 70 7061 79
rect 7009 36 7018 70
rect 7018 36 7052 70
rect 7052 36 7061 70
rect 7009 27 7061 36
rect 6909 -60 6961 -15
rect 6909 -67 6918 -60
rect 6918 -67 6952 -60
rect 6952 -67 6961 -60
rect 6709 -166 6718 -143
rect 6718 -166 6752 -143
rect 6752 -166 6761 -143
rect 6709 -195 6761 -166
rect 6725 -248 6777 -239
rect 6725 -282 6734 -248
rect 6734 -282 6768 -248
rect 6768 -282 6777 -248
rect 6725 -291 6777 -282
rect 6709 -363 6761 -326
rect 6709 -378 6718 -363
rect 6718 -378 6752 -363
rect 6752 -378 6761 -363
rect 6709 -397 6718 -390
rect 6718 -397 6752 -390
rect 6752 -397 6761 -390
rect 6709 -435 6761 -397
rect 6709 -442 6718 -435
rect 6718 -442 6752 -435
rect 6752 -442 6761 -435
rect 6709 -469 6718 -454
rect 6718 -469 6752 -454
rect 6752 -469 6761 -454
rect 6709 -506 6761 -469
rect 6909 -94 6918 -79
rect 6918 -94 6952 -79
rect 6952 -94 6961 -79
rect 6909 -131 6961 -94
rect 7009 -74 7061 -22
rect 7209 143 7218 151
rect 7218 143 7252 151
rect 7252 143 7261 151
rect 7209 99 7261 143
rect 7409 317 7461 361
rect 7409 309 7418 317
rect 7418 309 7452 317
rect 7452 309 7461 317
rect 7609 423 7618 431
rect 7618 423 7652 431
rect 7652 423 7661 431
rect 7609 379 7661 423
rect 7809 597 7861 641
rect 7809 589 7818 597
rect 7818 589 7852 597
rect 7852 589 7861 597
rect 8009 703 8018 711
rect 8018 703 8052 711
rect 8052 703 8061 711
rect 8009 659 8061 703
rect 8209 877 8261 921
rect 8209 869 8218 877
rect 8218 869 8252 877
rect 8252 869 8261 877
rect 8409 983 8418 991
rect 8418 983 8452 991
rect 8452 983 8461 991
rect 8409 939 8461 983
rect 8609 1157 8661 1201
rect 8609 1149 8618 1157
rect 8618 1149 8652 1157
rect 8652 1149 8661 1157
rect 8809 1353 8818 1361
rect 8818 1353 8852 1361
rect 8852 1353 8861 1361
rect 8809 1309 8861 1353
rect 9009 1527 9061 1571
rect 9009 1519 9018 1527
rect 9018 1519 9052 1527
rect 9052 1519 9061 1527
rect 9209 1633 9218 1641
rect 9218 1633 9252 1641
rect 9252 1633 9261 1641
rect 9209 1589 9261 1633
rect 9409 1807 9461 1851
rect 9409 1799 9418 1807
rect 9418 1799 9452 1807
rect 9452 1799 9461 1807
rect 9609 1913 9618 1921
rect 9618 1913 9652 1921
rect 9652 1913 9661 1921
rect 9609 1869 9661 1913
rect 9809 2087 9861 2131
rect 9809 2079 9818 2087
rect 9818 2079 9852 2087
rect 9852 2079 9861 2087
rect 10009 2193 10018 2201
rect 10018 2193 10052 2201
rect 10052 2193 10061 2201
rect 10009 2149 10061 2193
rect 10209 2367 10261 2411
rect 10209 2359 10218 2367
rect 10218 2359 10252 2367
rect 10252 2359 10261 2367
rect 10409 2563 10418 2571
rect 10418 2563 10452 2571
rect 10452 2563 10461 2571
rect 10409 2519 10461 2563
rect 10609 2737 10661 2781
rect 10609 2729 10618 2737
rect 10618 2729 10652 2737
rect 10652 2729 10661 2737
rect 10809 2843 10818 2851
rect 10818 2843 10852 2851
rect 10852 2843 10861 2851
rect 10809 2799 10861 2843
rect 11009 3017 11061 3061
rect 11009 3009 11018 3017
rect 11018 3009 11052 3017
rect 11052 3009 11061 3017
rect 11209 3123 11218 3131
rect 11218 3123 11252 3131
rect 11252 3123 11261 3131
rect 11209 3079 11261 3123
rect 11409 3297 11461 3341
rect 11409 3289 11418 3297
rect 11418 3289 11452 3297
rect 11452 3289 11461 3297
rect 11609 3403 11618 3411
rect 11618 3403 11652 3411
rect 11652 3403 11661 3411
rect 11609 3359 11661 3403
rect 11809 3577 11861 3621
rect 11809 3569 11818 3577
rect 11818 3569 11852 3577
rect 11852 3569 11861 3577
rect 12009 3773 12018 3781
rect 12018 3773 12052 3781
rect 12052 3773 12061 3781
rect 12009 3729 12061 3773
rect 12209 3947 12261 3991
rect 12209 3939 12218 3947
rect 12218 3939 12252 3947
rect 12252 3939 12261 3947
rect 12409 4053 12418 4061
rect 12418 4053 12452 4061
rect 12452 4053 12461 4061
rect 12409 4009 12461 4053
rect 12609 4227 12661 4271
rect 12609 4219 12618 4227
rect 12618 4219 12652 4227
rect 12652 4219 12661 4227
rect 12809 4333 12818 4341
rect 12818 4333 12852 4341
rect 12852 4333 12861 4341
rect 12809 4289 12861 4333
rect 12907 4289 12959 4341
rect 12009 3684 12061 3693
rect 12009 3650 12018 3684
rect 12018 3650 12052 3684
rect 12052 3650 12061 3684
rect 12009 3641 12061 3650
rect 10409 2474 10461 2483
rect 10409 2440 10418 2474
rect 10418 2440 10452 2474
rect 10452 2440 10461 2474
rect 10409 2431 10461 2440
rect 8809 1264 8861 1273
rect 8809 1230 8818 1264
rect 8818 1230 8852 1264
rect 8852 1230 8861 1264
rect 8809 1221 8861 1230
rect 7209 54 7261 63
rect 7209 20 7218 54
rect 7218 20 7252 54
rect 7252 20 7261 54
rect 7209 11 7261 20
rect 7109 -60 7161 -15
rect 7109 -67 7118 -60
rect 7118 -67 7152 -60
rect 7152 -67 7161 -60
rect 6909 -166 6918 -143
rect 6918 -166 6952 -143
rect 6952 -166 6961 -143
rect 6909 -195 6961 -166
rect 6925 -248 6977 -239
rect 6925 -282 6934 -248
rect 6934 -282 6968 -248
rect 6968 -282 6977 -248
rect 6925 -291 6977 -282
rect 6909 -363 6961 -326
rect 6909 -378 6918 -363
rect 6918 -378 6952 -363
rect 6952 -378 6961 -363
rect 6909 -397 6918 -390
rect 6918 -397 6952 -390
rect 6952 -397 6961 -390
rect 6909 -435 6961 -397
rect 6909 -442 6918 -435
rect 6918 -442 6952 -435
rect 6952 -442 6961 -435
rect 6909 -469 6918 -454
rect 6918 -469 6952 -454
rect 6952 -469 6961 -454
rect 6909 -506 6961 -469
rect 7109 -94 7118 -79
rect 7118 -94 7152 -79
rect 7152 -94 7161 -79
rect 7109 -131 7161 -94
rect 7209 -74 7261 -22
rect 7409 177 7461 221
rect 7409 169 7418 177
rect 7418 169 7452 177
rect 7452 169 7461 177
rect 7609 283 7618 291
rect 7618 283 7652 291
rect 7652 283 7661 291
rect 7609 239 7661 283
rect 7809 457 7861 501
rect 7809 449 7818 457
rect 7818 449 7852 457
rect 7852 449 7861 457
rect 8009 563 8018 571
rect 8018 563 8052 571
rect 8052 563 8061 571
rect 8009 519 8061 563
rect 8209 737 8261 781
rect 8209 729 8218 737
rect 8218 729 8252 737
rect 8252 729 8261 737
rect 8409 843 8418 851
rect 8418 843 8452 851
rect 8452 843 8461 851
rect 8409 799 8461 843
rect 8609 1017 8661 1061
rect 8609 1009 8618 1017
rect 8618 1009 8652 1017
rect 8652 1009 8661 1017
rect 8809 1123 8818 1131
rect 8818 1123 8852 1131
rect 8852 1123 8861 1131
rect 8809 1079 8861 1123
rect 9009 1387 9061 1431
rect 9009 1379 9018 1387
rect 9018 1379 9052 1387
rect 9052 1379 9061 1387
rect 9209 1493 9218 1501
rect 9218 1493 9252 1501
rect 9252 1493 9261 1501
rect 9209 1449 9261 1493
rect 9409 1667 9461 1711
rect 9409 1659 9418 1667
rect 9418 1659 9452 1667
rect 9452 1659 9461 1667
rect 9609 1773 9618 1781
rect 9618 1773 9652 1781
rect 9652 1773 9661 1781
rect 9609 1729 9661 1773
rect 9809 1947 9861 1991
rect 9809 1939 9818 1947
rect 9818 1939 9852 1947
rect 9852 1939 9861 1947
rect 10009 2053 10018 2061
rect 10018 2053 10052 2061
rect 10052 2053 10061 2061
rect 10009 2009 10061 2053
rect 10209 2227 10261 2271
rect 10209 2219 10218 2227
rect 10218 2219 10252 2227
rect 10252 2219 10261 2227
rect 10409 2333 10418 2341
rect 10418 2333 10452 2341
rect 10452 2333 10461 2341
rect 10409 2289 10461 2333
rect 10609 2597 10661 2641
rect 10609 2589 10618 2597
rect 10618 2589 10652 2597
rect 10652 2589 10661 2597
rect 10809 2703 10818 2711
rect 10818 2703 10852 2711
rect 10852 2703 10861 2711
rect 10809 2659 10861 2703
rect 11009 2877 11061 2921
rect 11009 2869 11018 2877
rect 11018 2869 11052 2877
rect 11052 2869 11061 2877
rect 11209 2983 11218 2991
rect 11218 2983 11252 2991
rect 11252 2983 11261 2991
rect 11209 2939 11261 2983
rect 11409 3157 11461 3201
rect 11409 3149 11418 3157
rect 11418 3149 11452 3157
rect 11452 3149 11461 3157
rect 11609 3263 11618 3271
rect 11618 3263 11652 3271
rect 11652 3263 11661 3271
rect 11609 3219 11661 3263
rect 11809 3437 11861 3481
rect 11809 3429 11818 3437
rect 11818 3429 11852 3437
rect 11852 3429 11861 3437
rect 12009 3543 12018 3551
rect 12018 3543 12052 3551
rect 12052 3543 12061 3551
rect 12009 3499 12061 3543
rect 12209 3807 12261 3851
rect 12209 3799 12218 3807
rect 12218 3799 12252 3807
rect 12252 3799 12261 3807
rect 12409 3913 12418 3921
rect 12418 3913 12452 3921
rect 12452 3913 12461 3921
rect 12409 3869 12461 3913
rect 12609 4087 12661 4131
rect 12609 4079 12618 4087
rect 12618 4079 12652 4087
rect 12652 4079 12661 4087
rect 12809 4193 12818 4201
rect 12818 4193 12852 4201
rect 12852 4193 12861 4201
rect 12809 4149 12861 4193
rect 12907 4149 12959 4201
rect 12209 3700 12261 3709
rect 12209 3666 12218 3700
rect 12218 3666 12252 3700
rect 12252 3666 12261 3700
rect 12209 3657 12261 3666
rect 10609 2490 10661 2499
rect 10609 2456 10618 2490
rect 10618 2456 10652 2490
rect 10652 2456 10661 2490
rect 10609 2447 10661 2456
rect 9009 1280 9061 1289
rect 9009 1246 9018 1280
rect 9018 1246 9052 1280
rect 9052 1246 9061 1280
rect 9009 1237 9061 1246
rect 7409 70 7461 79
rect 7409 36 7418 70
rect 7418 36 7452 70
rect 7452 36 7461 70
rect 7409 27 7461 36
rect 7309 -60 7361 -15
rect 7309 -67 7318 -60
rect 7318 -67 7352 -60
rect 7352 -67 7361 -60
rect 7109 -166 7118 -143
rect 7118 -166 7152 -143
rect 7152 -166 7161 -143
rect 7109 -195 7161 -166
rect 7125 -248 7177 -239
rect 7125 -282 7134 -248
rect 7134 -282 7168 -248
rect 7168 -282 7177 -248
rect 7125 -291 7177 -282
rect 7109 -363 7161 -326
rect 7109 -378 7118 -363
rect 7118 -378 7152 -363
rect 7152 -378 7161 -363
rect 7109 -397 7118 -390
rect 7118 -397 7152 -390
rect 7152 -397 7161 -390
rect 7109 -435 7161 -397
rect 7109 -442 7118 -435
rect 7118 -442 7152 -435
rect 7152 -442 7161 -435
rect 7109 -469 7118 -454
rect 7118 -469 7152 -454
rect 7152 -469 7161 -454
rect 7109 -506 7161 -469
rect 7309 -94 7318 -79
rect 7318 -94 7352 -79
rect 7352 -94 7361 -79
rect 7309 -131 7361 -94
rect 7409 -74 7461 -22
rect 7609 143 7618 151
rect 7618 143 7652 151
rect 7652 143 7661 151
rect 7609 99 7661 143
rect 7809 317 7861 361
rect 7809 309 7818 317
rect 7818 309 7852 317
rect 7852 309 7861 317
rect 8009 423 8018 431
rect 8018 423 8052 431
rect 8052 423 8061 431
rect 8009 379 8061 423
rect 8209 597 8261 641
rect 8209 589 8218 597
rect 8218 589 8252 597
rect 8252 589 8261 597
rect 8409 703 8418 711
rect 8418 703 8452 711
rect 8452 703 8461 711
rect 8409 659 8461 703
rect 8609 877 8661 921
rect 8609 869 8618 877
rect 8618 869 8652 877
rect 8652 869 8661 877
rect 8809 983 8818 991
rect 8818 983 8852 991
rect 8852 983 8861 991
rect 8809 939 8861 983
rect 9009 1157 9061 1201
rect 9009 1149 9018 1157
rect 9018 1149 9052 1157
rect 9052 1149 9061 1157
rect 9209 1353 9218 1361
rect 9218 1353 9252 1361
rect 9252 1353 9261 1361
rect 9209 1309 9261 1353
rect 9409 1527 9461 1571
rect 9409 1519 9418 1527
rect 9418 1519 9452 1527
rect 9452 1519 9461 1527
rect 9609 1633 9618 1641
rect 9618 1633 9652 1641
rect 9652 1633 9661 1641
rect 9609 1589 9661 1633
rect 9809 1807 9861 1851
rect 9809 1799 9818 1807
rect 9818 1799 9852 1807
rect 9852 1799 9861 1807
rect 10009 1913 10018 1921
rect 10018 1913 10052 1921
rect 10052 1913 10061 1921
rect 10009 1869 10061 1913
rect 10209 2087 10261 2131
rect 10209 2079 10218 2087
rect 10218 2079 10252 2087
rect 10252 2079 10261 2087
rect 10409 2193 10418 2201
rect 10418 2193 10452 2201
rect 10452 2193 10461 2201
rect 10409 2149 10461 2193
rect 10609 2367 10661 2411
rect 10609 2359 10618 2367
rect 10618 2359 10652 2367
rect 10652 2359 10661 2367
rect 10809 2563 10818 2571
rect 10818 2563 10852 2571
rect 10852 2563 10861 2571
rect 10809 2519 10861 2563
rect 11009 2737 11061 2781
rect 11009 2729 11018 2737
rect 11018 2729 11052 2737
rect 11052 2729 11061 2737
rect 11209 2843 11218 2851
rect 11218 2843 11252 2851
rect 11252 2843 11261 2851
rect 11209 2799 11261 2843
rect 11409 3017 11461 3061
rect 11409 3009 11418 3017
rect 11418 3009 11452 3017
rect 11452 3009 11461 3017
rect 11609 3123 11618 3131
rect 11618 3123 11652 3131
rect 11652 3123 11661 3131
rect 11609 3079 11661 3123
rect 11809 3297 11861 3341
rect 11809 3289 11818 3297
rect 11818 3289 11852 3297
rect 11852 3289 11861 3297
rect 12009 3403 12018 3411
rect 12018 3403 12052 3411
rect 12052 3403 12061 3411
rect 12009 3359 12061 3403
rect 12209 3577 12261 3621
rect 12209 3569 12218 3577
rect 12218 3569 12252 3577
rect 12252 3569 12261 3577
rect 12409 3773 12418 3781
rect 12418 3773 12452 3781
rect 12452 3773 12461 3781
rect 12409 3729 12461 3773
rect 12609 3947 12661 3991
rect 12609 3939 12618 3947
rect 12618 3939 12652 3947
rect 12652 3939 12661 3947
rect 12809 4053 12818 4061
rect 12818 4053 12852 4061
rect 12852 4053 12861 4061
rect 12809 4009 12861 4053
rect 12907 4009 12959 4061
rect 12409 3684 12461 3693
rect 12409 3650 12418 3684
rect 12418 3650 12452 3684
rect 12452 3650 12461 3684
rect 12409 3641 12461 3650
rect 10809 2474 10861 2483
rect 10809 2440 10818 2474
rect 10818 2440 10852 2474
rect 10852 2440 10861 2474
rect 10809 2431 10861 2440
rect 9209 1264 9261 1273
rect 9209 1230 9218 1264
rect 9218 1230 9252 1264
rect 9252 1230 9261 1264
rect 9209 1221 9261 1230
rect 7609 54 7661 63
rect 7609 20 7618 54
rect 7618 20 7652 54
rect 7652 20 7661 54
rect 7609 11 7661 20
rect 7509 -60 7561 -15
rect 7509 -67 7518 -60
rect 7518 -67 7552 -60
rect 7552 -67 7561 -60
rect 7309 -166 7318 -143
rect 7318 -166 7352 -143
rect 7352 -166 7361 -143
rect 7309 -195 7361 -166
rect 7325 -248 7377 -239
rect 7325 -282 7334 -248
rect 7334 -282 7368 -248
rect 7368 -282 7377 -248
rect 7325 -291 7377 -282
rect 7309 -363 7361 -326
rect 7309 -378 7318 -363
rect 7318 -378 7352 -363
rect 7352 -378 7361 -363
rect 7309 -397 7318 -390
rect 7318 -397 7352 -390
rect 7352 -397 7361 -390
rect 7309 -435 7361 -397
rect 7309 -442 7318 -435
rect 7318 -442 7352 -435
rect 7352 -442 7361 -435
rect 7309 -469 7318 -454
rect 7318 -469 7352 -454
rect 7352 -469 7361 -454
rect 7309 -506 7361 -469
rect 7509 -94 7518 -79
rect 7518 -94 7552 -79
rect 7552 -94 7561 -79
rect 7509 -131 7561 -94
rect 7609 -74 7661 -22
rect 7809 177 7861 221
rect 7809 169 7818 177
rect 7818 169 7852 177
rect 7852 169 7861 177
rect 8009 283 8018 291
rect 8018 283 8052 291
rect 8052 283 8061 291
rect 8009 239 8061 283
rect 8209 457 8261 501
rect 8209 449 8218 457
rect 8218 449 8252 457
rect 8252 449 8261 457
rect 8409 563 8418 571
rect 8418 563 8452 571
rect 8452 563 8461 571
rect 8409 519 8461 563
rect 8609 737 8661 781
rect 8609 729 8618 737
rect 8618 729 8652 737
rect 8652 729 8661 737
rect 8809 843 8818 851
rect 8818 843 8852 851
rect 8852 843 8861 851
rect 8809 799 8861 843
rect 9009 1017 9061 1061
rect 9009 1009 9018 1017
rect 9018 1009 9052 1017
rect 9052 1009 9061 1017
rect 9209 1123 9218 1131
rect 9218 1123 9252 1131
rect 9252 1123 9261 1131
rect 9209 1079 9261 1123
rect 9409 1387 9461 1431
rect 9409 1379 9418 1387
rect 9418 1379 9452 1387
rect 9452 1379 9461 1387
rect 9609 1493 9618 1501
rect 9618 1493 9652 1501
rect 9652 1493 9661 1501
rect 9609 1449 9661 1493
rect 9809 1667 9861 1711
rect 9809 1659 9818 1667
rect 9818 1659 9852 1667
rect 9852 1659 9861 1667
rect 10009 1773 10018 1781
rect 10018 1773 10052 1781
rect 10052 1773 10061 1781
rect 10009 1729 10061 1773
rect 10209 1947 10261 1991
rect 10209 1939 10218 1947
rect 10218 1939 10252 1947
rect 10252 1939 10261 1947
rect 10409 2053 10418 2061
rect 10418 2053 10452 2061
rect 10452 2053 10461 2061
rect 10409 2009 10461 2053
rect 10609 2227 10661 2271
rect 10609 2219 10618 2227
rect 10618 2219 10652 2227
rect 10652 2219 10661 2227
rect 10809 2333 10818 2341
rect 10818 2333 10852 2341
rect 10852 2333 10861 2341
rect 10809 2289 10861 2333
rect 11009 2597 11061 2641
rect 11009 2589 11018 2597
rect 11018 2589 11052 2597
rect 11052 2589 11061 2597
rect 11209 2703 11218 2711
rect 11218 2703 11252 2711
rect 11252 2703 11261 2711
rect 11209 2659 11261 2703
rect 11409 2877 11461 2921
rect 11409 2869 11418 2877
rect 11418 2869 11452 2877
rect 11452 2869 11461 2877
rect 11609 2983 11618 2991
rect 11618 2983 11652 2991
rect 11652 2983 11661 2991
rect 11609 2939 11661 2983
rect 11809 3157 11861 3201
rect 11809 3149 11818 3157
rect 11818 3149 11852 3157
rect 11852 3149 11861 3157
rect 12009 3263 12018 3271
rect 12018 3263 12052 3271
rect 12052 3263 12061 3271
rect 12009 3219 12061 3263
rect 12209 3437 12261 3481
rect 12209 3429 12218 3437
rect 12218 3429 12252 3437
rect 12252 3429 12261 3437
rect 12409 3543 12418 3551
rect 12418 3543 12452 3551
rect 12452 3543 12461 3551
rect 12409 3499 12461 3543
rect 12609 3807 12661 3851
rect 12609 3799 12618 3807
rect 12618 3799 12652 3807
rect 12652 3799 12661 3807
rect 12809 3913 12818 3921
rect 12818 3913 12852 3921
rect 12852 3913 12861 3921
rect 12809 3869 12861 3913
rect 12907 3869 12959 3921
rect 12609 3700 12661 3709
rect 12609 3666 12618 3700
rect 12618 3666 12652 3700
rect 12652 3666 12661 3700
rect 12609 3657 12661 3666
rect 11009 2490 11061 2499
rect 11009 2456 11018 2490
rect 11018 2456 11052 2490
rect 11052 2456 11061 2490
rect 11009 2447 11061 2456
rect 9409 1280 9461 1289
rect 9409 1246 9418 1280
rect 9418 1246 9452 1280
rect 9452 1246 9461 1280
rect 9409 1237 9461 1246
rect 7809 70 7861 79
rect 7809 36 7818 70
rect 7818 36 7852 70
rect 7852 36 7861 70
rect 7809 27 7861 36
rect 7709 -60 7761 -15
rect 7709 -67 7718 -60
rect 7718 -67 7752 -60
rect 7752 -67 7761 -60
rect 7509 -166 7518 -143
rect 7518 -166 7552 -143
rect 7552 -166 7561 -143
rect 7509 -195 7561 -166
rect 7525 -248 7577 -239
rect 7525 -282 7534 -248
rect 7534 -282 7568 -248
rect 7568 -282 7577 -248
rect 7525 -291 7577 -282
rect 7509 -363 7561 -326
rect 7509 -378 7518 -363
rect 7518 -378 7552 -363
rect 7552 -378 7561 -363
rect 7509 -397 7518 -390
rect 7518 -397 7552 -390
rect 7552 -397 7561 -390
rect 7509 -435 7561 -397
rect 7509 -442 7518 -435
rect 7518 -442 7552 -435
rect 7552 -442 7561 -435
rect 7509 -469 7518 -454
rect 7518 -469 7552 -454
rect 7552 -469 7561 -454
rect 7509 -506 7561 -469
rect 7709 -94 7718 -79
rect 7718 -94 7752 -79
rect 7752 -94 7761 -79
rect 7709 -131 7761 -94
rect 7809 -74 7861 -22
rect 8009 143 8018 151
rect 8018 143 8052 151
rect 8052 143 8061 151
rect 8009 99 8061 143
rect 8209 317 8261 361
rect 8209 309 8218 317
rect 8218 309 8252 317
rect 8252 309 8261 317
rect 8409 423 8418 431
rect 8418 423 8452 431
rect 8452 423 8461 431
rect 8409 379 8461 423
rect 8609 597 8661 641
rect 8609 589 8618 597
rect 8618 589 8652 597
rect 8652 589 8661 597
rect 8809 703 8818 711
rect 8818 703 8852 711
rect 8852 703 8861 711
rect 8809 659 8861 703
rect 9009 877 9061 921
rect 9009 869 9018 877
rect 9018 869 9052 877
rect 9052 869 9061 877
rect 9209 983 9218 991
rect 9218 983 9252 991
rect 9252 983 9261 991
rect 9209 939 9261 983
rect 9409 1157 9461 1201
rect 9409 1149 9418 1157
rect 9418 1149 9452 1157
rect 9452 1149 9461 1157
rect 9609 1353 9618 1361
rect 9618 1353 9652 1361
rect 9652 1353 9661 1361
rect 9609 1309 9661 1353
rect 9809 1527 9861 1571
rect 9809 1519 9818 1527
rect 9818 1519 9852 1527
rect 9852 1519 9861 1527
rect 10009 1633 10018 1641
rect 10018 1633 10052 1641
rect 10052 1633 10061 1641
rect 10009 1589 10061 1633
rect 10209 1807 10261 1851
rect 10209 1799 10218 1807
rect 10218 1799 10252 1807
rect 10252 1799 10261 1807
rect 10409 1913 10418 1921
rect 10418 1913 10452 1921
rect 10452 1913 10461 1921
rect 10409 1869 10461 1913
rect 10609 2087 10661 2131
rect 10609 2079 10618 2087
rect 10618 2079 10652 2087
rect 10652 2079 10661 2087
rect 10809 2193 10818 2201
rect 10818 2193 10852 2201
rect 10852 2193 10861 2201
rect 10809 2149 10861 2193
rect 11009 2367 11061 2411
rect 11009 2359 11018 2367
rect 11018 2359 11052 2367
rect 11052 2359 11061 2367
rect 11209 2563 11218 2571
rect 11218 2563 11252 2571
rect 11252 2563 11261 2571
rect 11209 2519 11261 2563
rect 11409 2737 11461 2781
rect 11409 2729 11418 2737
rect 11418 2729 11452 2737
rect 11452 2729 11461 2737
rect 11609 2843 11618 2851
rect 11618 2843 11652 2851
rect 11652 2843 11661 2851
rect 11609 2799 11661 2843
rect 11809 3017 11861 3061
rect 11809 3009 11818 3017
rect 11818 3009 11852 3017
rect 11852 3009 11861 3017
rect 12009 3123 12018 3131
rect 12018 3123 12052 3131
rect 12052 3123 12061 3131
rect 12009 3079 12061 3123
rect 12209 3297 12261 3341
rect 12209 3289 12218 3297
rect 12218 3289 12252 3297
rect 12252 3289 12261 3297
rect 12409 3403 12418 3411
rect 12418 3403 12452 3411
rect 12452 3403 12461 3411
rect 12409 3359 12461 3403
rect 12609 3577 12661 3621
rect 12609 3569 12618 3577
rect 12618 3569 12652 3577
rect 12652 3569 12661 3577
rect 12809 3773 12818 3781
rect 12818 3773 12852 3781
rect 12852 3773 12861 3781
rect 12809 3729 12861 3773
rect 12907 3729 12959 3781
rect 11209 2474 11261 2483
rect 11209 2440 11218 2474
rect 11218 2440 11252 2474
rect 11252 2440 11261 2474
rect 11209 2431 11261 2440
rect 9609 1264 9661 1273
rect 9609 1230 9618 1264
rect 9618 1230 9652 1264
rect 9652 1230 9661 1264
rect 9609 1221 9661 1230
rect 8009 54 8061 63
rect 8009 20 8018 54
rect 8018 20 8052 54
rect 8052 20 8061 54
rect 8009 11 8061 20
rect 7909 -60 7961 -15
rect 7909 -67 7918 -60
rect 7918 -67 7952 -60
rect 7952 -67 7961 -60
rect 7709 -166 7718 -143
rect 7718 -166 7752 -143
rect 7752 -166 7761 -143
rect 7709 -195 7761 -166
rect 7725 -248 7777 -239
rect 7725 -282 7734 -248
rect 7734 -282 7768 -248
rect 7768 -282 7777 -248
rect 7725 -291 7777 -282
rect 7709 -363 7761 -326
rect 7709 -378 7718 -363
rect 7718 -378 7752 -363
rect 7752 -378 7761 -363
rect 7709 -397 7718 -390
rect 7718 -397 7752 -390
rect 7752 -397 7761 -390
rect 7709 -435 7761 -397
rect 7709 -442 7718 -435
rect 7718 -442 7752 -435
rect 7752 -442 7761 -435
rect 7709 -469 7718 -454
rect 7718 -469 7752 -454
rect 7752 -469 7761 -454
rect 7709 -506 7761 -469
rect 7909 -94 7918 -79
rect 7918 -94 7952 -79
rect 7952 -94 7961 -79
rect 7909 -131 7961 -94
rect 8009 -74 8061 -22
rect 8209 177 8261 221
rect 8209 169 8218 177
rect 8218 169 8252 177
rect 8252 169 8261 177
rect 8409 283 8418 291
rect 8418 283 8452 291
rect 8452 283 8461 291
rect 8409 239 8461 283
rect 8609 457 8661 501
rect 8609 449 8618 457
rect 8618 449 8652 457
rect 8652 449 8661 457
rect 8809 563 8818 571
rect 8818 563 8852 571
rect 8852 563 8861 571
rect 8809 519 8861 563
rect 9009 737 9061 781
rect 9009 729 9018 737
rect 9018 729 9052 737
rect 9052 729 9061 737
rect 9209 843 9218 851
rect 9218 843 9252 851
rect 9252 843 9261 851
rect 9209 799 9261 843
rect 9409 1017 9461 1061
rect 9409 1009 9418 1017
rect 9418 1009 9452 1017
rect 9452 1009 9461 1017
rect 9609 1123 9618 1131
rect 9618 1123 9652 1131
rect 9652 1123 9661 1131
rect 9609 1079 9661 1123
rect 9809 1387 9861 1431
rect 9809 1379 9818 1387
rect 9818 1379 9852 1387
rect 9852 1379 9861 1387
rect 10009 1493 10018 1501
rect 10018 1493 10052 1501
rect 10052 1493 10061 1501
rect 10009 1449 10061 1493
rect 10209 1667 10261 1711
rect 10209 1659 10218 1667
rect 10218 1659 10252 1667
rect 10252 1659 10261 1667
rect 10409 1773 10418 1781
rect 10418 1773 10452 1781
rect 10452 1773 10461 1781
rect 10409 1729 10461 1773
rect 10609 1947 10661 1991
rect 10609 1939 10618 1947
rect 10618 1939 10652 1947
rect 10652 1939 10661 1947
rect 10809 2053 10818 2061
rect 10818 2053 10852 2061
rect 10852 2053 10861 2061
rect 10809 2009 10861 2053
rect 11009 2227 11061 2271
rect 11009 2219 11018 2227
rect 11018 2219 11052 2227
rect 11052 2219 11061 2227
rect 11209 2333 11218 2341
rect 11218 2333 11252 2341
rect 11252 2333 11261 2341
rect 11209 2289 11261 2333
rect 11409 2597 11461 2641
rect 11409 2589 11418 2597
rect 11418 2589 11452 2597
rect 11452 2589 11461 2597
rect 11609 2703 11618 2711
rect 11618 2703 11652 2711
rect 11652 2703 11661 2711
rect 11609 2659 11661 2703
rect 11809 2877 11861 2921
rect 11809 2869 11818 2877
rect 11818 2869 11852 2877
rect 11852 2869 11861 2877
rect 12009 2983 12018 2991
rect 12018 2983 12052 2991
rect 12052 2983 12061 2991
rect 12009 2939 12061 2983
rect 12209 3157 12261 3201
rect 12209 3149 12218 3157
rect 12218 3149 12252 3157
rect 12252 3149 12261 3157
rect 12409 3263 12418 3271
rect 12418 3263 12452 3271
rect 12452 3263 12461 3271
rect 12409 3219 12461 3263
rect 12609 3437 12661 3481
rect 12609 3429 12618 3437
rect 12618 3429 12652 3437
rect 12652 3429 12661 3437
rect 12809 3543 12818 3551
rect 12818 3543 12852 3551
rect 12852 3543 12861 3551
rect 12809 3499 12861 3543
rect 12907 3499 12959 3551
rect 11409 2490 11461 2499
rect 11409 2456 11418 2490
rect 11418 2456 11452 2490
rect 11452 2456 11461 2490
rect 11409 2447 11461 2456
rect 9809 1280 9861 1289
rect 9809 1246 9818 1280
rect 9818 1246 9852 1280
rect 9852 1246 9861 1280
rect 9809 1237 9861 1246
rect 8209 70 8261 79
rect 8209 36 8218 70
rect 8218 36 8252 70
rect 8252 36 8261 70
rect 8209 27 8261 36
rect 8109 -60 8161 -15
rect 8109 -67 8118 -60
rect 8118 -67 8152 -60
rect 8152 -67 8161 -60
rect 7909 -166 7918 -143
rect 7918 -166 7952 -143
rect 7952 -166 7961 -143
rect 7909 -195 7961 -166
rect 7925 -248 7977 -239
rect 7925 -282 7934 -248
rect 7934 -282 7968 -248
rect 7968 -282 7977 -248
rect 7925 -291 7977 -282
rect 7909 -363 7961 -326
rect 7909 -378 7918 -363
rect 7918 -378 7952 -363
rect 7952 -378 7961 -363
rect 7909 -397 7918 -390
rect 7918 -397 7952 -390
rect 7952 -397 7961 -390
rect 7909 -435 7961 -397
rect 7909 -442 7918 -435
rect 7918 -442 7952 -435
rect 7952 -442 7961 -435
rect 7909 -469 7918 -454
rect 7918 -469 7952 -454
rect 7952 -469 7961 -454
rect 7909 -506 7961 -469
rect 8109 -94 8118 -79
rect 8118 -94 8152 -79
rect 8152 -94 8161 -79
rect 8109 -131 8161 -94
rect 8209 -74 8261 -22
rect 8409 143 8418 151
rect 8418 143 8452 151
rect 8452 143 8461 151
rect 8409 99 8461 143
rect 8609 317 8661 361
rect 8609 309 8618 317
rect 8618 309 8652 317
rect 8652 309 8661 317
rect 8809 423 8818 431
rect 8818 423 8852 431
rect 8852 423 8861 431
rect 8809 379 8861 423
rect 9009 597 9061 641
rect 9009 589 9018 597
rect 9018 589 9052 597
rect 9052 589 9061 597
rect 9209 703 9218 711
rect 9218 703 9252 711
rect 9252 703 9261 711
rect 9209 659 9261 703
rect 9409 877 9461 921
rect 9409 869 9418 877
rect 9418 869 9452 877
rect 9452 869 9461 877
rect 9609 983 9618 991
rect 9618 983 9652 991
rect 9652 983 9661 991
rect 9609 939 9661 983
rect 9809 1157 9861 1201
rect 9809 1149 9818 1157
rect 9818 1149 9852 1157
rect 9852 1149 9861 1157
rect 10009 1353 10018 1361
rect 10018 1353 10052 1361
rect 10052 1353 10061 1361
rect 10009 1309 10061 1353
rect 10209 1527 10261 1571
rect 10209 1519 10218 1527
rect 10218 1519 10252 1527
rect 10252 1519 10261 1527
rect 10409 1633 10418 1641
rect 10418 1633 10452 1641
rect 10452 1633 10461 1641
rect 10409 1589 10461 1633
rect 10609 1807 10661 1851
rect 10609 1799 10618 1807
rect 10618 1799 10652 1807
rect 10652 1799 10661 1807
rect 10809 1913 10818 1921
rect 10818 1913 10852 1921
rect 10852 1913 10861 1921
rect 10809 1869 10861 1913
rect 11009 2087 11061 2131
rect 11009 2079 11018 2087
rect 11018 2079 11052 2087
rect 11052 2079 11061 2087
rect 11209 2193 11218 2201
rect 11218 2193 11252 2201
rect 11252 2193 11261 2201
rect 11209 2149 11261 2193
rect 11409 2367 11461 2411
rect 11409 2359 11418 2367
rect 11418 2359 11452 2367
rect 11452 2359 11461 2367
rect 11609 2563 11618 2571
rect 11618 2563 11652 2571
rect 11652 2563 11661 2571
rect 11609 2519 11661 2563
rect 11809 2737 11861 2781
rect 11809 2729 11818 2737
rect 11818 2729 11852 2737
rect 11852 2729 11861 2737
rect 12009 2843 12018 2851
rect 12018 2843 12052 2851
rect 12052 2843 12061 2851
rect 12009 2799 12061 2843
rect 12209 3017 12261 3061
rect 12209 3009 12218 3017
rect 12218 3009 12252 3017
rect 12252 3009 12261 3017
rect 12409 3123 12418 3131
rect 12418 3123 12452 3131
rect 12452 3123 12461 3131
rect 12409 3079 12461 3123
rect 12609 3297 12661 3341
rect 12609 3289 12618 3297
rect 12618 3289 12652 3297
rect 12652 3289 12661 3297
rect 12809 3403 12818 3411
rect 12818 3403 12852 3411
rect 12852 3403 12861 3411
rect 12809 3359 12861 3403
rect 12907 3359 12959 3411
rect 11609 2474 11661 2483
rect 11609 2440 11618 2474
rect 11618 2440 11652 2474
rect 11652 2440 11661 2474
rect 11609 2431 11661 2440
rect 10009 1264 10061 1273
rect 10009 1230 10018 1264
rect 10018 1230 10052 1264
rect 10052 1230 10061 1264
rect 10009 1221 10061 1230
rect 8409 54 8461 63
rect 8409 20 8418 54
rect 8418 20 8452 54
rect 8452 20 8461 54
rect 8409 11 8461 20
rect 8309 -60 8361 -15
rect 8309 -67 8318 -60
rect 8318 -67 8352 -60
rect 8352 -67 8361 -60
rect 8109 -166 8118 -143
rect 8118 -166 8152 -143
rect 8152 -166 8161 -143
rect 8109 -195 8161 -166
rect 8125 -248 8177 -239
rect 8125 -282 8134 -248
rect 8134 -282 8168 -248
rect 8168 -282 8177 -248
rect 8125 -291 8177 -282
rect 8109 -363 8161 -326
rect 8109 -378 8118 -363
rect 8118 -378 8152 -363
rect 8152 -378 8161 -363
rect 8109 -397 8118 -390
rect 8118 -397 8152 -390
rect 8152 -397 8161 -390
rect 8109 -435 8161 -397
rect 8109 -442 8118 -435
rect 8118 -442 8152 -435
rect 8152 -442 8161 -435
rect 8109 -469 8118 -454
rect 8118 -469 8152 -454
rect 8152 -469 8161 -454
rect 8109 -506 8161 -469
rect 8309 -94 8318 -79
rect 8318 -94 8352 -79
rect 8352 -94 8361 -79
rect 8309 -131 8361 -94
rect 8409 -74 8461 -22
rect 8609 177 8661 221
rect 8609 169 8618 177
rect 8618 169 8652 177
rect 8652 169 8661 177
rect 8809 283 8818 291
rect 8818 283 8852 291
rect 8852 283 8861 291
rect 8809 239 8861 283
rect 9009 457 9061 501
rect 9009 449 9018 457
rect 9018 449 9052 457
rect 9052 449 9061 457
rect 9209 563 9218 571
rect 9218 563 9252 571
rect 9252 563 9261 571
rect 9209 519 9261 563
rect 9409 737 9461 781
rect 9409 729 9418 737
rect 9418 729 9452 737
rect 9452 729 9461 737
rect 9609 843 9618 851
rect 9618 843 9652 851
rect 9652 843 9661 851
rect 9609 799 9661 843
rect 9809 1017 9861 1061
rect 9809 1009 9818 1017
rect 9818 1009 9852 1017
rect 9852 1009 9861 1017
rect 10009 1123 10018 1131
rect 10018 1123 10052 1131
rect 10052 1123 10061 1131
rect 10009 1079 10061 1123
rect 10209 1387 10261 1431
rect 10209 1379 10218 1387
rect 10218 1379 10252 1387
rect 10252 1379 10261 1387
rect 10409 1493 10418 1501
rect 10418 1493 10452 1501
rect 10452 1493 10461 1501
rect 10409 1449 10461 1493
rect 10609 1667 10661 1711
rect 10609 1659 10618 1667
rect 10618 1659 10652 1667
rect 10652 1659 10661 1667
rect 10809 1773 10818 1781
rect 10818 1773 10852 1781
rect 10852 1773 10861 1781
rect 10809 1729 10861 1773
rect 11009 1947 11061 1991
rect 11009 1939 11018 1947
rect 11018 1939 11052 1947
rect 11052 1939 11061 1947
rect 11209 2053 11218 2061
rect 11218 2053 11252 2061
rect 11252 2053 11261 2061
rect 11209 2009 11261 2053
rect 11409 2227 11461 2271
rect 11409 2219 11418 2227
rect 11418 2219 11452 2227
rect 11452 2219 11461 2227
rect 11609 2333 11618 2341
rect 11618 2333 11652 2341
rect 11652 2333 11661 2341
rect 11609 2289 11661 2333
rect 11809 2597 11861 2641
rect 11809 2589 11818 2597
rect 11818 2589 11852 2597
rect 11852 2589 11861 2597
rect 12009 2703 12018 2711
rect 12018 2703 12052 2711
rect 12052 2703 12061 2711
rect 12009 2659 12061 2703
rect 12209 2877 12261 2921
rect 12209 2869 12218 2877
rect 12218 2869 12252 2877
rect 12252 2869 12261 2877
rect 12409 2983 12418 2991
rect 12418 2983 12452 2991
rect 12452 2983 12461 2991
rect 12409 2939 12461 2983
rect 12609 3157 12661 3201
rect 12609 3149 12618 3157
rect 12618 3149 12652 3157
rect 12652 3149 12661 3157
rect 12809 3263 12818 3271
rect 12818 3263 12852 3271
rect 12852 3263 12861 3271
rect 12809 3219 12861 3263
rect 12907 3219 12959 3271
rect 11809 2490 11861 2499
rect 11809 2456 11818 2490
rect 11818 2456 11852 2490
rect 11852 2456 11861 2490
rect 11809 2447 11861 2456
rect 10209 1280 10261 1289
rect 10209 1246 10218 1280
rect 10218 1246 10252 1280
rect 10252 1246 10261 1280
rect 10209 1237 10261 1246
rect 8609 70 8661 79
rect 8609 36 8618 70
rect 8618 36 8652 70
rect 8652 36 8661 70
rect 8609 27 8661 36
rect 8509 -60 8561 -15
rect 8509 -67 8518 -60
rect 8518 -67 8552 -60
rect 8552 -67 8561 -60
rect 8309 -166 8318 -143
rect 8318 -166 8352 -143
rect 8352 -166 8361 -143
rect 8309 -195 8361 -166
rect 8325 -248 8377 -239
rect 8325 -282 8334 -248
rect 8334 -282 8368 -248
rect 8368 -282 8377 -248
rect 8325 -291 8377 -282
rect 8309 -363 8361 -326
rect 8309 -378 8318 -363
rect 8318 -378 8352 -363
rect 8352 -378 8361 -363
rect 8309 -397 8318 -390
rect 8318 -397 8352 -390
rect 8352 -397 8361 -390
rect 8309 -435 8361 -397
rect 8309 -442 8318 -435
rect 8318 -442 8352 -435
rect 8352 -442 8361 -435
rect 8309 -469 8318 -454
rect 8318 -469 8352 -454
rect 8352 -469 8361 -454
rect 8309 -506 8361 -469
rect 8509 -94 8518 -79
rect 8518 -94 8552 -79
rect 8552 -94 8561 -79
rect 8509 -131 8561 -94
rect 8609 -74 8661 -22
rect 8809 143 8818 151
rect 8818 143 8852 151
rect 8852 143 8861 151
rect 8809 99 8861 143
rect 9009 317 9061 361
rect 9009 309 9018 317
rect 9018 309 9052 317
rect 9052 309 9061 317
rect 9209 423 9218 431
rect 9218 423 9252 431
rect 9252 423 9261 431
rect 9209 379 9261 423
rect 9409 597 9461 641
rect 9409 589 9418 597
rect 9418 589 9452 597
rect 9452 589 9461 597
rect 9609 703 9618 711
rect 9618 703 9652 711
rect 9652 703 9661 711
rect 9609 659 9661 703
rect 9809 877 9861 921
rect 9809 869 9818 877
rect 9818 869 9852 877
rect 9852 869 9861 877
rect 10009 983 10018 991
rect 10018 983 10052 991
rect 10052 983 10061 991
rect 10009 939 10061 983
rect 10209 1157 10261 1201
rect 10209 1149 10218 1157
rect 10218 1149 10252 1157
rect 10252 1149 10261 1157
rect 10409 1353 10418 1361
rect 10418 1353 10452 1361
rect 10452 1353 10461 1361
rect 10409 1309 10461 1353
rect 10609 1527 10661 1571
rect 10609 1519 10618 1527
rect 10618 1519 10652 1527
rect 10652 1519 10661 1527
rect 10809 1633 10818 1641
rect 10818 1633 10852 1641
rect 10852 1633 10861 1641
rect 10809 1589 10861 1633
rect 11009 1807 11061 1851
rect 11009 1799 11018 1807
rect 11018 1799 11052 1807
rect 11052 1799 11061 1807
rect 11209 1913 11218 1921
rect 11218 1913 11252 1921
rect 11252 1913 11261 1921
rect 11209 1869 11261 1913
rect 11409 2087 11461 2131
rect 11409 2079 11418 2087
rect 11418 2079 11452 2087
rect 11452 2079 11461 2087
rect 11609 2193 11618 2201
rect 11618 2193 11652 2201
rect 11652 2193 11661 2201
rect 11609 2149 11661 2193
rect 11809 2367 11861 2411
rect 11809 2359 11818 2367
rect 11818 2359 11852 2367
rect 11852 2359 11861 2367
rect 12009 2563 12018 2571
rect 12018 2563 12052 2571
rect 12052 2563 12061 2571
rect 12009 2519 12061 2563
rect 12209 2737 12261 2781
rect 12209 2729 12218 2737
rect 12218 2729 12252 2737
rect 12252 2729 12261 2737
rect 12409 2843 12418 2851
rect 12418 2843 12452 2851
rect 12452 2843 12461 2851
rect 12409 2799 12461 2843
rect 12609 3017 12661 3061
rect 12609 3009 12618 3017
rect 12618 3009 12652 3017
rect 12652 3009 12661 3017
rect 12809 3123 12818 3131
rect 12818 3123 12852 3131
rect 12852 3123 12861 3131
rect 12809 3079 12861 3123
rect 12907 3079 12959 3131
rect 12009 2474 12061 2483
rect 12009 2440 12018 2474
rect 12018 2440 12052 2474
rect 12052 2440 12061 2474
rect 12009 2431 12061 2440
rect 10409 1264 10461 1273
rect 10409 1230 10418 1264
rect 10418 1230 10452 1264
rect 10452 1230 10461 1264
rect 10409 1221 10461 1230
rect 8809 54 8861 63
rect 8809 20 8818 54
rect 8818 20 8852 54
rect 8852 20 8861 54
rect 8809 11 8861 20
rect 8709 -60 8761 -15
rect 8709 -67 8718 -60
rect 8718 -67 8752 -60
rect 8752 -67 8761 -60
rect 8509 -166 8518 -143
rect 8518 -166 8552 -143
rect 8552 -166 8561 -143
rect 8509 -195 8561 -166
rect 8525 -248 8577 -239
rect 8525 -282 8534 -248
rect 8534 -282 8568 -248
rect 8568 -282 8577 -248
rect 8525 -291 8577 -282
rect 8509 -363 8561 -326
rect 8509 -378 8518 -363
rect 8518 -378 8552 -363
rect 8552 -378 8561 -363
rect 8509 -397 8518 -390
rect 8518 -397 8552 -390
rect 8552 -397 8561 -390
rect 8509 -435 8561 -397
rect 8509 -442 8518 -435
rect 8518 -442 8552 -435
rect 8552 -442 8561 -435
rect 8509 -469 8518 -454
rect 8518 -469 8552 -454
rect 8552 -469 8561 -454
rect 8509 -506 8561 -469
rect 8709 -94 8718 -79
rect 8718 -94 8752 -79
rect 8752 -94 8761 -79
rect 8709 -131 8761 -94
rect 8809 -74 8861 -22
rect 9009 177 9061 221
rect 9009 169 9018 177
rect 9018 169 9052 177
rect 9052 169 9061 177
rect 9209 283 9218 291
rect 9218 283 9252 291
rect 9252 283 9261 291
rect 9209 239 9261 283
rect 9409 457 9461 501
rect 9409 449 9418 457
rect 9418 449 9452 457
rect 9452 449 9461 457
rect 9609 563 9618 571
rect 9618 563 9652 571
rect 9652 563 9661 571
rect 9609 519 9661 563
rect 9809 737 9861 781
rect 9809 729 9818 737
rect 9818 729 9852 737
rect 9852 729 9861 737
rect 10009 843 10018 851
rect 10018 843 10052 851
rect 10052 843 10061 851
rect 10009 799 10061 843
rect 10209 1017 10261 1061
rect 10209 1009 10218 1017
rect 10218 1009 10252 1017
rect 10252 1009 10261 1017
rect 10409 1123 10418 1131
rect 10418 1123 10452 1131
rect 10452 1123 10461 1131
rect 10409 1079 10461 1123
rect 10609 1387 10661 1431
rect 10609 1379 10618 1387
rect 10618 1379 10652 1387
rect 10652 1379 10661 1387
rect 10809 1493 10818 1501
rect 10818 1493 10852 1501
rect 10852 1493 10861 1501
rect 10809 1449 10861 1493
rect 11009 1667 11061 1711
rect 11009 1659 11018 1667
rect 11018 1659 11052 1667
rect 11052 1659 11061 1667
rect 11209 1773 11218 1781
rect 11218 1773 11252 1781
rect 11252 1773 11261 1781
rect 11209 1729 11261 1773
rect 11409 1947 11461 1991
rect 11409 1939 11418 1947
rect 11418 1939 11452 1947
rect 11452 1939 11461 1947
rect 11609 2053 11618 2061
rect 11618 2053 11652 2061
rect 11652 2053 11661 2061
rect 11609 2009 11661 2053
rect 11809 2227 11861 2271
rect 11809 2219 11818 2227
rect 11818 2219 11852 2227
rect 11852 2219 11861 2227
rect 12009 2333 12018 2341
rect 12018 2333 12052 2341
rect 12052 2333 12061 2341
rect 12009 2289 12061 2333
rect 12209 2597 12261 2641
rect 12209 2589 12218 2597
rect 12218 2589 12252 2597
rect 12252 2589 12261 2597
rect 12409 2703 12418 2711
rect 12418 2703 12452 2711
rect 12452 2703 12461 2711
rect 12409 2659 12461 2703
rect 12609 2877 12661 2921
rect 12609 2869 12618 2877
rect 12618 2869 12652 2877
rect 12652 2869 12661 2877
rect 12809 2983 12818 2991
rect 12818 2983 12852 2991
rect 12852 2983 12861 2991
rect 12809 2939 12861 2983
rect 12907 2939 12959 2991
rect 12209 2490 12261 2499
rect 12209 2456 12218 2490
rect 12218 2456 12252 2490
rect 12252 2456 12261 2490
rect 12209 2447 12261 2456
rect 10609 1280 10661 1289
rect 10609 1246 10618 1280
rect 10618 1246 10652 1280
rect 10652 1246 10661 1280
rect 10609 1237 10661 1246
rect 9009 70 9061 79
rect 9009 36 9018 70
rect 9018 36 9052 70
rect 9052 36 9061 70
rect 9009 27 9061 36
rect 8909 -60 8961 -15
rect 8909 -67 8918 -60
rect 8918 -67 8952 -60
rect 8952 -67 8961 -60
rect 8709 -166 8718 -143
rect 8718 -166 8752 -143
rect 8752 -166 8761 -143
rect 8709 -195 8761 -166
rect 8725 -248 8777 -239
rect 8725 -282 8734 -248
rect 8734 -282 8768 -248
rect 8768 -282 8777 -248
rect 8725 -291 8777 -282
rect 8709 -363 8761 -326
rect 8709 -378 8718 -363
rect 8718 -378 8752 -363
rect 8752 -378 8761 -363
rect 8709 -397 8718 -390
rect 8718 -397 8752 -390
rect 8752 -397 8761 -390
rect 8709 -435 8761 -397
rect 8709 -442 8718 -435
rect 8718 -442 8752 -435
rect 8752 -442 8761 -435
rect 8709 -469 8718 -454
rect 8718 -469 8752 -454
rect 8752 -469 8761 -454
rect 8709 -506 8761 -469
rect 8909 -94 8918 -79
rect 8918 -94 8952 -79
rect 8952 -94 8961 -79
rect 8909 -131 8961 -94
rect 9009 -74 9061 -22
rect 9209 143 9218 151
rect 9218 143 9252 151
rect 9252 143 9261 151
rect 9209 99 9261 143
rect 9409 317 9461 361
rect 9409 309 9418 317
rect 9418 309 9452 317
rect 9452 309 9461 317
rect 9609 423 9618 431
rect 9618 423 9652 431
rect 9652 423 9661 431
rect 9609 379 9661 423
rect 9809 597 9861 641
rect 9809 589 9818 597
rect 9818 589 9852 597
rect 9852 589 9861 597
rect 10009 703 10018 711
rect 10018 703 10052 711
rect 10052 703 10061 711
rect 10009 659 10061 703
rect 10209 877 10261 921
rect 10209 869 10218 877
rect 10218 869 10252 877
rect 10252 869 10261 877
rect 10409 983 10418 991
rect 10418 983 10452 991
rect 10452 983 10461 991
rect 10409 939 10461 983
rect 10609 1157 10661 1201
rect 10609 1149 10618 1157
rect 10618 1149 10652 1157
rect 10652 1149 10661 1157
rect 10809 1353 10818 1361
rect 10818 1353 10852 1361
rect 10852 1353 10861 1361
rect 10809 1309 10861 1353
rect 11009 1527 11061 1571
rect 11009 1519 11018 1527
rect 11018 1519 11052 1527
rect 11052 1519 11061 1527
rect 11209 1633 11218 1641
rect 11218 1633 11252 1641
rect 11252 1633 11261 1641
rect 11209 1589 11261 1633
rect 11409 1807 11461 1851
rect 11409 1799 11418 1807
rect 11418 1799 11452 1807
rect 11452 1799 11461 1807
rect 11609 1913 11618 1921
rect 11618 1913 11652 1921
rect 11652 1913 11661 1921
rect 11609 1869 11661 1913
rect 11809 2087 11861 2131
rect 11809 2079 11818 2087
rect 11818 2079 11852 2087
rect 11852 2079 11861 2087
rect 12009 2193 12018 2201
rect 12018 2193 12052 2201
rect 12052 2193 12061 2201
rect 12009 2149 12061 2193
rect 12209 2367 12261 2411
rect 12209 2359 12218 2367
rect 12218 2359 12252 2367
rect 12252 2359 12261 2367
rect 12409 2563 12418 2571
rect 12418 2563 12452 2571
rect 12452 2563 12461 2571
rect 12409 2519 12461 2563
rect 12609 2737 12661 2781
rect 12609 2729 12618 2737
rect 12618 2729 12652 2737
rect 12652 2729 12661 2737
rect 12809 2843 12818 2851
rect 12818 2843 12852 2851
rect 12852 2843 12861 2851
rect 12809 2799 12861 2843
rect 12907 2799 12959 2851
rect 12409 2474 12461 2483
rect 12409 2440 12418 2474
rect 12418 2440 12452 2474
rect 12452 2440 12461 2474
rect 12409 2431 12461 2440
rect 10809 1264 10861 1273
rect 10809 1230 10818 1264
rect 10818 1230 10852 1264
rect 10852 1230 10861 1264
rect 10809 1221 10861 1230
rect 9209 54 9261 63
rect 9209 20 9218 54
rect 9218 20 9252 54
rect 9252 20 9261 54
rect 9209 11 9261 20
rect 9109 -60 9161 -15
rect 9109 -67 9118 -60
rect 9118 -67 9152 -60
rect 9152 -67 9161 -60
rect 8909 -166 8918 -143
rect 8918 -166 8952 -143
rect 8952 -166 8961 -143
rect 8909 -195 8961 -166
rect 8925 -248 8977 -239
rect 8925 -282 8934 -248
rect 8934 -282 8968 -248
rect 8968 -282 8977 -248
rect 8925 -291 8977 -282
rect 8909 -363 8961 -326
rect 8909 -378 8918 -363
rect 8918 -378 8952 -363
rect 8952 -378 8961 -363
rect 8909 -397 8918 -390
rect 8918 -397 8952 -390
rect 8952 -397 8961 -390
rect 8909 -435 8961 -397
rect 8909 -442 8918 -435
rect 8918 -442 8952 -435
rect 8952 -442 8961 -435
rect 8909 -469 8918 -454
rect 8918 -469 8952 -454
rect 8952 -469 8961 -454
rect 8909 -506 8961 -469
rect 9109 -94 9118 -79
rect 9118 -94 9152 -79
rect 9152 -94 9161 -79
rect 9109 -131 9161 -94
rect 9209 -74 9261 -22
rect 9409 177 9461 221
rect 9409 169 9418 177
rect 9418 169 9452 177
rect 9452 169 9461 177
rect 9609 283 9618 291
rect 9618 283 9652 291
rect 9652 283 9661 291
rect 9609 239 9661 283
rect 9809 457 9861 501
rect 9809 449 9818 457
rect 9818 449 9852 457
rect 9852 449 9861 457
rect 10009 563 10018 571
rect 10018 563 10052 571
rect 10052 563 10061 571
rect 10009 519 10061 563
rect 10209 737 10261 781
rect 10209 729 10218 737
rect 10218 729 10252 737
rect 10252 729 10261 737
rect 10409 843 10418 851
rect 10418 843 10452 851
rect 10452 843 10461 851
rect 10409 799 10461 843
rect 10609 1017 10661 1061
rect 10609 1009 10618 1017
rect 10618 1009 10652 1017
rect 10652 1009 10661 1017
rect 10809 1123 10818 1131
rect 10818 1123 10852 1131
rect 10852 1123 10861 1131
rect 10809 1079 10861 1123
rect 11009 1387 11061 1431
rect 11009 1379 11018 1387
rect 11018 1379 11052 1387
rect 11052 1379 11061 1387
rect 11209 1493 11218 1501
rect 11218 1493 11252 1501
rect 11252 1493 11261 1501
rect 11209 1449 11261 1493
rect 11409 1667 11461 1711
rect 11409 1659 11418 1667
rect 11418 1659 11452 1667
rect 11452 1659 11461 1667
rect 11609 1773 11618 1781
rect 11618 1773 11652 1781
rect 11652 1773 11661 1781
rect 11609 1729 11661 1773
rect 11809 1947 11861 1991
rect 11809 1939 11818 1947
rect 11818 1939 11852 1947
rect 11852 1939 11861 1947
rect 12009 2053 12018 2061
rect 12018 2053 12052 2061
rect 12052 2053 12061 2061
rect 12009 2009 12061 2053
rect 12209 2227 12261 2271
rect 12209 2219 12218 2227
rect 12218 2219 12252 2227
rect 12252 2219 12261 2227
rect 12409 2333 12418 2341
rect 12418 2333 12452 2341
rect 12452 2333 12461 2341
rect 12409 2289 12461 2333
rect 12609 2597 12661 2641
rect 12609 2589 12618 2597
rect 12618 2589 12652 2597
rect 12652 2589 12661 2597
rect 12809 2703 12818 2711
rect 12818 2703 12852 2711
rect 12852 2703 12861 2711
rect 12809 2659 12861 2703
rect 12907 2659 12959 2711
rect 12609 2490 12661 2499
rect 12609 2456 12618 2490
rect 12618 2456 12652 2490
rect 12652 2456 12661 2490
rect 12609 2447 12661 2456
rect 11009 1280 11061 1289
rect 11009 1246 11018 1280
rect 11018 1246 11052 1280
rect 11052 1246 11061 1280
rect 11009 1237 11061 1246
rect 9409 70 9461 79
rect 9409 36 9418 70
rect 9418 36 9452 70
rect 9452 36 9461 70
rect 9409 27 9461 36
rect 9309 -60 9361 -15
rect 9309 -67 9318 -60
rect 9318 -67 9352 -60
rect 9352 -67 9361 -60
rect 9109 -166 9118 -143
rect 9118 -166 9152 -143
rect 9152 -166 9161 -143
rect 9109 -195 9161 -166
rect 9125 -248 9177 -239
rect 9125 -282 9134 -248
rect 9134 -282 9168 -248
rect 9168 -282 9177 -248
rect 9125 -291 9177 -282
rect 9109 -363 9161 -326
rect 9109 -378 9118 -363
rect 9118 -378 9152 -363
rect 9152 -378 9161 -363
rect 9109 -397 9118 -390
rect 9118 -397 9152 -390
rect 9152 -397 9161 -390
rect 9109 -435 9161 -397
rect 9109 -442 9118 -435
rect 9118 -442 9152 -435
rect 9152 -442 9161 -435
rect 9109 -469 9118 -454
rect 9118 -469 9152 -454
rect 9152 -469 9161 -454
rect 9109 -506 9161 -469
rect 9309 -94 9318 -79
rect 9318 -94 9352 -79
rect 9352 -94 9361 -79
rect 9309 -131 9361 -94
rect 9409 -74 9461 -22
rect 9609 143 9618 151
rect 9618 143 9652 151
rect 9652 143 9661 151
rect 9609 99 9661 143
rect 9809 317 9861 361
rect 9809 309 9818 317
rect 9818 309 9852 317
rect 9852 309 9861 317
rect 10009 423 10018 431
rect 10018 423 10052 431
rect 10052 423 10061 431
rect 10009 379 10061 423
rect 10209 597 10261 641
rect 10209 589 10218 597
rect 10218 589 10252 597
rect 10252 589 10261 597
rect 10409 703 10418 711
rect 10418 703 10452 711
rect 10452 703 10461 711
rect 10409 659 10461 703
rect 10609 877 10661 921
rect 10609 869 10618 877
rect 10618 869 10652 877
rect 10652 869 10661 877
rect 10809 983 10818 991
rect 10818 983 10852 991
rect 10852 983 10861 991
rect 10809 939 10861 983
rect 11009 1157 11061 1201
rect 11009 1149 11018 1157
rect 11018 1149 11052 1157
rect 11052 1149 11061 1157
rect 11209 1353 11218 1361
rect 11218 1353 11252 1361
rect 11252 1353 11261 1361
rect 11209 1309 11261 1353
rect 11409 1527 11461 1571
rect 11409 1519 11418 1527
rect 11418 1519 11452 1527
rect 11452 1519 11461 1527
rect 11609 1633 11618 1641
rect 11618 1633 11652 1641
rect 11652 1633 11661 1641
rect 11609 1589 11661 1633
rect 11809 1807 11861 1851
rect 11809 1799 11818 1807
rect 11818 1799 11852 1807
rect 11852 1799 11861 1807
rect 12009 1913 12018 1921
rect 12018 1913 12052 1921
rect 12052 1913 12061 1921
rect 12009 1869 12061 1913
rect 12209 2087 12261 2131
rect 12209 2079 12218 2087
rect 12218 2079 12252 2087
rect 12252 2079 12261 2087
rect 12409 2193 12418 2201
rect 12418 2193 12452 2201
rect 12452 2193 12461 2201
rect 12409 2149 12461 2193
rect 12609 2367 12661 2411
rect 12609 2359 12618 2367
rect 12618 2359 12652 2367
rect 12652 2359 12661 2367
rect 12809 2563 12818 2571
rect 12818 2563 12852 2571
rect 12852 2563 12861 2571
rect 12809 2519 12861 2563
rect 12907 2519 12959 2571
rect 11209 1264 11261 1273
rect 11209 1230 11218 1264
rect 11218 1230 11252 1264
rect 11252 1230 11261 1264
rect 11209 1221 11261 1230
rect 9609 54 9661 63
rect 9609 20 9618 54
rect 9618 20 9652 54
rect 9652 20 9661 54
rect 9609 11 9661 20
rect 9509 -60 9561 -15
rect 9509 -67 9518 -60
rect 9518 -67 9552 -60
rect 9552 -67 9561 -60
rect 9309 -166 9318 -143
rect 9318 -166 9352 -143
rect 9352 -166 9361 -143
rect 9309 -195 9361 -166
rect 9325 -248 9377 -239
rect 9325 -282 9334 -248
rect 9334 -282 9368 -248
rect 9368 -282 9377 -248
rect 9325 -291 9377 -282
rect 9309 -363 9361 -326
rect 9309 -378 9318 -363
rect 9318 -378 9352 -363
rect 9352 -378 9361 -363
rect 9309 -397 9318 -390
rect 9318 -397 9352 -390
rect 9352 -397 9361 -390
rect 9309 -435 9361 -397
rect 9309 -442 9318 -435
rect 9318 -442 9352 -435
rect 9352 -442 9361 -435
rect 9309 -469 9318 -454
rect 9318 -469 9352 -454
rect 9352 -469 9361 -454
rect 9309 -506 9361 -469
rect 9509 -94 9518 -79
rect 9518 -94 9552 -79
rect 9552 -94 9561 -79
rect 9509 -131 9561 -94
rect 9609 -74 9661 -22
rect 9809 177 9861 221
rect 9809 169 9818 177
rect 9818 169 9852 177
rect 9852 169 9861 177
rect 10009 283 10018 291
rect 10018 283 10052 291
rect 10052 283 10061 291
rect 10009 239 10061 283
rect 10209 457 10261 501
rect 10209 449 10218 457
rect 10218 449 10252 457
rect 10252 449 10261 457
rect 10409 563 10418 571
rect 10418 563 10452 571
rect 10452 563 10461 571
rect 10409 519 10461 563
rect 10609 737 10661 781
rect 10609 729 10618 737
rect 10618 729 10652 737
rect 10652 729 10661 737
rect 10809 843 10818 851
rect 10818 843 10852 851
rect 10852 843 10861 851
rect 10809 799 10861 843
rect 11009 1017 11061 1061
rect 11009 1009 11018 1017
rect 11018 1009 11052 1017
rect 11052 1009 11061 1017
rect 11209 1123 11218 1131
rect 11218 1123 11252 1131
rect 11252 1123 11261 1131
rect 11209 1079 11261 1123
rect 11409 1387 11461 1431
rect 11409 1379 11418 1387
rect 11418 1379 11452 1387
rect 11452 1379 11461 1387
rect 11609 1493 11618 1501
rect 11618 1493 11652 1501
rect 11652 1493 11661 1501
rect 11609 1449 11661 1493
rect 11809 1667 11861 1711
rect 11809 1659 11818 1667
rect 11818 1659 11852 1667
rect 11852 1659 11861 1667
rect 12009 1773 12018 1781
rect 12018 1773 12052 1781
rect 12052 1773 12061 1781
rect 12009 1729 12061 1773
rect 12209 1947 12261 1991
rect 12209 1939 12218 1947
rect 12218 1939 12252 1947
rect 12252 1939 12261 1947
rect 12409 2053 12418 2061
rect 12418 2053 12452 2061
rect 12452 2053 12461 2061
rect 12409 2009 12461 2053
rect 12609 2227 12661 2271
rect 12609 2219 12618 2227
rect 12618 2219 12652 2227
rect 12652 2219 12661 2227
rect 12809 2333 12818 2341
rect 12818 2333 12852 2341
rect 12852 2333 12861 2341
rect 12809 2289 12861 2333
rect 12907 2289 12959 2341
rect 11409 1280 11461 1289
rect 11409 1246 11418 1280
rect 11418 1246 11452 1280
rect 11452 1246 11461 1280
rect 11409 1237 11461 1246
rect 9809 70 9861 79
rect 9809 36 9818 70
rect 9818 36 9852 70
rect 9852 36 9861 70
rect 9809 27 9861 36
rect 9709 -60 9761 -15
rect 9709 -67 9718 -60
rect 9718 -67 9752 -60
rect 9752 -67 9761 -60
rect 9509 -166 9518 -143
rect 9518 -166 9552 -143
rect 9552 -166 9561 -143
rect 9509 -195 9561 -166
rect 9525 -248 9577 -239
rect 9525 -282 9534 -248
rect 9534 -282 9568 -248
rect 9568 -282 9577 -248
rect 9525 -291 9577 -282
rect 9509 -363 9561 -326
rect 9509 -378 9518 -363
rect 9518 -378 9552 -363
rect 9552 -378 9561 -363
rect 9509 -397 9518 -390
rect 9518 -397 9552 -390
rect 9552 -397 9561 -390
rect 9509 -435 9561 -397
rect 9509 -442 9518 -435
rect 9518 -442 9552 -435
rect 9552 -442 9561 -435
rect 9509 -469 9518 -454
rect 9518 -469 9552 -454
rect 9552 -469 9561 -454
rect 9509 -506 9561 -469
rect 9709 -94 9718 -79
rect 9718 -94 9752 -79
rect 9752 -94 9761 -79
rect 9709 -131 9761 -94
rect 9809 -74 9861 -22
rect 10009 143 10018 151
rect 10018 143 10052 151
rect 10052 143 10061 151
rect 10009 99 10061 143
rect 10209 317 10261 361
rect 10209 309 10218 317
rect 10218 309 10252 317
rect 10252 309 10261 317
rect 10409 423 10418 431
rect 10418 423 10452 431
rect 10452 423 10461 431
rect 10409 379 10461 423
rect 10609 597 10661 641
rect 10609 589 10618 597
rect 10618 589 10652 597
rect 10652 589 10661 597
rect 10809 703 10818 711
rect 10818 703 10852 711
rect 10852 703 10861 711
rect 10809 659 10861 703
rect 11009 877 11061 921
rect 11009 869 11018 877
rect 11018 869 11052 877
rect 11052 869 11061 877
rect 11209 983 11218 991
rect 11218 983 11252 991
rect 11252 983 11261 991
rect 11209 939 11261 983
rect 11409 1157 11461 1201
rect 11409 1149 11418 1157
rect 11418 1149 11452 1157
rect 11452 1149 11461 1157
rect 11609 1353 11618 1361
rect 11618 1353 11652 1361
rect 11652 1353 11661 1361
rect 11609 1309 11661 1353
rect 11809 1527 11861 1571
rect 11809 1519 11818 1527
rect 11818 1519 11852 1527
rect 11852 1519 11861 1527
rect 12009 1633 12018 1641
rect 12018 1633 12052 1641
rect 12052 1633 12061 1641
rect 12009 1589 12061 1633
rect 12209 1807 12261 1851
rect 12209 1799 12218 1807
rect 12218 1799 12252 1807
rect 12252 1799 12261 1807
rect 12409 1913 12418 1921
rect 12418 1913 12452 1921
rect 12452 1913 12461 1921
rect 12409 1869 12461 1913
rect 12609 2087 12661 2131
rect 12609 2079 12618 2087
rect 12618 2079 12652 2087
rect 12652 2079 12661 2087
rect 12809 2193 12818 2201
rect 12818 2193 12852 2201
rect 12852 2193 12861 2201
rect 12809 2149 12861 2193
rect 12907 2149 12959 2201
rect 11609 1264 11661 1273
rect 11609 1230 11618 1264
rect 11618 1230 11652 1264
rect 11652 1230 11661 1264
rect 11609 1221 11661 1230
rect 10009 54 10061 63
rect 10009 20 10018 54
rect 10018 20 10052 54
rect 10052 20 10061 54
rect 10009 11 10061 20
rect 9909 -60 9961 -15
rect 9909 -67 9918 -60
rect 9918 -67 9952 -60
rect 9952 -67 9961 -60
rect 9709 -166 9718 -143
rect 9718 -166 9752 -143
rect 9752 -166 9761 -143
rect 9709 -195 9761 -166
rect 9725 -248 9777 -239
rect 9725 -282 9734 -248
rect 9734 -282 9768 -248
rect 9768 -282 9777 -248
rect 9725 -291 9777 -282
rect 9709 -363 9761 -326
rect 9709 -378 9718 -363
rect 9718 -378 9752 -363
rect 9752 -378 9761 -363
rect 9709 -397 9718 -390
rect 9718 -397 9752 -390
rect 9752 -397 9761 -390
rect 9709 -435 9761 -397
rect 9709 -442 9718 -435
rect 9718 -442 9752 -435
rect 9752 -442 9761 -435
rect 9709 -469 9718 -454
rect 9718 -469 9752 -454
rect 9752 -469 9761 -454
rect 9709 -506 9761 -469
rect 9909 -94 9918 -79
rect 9918 -94 9952 -79
rect 9952 -94 9961 -79
rect 9909 -131 9961 -94
rect 10009 -74 10061 -22
rect 10209 177 10261 221
rect 10209 169 10218 177
rect 10218 169 10252 177
rect 10252 169 10261 177
rect 10409 283 10418 291
rect 10418 283 10452 291
rect 10452 283 10461 291
rect 10409 239 10461 283
rect 10609 457 10661 501
rect 10609 449 10618 457
rect 10618 449 10652 457
rect 10652 449 10661 457
rect 10809 563 10818 571
rect 10818 563 10852 571
rect 10852 563 10861 571
rect 10809 519 10861 563
rect 11009 737 11061 781
rect 11009 729 11018 737
rect 11018 729 11052 737
rect 11052 729 11061 737
rect 11209 843 11218 851
rect 11218 843 11252 851
rect 11252 843 11261 851
rect 11209 799 11261 843
rect 11409 1017 11461 1061
rect 11409 1009 11418 1017
rect 11418 1009 11452 1017
rect 11452 1009 11461 1017
rect 11609 1123 11618 1131
rect 11618 1123 11652 1131
rect 11652 1123 11661 1131
rect 11609 1079 11661 1123
rect 11809 1387 11861 1431
rect 11809 1379 11818 1387
rect 11818 1379 11852 1387
rect 11852 1379 11861 1387
rect 12009 1493 12018 1501
rect 12018 1493 12052 1501
rect 12052 1493 12061 1501
rect 12009 1449 12061 1493
rect 12209 1667 12261 1711
rect 12209 1659 12218 1667
rect 12218 1659 12252 1667
rect 12252 1659 12261 1667
rect 12409 1773 12418 1781
rect 12418 1773 12452 1781
rect 12452 1773 12461 1781
rect 12409 1729 12461 1773
rect 12609 1947 12661 1991
rect 12609 1939 12618 1947
rect 12618 1939 12652 1947
rect 12652 1939 12661 1947
rect 12809 2053 12818 2061
rect 12818 2053 12852 2061
rect 12852 2053 12861 2061
rect 12809 2009 12861 2053
rect 12907 2009 12959 2061
rect 11809 1280 11861 1289
rect 11809 1246 11818 1280
rect 11818 1246 11852 1280
rect 11852 1246 11861 1280
rect 11809 1237 11861 1246
rect 10209 70 10261 79
rect 10209 36 10218 70
rect 10218 36 10252 70
rect 10252 36 10261 70
rect 10209 27 10261 36
rect 10109 -60 10161 -15
rect 10109 -67 10118 -60
rect 10118 -67 10152 -60
rect 10152 -67 10161 -60
rect 9909 -166 9918 -143
rect 9918 -166 9952 -143
rect 9952 -166 9961 -143
rect 9909 -195 9961 -166
rect 9925 -248 9977 -239
rect 9925 -282 9934 -248
rect 9934 -282 9968 -248
rect 9968 -282 9977 -248
rect 9925 -291 9977 -282
rect 9909 -363 9961 -326
rect 9909 -378 9918 -363
rect 9918 -378 9952 -363
rect 9952 -378 9961 -363
rect 9909 -397 9918 -390
rect 9918 -397 9952 -390
rect 9952 -397 9961 -390
rect 9909 -435 9961 -397
rect 9909 -442 9918 -435
rect 9918 -442 9952 -435
rect 9952 -442 9961 -435
rect 9909 -469 9918 -454
rect 9918 -469 9952 -454
rect 9952 -469 9961 -454
rect 9909 -506 9961 -469
rect 10109 -94 10118 -79
rect 10118 -94 10152 -79
rect 10152 -94 10161 -79
rect 10109 -131 10161 -94
rect 10209 -74 10261 -22
rect 10409 143 10418 151
rect 10418 143 10452 151
rect 10452 143 10461 151
rect 10409 99 10461 143
rect 10609 317 10661 361
rect 10609 309 10618 317
rect 10618 309 10652 317
rect 10652 309 10661 317
rect 10809 423 10818 431
rect 10818 423 10852 431
rect 10852 423 10861 431
rect 10809 379 10861 423
rect 11009 597 11061 641
rect 11009 589 11018 597
rect 11018 589 11052 597
rect 11052 589 11061 597
rect 11209 703 11218 711
rect 11218 703 11252 711
rect 11252 703 11261 711
rect 11209 659 11261 703
rect 11409 877 11461 921
rect 11409 869 11418 877
rect 11418 869 11452 877
rect 11452 869 11461 877
rect 11609 983 11618 991
rect 11618 983 11652 991
rect 11652 983 11661 991
rect 11609 939 11661 983
rect 11809 1157 11861 1201
rect 11809 1149 11818 1157
rect 11818 1149 11852 1157
rect 11852 1149 11861 1157
rect 12009 1353 12018 1361
rect 12018 1353 12052 1361
rect 12052 1353 12061 1361
rect 12009 1309 12061 1353
rect 12209 1527 12261 1571
rect 12209 1519 12218 1527
rect 12218 1519 12252 1527
rect 12252 1519 12261 1527
rect 12409 1633 12418 1641
rect 12418 1633 12452 1641
rect 12452 1633 12461 1641
rect 12409 1589 12461 1633
rect 12609 1807 12661 1851
rect 12609 1799 12618 1807
rect 12618 1799 12652 1807
rect 12652 1799 12661 1807
rect 12809 1913 12818 1921
rect 12818 1913 12852 1921
rect 12852 1913 12861 1921
rect 12809 1869 12861 1913
rect 12907 1869 12959 1921
rect 12009 1264 12061 1273
rect 12009 1230 12018 1264
rect 12018 1230 12052 1264
rect 12052 1230 12061 1264
rect 12009 1221 12061 1230
rect 10409 54 10461 63
rect 10409 20 10418 54
rect 10418 20 10452 54
rect 10452 20 10461 54
rect 10409 11 10461 20
rect 10309 -60 10361 -15
rect 10309 -67 10318 -60
rect 10318 -67 10352 -60
rect 10352 -67 10361 -60
rect 10109 -166 10118 -143
rect 10118 -166 10152 -143
rect 10152 -166 10161 -143
rect 10109 -195 10161 -166
rect 10125 -248 10177 -239
rect 10125 -282 10134 -248
rect 10134 -282 10168 -248
rect 10168 -282 10177 -248
rect 10125 -291 10177 -282
rect 10109 -363 10161 -326
rect 10109 -378 10118 -363
rect 10118 -378 10152 -363
rect 10152 -378 10161 -363
rect 10109 -397 10118 -390
rect 10118 -397 10152 -390
rect 10152 -397 10161 -390
rect 10109 -435 10161 -397
rect 10109 -442 10118 -435
rect 10118 -442 10152 -435
rect 10152 -442 10161 -435
rect 10109 -469 10118 -454
rect 10118 -469 10152 -454
rect 10152 -469 10161 -454
rect 10109 -506 10161 -469
rect 10309 -94 10318 -79
rect 10318 -94 10352 -79
rect 10352 -94 10361 -79
rect 10309 -131 10361 -94
rect 10409 -74 10461 -22
rect 10609 177 10661 221
rect 10609 169 10618 177
rect 10618 169 10652 177
rect 10652 169 10661 177
rect 10809 283 10818 291
rect 10818 283 10852 291
rect 10852 283 10861 291
rect 10809 239 10861 283
rect 11009 457 11061 501
rect 11009 449 11018 457
rect 11018 449 11052 457
rect 11052 449 11061 457
rect 11209 563 11218 571
rect 11218 563 11252 571
rect 11252 563 11261 571
rect 11209 519 11261 563
rect 11409 737 11461 781
rect 11409 729 11418 737
rect 11418 729 11452 737
rect 11452 729 11461 737
rect 11609 843 11618 851
rect 11618 843 11652 851
rect 11652 843 11661 851
rect 11609 799 11661 843
rect 11809 1017 11861 1061
rect 11809 1009 11818 1017
rect 11818 1009 11852 1017
rect 11852 1009 11861 1017
rect 12009 1123 12018 1131
rect 12018 1123 12052 1131
rect 12052 1123 12061 1131
rect 12009 1079 12061 1123
rect 12209 1387 12261 1431
rect 12209 1379 12218 1387
rect 12218 1379 12252 1387
rect 12252 1379 12261 1387
rect 12409 1493 12418 1501
rect 12418 1493 12452 1501
rect 12452 1493 12461 1501
rect 12409 1449 12461 1493
rect 12609 1667 12661 1711
rect 12609 1659 12618 1667
rect 12618 1659 12652 1667
rect 12652 1659 12661 1667
rect 12809 1773 12818 1781
rect 12818 1773 12852 1781
rect 12852 1773 12861 1781
rect 12809 1729 12861 1773
rect 12907 1729 12959 1781
rect 12209 1280 12261 1289
rect 12209 1246 12218 1280
rect 12218 1246 12252 1280
rect 12252 1246 12261 1280
rect 12209 1237 12261 1246
rect 10609 70 10661 79
rect 10609 36 10618 70
rect 10618 36 10652 70
rect 10652 36 10661 70
rect 10609 27 10661 36
rect 10509 -60 10561 -15
rect 10509 -67 10518 -60
rect 10518 -67 10552 -60
rect 10552 -67 10561 -60
rect 10309 -166 10318 -143
rect 10318 -166 10352 -143
rect 10352 -166 10361 -143
rect 10309 -195 10361 -166
rect 10325 -248 10377 -239
rect 10325 -282 10334 -248
rect 10334 -282 10368 -248
rect 10368 -282 10377 -248
rect 10325 -291 10377 -282
rect 10309 -363 10361 -326
rect 10309 -378 10318 -363
rect 10318 -378 10352 -363
rect 10352 -378 10361 -363
rect 10309 -397 10318 -390
rect 10318 -397 10352 -390
rect 10352 -397 10361 -390
rect 10309 -435 10361 -397
rect 10309 -442 10318 -435
rect 10318 -442 10352 -435
rect 10352 -442 10361 -435
rect 10309 -469 10318 -454
rect 10318 -469 10352 -454
rect 10352 -469 10361 -454
rect 10309 -506 10361 -469
rect 10509 -94 10518 -79
rect 10518 -94 10552 -79
rect 10552 -94 10561 -79
rect 10509 -131 10561 -94
rect 10609 -74 10661 -22
rect 10809 143 10818 151
rect 10818 143 10852 151
rect 10852 143 10861 151
rect 10809 99 10861 143
rect 11009 317 11061 361
rect 11009 309 11018 317
rect 11018 309 11052 317
rect 11052 309 11061 317
rect 11209 423 11218 431
rect 11218 423 11252 431
rect 11252 423 11261 431
rect 11209 379 11261 423
rect 11409 597 11461 641
rect 11409 589 11418 597
rect 11418 589 11452 597
rect 11452 589 11461 597
rect 11609 703 11618 711
rect 11618 703 11652 711
rect 11652 703 11661 711
rect 11609 659 11661 703
rect 11809 877 11861 921
rect 11809 869 11818 877
rect 11818 869 11852 877
rect 11852 869 11861 877
rect 12009 983 12018 991
rect 12018 983 12052 991
rect 12052 983 12061 991
rect 12009 939 12061 983
rect 12209 1157 12261 1201
rect 12209 1149 12218 1157
rect 12218 1149 12252 1157
rect 12252 1149 12261 1157
rect 12409 1353 12418 1361
rect 12418 1353 12452 1361
rect 12452 1353 12461 1361
rect 12409 1309 12461 1353
rect 12609 1527 12661 1571
rect 12609 1519 12618 1527
rect 12618 1519 12652 1527
rect 12652 1519 12661 1527
rect 12809 1633 12818 1641
rect 12818 1633 12852 1641
rect 12852 1633 12861 1641
rect 12809 1589 12861 1633
rect 12907 1589 12959 1641
rect 12409 1264 12461 1273
rect 12409 1230 12418 1264
rect 12418 1230 12452 1264
rect 12452 1230 12461 1264
rect 12409 1221 12461 1230
rect 10809 54 10861 63
rect 10809 20 10818 54
rect 10818 20 10852 54
rect 10852 20 10861 54
rect 10809 11 10861 20
rect 10709 -60 10761 -15
rect 10709 -67 10718 -60
rect 10718 -67 10752 -60
rect 10752 -67 10761 -60
rect 10509 -166 10518 -143
rect 10518 -166 10552 -143
rect 10552 -166 10561 -143
rect 10509 -195 10561 -166
rect 10525 -248 10577 -239
rect 10525 -282 10534 -248
rect 10534 -282 10568 -248
rect 10568 -282 10577 -248
rect 10525 -291 10577 -282
rect 10509 -363 10561 -326
rect 10509 -378 10518 -363
rect 10518 -378 10552 -363
rect 10552 -378 10561 -363
rect 10509 -397 10518 -390
rect 10518 -397 10552 -390
rect 10552 -397 10561 -390
rect 10509 -435 10561 -397
rect 10509 -442 10518 -435
rect 10518 -442 10552 -435
rect 10552 -442 10561 -435
rect 10509 -469 10518 -454
rect 10518 -469 10552 -454
rect 10552 -469 10561 -454
rect 10509 -506 10561 -469
rect 10709 -94 10718 -79
rect 10718 -94 10752 -79
rect 10752 -94 10761 -79
rect 10709 -131 10761 -94
rect 10809 -74 10861 -22
rect 11009 177 11061 221
rect 11009 169 11018 177
rect 11018 169 11052 177
rect 11052 169 11061 177
rect 11209 283 11218 291
rect 11218 283 11252 291
rect 11252 283 11261 291
rect 11209 239 11261 283
rect 11409 457 11461 501
rect 11409 449 11418 457
rect 11418 449 11452 457
rect 11452 449 11461 457
rect 11609 563 11618 571
rect 11618 563 11652 571
rect 11652 563 11661 571
rect 11609 519 11661 563
rect 11809 737 11861 781
rect 11809 729 11818 737
rect 11818 729 11852 737
rect 11852 729 11861 737
rect 12009 843 12018 851
rect 12018 843 12052 851
rect 12052 843 12061 851
rect 12009 799 12061 843
rect 12209 1017 12261 1061
rect 12209 1009 12218 1017
rect 12218 1009 12252 1017
rect 12252 1009 12261 1017
rect 12409 1123 12418 1131
rect 12418 1123 12452 1131
rect 12452 1123 12461 1131
rect 12409 1079 12461 1123
rect 12609 1387 12661 1431
rect 12609 1379 12618 1387
rect 12618 1379 12652 1387
rect 12652 1379 12661 1387
rect 12809 1493 12818 1501
rect 12818 1493 12852 1501
rect 12852 1493 12861 1501
rect 12809 1449 12861 1493
rect 12907 1449 12959 1501
rect 12609 1280 12661 1289
rect 12609 1246 12618 1280
rect 12618 1246 12652 1280
rect 12652 1246 12661 1280
rect 12609 1237 12661 1246
rect 11009 70 11061 79
rect 11009 36 11018 70
rect 11018 36 11052 70
rect 11052 36 11061 70
rect 11009 27 11061 36
rect 10909 -60 10961 -15
rect 10909 -67 10918 -60
rect 10918 -67 10952 -60
rect 10952 -67 10961 -60
rect 10709 -166 10718 -143
rect 10718 -166 10752 -143
rect 10752 -166 10761 -143
rect 10709 -195 10761 -166
rect 10725 -248 10777 -239
rect 10725 -282 10734 -248
rect 10734 -282 10768 -248
rect 10768 -282 10777 -248
rect 10725 -291 10777 -282
rect 10709 -363 10761 -326
rect 10709 -378 10718 -363
rect 10718 -378 10752 -363
rect 10752 -378 10761 -363
rect 10709 -397 10718 -390
rect 10718 -397 10752 -390
rect 10752 -397 10761 -390
rect 10709 -435 10761 -397
rect 10709 -442 10718 -435
rect 10718 -442 10752 -435
rect 10752 -442 10761 -435
rect 10709 -469 10718 -454
rect 10718 -469 10752 -454
rect 10752 -469 10761 -454
rect 10709 -506 10761 -469
rect 10909 -94 10918 -79
rect 10918 -94 10952 -79
rect 10952 -94 10961 -79
rect 10909 -131 10961 -94
rect 11009 -74 11061 -22
rect 11209 143 11218 151
rect 11218 143 11252 151
rect 11252 143 11261 151
rect 11209 99 11261 143
rect 11409 317 11461 361
rect 11409 309 11418 317
rect 11418 309 11452 317
rect 11452 309 11461 317
rect 11609 423 11618 431
rect 11618 423 11652 431
rect 11652 423 11661 431
rect 11609 379 11661 423
rect 11809 597 11861 641
rect 11809 589 11818 597
rect 11818 589 11852 597
rect 11852 589 11861 597
rect 12009 703 12018 711
rect 12018 703 12052 711
rect 12052 703 12061 711
rect 12009 659 12061 703
rect 12209 877 12261 921
rect 12209 869 12218 877
rect 12218 869 12252 877
rect 12252 869 12261 877
rect 12409 983 12418 991
rect 12418 983 12452 991
rect 12452 983 12461 991
rect 12409 939 12461 983
rect 12609 1157 12661 1201
rect 12609 1149 12618 1157
rect 12618 1149 12652 1157
rect 12652 1149 12661 1157
rect 12809 1353 12818 1361
rect 12818 1353 12852 1361
rect 12852 1353 12861 1361
rect 12809 1309 12861 1353
rect 12907 1309 12959 1361
rect 11209 54 11261 63
rect 11209 20 11218 54
rect 11218 20 11252 54
rect 11252 20 11261 54
rect 11209 11 11261 20
rect 11109 -60 11161 -15
rect 11109 -67 11118 -60
rect 11118 -67 11152 -60
rect 11152 -67 11161 -60
rect 10909 -166 10918 -143
rect 10918 -166 10952 -143
rect 10952 -166 10961 -143
rect 10909 -195 10961 -166
rect 10925 -248 10977 -239
rect 10925 -282 10934 -248
rect 10934 -282 10968 -248
rect 10968 -282 10977 -248
rect 10925 -291 10977 -282
rect 10909 -363 10961 -326
rect 10909 -378 10918 -363
rect 10918 -378 10952 -363
rect 10952 -378 10961 -363
rect 10909 -397 10918 -390
rect 10918 -397 10952 -390
rect 10952 -397 10961 -390
rect 10909 -435 10961 -397
rect 10909 -442 10918 -435
rect 10918 -442 10952 -435
rect 10952 -442 10961 -435
rect 10909 -469 10918 -454
rect 10918 -469 10952 -454
rect 10952 -469 10961 -454
rect 10909 -506 10961 -469
rect 11109 -94 11118 -79
rect 11118 -94 11152 -79
rect 11152 -94 11161 -79
rect 11109 -131 11161 -94
rect 11209 -74 11261 -22
rect 11409 177 11461 221
rect 11409 169 11418 177
rect 11418 169 11452 177
rect 11452 169 11461 177
rect 11609 283 11618 291
rect 11618 283 11652 291
rect 11652 283 11661 291
rect 11609 239 11661 283
rect 11809 457 11861 501
rect 11809 449 11818 457
rect 11818 449 11852 457
rect 11852 449 11861 457
rect 12009 563 12018 571
rect 12018 563 12052 571
rect 12052 563 12061 571
rect 12009 519 12061 563
rect 12209 737 12261 781
rect 12209 729 12218 737
rect 12218 729 12252 737
rect 12252 729 12261 737
rect 12409 843 12418 851
rect 12418 843 12452 851
rect 12452 843 12461 851
rect 12409 799 12461 843
rect 12609 1017 12661 1061
rect 12609 1009 12618 1017
rect 12618 1009 12652 1017
rect 12652 1009 12661 1017
rect 12809 1123 12818 1131
rect 12818 1123 12852 1131
rect 12852 1123 12861 1131
rect 12809 1079 12861 1123
rect 12907 1079 12959 1131
rect 11409 70 11461 79
rect 11409 36 11418 70
rect 11418 36 11452 70
rect 11452 36 11461 70
rect 11409 27 11461 36
rect 11309 -60 11361 -15
rect 11309 -67 11318 -60
rect 11318 -67 11352 -60
rect 11352 -67 11361 -60
rect 11109 -166 11118 -143
rect 11118 -166 11152 -143
rect 11152 -166 11161 -143
rect 11109 -195 11161 -166
rect 11125 -248 11177 -239
rect 11125 -282 11134 -248
rect 11134 -282 11168 -248
rect 11168 -282 11177 -248
rect 11125 -291 11177 -282
rect 11109 -363 11161 -326
rect 11109 -378 11118 -363
rect 11118 -378 11152 -363
rect 11152 -378 11161 -363
rect 11109 -397 11118 -390
rect 11118 -397 11152 -390
rect 11152 -397 11161 -390
rect 11109 -435 11161 -397
rect 11109 -442 11118 -435
rect 11118 -442 11152 -435
rect 11152 -442 11161 -435
rect 11109 -469 11118 -454
rect 11118 -469 11152 -454
rect 11152 -469 11161 -454
rect 11109 -506 11161 -469
rect 11309 -94 11318 -79
rect 11318 -94 11352 -79
rect 11352 -94 11361 -79
rect 11309 -131 11361 -94
rect 11409 -74 11461 -22
rect 11609 143 11618 151
rect 11618 143 11652 151
rect 11652 143 11661 151
rect 11609 99 11661 143
rect 11809 317 11861 361
rect 11809 309 11818 317
rect 11818 309 11852 317
rect 11852 309 11861 317
rect 12009 423 12018 431
rect 12018 423 12052 431
rect 12052 423 12061 431
rect 12009 379 12061 423
rect 12209 597 12261 641
rect 12209 589 12218 597
rect 12218 589 12252 597
rect 12252 589 12261 597
rect 12409 703 12418 711
rect 12418 703 12452 711
rect 12452 703 12461 711
rect 12409 659 12461 703
rect 12609 877 12661 921
rect 12609 869 12618 877
rect 12618 869 12652 877
rect 12652 869 12661 877
rect 12809 983 12818 991
rect 12818 983 12852 991
rect 12852 983 12861 991
rect 12809 939 12861 983
rect 12907 939 12959 991
rect 11609 54 11661 63
rect 11609 20 11618 54
rect 11618 20 11652 54
rect 11652 20 11661 54
rect 11609 11 11661 20
rect 11509 -60 11561 -15
rect 11509 -67 11518 -60
rect 11518 -67 11552 -60
rect 11552 -67 11561 -60
rect 11309 -166 11318 -143
rect 11318 -166 11352 -143
rect 11352 -166 11361 -143
rect 11309 -195 11361 -166
rect 11325 -248 11377 -239
rect 11325 -282 11334 -248
rect 11334 -282 11368 -248
rect 11368 -282 11377 -248
rect 11325 -291 11377 -282
rect 11309 -363 11361 -326
rect 11309 -378 11318 -363
rect 11318 -378 11352 -363
rect 11352 -378 11361 -363
rect 11309 -397 11318 -390
rect 11318 -397 11352 -390
rect 11352 -397 11361 -390
rect 11309 -435 11361 -397
rect 11309 -442 11318 -435
rect 11318 -442 11352 -435
rect 11352 -442 11361 -435
rect 11309 -469 11318 -454
rect 11318 -469 11352 -454
rect 11352 -469 11361 -454
rect 11309 -506 11361 -469
rect 11509 -94 11518 -79
rect 11518 -94 11552 -79
rect 11552 -94 11561 -79
rect 11509 -131 11561 -94
rect 11609 -74 11661 -22
rect 11809 177 11861 221
rect 11809 169 11818 177
rect 11818 169 11852 177
rect 11852 169 11861 177
rect 12009 283 12018 291
rect 12018 283 12052 291
rect 12052 283 12061 291
rect 12009 239 12061 283
rect 12209 457 12261 501
rect 12209 449 12218 457
rect 12218 449 12252 457
rect 12252 449 12261 457
rect 12409 563 12418 571
rect 12418 563 12452 571
rect 12452 563 12461 571
rect 12409 519 12461 563
rect 12609 737 12661 781
rect 12609 729 12618 737
rect 12618 729 12652 737
rect 12652 729 12661 737
rect 12809 843 12818 851
rect 12818 843 12852 851
rect 12852 843 12861 851
rect 12809 799 12861 843
rect 12907 799 12959 851
rect 11809 70 11861 79
rect 11809 36 11818 70
rect 11818 36 11852 70
rect 11852 36 11861 70
rect 11809 27 11861 36
rect 11709 -60 11761 -15
rect 11709 -67 11718 -60
rect 11718 -67 11752 -60
rect 11752 -67 11761 -60
rect 11509 -166 11518 -143
rect 11518 -166 11552 -143
rect 11552 -166 11561 -143
rect 11509 -195 11561 -166
rect 11525 -248 11577 -239
rect 11525 -282 11534 -248
rect 11534 -282 11568 -248
rect 11568 -282 11577 -248
rect 11525 -291 11577 -282
rect 11509 -363 11561 -326
rect 11509 -378 11518 -363
rect 11518 -378 11552 -363
rect 11552 -378 11561 -363
rect 11509 -397 11518 -390
rect 11518 -397 11552 -390
rect 11552 -397 11561 -390
rect 11509 -435 11561 -397
rect 11509 -442 11518 -435
rect 11518 -442 11552 -435
rect 11552 -442 11561 -435
rect 11509 -469 11518 -454
rect 11518 -469 11552 -454
rect 11552 -469 11561 -454
rect 11509 -506 11561 -469
rect 11709 -94 11718 -79
rect 11718 -94 11752 -79
rect 11752 -94 11761 -79
rect 11709 -131 11761 -94
rect 11809 -74 11861 -22
rect 12009 143 12018 151
rect 12018 143 12052 151
rect 12052 143 12061 151
rect 12009 99 12061 143
rect 12209 317 12261 361
rect 12209 309 12218 317
rect 12218 309 12252 317
rect 12252 309 12261 317
rect 12409 423 12418 431
rect 12418 423 12452 431
rect 12452 423 12461 431
rect 12409 379 12461 423
rect 12609 597 12661 641
rect 12609 589 12618 597
rect 12618 589 12652 597
rect 12652 589 12661 597
rect 12809 703 12818 711
rect 12818 703 12852 711
rect 12852 703 12861 711
rect 12809 659 12861 703
rect 12907 659 12959 711
rect 12009 54 12061 63
rect 12009 20 12018 54
rect 12018 20 12052 54
rect 12052 20 12061 54
rect 12009 11 12061 20
rect 11909 -60 11961 -15
rect 11909 -67 11918 -60
rect 11918 -67 11952 -60
rect 11952 -67 11961 -60
rect 11709 -166 11718 -143
rect 11718 -166 11752 -143
rect 11752 -166 11761 -143
rect 11709 -195 11761 -166
rect 11725 -248 11777 -239
rect 11725 -282 11734 -248
rect 11734 -282 11768 -248
rect 11768 -282 11777 -248
rect 11725 -291 11777 -282
rect 11709 -363 11761 -326
rect 11709 -378 11718 -363
rect 11718 -378 11752 -363
rect 11752 -378 11761 -363
rect 11709 -397 11718 -390
rect 11718 -397 11752 -390
rect 11752 -397 11761 -390
rect 11709 -435 11761 -397
rect 11709 -442 11718 -435
rect 11718 -442 11752 -435
rect 11752 -442 11761 -435
rect 11709 -469 11718 -454
rect 11718 -469 11752 -454
rect 11752 -469 11761 -454
rect 11709 -506 11761 -469
rect 11909 -94 11918 -79
rect 11918 -94 11952 -79
rect 11952 -94 11961 -79
rect 11909 -131 11961 -94
rect 12009 -74 12061 -22
rect 12209 177 12261 221
rect 12209 169 12218 177
rect 12218 169 12252 177
rect 12252 169 12261 177
rect 12409 283 12418 291
rect 12418 283 12452 291
rect 12452 283 12461 291
rect 12409 239 12461 283
rect 12609 457 12661 501
rect 12609 449 12618 457
rect 12618 449 12652 457
rect 12652 449 12661 457
rect 12809 563 12818 571
rect 12818 563 12852 571
rect 12852 563 12861 571
rect 12809 519 12861 563
rect 12907 519 12959 571
rect 12209 70 12261 79
rect 12209 36 12218 70
rect 12218 36 12252 70
rect 12252 36 12261 70
rect 12209 27 12261 36
rect 12109 -60 12161 -15
rect 12109 -67 12118 -60
rect 12118 -67 12152 -60
rect 12152 -67 12161 -60
rect 11909 -166 11918 -143
rect 11918 -166 11952 -143
rect 11952 -166 11961 -143
rect 11909 -195 11961 -166
rect 11925 -248 11977 -239
rect 11925 -282 11934 -248
rect 11934 -282 11968 -248
rect 11968 -282 11977 -248
rect 11925 -291 11977 -282
rect 11909 -363 11961 -326
rect 11909 -378 11918 -363
rect 11918 -378 11952 -363
rect 11952 -378 11961 -363
rect 11909 -397 11918 -390
rect 11918 -397 11952 -390
rect 11952 -397 11961 -390
rect 11909 -435 11961 -397
rect 11909 -442 11918 -435
rect 11918 -442 11952 -435
rect 11952 -442 11961 -435
rect 11909 -469 11918 -454
rect 11918 -469 11952 -454
rect 11952 -469 11961 -454
rect 11909 -506 11961 -469
rect 12109 -94 12118 -79
rect 12118 -94 12152 -79
rect 12152 -94 12161 -79
rect 12109 -131 12161 -94
rect 12209 -74 12261 -22
rect 12409 143 12418 151
rect 12418 143 12452 151
rect 12452 143 12461 151
rect 12409 99 12461 143
rect 12609 317 12661 361
rect 12609 309 12618 317
rect 12618 309 12652 317
rect 12652 309 12661 317
rect 12809 423 12818 431
rect 12818 423 12852 431
rect 12852 423 12861 431
rect 12809 379 12861 423
rect 12907 379 12959 431
rect 12409 54 12461 63
rect 12409 20 12418 54
rect 12418 20 12452 54
rect 12452 20 12461 54
rect 12409 11 12461 20
rect 12309 -60 12361 -15
rect 12309 -67 12318 -60
rect 12318 -67 12352 -60
rect 12352 -67 12361 -60
rect 12109 -166 12118 -143
rect 12118 -166 12152 -143
rect 12152 -166 12161 -143
rect 12109 -195 12161 -166
rect 12125 -248 12177 -239
rect 12125 -282 12134 -248
rect 12134 -282 12168 -248
rect 12168 -282 12177 -248
rect 12125 -291 12177 -282
rect 12109 -363 12161 -326
rect 12109 -378 12118 -363
rect 12118 -378 12152 -363
rect 12152 -378 12161 -363
rect 12109 -397 12118 -390
rect 12118 -397 12152 -390
rect 12152 -397 12161 -390
rect 12109 -435 12161 -397
rect 12109 -442 12118 -435
rect 12118 -442 12152 -435
rect 12152 -442 12161 -435
rect 12109 -469 12118 -454
rect 12118 -469 12152 -454
rect 12152 -469 12161 -454
rect 12109 -506 12161 -469
rect 12309 -94 12318 -79
rect 12318 -94 12352 -79
rect 12352 -94 12361 -79
rect 12309 -131 12361 -94
rect 12409 -74 12461 -22
rect 12609 177 12661 221
rect 12609 169 12618 177
rect 12618 169 12652 177
rect 12652 169 12661 177
rect 12809 283 12818 291
rect 12818 283 12852 291
rect 12852 283 12861 291
rect 12809 239 12861 283
rect 12907 239 12959 291
rect 12609 70 12661 79
rect 12609 36 12618 70
rect 12618 36 12652 70
rect 12652 36 12661 70
rect 12609 27 12661 36
rect 12509 -60 12561 -15
rect 12509 -67 12518 -60
rect 12518 -67 12552 -60
rect 12552 -67 12561 -60
rect 12309 -166 12318 -143
rect 12318 -166 12352 -143
rect 12352 -166 12361 -143
rect 12309 -195 12361 -166
rect 12325 -248 12377 -239
rect 12325 -282 12334 -248
rect 12334 -282 12368 -248
rect 12368 -282 12377 -248
rect 12325 -291 12377 -282
rect 12309 -363 12361 -326
rect 12309 -378 12318 -363
rect 12318 -378 12352 -363
rect 12352 -378 12361 -363
rect 12309 -397 12318 -390
rect 12318 -397 12352 -390
rect 12352 -397 12361 -390
rect 12309 -435 12361 -397
rect 12309 -442 12318 -435
rect 12318 -442 12352 -435
rect 12352 -442 12361 -435
rect 12309 -469 12318 -454
rect 12318 -469 12352 -454
rect 12352 -469 12361 -454
rect 12309 -506 12361 -469
rect 12509 -94 12518 -79
rect 12518 -94 12552 -79
rect 12552 -94 12561 -79
rect 12509 -131 12561 -94
rect 12609 -74 12661 -22
rect 12809 143 12818 151
rect 12818 143 12852 151
rect 12852 143 12861 151
rect 12809 99 12861 143
rect 12907 99 12959 151
rect 13111 4779 13163 4831
rect 13111 4639 13163 4691
rect 13111 4499 13163 4551
rect 13111 4359 13163 4411
rect 13111 4219 13163 4271
rect 13111 4079 13163 4131
rect 13111 3939 13163 3991
rect 13111 3799 13163 3851
rect 13111 3569 13163 3621
rect 13111 3429 13163 3481
rect 13111 3289 13163 3341
rect 13111 3149 13163 3201
rect 13111 3009 13163 3061
rect 13111 2869 13163 2921
rect 13111 2729 13163 2781
rect 13111 2589 13163 2641
rect 13111 2359 13163 2411
rect 13111 2219 13163 2271
rect 13111 2079 13163 2131
rect 13111 1939 13163 1991
rect 13111 1799 13163 1851
rect 13111 1659 13163 1711
rect 13111 1519 13163 1571
rect 13111 1379 13163 1431
rect 13111 1149 13163 1201
rect 13111 1009 13163 1061
rect 13111 869 13163 921
rect 13111 729 13163 781
rect 13111 589 13163 641
rect 13111 449 13163 501
rect 13111 309 13163 361
rect 13111 169 13163 221
rect 12709 -60 12761 -15
rect 12709 -67 12718 -60
rect 12718 -67 12752 -60
rect 12752 -67 12761 -60
rect 12509 -166 12518 -143
rect 12518 -166 12552 -143
rect 12552 -166 12561 -143
rect 12509 -195 12561 -166
rect 12525 -248 12577 -239
rect 12525 -282 12534 -248
rect 12534 -282 12568 -248
rect 12568 -282 12577 -248
rect 12525 -291 12577 -282
rect 12509 -363 12561 -326
rect 12509 -378 12518 -363
rect 12518 -378 12552 -363
rect 12552 -378 12561 -363
rect 12509 -397 12518 -390
rect 12518 -397 12552 -390
rect 12552 -397 12561 -390
rect 12509 -435 12561 -397
rect 12509 -442 12518 -435
rect 12518 -442 12552 -435
rect 12552 -442 12561 -435
rect 12509 -469 12518 -454
rect 12518 -469 12552 -454
rect 12552 -469 12561 -454
rect 12509 -506 12561 -469
rect 12709 -94 12718 -79
rect 12718 -94 12752 -79
rect 12752 -94 12761 -79
rect 12709 -131 12761 -94
rect 12709 -166 12718 -143
rect 12718 -166 12752 -143
rect 12752 -166 12761 -143
rect 12709 -195 12761 -166
rect 14553 -208 14605 -199
rect 14553 -242 14558 -208
rect 14558 -242 14592 -208
rect 14592 -242 14605 -208
rect 14553 -251 14605 -242
rect 14617 -208 14669 -199
rect 14617 -242 14630 -208
rect 14630 -242 14664 -208
rect 14664 -242 14669 -208
rect 14617 -251 14669 -242
rect 14816 -208 14868 -199
rect 14880 -208 14932 -199
rect 14944 -208 14996 -199
rect 15008 -208 15060 -199
rect 15072 -208 15124 -199
rect 14816 -242 14842 -208
rect 14842 -242 14868 -208
rect 14880 -242 14914 -208
rect 14914 -242 14932 -208
rect 14944 -242 14948 -208
rect 14948 -242 14986 -208
rect 14986 -242 14996 -208
rect 15008 -242 15020 -208
rect 15020 -242 15058 -208
rect 15058 -242 15060 -208
rect 15072 -242 15092 -208
rect 15092 -242 15124 -208
rect 14816 -251 14868 -242
rect 14880 -251 14932 -242
rect 14944 -251 14996 -242
rect 15008 -251 15060 -242
rect 15072 -251 15124 -242
rect 15217 -208 15269 -199
rect 15281 -208 15333 -199
rect 15345 -208 15397 -199
rect 15409 -208 15461 -199
rect 15473 -208 15525 -199
rect 15217 -242 15249 -208
rect 15249 -242 15269 -208
rect 15281 -242 15283 -208
rect 15283 -242 15321 -208
rect 15321 -242 15333 -208
rect 15345 -242 15355 -208
rect 15355 -242 15393 -208
rect 15393 -242 15397 -208
rect 15409 -242 15427 -208
rect 15427 -242 15461 -208
rect 15473 -242 15499 -208
rect 15499 -242 15525 -208
rect 15217 -251 15269 -242
rect 15281 -251 15333 -242
rect 15345 -251 15397 -242
rect 15409 -251 15461 -242
rect 15473 -251 15525 -242
rect 15672 -208 15724 -199
rect 15672 -242 15677 -208
rect 15677 -242 15711 -208
rect 15711 -242 15724 -208
rect 15672 -251 15724 -242
rect 15736 -208 15788 -199
rect 15736 -242 15749 -208
rect 15749 -242 15783 -208
rect 15783 -242 15788 -208
rect 15736 -251 15788 -242
rect 12709 -363 12761 -326
rect 15212 -308 15264 -299
rect 15212 -342 15251 -308
rect 15251 -342 15264 -308
rect 15212 -351 15264 -342
rect 12709 -378 12718 -363
rect 12718 -378 12752 -363
rect 12752 -378 12761 -363
rect 12709 -397 12718 -390
rect 12718 -397 12752 -390
rect 12752 -397 12761 -390
rect 12709 -435 12761 -397
rect 12709 -442 12718 -435
rect 12718 -442 12752 -435
rect 12752 -442 12761 -435
rect 14440 -451 14492 -399
rect 14553 -408 14605 -399
rect 14553 -442 14558 -408
rect 14558 -442 14592 -408
rect 14592 -442 14605 -408
rect 14553 -451 14605 -442
rect 14617 -408 14669 -399
rect 14617 -442 14630 -408
rect 14630 -442 14664 -408
rect 14664 -442 14669 -408
rect 14617 -451 14669 -442
rect 12709 -469 12718 -454
rect 12718 -469 12752 -454
rect 12752 -469 12761 -454
rect 14725 -408 14777 -399
rect 14725 -442 14734 -408
rect 14734 -442 14768 -408
rect 14768 -442 14777 -408
rect 14725 -451 14777 -442
rect 14816 -408 14868 -399
rect 14880 -408 14932 -399
rect 14944 -408 14996 -399
rect 15008 -408 15060 -399
rect 15072 -408 15124 -399
rect 14816 -442 14842 -408
rect 14842 -442 14868 -408
rect 14880 -442 14914 -408
rect 14914 -442 14932 -408
rect 14944 -442 14948 -408
rect 14948 -442 14986 -408
rect 14986 -442 14996 -408
rect 15008 -442 15020 -408
rect 15020 -442 15058 -408
rect 15058 -442 15060 -408
rect 15072 -442 15092 -408
rect 15092 -442 15124 -408
rect 14816 -451 14868 -442
rect 14880 -451 14932 -442
rect 14944 -451 14996 -442
rect 15008 -451 15060 -442
rect 15072 -451 15124 -442
rect 15217 -408 15269 -399
rect 15281 -408 15333 -399
rect 15345 -408 15397 -399
rect 15409 -408 15461 -399
rect 15473 -408 15525 -399
rect 15217 -442 15249 -408
rect 15249 -442 15269 -408
rect 15281 -442 15283 -408
rect 15283 -442 15321 -408
rect 15321 -442 15333 -408
rect 15345 -442 15355 -408
rect 15355 -442 15393 -408
rect 15393 -442 15397 -408
rect 15409 -442 15427 -408
rect 15427 -442 15461 -408
rect 15473 -442 15499 -408
rect 15499 -442 15525 -408
rect 15217 -451 15269 -442
rect 15281 -451 15333 -442
rect 15345 -451 15397 -442
rect 15409 -451 15461 -442
rect 15473 -451 15525 -442
rect 15565 -408 15617 -399
rect 15565 -442 15574 -408
rect 15574 -442 15608 -408
rect 15608 -442 15617 -408
rect 15565 -451 15617 -442
rect 15672 -408 15724 -399
rect 15672 -442 15677 -408
rect 15677 -442 15711 -408
rect 15711 -442 15724 -408
rect 15672 -451 15724 -442
rect 15736 -408 15788 -399
rect 15736 -442 15749 -408
rect 15749 -442 15783 -408
rect 15783 -442 15788 -408
rect 15736 -451 15788 -442
rect 12709 -506 12761 -469
rect 15212 -508 15264 -499
rect 15212 -542 15251 -508
rect 15251 -542 15264 -508
rect 15212 -551 15264 -542
rect 14440 -651 14492 -599
rect 14553 -608 14605 -599
rect 14553 -642 14558 -608
rect 14558 -642 14592 -608
rect 14592 -642 14605 -608
rect 14553 -651 14605 -642
rect 14617 -608 14669 -599
rect 14617 -642 14630 -608
rect 14630 -642 14664 -608
rect 14664 -642 14669 -608
rect 14617 -651 14669 -642
rect 14725 -608 14777 -599
rect 14725 -642 14734 -608
rect 14734 -642 14768 -608
rect 14768 -642 14777 -608
rect 14725 -651 14777 -642
rect 14816 -608 14868 -599
rect 14880 -608 14932 -599
rect 14944 -608 14996 -599
rect 15008 -608 15060 -599
rect 15072 -608 15124 -599
rect 14816 -642 14842 -608
rect 14842 -642 14868 -608
rect 14880 -642 14914 -608
rect 14914 -642 14932 -608
rect 14944 -642 14948 -608
rect 14948 -642 14986 -608
rect 14986 -642 14996 -608
rect 15008 -642 15020 -608
rect 15020 -642 15058 -608
rect 15058 -642 15060 -608
rect 15072 -642 15092 -608
rect 15092 -642 15124 -608
rect 14816 -651 14868 -642
rect 14880 -651 14932 -642
rect 14944 -651 14996 -642
rect 15008 -651 15060 -642
rect 15072 -651 15124 -642
rect 15217 -608 15269 -599
rect 15281 -608 15333 -599
rect 15345 -608 15397 -599
rect 15409 -608 15461 -599
rect 15473 -608 15525 -599
rect 15217 -642 15249 -608
rect 15249 -642 15269 -608
rect 15281 -642 15283 -608
rect 15283 -642 15321 -608
rect 15321 -642 15333 -608
rect 15345 -642 15355 -608
rect 15355 -642 15393 -608
rect 15393 -642 15397 -608
rect 15409 -642 15427 -608
rect 15427 -642 15461 -608
rect 15473 -642 15499 -608
rect 15499 -642 15525 -608
rect 15217 -651 15269 -642
rect 15281 -651 15333 -642
rect 15345 -651 15397 -642
rect 15409 -651 15461 -642
rect 15473 -651 15525 -642
rect 15565 -608 15617 -599
rect 15565 -642 15574 -608
rect 15574 -642 15608 -608
rect 15608 -642 15617 -608
rect 15565 -651 15617 -642
rect 15672 -608 15724 -599
rect 15672 -642 15677 -608
rect 15677 -642 15711 -608
rect 15711 -642 15724 -608
rect 15672 -651 15724 -642
rect 15736 -608 15788 -599
rect 15736 -642 15749 -608
rect 15749 -642 15783 -608
rect 15783 -642 15788 -608
rect 15736 -651 15788 -642
rect 15212 -708 15264 -699
rect 15212 -742 15251 -708
rect 15251 -742 15264 -708
rect 15212 -751 15264 -742
rect -9 -837 43 -828
rect -9 -871 -4 -837
rect -4 -871 30 -837
rect 30 -871 43 -837
rect -9 -880 43 -871
rect 55 -837 107 -828
rect 55 -871 68 -837
rect 68 -871 102 -837
rect 102 -871 107 -837
rect 55 -880 107 -871
rect 163 -837 215 -828
rect 163 -871 168 -837
rect 168 -871 202 -837
rect 202 -871 215 -837
rect 163 -880 215 -871
rect 227 -837 279 -828
rect 227 -871 240 -837
rect 240 -871 274 -837
rect 274 -871 279 -837
rect 227 -880 279 -871
rect 391 -837 443 -828
rect 391 -871 396 -837
rect 396 -871 430 -837
rect 430 -871 443 -837
rect 391 -880 443 -871
rect 455 -837 507 -828
rect 455 -871 468 -837
rect 468 -871 502 -837
rect 502 -871 507 -837
rect 455 -880 507 -871
rect 563 -837 615 -828
rect 563 -871 568 -837
rect 568 -871 602 -837
rect 602 -871 615 -837
rect 563 -880 615 -871
rect 627 -837 679 -828
rect 627 -871 640 -837
rect 640 -871 674 -837
rect 674 -871 679 -837
rect 627 -880 679 -871
rect 791 -837 843 -828
rect 791 -871 796 -837
rect 796 -871 830 -837
rect 830 -871 843 -837
rect 791 -880 843 -871
rect 855 -837 907 -828
rect 855 -871 868 -837
rect 868 -871 902 -837
rect 902 -871 907 -837
rect 855 -880 907 -871
rect 963 -837 1015 -828
rect 963 -871 968 -837
rect 968 -871 1002 -837
rect 1002 -871 1015 -837
rect 963 -880 1015 -871
rect 1027 -837 1079 -828
rect 1027 -871 1040 -837
rect 1040 -871 1074 -837
rect 1074 -871 1079 -837
rect 1027 -880 1079 -871
rect 1191 -837 1243 -828
rect 1191 -871 1196 -837
rect 1196 -871 1230 -837
rect 1230 -871 1243 -837
rect 1191 -880 1243 -871
rect 1255 -837 1307 -828
rect 1255 -871 1268 -837
rect 1268 -871 1302 -837
rect 1302 -871 1307 -837
rect 1255 -880 1307 -871
rect 1363 -837 1415 -828
rect 1363 -871 1368 -837
rect 1368 -871 1402 -837
rect 1402 -871 1415 -837
rect 1363 -880 1415 -871
rect 1427 -837 1479 -828
rect 1427 -871 1440 -837
rect 1440 -871 1474 -837
rect 1474 -871 1479 -837
rect 1427 -880 1479 -871
rect 1591 -837 1643 -828
rect 1591 -871 1596 -837
rect 1596 -871 1630 -837
rect 1630 -871 1643 -837
rect 1591 -880 1643 -871
rect 1655 -837 1707 -828
rect 1655 -871 1668 -837
rect 1668 -871 1702 -837
rect 1702 -871 1707 -837
rect 1655 -880 1707 -871
rect 1763 -837 1815 -828
rect 1763 -871 1768 -837
rect 1768 -871 1802 -837
rect 1802 -871 1815 -837
rect 1763 -880 1815 -871
rect 1827 -837 1879 -828
rect 1827 -871 1840 -837
rect 1840 -871 1874 -837
rect 1874 -871 1879 -837
rect 1827 -880 1879 -871
rect 1991 -837 2043 -828
rect 1991 -871 1996 -837
rect 1996 -871 2030 -837
rect 2030 -871 2043 -837
rect 1991 -880 2043 -871
rect 2055 -837 2107 -828
rect 2055 -871 2068 -837
rect 2068 -871 2102 -837
rect 2102 -871 2107 -837
rect 2055 -880 2107 -871
rect 2163 -837 2215 -828
rect 2163 -871 2168 -837
rect 2168 -871 2202 -837
rect 2202 -871 2215 -837
rect 2163 -880 2215 -871
rect 2227 -837 2279 -828
rect 2227 -871 2240 -837
rect 2240 -871 2274 -837
rect 2274 -871 2279 -837
rect 2227 -880 2279 -871
rect 2391 -837 2443 -828
rect 2391 -871 2396 -837
rect 2396 -871 2430 -837
rect 2430 -871 2443 -837
rect 2391 -880 2443 -871
rect 2455 -837 2507 -828
rect 2455 -871 2468 -837
rect 2468 -871 2502 -837
rect 2502 -871 2507 -837
rect 2455 -880 2507 -871
rect 2563 -837 2615 -828
rect 2563 -871 2568 -837
rect 2568 -871 2602 -837
rect 2602 -871 2615 -837
rect 2563 -880 2615 -871
rect 2627 -837 2679 -828
rect 2627 -871 2640 -837
rect 2640 -871 2674 -837
rect 2674 -871 2679 -837
rect 2627 -880 2679 -871
rect 2791 -837 2843 -828
rect 2791 -871 2796 -837
rect 2796 -871 2830 -837
rect 2830 -871 2843 -837
rect 2791 -880 2843 -871
rect 2855 -837 2907 -828
rect 2855 -871 2868 -837
rect 2868 -871 2902 -837
rect 2902 -871 2907 -837
rect 2855 -880 2907 -871
rect 2963 -837 3015 -828
rect 2963 -871 2968 -837
rect 2968 -871 3002 -837
rect 3002 -871 3015 -837
rect 2963 -880 3015 -871
rect 3027 -837 3079 -828
rect 3027 -871 3040 -837
rect 3040 -871 3074 -837
rect 3074 -871 3079 -837
rect 3027 -880 3079 -871
rect 3191 -837 3243 -828
rect 3191 -871 3196 -837
rect 3196 -871 3230 -837
rect 3230 -871 3243 -837
rect 3191 -880 3243 -871
rect 3255 -837 3307 -828
rect 3255 -871 3268 -837
rect 3268 -871 3302 -837
rect 3302 -871 3307 -837
rect 3255 -880 3307 -871
rect 3363 -837 3415 -828
rect 3363 -871 3368 -837
rect 3368 -871 3402 -837
rect 3402 -871 3415 -837
rect 3363 -880 3415 -871
rect 3427 -837 3479 -828
rect 3427 -871 3440 -837
rect 3440 -871 3474 -837
rect 3474 -871 3479 -837
rect 3427 -880 3479 -871
rect 3591 -837 3643 -828
rect 3591 -871 3596 -837
rect 3596 -871 3630 -837
rect 3630 -871 3643 -837
rect 3591 -880 3643 -871
rect 3655 -837 3707 -828
rect 3655 -871 3668 -837
rect 3668 -871 3702 -837
rect 3702 -871 3707 -837
rect 3655 -880 3707 -871
rect 3763 -837 3815 -828
rect 3763 -871 3768 -837
rect 3768 -871 3802 -837
rect 3802 -871 3815 -837
rect 3763 -880 3815 -871
rect 3827 -837 3879 -828
rect 3827 -871 3840 -837
rect 3840 -871 3874 -837
rect 3874 -871 3879 -837
rect 3827 -880 3879 -871
rect 3991 -837 4043 -828
rect 3991 -871 3996 -837
rect 3996 -871 4030 -837
rect 4030 -871 4043 -837
rect 3991 -880 4043 -871
rect 4055 -837 4107 -828
rect 4055 -871 4068 -837
rect 4068 -871 4102 -837
rect 4102 -871 4107 -837
rect 4055 -880 4107 -871
rect 4163 -837 4215 -828
rect 4163 -871 4168 -837
rect 4168 -871 4202 -837
rect 4202 -871 4215 -837
rect 4163 -880 4215 -871
rect 4227 -837 4279 -828
rect 4227 -871 4240 -837
rect 4240 -871 4274 -837
rect 4274 -871 4279 -837
rect 4227 -880 4279 -871
rect 4391 -837 4443 -828
rect 4391 -871 4396 -837
rect 4396 -871 4430 -837
rect 4430 -871 4443 -837
rect 4391 -880 4443 -871
rect 4455 -837 4507 -828
rect 4455 -871 4468 -837
rect 4468 -871 4502 -837
rect 4502 -871 4507 -837
rect 4455 -880 4507 -871
rect 4563 -837 4615 -828
rect 4563 -871 4568 -837
rect 4568 -871 4602 -837
rect 4602 -871 4615 -837
rect 4563 -880 4615 -871
rect 4627 -837 4679 -828
rect 4627 -871 4640 -837
rect 4640 -871 4674 -837
rect 4674 -871 4679 -837
rect 4627 -880 4679 -871
rect 4791 -837 4843 -828
rect 4791 -871 4796 -837
rect 4796 -871 4830 -837
rect 4830 -871 4843 -837
rect 4791 -880 4843 -871
rect 4855 -837 4907 -828
rect 4855 -871 4868 -837
rect 4868 -871 4902 -837
rect 4902 -871 4907 -837
rect 4855 -880 4907 -871
rect 4963 -837 5015 -828
rect 4963 -871 4968 -837
rect 4968 -871 5002 -837
rect 5002 -871 5015 -837
rect 4963 -880 5015 -871
rect 5027 -837 5079 -828
rect 5027 -871 5040 -837
rect 5040 -871 5074 -837
rect 5074 -871 5079 -837
rect 5027 -880 5079 -871
rect 5191 -837 5243 -828
rect 5191 -871 5196 -837
rect 5196 -871 5230 -837
rect 5230 -871 5243 -837
rect 5191 -880 5243 -871
rect 5255 -837 5307 -828
rect 5255 -871 5268 -837
rect 5268 -871 5302 -837
rect 5302 -871 5307 -837
rect 5255 -880 5307 -871
rect 5363 -837 5415 -828
rect 5363 -871 5368 -837
rect 5368 -871 5402 -837
rect 5402 -871 5415 -837
rect 5363 -880 5415 -871
rect 5427 -837 5479 -828
rect 5427 -871 5440 -837
rect 5440 -871 5474 -837
rect 5474 -871 5479 -837
rect 5427 -880 5479 -871
rect 5591 -837 5643 -828
rect 5591 -871 5596 -837
rect 5596 -871 5630 -837
rect 5630 -871 5643 -837
rect 5591 -880 5643 -871
rect 5655 -837 5707 -828
rect 5655 -871 5668 -837
rect 5668 -871 5702 -837
rect 5702 -871 5707 -837
rect 5655 -880 5707 -871
rect 5763 -837 5815 -828
rect 5763 -871 5768 -837
rect 5768 -871 5802 -837
rect 5802 -871 5815 -837
rect 5763 -880 5815 -871
rect 5827 -837 5879 -828
rect 5827 -871 5840 -837
rect 5840 -871 5874 -837
rect 5874 -871 5879 -837
rect 5827 -880 5879 -871
rect 5991 -837 6043 -828
rect 5991 -871 5996 -837
rect 5996 -871 6030 -837
rect 6030 -871 6043 -837
rect 5991 -880 6043 -871
rect 6055 -837 6107 -828
rect 6055 -871 6068 -837
rect 6068 -871 6102 -837
rect 6102 -871 6107 -837
rect 6055 -880 6107 -871
rect 6163 -837 6215 -828
rect 6163 -871 6168 -837
rect 6168 -871 6202 -837
rect 6202 -871 6215 -837
rect 6163 -880 6215 -871
rect 6227 -837 6279 -828
rect 6227 -871 6240 -837
rect 6240 -871 6274 -837
rect 6274 -871 6279 -837
rect 6227 -880 6279 -871
rect 6391 -837 6443 -828
rect 6391 -871 6396 -837
rect 6396 -871 6430 -837
rect 6430 -871 6443 -837
rect 6391 -880 6443 -871
rect 6455 -837 6507 -828
rect 6455 -871 6468 -837
rect 6468 -871 6502 -837
rect 6502 -871 6507 -837
rect 6455 -880 6507 -871
rect 6563 -837 6615 -828
rect 6563 -871 6568 -837
rect 6568 -871 6602 -837
rect 6602 -871 6615 -837
rect 6563 -880 6615 -871
rect 6627 -837 6679 -828
rect 6627 -871 6640 -837
rect 6640 -871 6674 -837
rect 6674 -871 6679 -837
rect 6627 -880 6679 -871
rect 6791 -837 6843 -828
rect 6791 -871 6796 -837
rect 6796 -871 6830 -837
rect 6830 -871 6843 -837
rect 6791 -880 6843 -871
rect 6855 -837 6907 -828
rect 6855 -871 6868 -837
rect 6868 -871 6902 -837
rect 6902 -871 6907 -837
rect 6855 -880 6907 -871
rect 6963 -837 7015 -828
rect 6963 -871 6968 -837
rect 6968 -871 7002 -837
rect 7002 -871 7015 -837
rect 6963 -880 7015 -871
rect 7027 -837 7079 -828
rect 7027 -871 7040 -837
rect 7040 -871 7074 -837
rect 7074 -871 7079 -837
rect 7027 -880 7079 -871
rect 7191 -837 7243 -828
rect 7191 -871 7196 -837
rect 7196 -871 7230 -837
rect 7230 -871 7243 -837
rect 7191 -880 7243 -871
rect 7255 -837 7307 -828
rect 7255 -871 7268 -837
rect 7268 -871 7302 -837
rect 7302 -871 7307 -837
rect 7255 -880 7307 -871
rect 7363 -837 7415 -828
rect 7363 -871 7368 -837
rect 7368 -871 7402 -837
rect 7402 -871 7415 -837
rect 7363 -880 7415 -871
rect 7427 -837 7479 -828
rect 7427 -871 7440 -837
rect 7440 -871 7474 -837
rect 7474 -871 7479 -837
rect 7427 -880 7479 -871
rect 7591 -837 7643 -828
rect 7591 -871 7596 -837
rect 7596 -871 7630 -837
rect 7630 -871 7643 -837
rect 7591 -880 7643 -871
rect 7655 -837 7707 -828
rect 7655 -871 7668 -837
rect 7668 -871 7702 -837
rect 7702 -871 7707 -837
rect 7655 -880 7707 -871
rect 7763 -837 7815 -828
rect 7763 -871 7768 -837
rect 7768 -871 7802 -837
rect 7802 -871 7815 -837
rect 7763 -880 7815 -871
rect 7827 -837 7879 -828
rect 7827 -871 7840 -837
rect 7840 -871 7874 -837
rect 7874 -871 7879 -837
rect 7827 -880 7879 -871
rect 7991 -837 8043 -828
rect 7991 -871 7996 -837
rect 7996 -871 8030 -837
rect 8030 -871 8043 -837
rect 7991 -880 8043 -871
rect 8055 -837 8107 -828
rect 8055 -871 8068 -837
rect 8068 -871 8102 -837
rect 8102 -871 8107 -837
rect 8055 -880 8107 -871
rect 8163 -837 8215 -828
rect 8163 -871 8168 -837
rect 8168 -871 8202 -837
rect 8202 -871 8215 -837
rect 8163 -880 8215 -871
rect 8227 -837 8279 -828
rect 8227 -871 8240 -837
rect 8240 -871 8274 -837
rect 8274 -871 8279 -837
rect 8227 -880 8279 -871
rect 8391 -837 8443 -828
rect 8391 -871 8396 -837
rect 8396 -871 8430 -837
rect 8430 -871 8443 -837
rect 8391 -880 8443 -871
rect 8455 -837 8507 -828
rect 8455 -871 8468 -837
rect 8468 -871 8502 -837
rect 8502 -871 8507 -837
rect 8455 -880 8507 -871
rect 8563 -837 8615 -828
rect 8563 -871 8568 -837
rect 8568 -871 8602 -837
rect 8602 -871 8615 -837
rect 8563 -880 8615 -871
rect 8627 -837 8679 -828
rect 8627 -871 8640 -837
rect 8640 -871 8674 -837
rect 8674 -871 8679 -837
rect 8627 -880 8679 -871
rect 8791 -837 8843 -828
rect 8791 -871 8796 -837
rect 8796 -871 8830 -837
rect 8830 -871 8843 -837
rect 8791 -880 8843 -871
rect 8855 -837 8907 -828
rect 8855 -871 8868 -837
rect 8868 -871 8902 -837
rect 8902 -871 8907 -837
rect 8855 -880 8907 -871
rect 8963 -837 9015 -828
rect 8963 -871 8968 -837
rect 8968 -871 9002 -837
rect 9002 -871 9015 -837
rect 8963 -880 9015 -871
rect 9027 -837 9079 -828
rect 9027 -871 9040 -837
rect 9040 -871 9074 -837
rect 9074 -871 9079 -837
rect 9027 -880 9079 -871
rect 9191 -837 9243 -828
rect 9191 -871 9196 -837
rect 9196 -871 9230 -837
rect 9230 -871 9243 -837
rect 9191 -880 9243 -871
rect 9255 -837 9307 -828
rect 9255 -871 9268 -837
rect 9268 -871 9302 -837
rect 9302 -871 9307 -837
rect 9255 -880 9307 -871
rect 9363 -837 9415 -828
rect 9363 -871 9368 -837
rect 9368 -871 9402 -837
rect 9402 -871 9415 -837
rect 9363 -880 9415 -871
rect 9427 -837 9479 -828
rect 9427 -871 9440 -837
rect 9440 -871 9474 -837
rect 9474 -871 9479 -837
rect 9427 -880 9479 -871
rect 9591 -837 9643 -828
rect 9591 -871 9596 -837
rect 9596 -871 9630 -837
rect 9630 -871 9643 -837
rect 9591 -880 9643 -871
rect 9655 -837 9707 -828
rect 9655 -871 9668 -837
rect 9668 -871 9702 -837
rect 9702 -871 9707 -837
rect 9655 -880 9707 -871
rect 9763 -837 9815 -828
rect 9763 -871 9768 -837
rect 9768 -871 9802 -837
rect 9802 -871 9815 -837
rect 9763 -880 9815 -871
rect 9827 -837 9879 -828
rect 9827 -871 9840 -837
rect 9840 -871 9874 -837
rect 9874 -871 9879 -837
rect 9827 -880 9879 -871
rect 9991 -837 10043 -828
rect 9991 -871 9996 -837
rect 9996 -871 10030 -837
rect 10030 -871 10043 -837
rect 9991 -880 10043 -871
rect 10055 -837 10107 -828
rect 10055 -871 10068 -837
rect 10068 -871 10102 -837
rect 10102 -871 10107 -837
rect 10055 -880 10107 -871
rect 10163 -837 10215 -828
rect 10163 -871 10168 -837
rect 10168 -871 10202 -837
rect 10202 -871 10215 -837
rect 10163 -880 10215 -871
rect 10227 -837 10279 -828
rect 10227 -871 10240 -837
rect 10240 -871 10274 -837
rect 10274 -871 10279 -837
rect 10227 -880 10279 -871
rect 10391 -837 10443 -828
rect 10391 -871 10396 -837
rect 10396 -871 10430 -837
rect 10430 -871 10443 -837
rect 10391 -880 10443 -871
rect 10455 -837 10507 -828
rect 10455 -871 10468 -837
rect 10468 -871 10502 -837
rect 10502 -871 10507 -837
rect 10455 -880 10507 -871
rect 10563 -837 10615 -828
rect 10563 -871 10568 -837
rect 10568 -871 10602 -837
rect 10602 -871 10615 -837
rect 10563 -880 10615 -871
rect 10627 -837 10679 -828
rect 10627 -871 10640 -837
rect 10640 -871 10674 -837
rect 10674 -871 10679 -837
rect 10627 -880 10679 -871
rect 10791 -837 10843 -828
rect 10791 -871 10796 -837
rect 10796 -871 10830 -837
rect 10830 -871 10843 -837
rect 10791 -880 10843 -871
rect 10855 -837 10907 -828
rect 10855 -871 10868 -837
rect 10868 -871 10902 -837
rect 10902 -871 10907 -837
rect 10855 -880 10907 -871
rect 10963 -837 11015 -828
rect 10963 -871 10968 -837
rect 10968 -871 11002 -837
rect 11002 -871 11015 -837
rect 10963 -880 11015 -871
rect 11027 -837 11079 -828
rect 11027 -871 11040 -837
rect 11040 -871 11074 -837
rect 11074 -871 11079 -837
rect 11027 -880 11079 -871
rect 11191 -837 11243 -828
rect 11191 -871 11196 -837
rect 11196 -871 11230 -837
rect 11230 -871 11243 -837
rect 11191 -880 11243 -871
rect 11255 -837 11307 -828
rect 11255 -871 11268 -837
rect 11268 -871 11302 -837
rect 11302 -871 11307 -837
rect 11255 -880 11307 -871
rect 11363 -837 11415 -828
rect 11363 -871 11368 -837
rect 11368 -871 11402 -837
rect 11402 -871 11415 -837
rect 11363 -880 11415 -871
rect 11427 -837 11479 -828
rect 11427 -871 11440 -837
rect 11440 -871 11474 -837
rect 11474 -871 11479 -837
rect 11427 -880 11479 -871
rect 11591 -837 11643 -828
rect 11591 -871 11596 -837
rect 11596 -871 11630 -837
rect 11630 -871 11643 -837
rect 11591 -880 11643 -871
rect 11655 -837 11707 -828
rect 11655 -871 11668 -837
rect 11668 -871 11702 -837
rect 11702 -871 11707 -837
rect 11655 -880 11707 -871
rect 11763 -837 11815 -828
rect 11763 -871 11768 -837
rect 11768 -871 11802 -837
rect 11802 -871 11815 -837
rect 11763 -880 11815 -871
rect 11827 -837 11879 -828
rect 11827 -871 11840 -837
rect 11840 -871 11874 -837
rect 11874 -871 11879 -837
rect 11827 -880 11879 -871
rect 11991 -837 12043 -828
rect 11991 -871 11996 -837
rect 11996 -871 12030 -837
rect 12030 -871 12043 -837
rect 11991 -880 12043 -871
rect 12055 -837 12107 -828
rect 12055 -871 12068 -837
rect 12068 -871 12102 -837
rect 12102 -871 12107 -837
rect 12055 -880 12107 -871
rect 12163 -837 12215 -828
rect 12163 -871 12168 -837
rect 12168 -871 12202 -837
rect 12202 -871 12215 -837
rect 12163 -880 12215 -871
rect 12227 -837 12279 -828
rect 12227 -871 12240 -837
rect 12240 -871 12274 -837
rect 12274 -871 12279 -837
rect 12227 -880 12279 -871
rect 12391 -837 12443 -828
rect 12391 -871 12396 -837
rect 12396 -871 12430 -837
rect 12430 -871 12443 -837
rect 12391 -880 12443 -871
rect 12455 -837 12507 -828
rect 12455 -871 12468 -837
rect 12468 -871 12502 -837
rect 12502 -871 12507 -837
rect 12455 -880 12507 -871
rect 12563 -837 12615 -828
rect 12563 -871 12568 -837
rect 12568 -871 12602 -837
rect 12602 -871 12615 -837
rect 12563 -880 12615 -871
rect 12627 -837 12679 -828
rect 12627 -871 12640 -837
rect 12640 -871 12674 -837
rect 12674 -871 12679 -837
rect 12627 -880 12679 -871
rect 14440 -851 14492 -799
rect 14553 -808 14605 -799
rect 14553 -842 14558 -808
rect 14558 -842 14592 -808
rect 14592 -842 14605 -808
rect 14553 -851 14605 -842
rect 14617 -808 14669 -799
rect 14617 -842 14630 -808
rect 14630 -842 14664 -808
rect 14664 -842 14669 -808
rect 14617 -851 14669 -842
rect 14725 -808 14777 -799
rect 14725 -842 14734 -808
rect 14734 -842 14768 -808
rect 14768 -842 14777 -808
rect 14725 -851 14777 -842
rect 14816 -808 14868 -799
rect 14880 -808 14932 -799
rect 14944 -808 14996 -799
rect 15008 -808 15060 -799
rect 15072 -808 15124 -799
rect 14816 -842 14842 -808
rect 14842 -842 14868 -808
rect 14880 -842 14914 -808
rect 14914 -842 14932 -808
rect 14944 -842 14948 -808
rect 14948 -842 14986 -808
rect 14986 -842 14996 -808
rect 15008 -842 15020 -808
rect 15020 -842 15058 -808
rect 15058 -842 15060 -808
rect 15072 -842 15092 -808
rect 15092 -842 15124 -808
rect 14816 -851 14868 -842
rect 14880 -851 14932 -842
rect 14944 -851 14996 -842
rect 15008 -851 15060 -842
rect 15072 -851 15124 -842
rect 15217 -808 15269 -799
rect 15281 -808 15333 -799
rect 15345 -808 15397 -799
rect 15409 -808 15461 -799
rect 15473 -808 15525 -799
rect 15217 -842 15249 -808
rect 15249 -842 15269 -808
rect 15281 -842 15283 -808
rect 15283 -842 15321 -808
rect 15321 -842 15333 -808
rect 15345 -842 15355 -808
rect 15355 -842 15393 -808
rect 15393 -842 15397 -808
rect 15409 -842 15427 -808
rect 15427 -842 15461 -808
rect 15473 -842 15499 -808
rect 15499 -842 15525 -808
rect 15217 -851 15269 -842
rect 15281 -851 15333 -842
rect 15345 -851 15397 -842
rect 15409 -851 15461 -842
rect 15473 -851 15525 -842
rect 15565 -808 15617 -799
rect 15565 -842 15574 -808
rect 15574 -842 15608 -808
rect 15608 -842 15617 -808
rect 15565 -851 15617 -842
rect 15672 -808 15724 -799
rect 15672 -842 15677 -808
rect 15677 -842 15711 -808
rect 15711 -842 15724 -808
rect 15672 -851 15724 -842
rect 15736 -808 15788 -799
rect 15736 -842 15749 -808
rect 15749 -842 15783 -808
rect 15783 -842 15788 -808
rect 15736 -851 15788 -842
rect 15212 -908 15264 -899
rect 15212 -942 15251 -908
rect 15251 -942 15264 -908
rect 15212 -951 15264 -942
rect 14440 -1051 14492 -999
rect 14553 -1008 14605 -999
rect 14553 -1042 14558 -1008
rect 14558 -1042 14592 -1008
rect 14592 -1042 14605 -1008
rect 14553 -1051 14605 -1042
rect 14617 -1008 14669 -999
rect 14617 -1042 14630 -1008
rect 14630 -1042 14664 -1008
rect 14664 -1042 14669 -1008
rect 14617 -1051 14669 -1042
rect 14725 -1008 14777 -999
rect 14725 -1042 14734 -1008
rect 14734 -1042 14768 -1008
rect 14768 -1042 14777 -1008
rect 14725 -1051 14777 -1042
rect 14816 -1008 14868 -999
rect 14880 -1008 14932 -999
rect 14944 -1008 14996 -999
rect 15008 -1008 15060 -999
rect 15072 -1008 15124 -999
rect 14816 -1042 14842 -1008
rect 14842 -1042 14868 -1008
rect 14880 -1042 14914 -1008
rect 14914 -1042 14932 -1008
rect 14944 -1042 14948 -1008
rect 14948 -1042 14986 -1008
rect 14986 -1042 14996 -1008
rect 15008 -1042 15020 -1008
rect 15020 -1042 15058 -1008
rect 15058 -1042 15060 -1008
rect 15072 -1042 15092 -1008
rect 15092 -1042 15124 -1008
rect 14816 -1051 14868 -1042
rect 14880 -1051 14932 -1042
rect 14944 -1051 14996 -1042
rect 15008 -1051 15060 -1042
rect 15072 -1051 15124 -1042
rect 15217 -1008 15269 -999
rect 15281 -1008 15333 -999
rect 15345 -1008 15397 -999
rect 15409 -1008 15461 -999
rect 15473 -1008 15525 -999
rect 15217 -1042 15249 -1008
rect 15249 -1042 15269 -1008
rect 15281 -1042 15283 -1008
rect 15283 -1042 15321 -1008
rect 15321 -1042 15333 -1008
rect 15345 -1042 15355 -1008
rect 15355 -1042 15393 -1008
rect 15393 -1042 15397 -1008
rect 15409 -1042 15427 -1008
rect 15427 -1042 15461 -1008
rect 15473 -1042 15499 -1008
rect 15499 -1042 15525 -1008
rect 15217 -1051 15269 -1042
rect 15281 -1051 15333 -1042
rect 15345 -1051 15397 -1042
rect 15409 -1051 15461 -1042
rect 15473 -1051 15525 -1042
rect 15565 -1008 15617 -999
rect 15565 -1042 15574 -1008
rect 15574 -1042 15608 -1008
rect 15608 -1042 15617 -1008
rect 15565 -1051 15617 -1042
rect 15672 -1008 15724 -999
rect 15672 -1042 15677 -1008
rect 15677 -1042 15711 -1008
rect 15711 -1042 15724 -1008
rect 15672 -1051 15724 -1042
rect 15736 -1008 15788 -999
rect 15736 -1042 15749 -1008
rect 15749 -1042 15783 -1008
rect 15783 -1042 15788 -1008
rect 15736 -1051 15788 -1042
rect 15212 -1108 15264 -1099
rect 15212 -1142 15251 -1108
rect 15251 -1142 15264 -1108
rect 15212 -1151 15264 -1142
rect 14440 -1251 14492 -1199
rect 14553 -1208 14605 -1199
rect 14553 -1242 14558 -1208
rect 14558 -1242 14592 -1208
rect 14592 -1242 14605 -1208
rect 14553 -1251 14605 -1242
rect 14617 -1208 14669 -1199
rect 14617 -1242 14630 -1208
rect 14630 -1242 14664 -1208
rect 14664 -1242 14669 -1208
rect 14617 -1251 14669 -1242
rect 14725 -1208 14777 -1199
rect 14725 -1242 14734 -1208
rect 14734 -1242 14768 -1208
rect 14768 -1242 14777 -1208
rect 14725 -1251 14777 -1242
rect 14816 -1208 14868 -1199
rect 14880 -1208 14932 -1199
rect 14944 -1208 14996 -1199
rect 15008 -1208 15060 -1199
rect 15072 -1208 15124 -1199
rect 14816 -1242 14842 -1208
rect 14842 -1242 14868 -1208
rect 14880 -1242 14914 -1208
rect 14914 -1242 14932 -1208
rect 14944 -1242 14948 -1208
rect 14948 -1242 14986 -1208
rect 14986 -1242 14996 -1208
rect 15008 -1242 15020 -1208
rect 15020 -1242 15058 -1208
rect 15058 -1242 15060 -1208
rect 15072 -1242 15092 -1208
rect 15092 -1242 15124 -1208
rect 14816 -1251 14868 -1242
rect 14880 -1251 14932 -1242
rect 14944 -1251 14996 -1242
rect 15008 -1251 15060 -1242
rect 15072 -1251 15124 -1242
rect 15217 -1208 15269 -1199
rect 15281 -1208 15333 -1199
rect 15345 -1208 15397 -1199
rect 15409 -1208 15461 -1199
rect 15473 -1208 15525 -1199
rect 15217 -1242 15249 -1208
rect 15249 -1242 15269 -1208
rect 15281 -1242 15283 -1208
rect 15283 -1242 15321 -1208
rect 15321 -1242 15333 -1208
rect 15345 -1242 15355 -1208
rect 15355 -1242 15393 -1208
rect 15393 -1242 15397 -1208
rect 15409 -1242 15427 -1208
rect 15427 -1242 15461 -1208
rect 15473 -1242 15499 -1208
rect 15499 -1242 15525 -1208
rect 15217 -1251 15269 -1242
rect 15281 -1251 15333 -1242
rect 15345 -1251 15397 -1242
rect 15409 -1251 15461 -1242
rect 15473 -1251 15525 -1242
rect 15565 -1208 15617 -1199
rect 15565 -1242 15574 -1208
rect 15574 -1242 15608 -1208
rect 15608 -1242 15617 -1208
rect 15565 -1251 15617 -1242
rect 15672 -1208 15724 -1199
rect 15672 -1242 15677 -1208
rect 15677 -1242 15711 -1208
rect 15711 -1242 15724 -1208
rect 15672 -1251 15724 -1242
rect 15736 -1208 15788 -1199
rect 15736 -1242 15749 -1208
rect 15749 -1242 15783 -1208
rect 15783 -1242 15788 -1208
rect 15736 -1251 15788 -1242
rect 15212 -1308 15264 -1299
rect 15212 -1342 15251 -1308
rect 15251 -1342 15264 -1308
rect 15212 -1351 15264 -1342
rect 14440 -1451 14492 -1399
rect 14553 -1408 14605 -1399
rect 14553 -1442 14558 -1408
rect 14558 -1442 14592 -1408
rect 14592 -1442 14605 -1408
rect 14553 -1451 14605 -1442
rect 14617 -1408 14669 -1399
rect 14617 -1442 14630 -1408
rect 14630 -1442 14664 -1408
rect 14664 -1442 14669 -1408
rect 14617 -1451 14669 -1442
rect 14725 -1408 14777 -1399
rect 14725 -1442 14734 -1408
rect 14734 -1442 14768 -1408
rect 14768 -1442 14777 -1408
rect 14725 -1451 14777 -1442
rect 14816 -1408 14868 -1399
rect 14880 -1408 14932 -1399
rect 14944 -1408 14996 -1399
rect 15008 -1408 15060 -1399
rect 15072 -1408 15124 -1399
rect 14816 -1442 14842 -1408
rect 14842 -1442 14868 -1408
rect 14880 -1442 14914 -1408
rect 14914 -1442 14932 -1408
rect 14944 -1442 14948 -1408
rect 14948 -1442 14986 -1408
rect 14986 -1442 14996 -1408
rect 15008 -1442 15020 -1408
rect 15020 -1442 15058 -1408
rect 15058 -1442 15060 -1408
rect 15072 -1442 15092 -1408
rect 15092 -1442 15124 -1408
rect 14816 -1451 14868 -1442
rect 14880 -1451 14932 -1442
rect 14944 -1451 14996 -1442
rect 15008 -1451 15060 -1442
rect 15072 -1451 15124 -1442
rect 15217 -1408 15269 -1399
rect 15281 -1408 15333 -1399
rect 15345 -1408 15397 -1399
rect 15409 -1408 15461 -1399
rect 15473 -1408 15525 -1399
rect 15217 -1442 15249 -1408
rect 15249 -1442 15269 -1408
rect 15281 -1442 15283 -1408
rect 15283 -1442 15321 -1408
rect 15321 -1442 15333 -1408
rect 15345 -1442 15355 -1408
rect 15355 -1442 15393 -1408
rect 15393 -1442 15397 -1408
rect 15409 -1442 15427 -1408
rect 15427 -1442 15461 -1408
rect 15473 -1442 15499 -1408
rect 15499 -1442 15525 -1408
rect 15217 -1451 15269 -1442
rect 15281 -1451 15333 -1442
rect 15345 -1451 15397 -1442
rect 15409 -1451 15461 -1442
rect 15473 -1451 15525 -1442
rect 15565 -1408 15617 -1399
rect 15565 -1442 15574 -1408
rect 15574 -1442 15608 -1408
rect 15608 -1442 15617 -1408
rect 15565 -1451 15617 -1442
rect 15672 -1408 15724 -1399
rect 15672 -1442 15677 -1408
rect 15677 -1442 15711 -1408
rect 15711 -1442 15724 -1408
rect 15672 -1451 15724 -1442
rect 15736 -1408 15788 -1399
rect 15736 -1442 15749 -1408
rect 15749 -1442 15783 -1408
rect 15783 -1442 15788 -1408
rect 15736 -1451 15788 -1442
rect 15212 -1508 15264 -1499
rect 15212 -1542 15251 -1508
rect 15251 -1542 15264 -1508
rect 15212 -1551 15264 -1542
rect 14440 -1651 14492 -1599
rect 14553 -1608 14605 -1599
rect 14553 -1642 14558 -1608
rect 14558 -1642 14592 -1608
rect 14592 -1642 14605 -1608
rect 14553 -1651 14605 -1642
rect 14617 -1608 14669 -1599
rect 14617 -1642 14630 -1608
rect 14630 -1642 14664 -1608
rect 14664 -1642 14669 -1608
rect 14617 -1651 14669 -1642
rect 14725 -1608 14777 -1599
rect 14725 -1642 14734 -1608
rect 14734 -1642 14768 -1608
rect 14768 -1642 14777 -1608
rect 14725 -1651 14777 -1642
rect 14816 -1608 14868 -1599
rect 14880 -1608 14932 -1599
rect 14944 -1608 14996 -1599
rect 15008 -1608 15060 -1599
rect 15072 -1608 15124 -1599
rect 14816 -1642 14842 -1608
rect 14842 -1642 14868 -1608
rect 14880 -1642 14914 -1608
rect 14914 -1642 14932 -1608
rect 14944 -1642 14948 -1608
rect 14948 -1642 14986 -1608
rect 14986 -1642 14996 -1608
rect 15008 -1642 15020 -1608
rect 15020 -1642 15058 -1608
rect 15058 -1642 15060 -1608
rect 15072 -1642 15092 -1608
rect 15092 -1642 15124 -1608
rect 14816 -1651 14868 -1642
rect 14880 -1651 14932 -1642
rect 14944 -1651 14996 -1642
rect 15008 -1651 15060 -1642
rect 15072 -1651 15124 -1642
rect 15217 -1608 15269 -1599
rect 15281 -1608 15333 -1599
rect 15345 -1608 15397 -1599
rect 15409 -1608 15461 -1599
rect 15473 -1608 15525 -1599
rect 15217 -1642 15249 -1608
rect 15249 -1642 15269 -1608
rect 15281 -1642 15283 -1608
rect 15283 -1642 15321 -1608
rect 15321 -1642 15333 -1608
rect 15345 -1642 15355 -1608
rect 15355 -1642 15393 -1608
rect 15393 -1642 15397 -1608
rect 15409 -1642 15427 -1608
rect 15427 -1642 15461 -1608
rect 15473 -1642 15499 -1608
rect 15499 -1642 15525 -1608
rect 15217 -1651 15269 -1642
rect 15281 -1651 15333 -1642
rect 15345 -1651 15397 -1642
rect 15409 -1651 15461 -1642
rect 15473 -1651 15525 -1642
rect 15565 -1608 15617 -1599
rect 15565 -1642 15574 -1608
rect 15574 -1642 15608 -1608
rect 15608 -1642 15617 -1608
rect 15565 -1651 15617 -1642
rect 15672 -1608 15724 -1599
rect 15672 -1642 15677 -1608
rect 15677 -1642 15711 -1608
rect 15711 -1642 15724 -1608
rect 15672 -1651 15724 -1642
rect 15736 -1608 15788 -1599
rect 15736 -1642 15749 -1608
rect 15749 -1642 15783 -1608
rect 15783 -1642 15788 -1608
rect 15736 -1651 15788 -1642
rect 15212 -1708 15264 -1699
rect 15212 -1742 15251 -1708
rect 15251 -1742 15264 -1708
rect 15212 -1751 15264 -1742
rect 14440 -1851 14492 -1799
rect 14553 -1808 14605 -1799
rect 14553 -1842 14558 -1808
rect 14558 -1842 14592 -1808
rect 14592 -1842 14605 -1808
rect 14553 -1851 14605 -1842
rect 14617 -1808 14669 -1799
rect 14617 -1842 14630 -1808
rect 14630 -1842 14664 -1808
rect 14664 -1842 14669 -1808
rect 14617 -1851 14669 -1842
rect 14725 -1808 14777 -1799
rect 14725 -1842 14734 -1808
rect 14734 -1842 14768 -1808
rect 14768 -1842 14777 -1808
rect 14725 -1851 14777 -1842
rect 14816 -1808 14868 -1799
rect 14880 -1808 14932 -1799
rect 14944 -1808 14996 -1799
rect 15008 -1808 15060 -1799
rect 15072 -1808 15124 -1799
rect 14816 -1842 14842 -1808
rect 14842 -1842 14868 -1808
rect 14880 -1842 14914 -1808
rect 14914 -1842 14932 -1808
rect 14944 -1842 14948 -1808
rect 14948 -1842 14986 -1808
rect 14986 -1842 14996 -1808
rect 15008 -1842 15020 -1808
rect 15020 -1842 15058 -1808
rect 15058 -1842 15060 -1808
rect 15072 -1842 15092 -1808
rect 15092 -1842 15124 -1808
rect 14816 -1851 14868 -1842
rect 14880 -1851 14932 -1842
rect 14944 -1851 14996 -1842
rect 15008 -1851 15060 -1842
rect 15072 -1851 15124 -1842
rect 15217 -1808 15269 -1799
rect 15281 -1808 15333 -1799
rect 15345 -1808 15397 -1799
rect 15409 -1808 15461 -1799
rect 15473 -1808 15525 -1799
rect 15217 -1842 15249 -1808
rect 15249 -1842 15269 -1808
rect 15281 -1842 15283 -1808
rect 15283 -1842 15321 -1808
rect 15321 -1842 15333 -1808
rect 15345 -1842 15355 -1808
rect 15355 -1842 15393 -1808
rect 15393 -1842 15397 -1808
rect 15409 -1842 15427 -1808
rect 15427 -1842 15461 -1808
rect 15473 -1842 15499 -1808
rect 15499 -1842 15525 -1808
rect 15217 -1851 15269 -1842
rect 15281 -1851 15333 -1842
rect 15345 -1851 15397 -1842
rect 15409 -1851 15461 -1842
rect 15473 -1851 15525 -1842
rect 15565 -1808 15617 -1799
rect 15565 -1842 15574 -1808
rect 15574 -1842 15608 -1808
rect 15608 -1842 15617 -1808
rect 15565 -1851 15617 -1842
rect 15672 -1808 15724 -1799
rect 15672 -1842 15677 -1808
rect 15677 -1842 15711 -1808
rect 15711 -1842 15724 -1808
rect 15672 -1851 15724 -1842
rect 15736 -1808 15788 -1799
rect 15736 -1842 15749 -1808
rect 15749 -1842 15783 -1808
rect 15783 -1842 15788 -1808
rect 15736 -1851 15788 -1842
rect 15212 -1908 15264 -1899
rect 15212 -1942 15251 -1908
rect 15251 -1942 15264 -1908
rect 15212 -1951 15264 -1942
rect 14440 -2051 14492 -1999
rect 14553 -2008 14605 -1999
rect 14553 -2042 14558 -2008
rect 14558 -2042 14592 -2008
rect 14592 -2042 14605 -2008
rect 14553 -2051 14605 -2042
rect 14617 -2008 14669 -1999
rect 14617 -2042 14630 -2008
rect 14630 -2042 14664 -2008
rect 14664 -2042 14669 -2008
rect 14617 -2051 14669 -2042
rect 14725 -2008 14777 -1999
rect 14725 -2042 14734 -2008
rect 14734 -2042 14768 -2008
rect 14768 -2042 14777 -2008
rect 14725 -2051 14777 -2042
rect 14816 -2008 14868 -1999
rect 14880 -2008 14932 -1999
rect 14944 -2008 14996 -1999
rect 15008 -2008 15060 -1999
rect 15072 -2008 15124 -1999
rect 14816 -2042 14842 -2008
rect 14842 -2042 14868 -2008
rect 14880 -2042 14914 -2008
rect 14914 -2042 14932 -2008
rect 14944 -2042 14948 -2008
rect 14948 -2042 14986 -2008
rect 14986 -2042 14996 -2008
rect 15008 -2042 15020 -2008
rect 15020 -2042 15058 -2008
rect 15058 -2042 15060 -2008
rect 15072 -2042 15092 -2008
rect 15092 -2042 15124 -2008
rect 14816 -2051 14868 -2042
rect 14880 -2051 14932 -2042
rect 14944 -2051 14996 -2042
rect 15008 -2051 15060 -2042
rect 15072 -2051 15124 -2042
rect 15217 -2008 15269 -1999
rect 15281 -2008 15333 -1999
rect 15345 -2008 15397 -1999
rect 15409 -2008 15461 -1999
rect 15473 -2008 15525 -1999
rect 15217 -2042 15249 -2008
rect 15249 -2042 15269 -2008
rect 15281 -2042 15283 -2008
rect 15283 -2042 15321 -2008
rect 15321 -2042 15333 -2008
rect 15345 -2042 15355 -2008
rect 15355 -2042 15393 -2008
rect 15393 -2042 15397 -2008
rect 15409 -2042 15427 -2008
rect 15427 -2042 15461 -2008
rect 15473 -2042 15499 -2008
rect 15499 -2042 15525 -2008
rect 15217 -2051 15269 -2042
rect 15281 -2051 15333 -2042
rect 15345 -2051 15397 -2042
rect 15409 -2051 15461 -2042
rect 15473 -2051 15525 -2042
rect 15565 -2008 15617 -1999
rect 15565 -2042 15574 -2008
rect 15574 -2042 15608 -2008
rect 15608 -2042 15617 -2008
rect 15565 -2051 15617 -2042
rect 15672 -2008 15724 -1999
rect 15672 -2042 15677 -2008
rect 15677 -2042 15711 -2008
rect 15711 -2042 15724 -2008
rect 15672 -2051 15724 -2042
rect 15736 -2008 15788 -1999
rect 15736 -2042 15749 -2008
rect 15749 -2042 15783 -2008
rect 15783 -2042 15788 -2008
rect 15736 -2051 15788 -2042
<< metal2 >>
rect 196 4921 274 4922
rect -4 4905 74 4906
rect -4 4849 7 4905
rect 63 4849 74 4905
rect 196 4865 207 4921
rect 263 4865 274 4921
rect 596 4921 674 4922
rect 196 4864 274 4865
rect 396 4905 474 4906
rect -4 4848 74 4849
rect 396 4849 407 4905
rect 463 4849 474 4905
rect 596 4865 607 4921
rect 663 4865 674 4921
rect 996 4921 1074 4922
rect 596 4864 674 4865
rect 796 4905 874 4906
rect 396 4848 474 4849
rect 796 4849 807 4905
rect 863 4849 874 4905
rect 996 4865 1007 4921
rect 1063 4865 1074 4921
rect 1396 4921 1474 4922
rect 996 4864 1074 4865
rect 1196 4905 1274 4906
rect 796 4848 874 4849
rect 1196 4849 1207 4905
rect 1263 4849 1274 4905
rect 1396 4865 1407 4921
rect 1463 4865 1474 4921
rect 1796 4921 1874 4922
rect 1396 4864 1474 4865
rect 1596 4905 1674 4906
rect 1196 4848 1274 4849
rect 1596 4849 1607 4905
rect 1663 4849 1674 4905
rect 1796 4865 1807 4921
rect 1863 4865 1874 4921
rect 2196 4921 2274 4922
rect 1796 4864 1874 4865
rect 1996 4905 2074 4906
rect 1596 4848 1674 4849
rect 1996 4849 2007 4905
rect 2063 4849 2074 4905
rect 2196 4865 2207 4921
rect 2263 4865 2274 4921
rect 2596 4921 2674 4922
rect 2196 4864 2274 4865
rect 2396 4905 2474 4906
rect 1996 4848 2074 4849
rect 2396 4849 2407 4905
rect 2463 4849 2474 4905
rect 2596 4865 2607 4921
rect 2663 4865 2674 4921
rect 2996 4921 3074 4922
rect 2596 4864 2674 4865
rect 2796 4905 2874 4906
rect 2396 4848 2474 4849
rect 2796 4849 2807 4905
rect 2863 4849 2874 4905
rect 2996 4865 3007 4921
rect 3063 4865 3074 4921
rect 3396 4921 3474 4922
rect 2996 4864 3074 4865
rect 3196 4905 3274 4906
rect 2796 4848 2874 4849
rect 3196 4849 3207 4905
rect 3263 4849 3274 4905
rect 3396 4865 3407 4921
rect 3463 4865 3474 4921
rect 3796 4921 3874 4922
rect 3396 4864 3474 4865
rect 3596 4905 3674 4906
rect 3196 4848 3274 4849
rect 3596 4849 3607 4905
rect 3663 4849 3674 4905
rect 3796 4865 3807 4921
rect 3863 4865 3874 4921
rect 4196 4921 4274 4922
rect 3796 4864 3874 4865
rect 3996 4905 4074 4906
rect 3596 4848 3674 4849
rect 3996 4849 4007 4905
rect 4063 4849 4074 4905
rect 4196 4865 4207 4921
rect 4263 4865 4274 4921
rect 4596 4921 4674 4922
rect 4196 4864 4274 4865
rect 4396 4905 4474 4906
rect 3996 4848 4074 4849
rect 4396 4849 4407 4905
rect 4463 4849 4474 4905
rect 4596 4865 4607 4921
rect 4663 4865 4674 4921
rect 4996 4921 5074 4922
rect 4596 4864 4674 4865
rect 4796 4905 4874 4906
rect 4396 4848 4474 4849
rect 4796 4849 4807 4905
rect 4863 4849 4874 4905
rect 4996 4865 5007 4921
rect 5063 4865 5074 4921
rect 5396 4921 5474 4922
rect 4996 4864 5074 4865
rect 5196 4905 5274 4906
rect 4796 4848 4874 4849
rect 5196 4849 5207 4905
rect 5263 4849 5274 4905
rect 5396 4865 5407 4921
rect 5463 4865 5474 4921
rect 5796 4921 5874 4922
rect 5396 4864 5474 4865
rect 5596 4905 5674 4906
rect 5196 4848 5274 4849
rect 5596 4849 5607 4905
rect 5663 4849 5674 4905
rect 5796 4865 5807 4921
rect 5863 4865 5874 4921
rect 6196 4921 6274 4922
rect 5796 4864 5874 4865
rect 5996 4905 6074 4906
rect 5596 4848 5674 4849
rect 5996 4849 6007 4905
rect 6063 4849 6074 4905
rect 6196 4865 6207 4921
rect 6263 4865 6274 4921
rect 6596 4921 6674 4922
rect 6196 4864 6274 4865
rect 6396 4905 6474 4906
rect 5996 4848 6074 4849
rect 6396 4849 6407 4905
rect 6463 4849 6474 4905
rect 6596 4865 6607 4921
rect 6663 4865 6674 4921
rect 6996 4921 7074 4922
rect 6596 4864 6674 4865
rect 6796 4905 6874 4906
rect 6396 4848 6474 4849
rect 6796 4849 6807 4905
rect 6863 4849 6874 4905
rect 6996 4865 7007 4921
rect 7063 4865 7074 4921
rect 7396 4921 7474 4922
rect 6996 4864 7074 4865
rect 7196 4905 7274 4906
rect 6796 4848 6874 4849
rect 7196 4849 7207 4905
rect 7263 4849 7274 4905
rect 7396 4865 7407 4921
rect 7463 4865 7474 4921
rect 7796 4921 7874 4922
rect 7396 4864 7474 4865
rect 7596 4905 7674 4906
rect 7196 4848 7274 4849
rect 7596 4849 7607 4905
rect 7663 4849 7674 4905
rect 7796 4865 7807 4921
rect 7863 4865 7874 4921
rect 8196 4921 8274 4922
rect 7796 4864 7874 4865
rect 7996 4905 8074 4906
rect 7596 4848 7674 4849
rect 7996 4849 8007 4905
rect 8063 4849 8074 4905
rect 8196 4865 8207 4921
rect 8263 4865 8274 4921
rect 8596 4921 8674 4922
rect 8196 4864 8274 4865
rect 8396 4905 8474 4906
rect 7996 4848 8074 4849
rect 8396 4849 8407 4905
rect 8463 4849 8474 4905
rect 8596 4865 8607 4921
rect 8663 4865 8674 4921
rect 8996 4921 9074 4922
rect 8596 4864 8674 4865
rect 8796 4905 8874 4906
rect 8396 4848 8474 4849
rect 8796 4849 8807 4905
rect 8863 4849 8874 4905
rect 8996 4865 9007 4921
rect 9063 4865 9074 4921
rect 9396 4921 9474 4922
rect 8996 4864 9074 4865
rect 9196 4905 9274 4906
rect 8796 4848 8874 4849
rect 9196 4849 9207 4905
rect 9263 4849 9274 4905
rect 9396 4865 9407 4921
rect 9463 4865 9474 4921
rect 9796 4921 9874 4922
rect 9396 4864 9474 4865
rect 9596 4905 9674 4906
rect 9196 4848 9274 4849
rect 9596 4849 9607 4905
rect 9663 4849 9674 4905
rect 9796 4865 9807 4921
rect 9863 4865 9874 4921
rect 10196 4921 10274 4922
rect 9796 4864 9874 4865
rect 9996 4905 10074 4906
rect 9596 4848 9674 4849
rect 9996 4849 10007 4905
rect 10063 4849 10074 4905
rect 10196 4865 10207 4921
rect 10263 4865 10274 4921
rect 10596 4921 10674 4922
rect 10196 4864 10274 4865
rect 10396 4905 10474 4906
rect 9996 4848 10074 4849
rect 10396 4849 10407 4905
rect 10463 4849 10474 4905
rect 10596 4865 10607 4921
rect 10663 4865 10674 4921
rect 10996 4921 11074 4922
rect 10596 4864 10674 4865
rect 10796 4905 10874 4906
rect 10396 4848 10474 4849
rect 10796 4849 10807 4905
rect 10863 4849 10874 4905
rect 10996 4865 11007 4921
rect 11063 4865 11074 4921
rect 11396 4921 11474 4922
rect 10996 4864 11074 4865
rect 11196 4905 11274 4906
rect 10796 4848 10874 4849
rect 11196 4849 11207 4905
rect 11263 4849 11274 4905
rect 11396 4865 11407 4921
rect 11463 4865 11474 4921
rect 11796 4921 11874 4922
rect 11396 4864 11474 4865
rect 11596 4905 11674 4906
rect 11196 4848 11274 4849
rect 11596 4849 11607 4905
rect 11663 4849 11674 4905
rect 11796 4865 11807 4921
rect 11863 4865 11874 4921
rect 12196 4921 12274 4922
rect 11796 4864 11874 4865
rect 11996 4905 12074 4906
rect 11596 4848 11674 4849
rect 11996 4849 12007 4905
rect 12063 4849 12074 4905
rect 12196 4865 12207 4921
rect 12263 4865 12274 4921
rect 12596 4921 12674 4922
rect 12196 4864 12274 4865
rect 12396 4905 12474 4906
rect 11996 4848 12074 4849
rect 12396 4849 12407 4905
rect 12463 4849 12474 4905
rect 12596 4865 12607 4921
rect 12663 4865 12674 4921
rect 12596 4864 12674 4865
rect 12396 4848 12474 4849
rect 202 4831 268 4832
rect 202 4820 209 4831
rect 0 4790 209 4820
rect 202 4779 209 4790
rect 261 4820 268 4831
rect 602 4831 668 4832
rect 602 4820 609 4831
rect 261 4790 609 4820
rect 261 4779 268 4790
rect 202 4778 268 4779
rect 602 4779 609 4790
rect 661 4820 668 4831
rect 1002 4831 1068 4832
rect 1002 4820 1009 4831
rect 661 4790 1009 4820
rect 661 4779 668 4790
rect 602 4778 668 4779
rect 1002 4779 1009 4790
rect 1061 4820 1068 4831
rect 1402 4831 1468 4832
rect 1402 4820 1409 4831
rect 1061 4790 1409 4820
rect 1061 4779 1068 4790
rect 1002 4778 1068 4779
rect 1402 4779 1409 4790
rect 1461 4820 1468 4831
rect 1802 4831 1868 4832
rect 1802 4820 1809 4831
rect 1461 4790 1809 4820
rect 1461 4779 1468 4790
rect 1402 4778 1468 4779
rect 1802 4779 1809 4790
rect 1861 4820 1868 4831
rect 2202 4831 2268 4832
rect 2202 4820 2209 4831
rect 1861 4790 2209 4820
rect 1861 4779 1868 4790
rect 1802 4778 1868 4779
rect 2202 4779 2209 4790
rect 2261 4820 2268 4831
rect 2602 4831 2668 4832
rect 2602 4820 2609 4831
rect 2261 4790 2609 4820
rect 2261 4779 2268 4790
rect 2202 4778 2268 4779
rect 2602 4779 2609 4790
rect 2661 4820 2668 4831
rect 3002 4831 3068 4832
rect 3002 4820 3009 4831
rect 2661 4790 3009 4820
rect 2661 4779 2668 4790
rect 2602 4778 2668 4779
rect 3002 4779 3009 4790
rect 3061 4820 3068 4831
rect 3402 4831 3468 4832
rect 3402 4820 3409 4831
rect 3061 4790 3409 4820
rect 3061 4779 3068 4790
rect 3002 4778 3068 4779
rect 3402 4779 3409 4790
rect 3461 4820 3468 4831
rect 3802 4831 3868 4832
rect 3802 4820 3809 4831
rect 3461 4790 3809 4820
rect 3461 4779 3468 4790
rect 3402 4778 3468 4779
rect 3802 4779 3809 4790
rect 3861 4820 3868 4831
rect 4202 4831 4268 4832
rect 4202 4820 4209 4831
rect 3861 4790 4209 4820
rect 3861 4779 3868 4790
rect 3802 4778 3868 4779
rect 4202 4779 4209 4790
rect 4261 4820 4268 4831
rect 4602 4831 4668 4832
rect 4602 4820 4609 4831
rect 4261 4790 4609 4820
rect 4261 4779 4268 4790
rect 4202 4778 4268 4779
rect 4602 4779 4609 4790
rect 4661 4820 4668 4831
rect 5002 4831 5068 4832
rect 5002 4820 5009 4831
rect 4661 4790 5009 4820
rect 4661 4779 4668 4790
rect 4602 4778 4668 4779
rect 5002 4779 5009 4790
rect 5061 4820 5068 4831
rect 5402 4831 5468 4832
rect 5402 4820 5409 4831
rect 5061 4790 5409 4820
rect 5061 4779 5068 4790
rect 5002 4778 5068 4779
rect 5402 4779 5409 4790
rect 5461 4820 5468 4831
rect 5802 4831 5868 4832
rect 5802 4820 5809 4831
rect 5461 4790 5809 4820
rect 5461 4779 5468 4790
rect 5402 4778 5468 4779
rect 5802 4779 5809 4790
rect 5861 4820 5868 4831
rect 6202 4831 6268 4832
rect 6202 4820 6209 4831
rect 5861 4790 6209 4820
rect 5861 4779 5868 4790
rect 5802 4778 5868 4779
rect 6202 4779 6209 4790
rect 6261 4820 6268 4831
rect 6602 4831 6668 4832
rect 6602 4820 6609 4831
rect 6261 4790 6609 4820
rect 6261 4779 6268 4790
rect 6202 4778 6268 4779
rect 6602 4779 6609 4790
rect 6661 4820 6668 4831
rect 7002 4831 7068 4832
rect 7002 4820 7009 4831
rect 6661 4790 7009 4820
rect 6661 4779 6668 4790
rect 6602 4778 6668 4779
rect 7002 4779 7009 4790
rect 7061 4820 7068 4831
rect 7402 4831 7468 4832
rect 7402 4820 7409 4831
rect 7061 4790 7409 4820
rect 7061 4779 7068 4790
rect 7002 4778 7068 4779
rect 7402 4779 7409 4790
rect 7461 4820 7468 4831
rect 7802 4831 7868 4832
rect 7802 4820 7809 4831
rect 7461 4790 7809 4820
rect 7461 4779 7468 4790
rect 7402 4778 7468 4779
rect 7802 4779 7809 4790
rect 7861 4820 7868 4831
rect 8202 4831 8268 4832
rect 8202 4820 8209 4831
rect 7861 4790 8209 4820
rect 7861 4779 7868 4790
rect 7802 4778 7868 4779
rect 8202 4779 8209 4790
rect 8261 4820 8268 4831
rect 8602 4831 8668 4832
rect 8602 4820 8609 4831
rect 8261 4790 8609 4820
rect 8261 4779 8268 4790
rect 8202 4778 8268 4779
rect 8602 4779 8609 4790
rect 8661 4820 8668 4831
rect 9002 4831 9068 4832
rect 9002 4820 9009 4831
rect 8661 4790 9009 4820
rect 8661 4779 8668 4790
rect 8602 4778 8668 4779
rect 9002 4779 9009 4790
rect 9061 4820 9068 4831
rect 9402 4831 9468 4832
rect 9402 4820 9409 4831
rect 9061 4790 9409 4820
rect 9061 4779 9068 4790
rect 9002 4778 9068 4779
rect 9402 4779 9409 4790
rect 9461 4820 9468 4831
rect 9802 4831 9868 4832
rect 9802 4820 9809 4831
rect 9461 4790 9809 4820
rect 9461 4779 9468 4790
rect 9402 4778 9468 4779
rect 9802 4779 9809 4790
rect 9861 4820 9868 4831
rect 10202 4831 10268 4832
rect 10202 4820 10209 4831
rect 9861 4790 10209 4820
rect 9861 4779 9868 4790
rect 9802 4778 9868 4779
rect 10202 4779 10209 4790
rect 10261 4820 10268 4831
rect 10602 4831 10668 4832
rect 10602 4820 10609 4831
rect 10261 4790 10609 4820
rect 10261 4779 10268 4790
rect 10202 4778 10268 4779
rect 10602 4779 10609 4790
rect 10661 4820 10668 4831
rect 11002 4831 11068 4832
rect 11002 4820 11009 4831
rect 10661 4790 11009 4820
rect 10661 4779 10668 4790
rect 10602 4778 10668 4779
rect 11002 4779 11009 4790
rect 11061 4820 11068 4831
rect 11402 4831 11468 4832
rect 11402 4820 11409 4831
rect 11061 4790 11409 4820
rect 11061 4779 11068 4790
rect 11002 4778 11068 4779
rect 11402 4779 11409 4790
rect 11461 4820 11468 4831
rect 11802 4831 11868 4832
rect 11802 4820 11809 4831
rect 11461 4790 11809 4820
rect 11461 4779 11468 4790
rect 11402 4778 11468 4779
rect 11802 4779 11809 4790
rect 11861 4820 11868 4831
rect 12202 4831 12268 4832
rect 12202 4820 12209 4831
rect 11861 4790 12209 4820
rect 11861 4779 11868 4790
rect 11802 4778 11868 4779
rect 12202 4779 12209 4790
rect 12261 4820 12268 4831
rect 12602 4831 12668 4832
rect 12602 4820 12609 4831
rect 12261 4790 12609 4820
rect 12261 4779 12268 4790
rect 12202 4778 12268 4779
rect 12602 4779 12609 4790
rect 12661 4820 12668 4831
rect 13104 4831 13170 4832
rect 13104 4820 13111 4831
rect 12661 4790 13111 4820
rect 12661 4779 12668 4790
rect 12602 4778 12668 4779
rect 13104 4779 13111 4790
rect 13163 4779 13170 4831
rect 13104 4778 13170 4779
rect 2 4761 68 4762
rect 2 4750 9 4761
rect 0 4720 9 4750
rect 2 4709 9 4720
rect 61 4750 68 4761
rect 402 4761 468 4762
rect 402 4750 409 4761
rect 61 4720 409 4750
rect 61 4709 68 4720
rect 2 4708 68 4709
rect 402 4709 409 4720
rect 461 4750 468 4761
rect 802 4761 868 4762
rect 802 4750 809 4761
rect 461 4720 809 4750
rect 461 4709 468 4720
rect 402 4708 468 4709
rect 802 4709 809 4720
rect 861 4750 868 4761
rect 1202 4761 1268 4762
rect 1202 4750 1209 4761
rect 861 4720 1209 4750
rect 861 4709 868 4720
rect 802 4708 868 4709
rect 1202 4709 1209 4720
rect 1261 4750 1268 4761
rect 1602 4761 1668 4762
rect 1602 4750 1609 4761
rect 1261 4720 1609 4750
rect 1261 4709 1268 4720
rect 1202 4708 1268 4709
rect 1602 4709 1609 4720
rect 1661 4750 1668 4761
rect 2002 4761 2068 4762
rect 2002 4750 2009 4761
rect 1661 4720 2009 4750
rect 1661 4709 1668 4720
rect 1602 4708 1668 4709
rect 2002 4709 2009 4720
rect 2061 4750 2068 4761
rect 2402 4761 2468 4762
rect 2402 4750 2409 4761
rect 2061 4720 2409 4750
rect 2061 4709 2068 4720
rect 2002 4708 2068 4709
rect 2402 4709 2409 4720
rect 2461 4750 2468 4761
rect 2802 4761 2868 4762
rect 2802 4750 2809 4761
rect 2461 4720 2809 4750
rect 2461 4709 2468 4720
rect 2402 4708 2468 4709
rect 2802 4709 2809 4720
rect 2861 4750 2868 4761
rect 3202 4761 3268 4762
rect 3202 4750 3209 4761
rect 2861 4720 3209 4750
rect 2861 4709 2868 4720
rect 2802 4708 2868 4709
rect 3202 4709 3209 4720
rect 3261 4750 3268 4761
rect 3602 4761 3668 4762
rect 3602 4750 3609 4761
rect 3261 4720 3609 4750
rect 3261 4709 3268 4720
rect 3202 4708 3268 4709
rect 3602 4709 3609 4720
rect 3661 4750 3668 4761
rect 4002 4761 4068 4762
rect 4002 4750 4009 4761
rect 3661 4720 4009 4750
rect 3661 4709 3668 4720
rect 3602 4708 3668 4709
rect 4002 4709 4009 4720
rect 4061 4750 4068 4761
rect 4402 4761 4468 4762
rect 4402 4750 4409 4761
rect 4061 4720 4409 4750
rect 4061 4709 4068 4720
rect 4002 4708 4068 4709
rect 4402 4709 4409 4720
rect 4461 4750 4468 4761
rect 4802 4761 4868 4762
rect 4802 4750 4809 4761
rect 4461 4720 4809 4750
rect 4461 4709 4468 4720
rect 4402 4708 4468 4709
rect 4802 4709 4809 4720
rect 4861 4750 4868 4761
rect 5202 4761 5268 4762
rect 5202 4750 5209 4761
rect 4861 4720 5209 4750
rect 4861 4709 4868 4720
rect 4802 4708 4868 4709
rect 5202 4709 5209 4720
rect 5261 4750 5268 4761
rect 5602 4761 5668 4762
rect 5602 4750 5609 4761
rect 5261 4720 5609 4750
rect 5261 4709 5268 4720
rect 5202 4708 5268 4709
rect 5602 4709 5609 4720
rect 5661 4750 5668 4761
rect 6002 4761 6068 4762
rect 6002 4750 6009 4761
rect 5661 4720 6009 4750
rect 5661 4709 5668 4720
rect 5602 4708 5668 4709
rect 6002 4709 6009 4720
rect 6061 4750 6068 4761
rect 6402 4761 6468 4762
rect 6402 4750 6409 4761
rect 6061 4720 6409 4750
rect 6061 4709 6068 4720
rect 6002 4708 6068 4709
rect 6402 4709 6409 4720
rect 6461 4750 6468 4761
rect 6802 4761 6868 4762
rect 6802 4750 6809 4761
rect 6461 4720 6809 4750
rect 6461 4709 6468 4720
rect 6402 4708 6468 4709
rect 6802 4709 6809 4720
rect 6861 4750 6868 4761
rect 7202 4761 7268 4762
rect 7202 4750 7209 4761
rect 6861 4720 7209 4750
rect 6861 4709 6868 4720
rect 6802 4708 6868 4709
rect 7202 4709 7209 4720
rect 7261 4750 7268 4761
rect 7602 4761 7668 4762
rect 7602 4750 7609 4761
rect 7261 4720 7609 4750
rect 7261 4709 7268 4720
rect 7202 4708 7268 4709
rect 7602 4709 7609 4720
rect 7661 4750 7668 4761
rect 8002 4761 8068 4762
rect 8002 4750 8009 4761
rect 7661 4720 8009 4750
rect 7661 4709 7668 4720
rect 7602 4708 7668 4709
rect 8002 4709 8009 4720
rect 8061 4750 8068 4761
rect 8402 4761 8468 4762
rect 8402 4750 8409 4761
rect 8061 4720 8409 4750
rect 8061 4709 8068 4720
rect 8002 4708 8068 4709
rect 8402 4709 8409 4720
rect 8461 4750 8468 4761
rect 8802 4761 8868 4762
rect 8802 4750 8809 4761
rect 8461 4720 8809 4750
rect 8461 4709 8468 4720
rect 8402 4708 8468 4709
rect 8802 4709 8809 4720
rect 8861 4750 8868 4761
rect 9202 4761 9268 4762
rect 9202 4750 9209 4761
rect 8861 4720 9209 4750
rect 8861 4709 8868 4720
rect 8802 4708 8868 4709
rect 9202 4709 9209 4720
rect 9261 4750 9268 4761
rect 9602 4761 9668 4762
rect 9602 4750 9609 4761
rect 9261 4720 9609 4750
rect 9261 4709 9268 4720
rect 9202 4708 9268 4709
rect 9602 4709 9609 4720
rect 9661 4750 9668 4761
rect 10002 4761 10068 4762
rect 10002 4750 10009 4761
rect 9661 4720 10009 4750
rect 9661 4709 9668 4720
rect 9602 4708 9668 4709
rect 10002 4709 10009 4720
rect 10061 4750 10068 4761
rect 10402 4761 10468 4762
rect 10402 4750 10409 4761
rect 10061 4720 10409 4750
rect 10061 4709 10068 4720
rect 10002 4708 10068 4709
rect 10402 4709 10409 4720
rect 10461 4750 10468 4761
rect 10802 4761 10868 4762
rect 10802 4750 10809 4761
rect 10461 4720 10809 4750
rect 10461 4709 10468 4720
rect 10402 4708 10468 4709
rect 10802 4709 10809 4720
rect 10861 4750 10868 4761
rect 11202 4761 11268 4762
rect 11202 4750 11209 4761
rect 10861 4720 11209 4750
rect 10861 4709 10868 4720
rect 10802 4708 10868 4709
rect 11202 4709 11209 4720
rect 11261 4750 11268 4761
rect 11602 4761 11668 4762
rect 11602 4750 11609 4761
rect 11261 4720 11609 4750
rect 11261 4709 11268 4720
rect 11202 4708 11268 4709
rect 11602 4709 11609 4720
rect 11661 4750 11668 4761
rect 12002 4761 12068 4762
rect 12002 4750 12009 4761
rect 11661 4720 12009 4750
rect 11661 4709 11668 4720
rect 11602 4708 11668 4709
rect 12002 4709 12009 4720
rect 12061 4750 12068 4761
rect 12402 4761 12468 4762
rect 12402 4750 12409 4761
rect 12061 4720 12409 4750
rect 12061 4709 12068 4720
rect 12002 4708 12068 4709
rect 12402 4709 12409 4720
rect 12461 4750 12468 4761
rect 12802 4761 12868 4762
rect 12802 4750 12809 4761
rect 12461 4720 12809 4750
rect 12461 4709 12468 4720
rect 12402 4708 12468 4709
rect 12802 4709 12809 4720
rect 12861 4750 12868 4761
rect 12900 4761 12966 4762
rect 12900 4750 12907 4761
rect 12861 4720 12907 4750
rect 12861 4709 12868 4720
rect 12802 4708 12868 4709
rect 12900 4709 12907 4720
rect 12959 4709 12966 4761
rect 12900 4708 12966 4709
rect 202 4691 268 4692
rect 202 4680 209 4691
rect 0 4650 209 4680
rect 202 4639 209 4650
rect 261 4680 268 4691
rect 602 4691 668 4692
rect 602 4680 609 4691
rect 261 4650 609 4680
rect 261 4639 268 4650
rect 202 4638 268 4639
rect 602 4639 609 4650
rect 661 4680 668 4691
rect 1002 4691 1068 4692
rect 1002 4680 1009 4691
rect 661 4650 1009 4680
rect 661 4639 668 4650
rect 602 4638 668 4639
rect 1002 4639 1009 4650
rect 1061 4680 1068 4691
rect 1402 4691 1468 4692
rect 1402 4680 1409 4691
rect 1061 4650 1409 4680
rect 1061 4639 1068 4650
rect 1002 4638 1068 4639
rect 1402 4639 1409 4650
rect 1461 4680 1468 4691
rect 1802 4691 1868 4692
rect 1802 4680 1809 4691
rect 1461 4650 1809 4680
rect 1461 4639 1468 4650
rect 1402 4638 1468 4639
rect 1802 4639 1809 4650
rect 1861 4680 1868 4691
rect 2202 4691 2268 4692
rect 2202 4680 2209 4691
rect 1861 4650 2209 4680
rect 1861 4639 1868 4650
rect 1802 4638 1868 4639
rect 2202 4639 2209 4650
rect 2261 4680 2268 4691
rect 2602 4691 2668 4692
rect 2602 4680 2609 4691
rect 2261 4650 2609 4680
rect 2261 4639 2268 4650
rect 2202 4638 2268 4639
rect 2602 4639 2609 4650
rect 2661 4680 2668 4691
rect 3002 4691 3068 4692
rect 3002 4680 3009 4691
rect 2661 4650 3009 4680
rect 2661 4639 2668 4650
rect 2602 4638 2668 4639
rect 3002 4639 3009 4650
rect 3061 4680 3068 4691
rect 3402 4691 3468 4692
rect 3402 4680 3409 4691
rect 3061 4650 3409 4680
rect 3061 4639 3068 4650
rect 3002 4638 3068 4639
rect 3402 4639 3409 4650
rect 3461 4680 3468 4691
rect 3802 4691 3868 4692
rect 3802 4680 3809 4691
rect 3461 4650 3809 4680
rect 3461 4639 3468 4650
rect 3402 4638 3468 4639
rect 3802 4639 3809 4650
rect 3861 4680 3868 4691
rect 4202 4691 4268 4692
rect 4202 4680 4209 4691
rect 3861 4650 4209 4680
rect 3861 4639 3868 4650
rect 3802 4638 3868 4639
rect 4202 4639 4209 4650
rect 4261 4680 4268 4691
rect 4602 4691 4668 4692
rect 4602 4680 4609 4691
rect 4261 4650 4609 4680
rect 4261 4639 4268 4650
rect 4202 4638 4268 4639
rect 4602 4639 4609 4650
rect 4661 4680 4668 4691
rect 5002 4691 5068 4692
rect 5002 4680 5009 4691
rect 4661 4650 5009 4680
rect 4661 4639 4668 4650
rect 4602 4638 4668 4639
rect 5002 4639 5009 4650
rect 5061 4680 5068 4691
rect 5402 4691 5468 4692
rect 5402 4680 5409 4691
rect 5061 4650 5409 4680
rect 5061 4639 5068 4650
rect 5002 4638 5068 4639
rect 5402 4639 5409 4650
rect 5461 4680 5468 4691
rect 5802 4691 5868 4692
rect 5802 4680 5809 4691
rect 5461 4650 5809 4680
rect 5461 4639 5468 4650
rect 5402 4638 5468 4639
rect 5802 4639 5809 4650
rect 5861 4680 5868 4691
rect 6202 4691 6268 4692
rect 6202 4680 6209 4691
rect 5861 4650 6209 4680
rect 5861 4639 5868 4650
rect 5802 4638 5868 4639
rect 6202 4639 6209 4650
rect 6261 4680 6268 4691
rect 6602 4691 6668 4692
rect 6602 4680 6609 4691
rect 6261 4650 6609 4680
rect 6261 4639 6268 4650
rect 6202 4638 6268 4639
rect 6602 4639 6609 4650
rect 6661 4680 6668 4691
rect 7002 4691 7068 4692
rect 7002 4680 7009 4691
rect 6661 4650 7009 4680
rect 6661 4639 6668 4650
rect 6602 4638 6668 4639
rect 7002 4639 7009 4650
rect 7061 4680 7068 4691
rect 7402 4691 7468 4692
rect 7402 4680 7409 4691
rect 7061 4650 7409 4680
rect 7061 4639 7068 4650
rect 7002 4638 7068 4639
rect 7402 4639 7409 4650
rect 7461 4680 7468 4691
rect 7802 4691 7868 4692
rect 7802 4680 7809 4691
rect 7461 4650 7809 4680
rect 7461 4639 7468 4650
rect 7402 4638 7468 4639
rect 7802 4639 7809 4650
rect 7861 4680 7868 4691
rect 8202 4691 8268 4692
rect 8202 4680 8209 4691
rect 7861 4650 8209 4680
rect 7861 4639 7868 4650
rect 7802 4638 7868 4639
rect 8202 4639 8209 4650
rect 8261 4680 8268 4691
rect 8602 4691 8668 4692
rect 8602 4680 8609 4691
rect 8261 4650 8609 4680
rect 8261 4639 8268 4650
rect 8202 4638 8268 4639
rect 8602 4639 8609 4650
rect 8661 4680 8668 4691
rect 9002 4691 9068 4692
rect 9002 4680 9009 4691
rect 8661 4650 9009 4680
rect 8661 4639 8668 4650
rect 8602 4638 8668 4639
rect 9002 4639 9009 4650
rect 9061 4680 9068 4691
rect 9402 4691 9468 4692
rect 9402 4680 9409 4691
rect 9061 4650 9409 4680
rect 9061 4639 9068 4650
rect 9002 4638 9068 4639
rect 9402 4639 9409 4650
rect 9461 4680 9468 4691
rect 9802 4691 9868 4692
rect 9802 4680 9809 4691
rect 9461 4650 9809 4680
rect 9461 4639 9468 4650
rect 9402 4638 9468 4639
rect 9802 4639 9809 4650
rect 9861 4680 9868 4691
rect 10202 4691 10268 4692
rect 10202 4680 10209 4691
rect 9861 4650 10209 4680
rect 9861 4639 9868 4650
rect 9802 4638 9868 4639
rect 10202 4639 10209 4650
rect 10261 4680 10268 4691
rect 10602 4691 10668 4692
rect 10602 4680 10609 4691
rect 10261 4650 10609 4680
rect 10261 4639 10268 4650
rect 10202 4638 10268 4639
rect 10602 4639 10609 4650
rect 10661 4680 10668 4691
rect 11002 4691 11068 4692
rect 11002 4680 11009 4691
rect 10661 4650 11009 4680
rect 10661 4639 10668 4650
rect 10602 4638 10668 4639
rect 11002 4639 11009 4650
rect 11061 4680 11068 4691
rect 11402 4691 11468 4692
rect 11402 4680 11409 4691
rect 11061 4650 11409 4680
rect 11061 4639 11068 4650
rect 11002 4638 11068 4639
rect 11402 4639 11409 4650
rect 11461 4680 11468 4691
rect 11802 4691 11868 4692
rect 11802 4680 11809 4691
rect 11461 4650 11809 4680
rect 11461 4639 11468 4650
rect 11402 4638 11468 4639
rect 11802 4639 11809 4650
rect 11861 4680 11868 4691
rect 12202 4691 12268 4692
rect 12202 4680 12209 4691
rect 11861 4650 12209 4680
rect 11861 4639 11868 4650
rect 11802 4638 11868 4639
rect 12202 4639 12209 4650
rect 12261 4680 12268 4691
rect 12602 4691 12668 4692
rect 12602 4680 12609 4691
rect 12261 4650 12609 4680
rect 12261 4639 12268 4650
rect 12202 4638 12268 4639
rect 12602 4639 12609 4650
rect 12661 4680 12668 4691
rect 13104 4691 13170 4692
rect 13104 4680 13111 4691
rect 12661 4650 13111 4680
rect 12661 4639 12668 4650
rect 12602 4638 12668 4639
rect 13104 4639 13111 4650
rect 13163 4639 13170 4691
rect 13104 4638 13170 4639
rect 2 4621 68 4622
rect 2 4610 9 4621
rect 0 4580 9 4610
rect 2 4569 9 4580
rect 61 4610 68 4621
rect 402 4621 468 4622
rect 402 4610 409 4621
rect 61 4580 409 4610
rect 61 4569 68 4580
rect 2 4568 68 4569
rect 402 4569 409 4580
rect 461 4610 468 4621
rect 802 4621 868 4622
rect 802 4610 809 4621
rect 461 4580 809 4610
rect 461 4569 468 4580
rect 402 4568 468 4569
rect 802 4569 809 4580
rect 861 4610 868 4621
rect 1202 4621 1268 4622
rect 1202 4610 1209 4621
rect 861 4580 1209 4610
rect 861 4569 868 4580
rect 802 4568 868 4569
rect 1202 4569 1209 4580
rect 1261 4610 1268 4621
rect 1602 4621 1668 4622
rect 1602 4610 1609 4621
rect 1261 4580 1609 4610
rect 1261 4569 1268 4580
rect 1202 4568 1268 4569
rect 1602 4569 1609 4580
rect 1661 4610 1668 4621
rect 2002 4621 2068 4622
rect 2002 4610 2009 4621
rect 1661 4580 2009 4610
rect 1661 4569 1668 4580
rect 1602 4568 1668 4569
rect 2002 4569 2009 4580
rect 2061 4610 2068 4621
rect 2402 4621 2468 4622
rect 2402 4610 2409 4621
rect 2061 4580 2409 4610
rect 2061 4569 2068 4580
rect 2002 4568 2068 4569
rect 2402 4569 2409 4580
rect 2461 4610 2468 4621
rect 2802 4621 2868 4622
rect 2802 4610 2809 4621
rect 2461 4580 2809 4610
rect 2461 4569 2468 4580
rect 2402 4568 2468 4569
rect 2802 4569 2809 4580
rect 2861 4610 2868 4621
rect 3202 4621 3268 4622
rect 3202 4610 3209 4621
rect 2861 4580 3209 4610
rect 2861 4569 2868 4580
rect 2802 4568 2868 4569
rect 3202 4569 3209 4580
rect 3261 4610 3268 4621
rect 3602 4621 3668 4622
rect 3602 4610 3609 4621
rect 3261 4580 3609 4610
rect 3261 4569 3268 4580
rect 3202 4568 3268 4569
rect 3602 4569 3609 4580
rect 3661 4610 3668 4621
rect 4002 4621 4068 4622
rect 4002 4610 4009 4621
rect 3661 4580 4009 4610
rect 3661 4569 3668 4580
rect 3602 4568 3668 4569
rect 4002 4569 4009 4580
rect 4061 4610 4068 4621
rect 4402 4621 4468 4622
rect 4402 4610 4409 4621
rect 4061 4580 4409 4610
rect 4061 4569 4068 4580
rect 4002 4568 4068 4569
rect 4402 4569 4409 4580
rect 4461 4610 4468 4621
rect 4802 4621 4868 4622
rect 4802 4610 4809 4621
rect 4461 4580 4809 4610
rect 4461 4569 4468 4580
rect 4402 4568 4468 4569
rect 4802 4569 4809 4580
rect 4861 4610 4868 4621
rect 5202 4621 5268 4622
rect 5202 4610 5209 4621
rect 4861 4580 5209 4610
rect 4861 4569 4868 4580
rect 4802 4568 4868 4569
rect 5202 4569 5209 4580
rect 5261 4610 5268 4621
rect 5602 4621 5668 4622
rect 5602 4610 5609 4621
rect 5261 4580 5609 4610
rect 5261 4569 5268 4580
rect 5202 4568 5268 4569
rect 5602 4569 5609 4580
rect 5661 4610 5668 4621
rect 6002 4621 6068 4622
rect 6002 4610 6009 4621
rect 5661 4580 6009 4610
rect 5661 4569 5668 4580
rect 5602 4568 5668 4569
rect 6002 4569 6009 4580
rect 6061 4610 6068 4621
rect 6402 4621 6468 4622
rect 6402 4610 6409 4621
rect 6061 4580 6409 4610
rect 6061 4569 6068 4580
rect 6002 4568 6068 4569
rect 6402 4569 6409 4580
rect 6461 4610 6468 4621
rect 6802 4621 6868 4622
rect 6802 4610 6809 4621
rect 6461 4580 6809 4610
rect 6461 4569 6468 4580
rect 6402 4568 6468 4569
rect 6802 4569 6809 4580
rect 6861 4610 6868 4621
rect 7202 4621 7268 4622
rect 7202 4610 7209 4621
rect 6861 4580 7209 4610
rect 6861 4569 6868 4580
rect 6802 4568 6868 4569
rect 7202 4569 7209 4580
rect 7261 4610 7268 4621
rect 7602 4621 7668 4622
rect 7602 4610 7609 4621
rect 7261 4580 7609 4610
rect 7261 4569 7268 4580
rect 7202 4568 7268 4569
rect 7602 4569 7609 4580
rect 7661 4610 7668 4621
rect 8002 4621 8068 4622
rect 8002 4610 8009 4621
rect 7661 4580 8009 4610
rect 7661 4569 7668 4580
rect 7602 4568 7668 4569
rect 8002 4569 8009 4580
rect 8061 4610 8068 4621
rect 8402 4621 8468 4622
rect 8402 4610 8409 4621
rect 8061 4580 8409 4610
rect 8061 4569 8068 4580
rect 8002 4568 8068 4569
rect 8402 4569 8409 4580
rect 8461 4610 8468 4621
rect 8802 4621 8868 4622
rect 8802 4610 8809 4621
rect 8461 4580 8809 4610
rect 8461 4569 8468 4580
rect 8402 4568 8468 4569
rect 8802 4569 8809 4580
rect 8861 4610 8868 4621
rect 9202 4621 9268 4622
rect 9202 4610 9209 4621
rect 8861 4580 9209 4610
rect 8861 4569 8868 4580
rect 8802 4568 8868 4569
rect 9202 4569 9209 4580
rect 9261 4610 9268 4621
rect 9602 4621 9668 4622
rect 9602 4610 9609 4621
rect 9261 4580 9609 4610
rect 9261 4569 9268 4580
rect 9202 4568 9268 4569
rect 9602 4569 9609 4580
rect 9661 4610 9668 4621
rect 10002 4621 10068 4622
rect 10002 4610 10009 4621
rect 9661 4580 10009 4610
rect 9661 4569 9668 4580
rect 9602 4568 9668 4569
rect 10002 4569 10009 4580
rect 10061 4610 10068 4621
rect 10402 4621 10468 4622
rect 10402 4610 10409 4621
rect 10061 4580 10409 4610
rect 10061 4569 10068 4580
rect 10002 4568 10068 4569
rect 10402 4569 10409 4580
rect 10461 4610 10468 4621
rect 10802 4621 10868 4622
rect 10802 4610 10809 4621
rect 10461 4580 10809 4610
rect 10461 4569 10468 4580
rect 10402 4568 10468 4569
rect 10802 4569 10809 4580
rect 10861 4610 10868 4621
rect 11202 4621 11268 4622
rect 11202 4610 11209 4621
rect 10861 4580 11209 4610
rect 10861 4569 10868 4580
rect 10802 4568 10868 4569
rect 11202 4569 11209 4580
rect 11261 4610 11268 4621
rect 11602 4621 11668 4622
rect 11602 4610 11609 4621
rect 11261 4580 11609 4610
rect 11261 4569 11268 4580
rect 11202 4568 11268 4569
rect 11602 4569 11609 4580
rect 11661 4610 11668 4621
rect 12002 4621 12068 4622
rect 12002 4610 12009 4621
rect 11661 4580 12009 4610
rect 11661 4569 11668 4580
rect 11602 4568 11668 4569
rect 12002 4569 12009 4580
rect 12061 4610 12068 4621
rect 12402 4621 12468 4622
rect 12402 4610 12409 4621
rect 12061 4580 12409 4610
rect 12061 4569 12068 4580
rect 12002 4568 12068 4569
rect 12402 4569 12409 4580
rect 12461 4610 12468 4621
rect 12802 4621 12868 4622
rect 12802 4610 12809 4621
rect 12461 4580 12809 4610
rect 12461 4569 12468 4580
rect 12402 4568 12468 4569
rect 12802 4569 12809 4580
rect 12861 4610 12868 4621
rect 12900 4621 12966 4622
rect 12900 4610 12907 4621
rect 12861 4580 12907 4610
rect 12861 4569 12868 4580
rect 12802 4568 12868 4569
rect 12900 4569 12907 4580
rect 12959 4569 12966 4621
rect 12900 4568 12966 4569
rect 202 4551 268 4552
rect 202 4540 209 4551
rect 0 4510 209 4540
rect 202 4499 209 4510
rect 261 4540 268 4551
rect 602 4551 668 4552
rect 602 4540 609 4551
rect 261 4510 609 4540
rect 261 4499 268 4510
rect 202 4498 268 4499
rect 602 4499 609 4510
rect 661 4540 668 4551
rect 1002 4551 1068 4552
rect 1002 4540 1009 4551
rect 661 4510 1009 4540
rect 661 4499 668 4510
rect 602 4498 668 4499
rect 1002 4499 1009 4510
rect 1061 4540 1068 4551
rect 1402 4551 1468 4552
rect 1402 4540 1409 4551
rect 1061 4510 1409 4540
rect 1061 4499 1068 4510
rect 1002 4498 1068 4499
rect 1402 4499 1409 4510
rect 1461 4540 1468 4551
rect 1802 4551 1868 4552
rect 1802 4540 1809 4551
rect 1461 4510 1809 4540
rect 1461 4499 1468 4510
rect 1402 4498 1468 4499
rect 1802 4499 1809 4510
rect 1861 4540 1868 4551
rect 2202 4551 2268 4552
rect 2202 4540 2209 4551
rect 1861 4510 2209 4540
rect 1861 4499 1868 4510
rect 1802 4498 1868 4499
rect 2202 4499 2209 4510
rect 2261 4540 2268 4551
rect 2602 4551 2668 4552
rect 2602 4540 2609 4551
rect 2261 4510 2609 4540
rect 2261 4499 2268 4510
rect 2202 4498 2268 4499
rect 2602 4499 2609 4510
rect 2661 4540 2668 4551
rect 3002 4551 3068 4552
rect 3002 4540 3009 4551
rect 2661 4510 3009 4540
rect 2661 4499 2668 4510
rect 2602 4498 2668 4499
rect 3002 4499 3009 4510
rect 3061 4540 3068 4551
rect 3402 4551 3468 4552
rect 3402 4540 3409 4551
rect 3061 4510 3409 4540
rect 3061 4499 3068 4510
rect 3002 4498 3068 4499
rect 3402 4499 3409 4510
rect 3461 4540 3468 4551
rect 3802 4551 3868 4552
rect 3802 4540 3809 4551
rect 3461 4510 3809 4540
rect 3461 4499 3468 4510
rect 3402 4498 3468 4499
rect 3802 4499 3809 4510
rect 3861 4540 3868 4551
rect 4202 4551 4268 4552
rect 4202 4540 4209 4551
rect 3861 4510 4209 4540
rect 3861 4499 3868 4510
rect 3802 4498 3868 4499
rect 4202 4499 4209 4510
rect 4261 4540 4268 4551
rect 4602 4551 4668 4552
rect 4602 4540 4609 4551
rect 4261 4510 4609 4540
rect 4261 4499 4268 4510
rect 4202 4498 4268 4499
rect 4602 4499 4609 4510
rect 4661 4540 4668 4551
rect 5002 4551 5068 4552
rect 5002 4540 5009 4551
rect 4661 4510 5009 4540
rect 4661 4499 4668 4510
rect 4602 4498 4668 4499
rect 5002 4499 5009 4510
rect 5061 4540 5068 4551
rect 5402 4551 5468 4552
rect 5402 4540 5409 4551
rect 5061 4510 5409 4540
rect 5061 4499 5068 4510
rect 5002 4498 5068 4499
rect 5402 4499 5409 4510
rect 5461 4540 5468 4551
rect 5802 4551 5868 4552
rect 5802 4540 5809 4551
rect 5461 4510 5809 4540
rect 5461 4499 5468 4510
rect 5402 4498 5468 4499
rect 5802 4499 5809 4510
rect 5861 4540 5868 4551
rect 6202 4551 6268 4552
rect 6202 4540 6209 4551
rect 5861 4510 6209 4540
rect 5861 4499 5868 4510
rect 5802 4498 5868 4499
rect 6202 4499 6209 4510
rect 6261 4540 6268 4551
rect 6602 4551 6668 4552
rect 6602 4540 6609 4551
rect 6261 4510 6609 4540
rect 6261 4499 6268 4510
rect 6202 4498 6268 4499
rect 6602 4499 6609 4510
rect 6661 4540 6668 4551
rect 7002 4551 7068 4552
rect 7002 4540 7009 4551
rect 6661 4510 7009 4540
rect 6661 4499 6668 4510
rect 6602 4498 6668 4499
rect 7002 4499 7009 4510
rect 7061 4540 7068 4551
rect 7402 4551 7468 4552
rect 7402 4540 7409 4551
rect 7061 4510 7409 4540
rect 7061 4499 7068 4510
rect 7002 4498 7068 4499
rect 7402 4499 7409 4510
rect 7461 4540 7468 4551
rect 7802 4551 7868 4552
rect 7802 4540 7809 4551
rect 7461 4510 7809 4540
rect 7461 4499 7468 4510
rect 7402 4498 7468 4499
rect 7802 4499 7809 4510
rect 7861 4540 7868 4551
rect 8202 4551 8268 4552
rect 8202 4540 8209 4551
rect 7861 4510 8209 4540
rect 7861 4499 7868 4510
rect 7802 4498 7868 4499
rect 8202 4499 8209 4510
rect 8261 4540 8268 4551
rect 8602 4551 8668 4552
rect 8602 4540 8609 4551
rect 8261 4510 8609 4540
rect 8261 4499 8268 4510
rect 8202 4498 8268 4499
rect 8602 4499 8609 4510
rect 8661 4540 8668 4551
rect 9002 4551 9068 4552
rect 9002 4540 9009 4551
rect 8661 4510 9009 4540
rect 8661 4499 8668 4510
rect 8602 4498 8668 4499
rect 9002 4499 9009 4510
rect 9061 4540 9068 4551
rect 9402 4551 9468 4552
rect 9402 4540 9409 4551
rect 9061 4510 9409 4540
rect 9061 4499 9068 4510
rect 9002 4498 9068 4499
rect 9402 4499 9409 4510
rect 9461 4540 9468 4551
rect 9802 4551 9868 4552
rect 9802 4540 9809 4551
rect 9461 4510 9809 4540
rect 9461 4499 9468 4510
rect 9402 4498 9468 4499
rect 9802 4499 9809 4510
rect 9861 4540 9868 4551
rect 10202 4551 10268 4552
rect 10202 4540 10209 4551
rect 9861 4510 10209 4540
rect 9861 4499 9868 4510
rect 9802 4498 9868 4499
rect 10202 4499 10209 4510
rect 10261 4540 10268 4551
rect 10602 4551 10668 4552
rect 10602 4540 10609 4551
rect 10261 4510 10609 4540
rect 10261 4499 10268 4510
rect 10202 4498 10268 4499
rect 10602 4499 10609 4510
rect 10661 4540 10668 4551
rect 11002 4551 11068 4552
rect 11002 4540 11009 4551
rect 10661 4510 11009 4540
rect 10661 4499 10668 4510
rect 10602 4498 10668 4499
rect 11002 4499 11009 4510
rect 11061 4540 11068 4551
rect 11402 4551 11468 4552
rect 11402 4540 11409 4551
rect 11061 4510 11409 4540
rect 11061 4499 11068 4510
rect 11002 4498 11068 4499
rect 11402 4499 11409 4510
rect 11461 4540 11468 4551
rect 11802 4551 11868 4552
rect 11802 4540 11809 4551
rect 11461 4510 11809 4540
rect 11461 4499 11468 4510
rect 11402 4498 11468 4499
rect 11802 4499 11809 4510
rect 11861 4540 11868 4551
rect 12202 4551 12268 4552
rect 12202 4540 12209 4551
rect 11861 4510 12209 4540
rect 11861 4499 11868 4510
rect 11802 4498 11868 4499
rect 12202 4499 12209 4510
rect 12261 4540 12268 4551
rect 12602 4551 12668 4552
rect 12602 4540 12609 4551
rect 12261 4510 12609 4540
rect 12261 4499 12268 4510
rect 12202 4498 12268 4499
rect 12602 4499 12609 4510
rect 12661 4540 12668 4551
rect 13104 4551 13170 4552
rect 13104 4540 13111 4551
rect 12661 4510 13111 4540
rect 12661 4499 12668 4510
rect 12602 4498 12668 4499
rect 13104 4499 13111 4510
rect 13163 4499 13170 4551
rect 13104 4498 13170 4499
rect 2 4481 68 4482
rect 2 4470 9 4481
rect 0 4440 9 4470
rect 2 4429 9 4440
rect 61 4470 68 4481
rect 402 4481 468 4482
rect 402 4470 409 4481
rect 61 4440 409 4470
rect 61 4429 68 4440
rect 2 4428 68 4429
rect 402 4429 409 4440
rect 461 4470 468 4481
rect 802 4481 868 4482
rect 802 4470 809 4481
rect 461 4440 809 4470
rect 461 4429 468 4440
rect 402 4428 468 4429
rect 802 4429 809 4440
rect 861 4470 868 4481
rect 1202 4481 1268 4482
rect 1202 4470 1209 4481
rect 861 4440 1209 4470
rect 861 4429 868 4440
rect 802 4428 868 4429
rect 1202 4429 1209 4440
rect 1261 4470 1268 4481
rect 1602 4481 1668 4482
rect 1602 4470 1609 4481
rect 1261 4440 1609 4470
rect 1261 4429 1268 4440
rect 1202 4428 1268 4429
rect 1602 4429 1609 4440
rect 1661 4470 1668 4481
rect 2002 4481 2068 4482
rect 2002 4470 2009 4481
rect 1661 4440 2009 4470
rect 1661 4429 1668 4440
rect 1602 4428 1668 4429
rect 2002 4429 2009 4440
rect 2061 4470 2068 4481
rect 2402 4481 2468 4482
rect 2402 4470 2409 4481
rect 2061 4440 2409 4470
rect 2061 4429 2068 4440
rect 2002 4428 2068 4429
rect 2402 4429 2409 4440
rect 2461 4470 2468 4481
rect 2802 4481 2868 4482
rect 2802 4470 2809 4481
rect 2461 4440 2809 4470
rect 2461 4429 2468 4440
rect 2402 4428 2468 4429
rect 2802 4429 2809 4440
rect 2861 4470 2868 4481
rect 3202 4481 3268 4482
rect 3202 4470 3209 4481
rect 2861 4440 3209 4470
rect 2861 4429 2868 4440
rect 2802 4428 2868 4429
rect 3202 4429 3209 4440
rect 3261 4470 3268 4481
rect 3602 4481 3668 4482
rect 3602 4470 3609 4481
rect 3261 4440 3609 4470
rect 3261 4429 3268 4440
rect 3202 4428 3268 4429
rect 3602 4429 3609 4440
rect 3661 4470 3668 4481
rect 4002 4481 4068 4482
rect 4002 4470 4009 4481
rect 3661 4440 4009 4470
rect 3661 4429 3668 4440
rect 3602 4428 3668 4429
rect 4002 4429 4009 4440
rect 4061 4470 4068 4481
rect 4402 4481 4468 4482
rect 4402 4470 4409 4481
rect 4061 4440 4409 4470
rect 4061 4429 4068 4440
rect 4002 4428 4068 4429
rect 4402 4429 4409 4440
rect 4461 4470 4468 4481
rect 4802 4481 4868 4482
rect 4802 4470 4809 4481
rect 4461 4440 4809 4470
rect 4461 4429 4468 4440
rect 4402 4428 4468 4429
rect 4802 4429 4809 4440
rect 4861 4470 4868 4481
rect 5202 4481 5268 4482
rect 5202 4470 5209 4481
rect 4861 4440 5209 4470
rect 4861 4429 4868 4440
rect 4802 4428 4868 4429
rect 5202 4429 5209 4440
rect 5261 4470 5268 4481
rect 5602 4481 5668 4482
rect 5602 4470 5609 4481
rect 5261 4440 5609 4470
rect 5261 4429 5268 4440
rect 5202 4428 5268 4429
rect 5602 4429 5609 4440
rect 5661 4470 5668 4481
rect 6002 4481 6068 4482
rect 6002 4470 6009 4481
rect 5661 4440 6009 4470
rect 5661 4429 5668 4440
rect 5602 4428 5668 4429
rect 6002 4429 6009 4440
rect 6061 4470 6068 4481
rect 6402 4481 6468 4482
rect 6402 4470 6409 4481
rect 6061 4440 6409 4470
rect 6061 4429 6068 4440
rect 6002 4428 6068 4429
rect 6402 4429 6409 4440
rect 6461 4470 6468 4481
rect 6802 4481 6868 4482
rect 6802 4470 6809 4481
rect 6461 4440 6809 4470
rect 6461 4429 6468 4440
rect 6402 4428 6468 4429
rect 6802 4429 6809 4440
rect 6861 4470 6868 4481
rect 7202 4481 7268 4482
rect 7202 4470 7209 4481
rect 6861 4440 7209 4470
rect 6861 4429 6868 4440
rect 6802 4428 6868 4429
rect 7202 4429 7209 4440
rect 7261 4470 7268 4481
rect 7602 4481 7668 4482
rect 7602 4470 7609 4481
rect 7261 4440 7609 4470
rect 7261 4429 7268 4440
rect 7202 4428 7268 4429
rect 7602 4429 7609 4440
rect 7661 4470 7668 4481
rect 8002 4481 8068 4482
rect 8002 4470 8009 4481
rect 7661 4440 8009 4470
rect 7661 4429 7668 4440
rect 7602 4428 7668 4429
rect 8002 4429 8009 4440
rect 8061 4470 8068 4481
rect 8402 4481 8468 4482
rect 8402 4470 8409 4481
rect 8061 4440 8409 4470
rect 8061 4429 8068 4440
rect 8002 4428 8068 4429
rect 8402 4429 8409 4440
rect 8461 4470 8468 4481
rect 8802 4481 8868 4482
rect 8802 4470 8809 4481
rect 8461 4440 8809 4470
rect 8461 4429 8468 4440
rect 8402 4428 8468 4429
rect 8802 4429 8809 4440
rect 8861 4470 8868 4481
rect 9202 4481 9268 4482
rect 9202 4470 9209 4481
rect 8861 4440 9209 4470
rect 8861 4429 8868 4440
rect 8802 4428 8868 4429
rect 9202 4429 9209 4440
rect 9261 4470 9268 4481
rect 9602 4481 9668 4482
rect 9602 4470 9609 4481
rect 9261 4440 9609 4470
rect 9261 4429 9268 4440
rect 9202 4428 9268 4429
rect 9602 4429 9609 4440
rect 9661 4470 9668 4481
rect 10002 4481 10068 4482
rect 10002 4470 10009 4481
rect 9661 4440 10009 4470
rect 9661 4429 9668 4440
rect 9602 4428 9668 4429
rect 10002 4429 10009 4440
rect 10061 4470 10068 4481
rect 10402 4481 10468 4482
rect 10402 4470 10409 4481
rect 10061 4440 10409 4470
rect 10061 4429 10068 4440
rect 10002 4428 10068 4429
rect 10402 4429 10409 4440
rect 10461 4470 10468 4481
rect 10802 4481 10868 4482
rect 10802 4470 10809 4481
rect 10461 4440 10809 4470
rect 10461 4429 10468 4440
rect 10402 4428 10468 4429
rect 10802 4429 10809 4440
rect 10861 4470 10868 4481
rect 11202 4481 11268 4482
rect 11202 4470 11209 4481
rect 10861 4440 11209 4470
rect 10861 4429 10868 4440
rect 10802 4428 10868 4429
rect 11202 4429 11209 4440
rect 11261 4470 11268 4481
rect 11602 4481 11668 4482
rect 11602 4470 11609 4481
rect 11261 4440 11609 4470
rect 11261 4429 11268 4440
rect 11202 4428 11268 4429
rect 11602 4429 11609 4440
rect 11661 4470 11668 4481
rect 12002 4481 12068 4482
rect 12002 4470 12009 4481
rect 11661 4440 12009 4470
rect 11661 4429 11668 4440
rect 11602 4428 11668 4429
rect 12002 4429 12009 4440
rect 12061 4470 12068 4481
rect 12402 4481 12468 4482
rect 12402 4470 12409 4481
rect 12061 4440 12409 4470
rect 12061 4429 12068 4440
rect 12002 4428 12068 4429
rect 12402 4429 12409 4440
rect 12461 4470 12468 4481
rect 12802 4481 12868 4482
rect 12802 4470 12809 4481
rect 12461 4440 12809 4470
rect 12461 4429 12468 4440
rect 12402 4428 12468 4429
rect 12802 4429 12809 4440
rect 12861 4470 12868 4481
rect 12900 4481 12966 4482
rect 12900 4470 12907 4481
rect 12861 4440 12907 4470
rect 12861 4429 12868 4440
rect 12802 4428 12868 4429
rect 12900 4429 12907 4440
rect 12959 4429 12966 4481
rect 12900 4428 12966 4429
rect 202 4411 268 4412
rect 202 4400 209 4411
rect 0 4370 209 4400
rect 202 4359 209 4370
rect 261 4400 268 4411
rect 602 4411 668 4412
rect 602 4400 609 4411
rect 261 4370 609 4400
rect 261 4359 268 4370
rect 202 4358 268 4359
rect 602 4359 609 4370
rect 661 4400 668 4411
rect 1002 4411 1068 4412
rect 1002 4400 1009 4411
rect 661 4370 1009 4400
rect 661 4359 668 4370
rect 602 4358 668 4359
rect 1002 4359 1009 4370
rect 1061 4400 1068 4411
rect 1402 4411 1468 4412
rect 1402 4400 1409 4411
rect 1061 4370 1409 4400
rect 1061 4359 1068 4370
rect 1002 4358 1068 4359
rect 1402 4359 1409 4370
rect 1461 4400 1468 4411
rect 1802 4411 1868 4412
rect 1802 4400 1809 4411
rect 1461 4370 1809 4400
rect 1461 4359 1468 4370
rect 1402 4358 1468 4359
rect 1802 4359 1809 4370
rect 1861 4400 1868 4411
rect 2202 4411 2268 4412
rect 2202 4400 2209 4411
rect 1861 4370 2209 4400
rect 1861 4359 1868 4370
rect 1802 4358 1868 4359
rect 2202 4359 2209 4370
rect 2261 4400 2268 4411
rect 2602 4411 2668 4412
rect 2602 4400 2609 4411
rect 2261 4370 2609 4400
rect 2261 4359 2268 4370
rect 2202 4358 2268 4359
rect 2602 4359 2609 4370
rect 2661 4400 2668 4411
rect 3002 4411 3068 4412
rect 3002 4400 3009 4411
rect 2661 4370 3009 4400
rect 2661 4359 2668 4370
rect 2602 4358 2668 4359
rect 3002 4359 3009 4370
rect 3061 4400 3068 4411
rect 3402 4411 3468 4412
rect 3402 4400 3409 4411
rect 3061 4370 3409 4400
rect 3061 4359 3068 4370
rect 3002 4358 3068 4359
rect 3402 4359 3409 4370
rect 3461 4400 3468 4411
rect 3802 4411 3868 4412
rect 3802 4400 3809 4411
rect 3461 4370 3809 4400
rect 3461 4359 3468 4370
rect 3402 4358 3468 4359
rect 3802 4359 3809 4370
rect 3861 4400 3868 4411
rect 4202 4411 4268 4412
rect 4202 4400 4209 4411
rect 3861 4370 4209 4400
rect 3861 4359 3868 4370
rect 3802 4358 3868 4359
rect 4202 4359 4209 4370
rect 4261 4400 4268 4411
rect 4602 4411 4668 4412
rect 4602 4400 4609 4411
rect 4261 4370 4609 4400
rect 4261 4359 4268 4370
rect 4202 4358 4268 4359
rect 4602 4359 4609 4370
rect 4661 4400 4668 4411
rect 5002 4411 5068 4412
rect 5002 4400 5009 4411
rect 4661 4370 5009 4400
rect 4661 4359 4668 4370
rect 4602 4358 4668 4359
rect 5002 4359 5009 4370
rect 5061 4400 5068 4411
rect 5402 4411 5468 4412
rect 5402 4400 5409 4411
rect 5061 4370 5409 4400
rect 5061 4359 5068 4370
rect 5002 4358 5068 4359
rect 5402 4359 5409 4370
rect 5461 4400 5468 4411
rect 5802 4411 5868 4412
rect 5802 4400 5809 4411
rect 5461 4370 5809 4400
rect 5461 4359 5468 4370
rect 5402 4358 5468 4359
rect 5802 4359 5809 4370
rect 5861 4400 5868 4411
rect 6202 4411 6268 4412
rect 6202 4400 6209 4411
rect 5861 4370 6209 4400
rect 5861 4359 5868 4370
rect 5802 4358 5868 4359
rect 6202 4359 6209 4370
rect 6261 4400 6268 4411
rect 6602 4411 6668 4412
rect 6602 4400 6609 4411
rect 6261 4370 6609 4400
rect 6261 4359 6268 4370
rect 6202 4358 6268 4359
rect 6602 4359 6609 4370
rect 6661 4400 6668 4411
rect 7002 4411 7068 4412
rect 7002 4400 7009 4411
rect 6661 4370 7009 4400
rect 6661 4359 6668 4370
rect 6602 4358 6668 4359
rect 7002 4359 7009 4370
rect 7061 4400 7068 4411
rect 7402 4411 7468 4412
rect 7402 4400 7409 4411
rect 7061 4370 7409 4400
rect 7061 4359 7068 4370
rect 7002 4358 7068 4359
rect 7402 4359 7409 4370
rect 7461 4400 7468 4411
rect 7802 4411 7868 4412
rect 7802 4400 7809 4411
rect 7461 4370 7809 4400
rect 7461 4359 7468 4370
rect 7402 4358 7468 4359
rect 7802 4359 7809 4370
rect 7861 4400 7868 4411
rect 8202 4411 8268 4412
rect 8202 4400 8209 4411
rect 7861 4370 8209 4400
rect 7861 4359 7868 4370
rect 7802 4358 7868 4359
rect 8202 4359 8209 4370
rect 8261 4400 8268 4411
rect 8602 4411 8668 4412
rect 8602 4400 8609 4411
rect 8261 4370 8609 4400
rect 8261 4359 8268 4370
rect 8202 4358 8268 4359
rect 8602 4359 8609 4370
rect 8661 4400 8668 4411
rect 9002 4411 9068 4412
rect 9002 4400 9009 4411
rect 8661 4370 9009 4400
rect 8661 4359 8668 4370
rect 8602 4358 8668 4359
rect 9002 4359 9009 4370
rect 9061 4400 9068 4411
rect 9402 4411 9468 4412
rect 9402 4400 9409 4411
rect 9061 4370 9409 4400
rect 9061 4359 9068 4370
rect 9002 4358 9068 4359
rect 9402 4359 9409 4370
rect 9461 4400 9468 4411
rect 9802 4411 9868 4412
rect 9802 4400 9809 4411
rect 9461 4370 9809 4400
rect 9461 4359 9468 4370
rect 9402 4358 9468 4359
rect 9802 4359 9809 4370
rect 9861 4400 9868 4411
rect 10202 4411 10268 4412
rect 10202 4400 10209 4411
rect 9861 4370 10209 4400
rect 9861 4359 9868 4370
rect 9802 4358 9868 4359
rect 10202 4359 10209 4370
rect 10261 4400 10268 4411
rect 10602 4411 10668 4412
rect 10602 4400 10609 4411
rect 10261 4370 10609 4400
rect 10261 4359 10268 4370
rect 10202 4358 10268 4359
rect 10602 4359 10609 4370
rect 10661 4400 10668 4411
rect 11002 4411 11068 4412
rect 11002 4400 11009 4411
rect 10661 4370 11009 4400
rect 10661 4359 10668 4370
rect 10602 4358 10668 4359
rect 11002 4359 11009 4370
rect 11061 4400 11068 4411
rect 11402 4411 11468 4412
rect 11402 4400 11409 4411
rect 11061 4370 11409 4400
rect 11061 4359 11068 4370
rect 11002 4358 11068 4359
rect 11402 4359 11409 4370
rect 11461 4400 11468 4411
rect 11802 4411 11868 4412
rect 11802 4400 11809 4411
rect 11461 4370 11809 4400
rect 11461 4359 11468 4370
rect 11402 4358 11468 4359
rect 11802 4359 11809 4370
rect 11861 4400 11868 4411
rect 12202 4411 12268 4412
rect 12202 4400 12209 4411
rect 11861 4370 12209 4400
rect 11861 4359 11868 4370
rect 11802 4358 11868 4359
rect 12202 4359 12209 4370
rect 12261 4400 12268 4411
rect 12602 4411 12668 4412
rect 12602 4400 12609 4411
rect 12261 4370 12609 4400
rect 12261 4359 12268 4370
rect 12202 4358 12268 4359
rect 12602 4359 12609 4370
rect 12661 4400 12668 4411
rect 13104 4411 13170 4412
rect 13104 4400 13111 4411
rect 12661 4370 13111 4400
rect 12661 4359 12668 4370
rect 12602 4358 12668 4359
rect 13104 4359 13111 4370
rect 13163 4359 13170 4411
rect 13104 4358 13170 4359
rect 2 4341 68 4342
rect 2 4330 9 4341
rect 0 4300 9 4330
rect 2 4289 9 4300
rect 61 4330 68 4341
rect 402 4341 468 4342
rect 402 4330 409 4341
rect 61 4300 409 4330
rect 61 4289 68 4300
rect 2 4288 68 4289
rect 402 4289 409 4300
rect 461 4330 468 4341
rect 802 4341 868 4342
rect 802 4330 809 4341
rect 461 4300 809 4330
rect 461 4289 468 4300
rect 402 4288 468 4289
rect 802 4289 809 4300
rect 861 4330 868 4341
rect 1202 4341 1268 4342
rect 1202 4330 1209 4341
rect 861 4300 1209 4330
rect 861 4289 868 4300
rect 802 4288 868 4289
rect 1202 4289 1209 4300
rect 1261 4330 1268 4341
rect 1602 4341 1668 4342
rect 1602 4330 1609 4341
rect 1261 4300 1609 4330
rect 1261 4289 1268 4300
rect 1202 4288 1268 4289
rect 1602 4289 1609 4300
rect 1661 4330 1668 4341
rect 2002 4341 2068 4342
rect 2002 4330 2009 4341
rect 1661 4300 2009 4330
rect 1661 4289 1668 4300
rect 1602 4288 1668 4289
rect 2002 4289 2009 4300
rect 2061 4330 2068 4341
rect 2402 4341 2468 4342
rect 2402 4330 2409 4341
rect 2061 4300 2409 4330
rect 2061 4289 2068 4300
rect 2002 4288 2068 4289
rect 2402 4289 2409 4300
rect 2461 4330 2468 4341
rect 2802 4341 2868 4342
rect 2802 4330 2809 4341
rect 2461 4300 2809 4330
rect 2461 4289 2468 4300
rect 2402 4288 2468 4289
rect 2802 4289 2809 4300
rect 2861 4330 2868 4341
rect 3202 4341 3268 4342
rect 3202 4330 3209 4341
rect 2861 4300 3209 4330
rect 2861 4289 2868 4300
rect 2802 4288 2868 4289
rect 3202 4289 3209 4300
rect 3261 4330 3268 4341
rect 3602 4341 3668 4342
rect 3602 4330 3609 4341
rect 3261 4300 3609 4330
rect 3261 4289 3268 4300
rect 3202 4288 3268 4289
rect 3602 4289 3609 4300
rect 3661 4330 3668 4341
rect 4002 4341 4068 4342
rect 4002 4330 4009 4341
rect 3661 4300 4009 4330
rect 3661 4289 3668 4300
rect 3602 4288 3668 4289
rect 4002 4289 4009 4300
rect 4061 4330 4068 4341
rect 4402 4341 4468 4342
rect 4402 4330 4409 4341
rect 4061 4300 4409 4330
rect 4061 4289 4068 4300
rect 4002 4288 4068 4289
rect 4402 4289 4409 4300
rect 4461 4330 4468 4341
rect 4802 4341 4868 4342
rect 4802 4330 4809 4341
rect 4461 4300 4809 4330
rect 4461 4289 4468 4300
rect 4402 4288 4468 4289
rect 4802 4289 4809 4300
rect 4861 4330 4868 4341
rect 5202 4341 5268 4342
rect 5202 4330 5209 4341
rect 4861 4300 5209 4330
rect 4861 4289 4868 4300
rect 4802 4288 4868 4289
rect 5202 4289 5209 4300
rect 5261 4330 5268 4341
rect 5602 4341 5668 4342
rect 5602 4330 5609 4341
rect 5261 4300 5609 4330
rect 5261 4289 5268 4300
rect 5202 4288 5268 4289
rect 5602 4289 5609 4300
rect 5661 4330 5668 4341
rect 6002 4341 6068 4342
rect 6002 4330 6009 4341
rect 5661 4300 6009 4330
rect 5661 4289 5668 4300
rect 5602 4288 5668 4289
rect 6002 4289 6009 4300
rect 6061 4330 6068 4341
rect 6402 4341 6468 4342
rect 6402 4330 6409 4341
rect 6061 4300 6409 4330
rect 6061 4289 6068 4300
rect 6002 4288 6068 4289
rect 6402 4289 6409 4300
rect 6461 4330 6468 4341
rect 6802 4341 6868 4342
rect 6802 4330 6809 4341
rect 6461 4300 6809 4330
rect 6461 4289 6468 4300
rect 6402 4288 6468 4289
rect 6802 4289 6809 4300
rect 6861 4330 6868 4341
rect 7202 4341 7268 4342
rect 7202 4330 7209 4341
rect 6861 4300 7209 4330
rect 6861 4289 6868 4300
rect 6802 4288 6868 4289
rect 7202 4289 7209 4300
rect 7261 4330 7268 4341
rect 7602 4341 7668 4342
rect 7602 4330 7609 4341
rect 7261 4300 7609 4330
rect 7261 4289 7268 4300
rect 7202 4288 7268 4289
rect 7602 4289 7609 4300
rect 7661 4330 7668 4341
rect 8002 4341 8068 4342
rect 8002 4330 8009 4341
rect 7661 4300 8009 4330
rect 7661 4289 7668 4300
rect 7602 4288 7668 4289
rect 8002 4289 8009 4300
rect 8061 4330 8068 4341
rect 8402 4341 8468 4342
rect 8402 4330 8409 4341
rect 8061 4300 8409 4330
rect 8061 4289 8068 4300
rect 8002 4288 8068 4289
rect 8402 4289 8409 4300
rect 8461 4330 8468 4341
rect 8802 4341 8868 4342
rect 8802 4330 8809 4341
rect 8461 4300 8809 4330
rect 8461 4289 8468 4300
rect 8402 4288 8468 4289
rect 8802 4289 8809 4300
rect 8861 4330 8868 4341
rect 9202 4341 9268 4342
rect 9202 4330 9209 4341
rect 8861 4300 9209 4330
rect 8861 4289 8868 4300
rect 8802 4288 8868 4289
rect 9202 4289 9209 4300
rect 9261 4330 9268 4341
rect 9602 4341 9668 4342
rect 9602 4330 9609 4341
rect 9261 4300 9609 4330
rect 9261 4289 9268 4300
rect 9202 4288 9268 4289
rect 9602 4289 9609 4300
rect 9661 4330 9668 4341
rect 10002 4341 10068 4342
rect 10002 4330 10009 4341
rect 9661 4300 10009 4330
rect 9661 4289 9668 4300
rect 9602 4288 9668 4289
rect 10002 4289 10009 4300
rect 10061 4330 10068 4341
rect 10402 4341 10468 4342
rect 10402 4330 10409 4341
rect 10061 4300 10409 4330
rect 10061 4289 10068 4300
rect 10002 4288 10068 4289
rect 10402 4289 10409 4300
rect 10461 4330 10468 4341
rect 10802 4341 10868 4342
rect 10802 4330 10809 4341
rect 10461 4300 10809 4330
rect 10461 4289 10468 4300
rect 10402 4288 10468 4289
rect 10802 4289 10809 4300
rect 10861 4330 10868 4341
rect 11202 4341 11268 4342
rect 11202 4330 11209 4341
rect 10861 4300 11209 4330
rect 10861 4289 10868 4300
rect 10802 4288 10868 4289
rect 11202 4289 11209 4300
rect 11261 4330 11268 4341
rect 11602 4341 11668 4342
rect 11602 4330 11609 4341
rect 11261 4300 11609 4330
rect 11261 4289 11268 4300
rect 11202 4288 11268 4289
rect 11602 4289 11609 4300
rect 11661 4330 11668 4341
rect 12002 4341 12068 4342
rect 12002 4330 12009 4341
rect 11661 4300 12009 4330
rect 11661 4289 11668 4300
rect 11602 4288 11668 4289
rect 12002 4289 12009 4300
rect 12061 4330 12068 4341
rect 12402 4341 12468 4342
rect 12402 4330 12409 4341
rect 12061 4300 12409 4330
rect 12061 4289 12068 4300
rect 12002 4288 12068 4289
rect 12402 4289 12409 4300
rect 12461 4330 12468 4341
rect 12802 4341 12868 4342
rect 12802 4330 12809 4341
rect 12461 4300 12809 4330
rect 12461 4289 12468 4300
rect 12402 4288 12468 4289
rect 12802 4289 12809 4300
rect 12861 4330 12868 4341
rect 12900 4341 12966 4342
rect 12900 4330 12907 4341
rect 12861 4300 12907 4330
rect 12861 4289 12868 4300
rect 12802 4288 12868 4289
rect 12900 4289 12907 4300
rect 12959 4289 12966 4341
rect 12900 4288 12966 4289
rect 202 4271 268 4272
rect 202 4260 209 4271
rect 0 4230 209 4260
rect 202 4219 209 4230
rect 261 4260 268 4271
rect 602 4271 668 4272
rect 602 4260 609 4271
rect 261 4230 609 4260
rect 261 4219 268 4230
rect 202 4218 268 4219
rect 602 4219 609 4230
rect 661 4260 668 4271
rect 1002 4271 1068 4272
rect 1002 4260 1009 4271
rect 661 4230 1009 4260
rect 661 4219 668 4230
rect 602 4218 668 4219
rect 1002 4219 1009 4230
rect 1061 4260 1068 4271
rect 1402 4271 1468 4272
rect 1402 4260 1409 4271
rect 1061 4230 1409 4260
rect 1061 4219 1068 4230
rect 1002 4218 1068 4219
rect 1402 4219 1409 4230
rect 1461 4260 1468 4271
rect 1802 4271 1868 4272
rect 1802 4260 1809 4271
rect 1461 4230 1809 4260
rect 1461 4219 1468 4230
rect 1402 4218 1468 4219
rect 1802 4219 1809 4230
rect 1861 4260 1868 4271
rect 2202 4271 2268 4272
rect 2202 4260 2209 4271
rect 1861 4230 2209 4260
rect 1861 4219 1868 4230
rect 1802 4218 1868 4219
rect 2202 4219 2209 4230
rect 2261 4260 2268 4271
rect 2602 4271 2668 4272
rect 2602 4260 2609 4271
rect 2261 4230 2609 4260
rect 2261 4219 2268 4230
rect 2202 4218 2268 4219
rect 2602 4219 2609 4230
rect 2661 4260 2668 4271
rect 3002 4271 3068 4272
rect 3002 4260 3009 4271
rect 2661 4230 3009 4260
rect 2661 4219 2668 4230
rect 2602 4218 2668 4219
rect 3002 4219 3009 4230
rect 3061 4260 3068 4271
rect 3402 4271 3468 4272
rect 3402 4260 3409 4271
rect 3061 4230 3409 4260
rect 3061 4219 3068 4230
rect 3002 4218 3068 4219
rect 3402 4219 3409 4230
rect 3461 4260 3468 4271
rect 3802 4271 3868 4272
rect 3802 4260 3809 4271
rect 3461 4230 3809 4260
rect 3461 4219 3468 4230
rect 3402 4218 3468 4219
rect 3802 4219 3809 4230
rect 3861 4260 3868 4271
rect 4202 4271 4268 4272
rect 4202 4260 4209 4271
rect 3861 4230 4209 4260
rect 3861 4219 3868 4230
rect 3802 4218 3868 4219
rect 4202 4219 4209 4230
rect 4261 4260 4268 4271
rect 4602 4271 4668 4272
rect 4602 4260 4609 4271
rect 4261 4230 4609 4260
rect 4261 4219 4268 4230
rect 4202 4218 4268 4219
rect 4602 4219 4609 4230
rect 4661 4260 4668 4271
rect 5002 4271 5068 4272
rect 5002 4260 5009 4271
rect 4661 4230 5009 4260
rect 4661 4219 4668 4230
rect 4602 4218 4668 4219
rect 5002 4219 5009 4230
rect 5061 4260 5068 4271
rect 5402 4271 5468 4272
rect 5402 4260 5409 4271
rect 5061 4230 5409 4260
rect 5061 4219 5068 4230
rect 5002 4218 5068 4219
rect 5402 4219 5409 4230
rect 5461 4260 5468 4271
rect 5802 4271 5868 4272
rect 5802 4260 5809 4271
rect 5461 4230 5809 4260
rect 5461 4219 5468 4230
rect 5402 4218 5468 4219
rect 5802 4219 5809 4230
rect 5861 4260 5868 4271
rect 6202 4271 6268 4272
rect 6202 4260 6209 4271
rect 5861 4230 6209 4260
rect 5861 4219 5868 4230
rect 5802 4218 5868 4219
rect 6202 4219 6209 4230
rect 6261 4260 6268 4271
rect 6602 4271 6668 4272
rect 6602 4260 6609 4271
rect 6261 4230 6609 4260
rect 6261 4219 6268 4230
rect 6202 4218 6268 4219
rect 6602 4219 6609 4230
rect 6661 4260 6668 4271
rect 7002 4271 7068 4272
rect 7002 4260 7009 4271
rect 6661 4230 7009 4260
rect 6661 4219 6668 4230
rect 6602 4218 6668 4219
rect 7002 4219 7009 4230
rect 7061 4260 7068 4271
rect 7402 4271 7468 4272
rect 7402 4260 7409 4271
rect 7061 4230 7409 4260
rect 7061 4219 7068 4230
rect 7002 4218 7068 4219
rect 7402 4219 7409 4230
rect 7461 4260 7468 4271
rect 7802 4271 7868 4272
rect 7802 4260 7809 4271
rect 7461 4230 7809 4260
rect 7461 4219 7468 4230
rect 7402 4218 7468 4219
rect 7802 4219 7809 4230
rect 7861 4260 7868 4271
rect 8202 4271 8268 4272
rect 8202 4260 8209 4271
rect 7861 4230 8209 4260
rect 7861 4219 7868 4230
rect 7802 4218 7868 4219
rect 8202 4219 8209 4230
rect 8261 4260 8268 4271
rect 8602 4271 8668 4272
rect 8602 4260 8609 4271
rect 8261 4230 8609 4260
rect 8261 4219 8268 4230
rect 8202 4218 8268 4219
rect 8602 4219 8609 4230
rect 8661 4260 8668 4271
rect 9002 4271 9068 4272
rect 9002 4260 9009 4271
rect 8661 4230 9009 4260
rect 8661 4219 8668 4230
rect 8602 4218 8668 4219
rect 9002 4219 9009 4230
rect 9061 4260 9068 4271
rect 9402 4271 9468 4272
rect 9402 4260 9409 4271
rect 9061 4230 9409 4260
rect 9061 4219 9068 4230
rect 9002 4218 9068 4219
rect 9402 4219 9409 4230
rect 9461 4260 9468 4271
rect 9802 4271 9868 4272
rect 9802 4260 9809 4271
rect 9461 4230 9809 4260
rect 9461 4219 9468 4230
rect 9402 4218 9468 4219
rect 9802 4219 9809 4230
rect 9861 4260 9868 4271
rect 10202 4271 10268 4272
rect 10202 4260 10209 4271
rect 9861 4230 10209 4260
rect 9861 4219 9868 4230
rect 9802 4218 9868 4219
rect 10202 4219 10209 4230
rect 10261 4260 10268 4271
rect 10602 4271 10668 4272
rect 10602 4260 10609 4271
rect 10261 4230 10609 4260
rect 10261 4219 10268 4230
rect 10202 4218 10268 4219
rect 10602 4219 10609 4230
rect 10661 4260 10668 4271
rect 11002 4271 11068 4272
rect 11002 4260 11009 4271
rect 10661 4230 11009 4260
rect 10661 4219 10668 4230
rect 10602 4218 10668 4219
rect 11002 4219 11009 4230
rect 11061 4260 11068 4271
rect 11402 4271 11468 4272
rect 11402 4260 11409 4271
rect 11061 4230 11409 4260
rect 11061 4219 11068 4230
rect 11002 4218 11068 4219
rect 11402 4219 11409 4230
rect 11461 4260 11468 4271
rect 11802 4271 11868 4272
rect 11802 4260 11809 4271
rect 11461 4230 11809 4260
rect 11461 4219 11468 4230
rect 11402 4218 11468 4219
rect 11802 4219 11809 4230
rect 11861 4260 11868 4271
rect 12202 4271 12268 4272
rect 12202 4260 12209 4271
rect 11861 4230 12209 4260
rect 11861 4219 11868 4230
rect 11802 4218 11868 4219
rect 12202 4219 12209 4230
rect 12261 4260 12268 4271
rect 12602 4271 12668 4272
rect 12602 4260 12609 4271
rect 12261 4230 12609 4260
rect 12261 4219 12268 4230
rect 12202 4218 12268 4219
rect 12602 4219 12609 4230
rect 12661 4260 12668 4271
rect 13104 4271 13170 4272
rect 13104 4260 13111 4271
rect 12661 4230 13111 4260
rect 12661 4219 12668 4230
rect 12602 4218 12668 4219
rect 13104 4219 13111 4230
rect 13163 4219 13170 4271
rect 13104 4218 13170 4219
rect 2 4201 68 4202
rect 2 4190 9 4201
rect 0 4160 9 4190
rect 2 4149 9 4160
rect 61 4190 68 4201
rect 402 4201 468 4202
rect 402 4190 409 4201
rect 61 4160 409 4190
rect 61 4149 68 4160
rect 2 4148 68 4149
rect 402 4149 409 4160
rect 461 4190 468 4201
rect 802 4201 868 4202
rect 802 4190 809 4201
rect 461 4160 809 4190
rect 461 4149 468 4160
rect 402 4148 468 4149
rect 802 4149 809 4160
rect 861 4190 868 4201
rect 1202 4201 1268 4202
rect 1202 4190 1209 4201
rect 861 4160 1209 4190
rect 861 4149 868 4160
rect 802 4148 868 4149
rect 1202 4149 1209 4160
rect 1261 4190 1268 4201
rect 1602 4201 1668 4202
rect 1602 4190 1609 4201
rect 1261 4160 1609 4190
rect 1261 4149 1268 4160
rect 1202 4148 1268 4149
rect 1602 4149 1609 4160
rect 1661 4190 1668 4201
rect 2002 4201 2068 4202
rect 2002 4190 2009 4201
rect 1661 4160 2009 4190
rect 1661 4149 1668 4160
rect 1602 4148 1668 4149
rect 2002 4149 2009 4160
rect 2061 4190 2068 4201
rect 2402 4201 2468 4202
rect 2402 4190 2409 4201
rect 2061 4160 2409 4190
rect 2061 4149 2068 4160
rect 2002 4148 2068 4149
rect 2402 4149 2409 4160
rect 2461 4190 2468 4201
rect 2802 4201 2868 4202
rect 2802 4190 2809 4201
rect 2461 4160 2809 4190
rect 2461 4149 2468 4160
rect 2402 4148 2468 4149
rect 2802 4149 2809 4160
rect 2861 4190 2868 4201
rect 3202 4201 3268 4202
rect 3202 4190 3209 4201
rect 2861 4160 3209 4190
rect 2861 4149 2868 4160
rect 2802 4148 2868 4149
rect 3202 4149 3209 4160
rect 3261 4190 3268 4201
rect 3602 4201 3668 4202
rect 3602 4190 3609 4201
rect 3261 4160 3609 4190
rect 3261 4149 3268 4160
rect 3202 4148 3268 4149
rect 3602 4149 3609 4160
rect 3661 4190 3668 4201
rect 4002 4201 4068 4202
rect 4002 4190 4009 4201
rect 3661 4160 4009 4190
rect 3661 4149 3668 4160
rect 3602 4148 3668 4149
rect 4002 4149 4009 4160
rect 4061 4190 4068 4201
rect 4402 4201 4468 4202
rect 4402 4190 4409 4201
rect 4061 4160 4409 4190
rect 4061 4149 4068 4160
rect 4002 4148 4068 4149
rect 4402 4149 4409 4160
rect 4461 4190 4468 4201
rect 4802 4201 4868 4202
rect 4802 4190 4809 4201
rect 4461 4160 4809 4190
rect 4461 4149 4468 4160
rect 4402 4148 4468 4149
rect 4802 4149 4809 4160
rect 4861 4190 4868 4201
rect 5202 4201 5268 4202
rect 5202 4190 5209 4201
rect 4861 4160 5209 4190
rect 4861 4149 4868 4160
rect 4802 4148 4868 4149
rect 5202 4149 5209 4160
rect 5261 4190 5268 4201
rect 5602 4201 5668 4202
rect 5602 4190 5609 4201
rect 5261 4160 5609 4190
rect 5261 4149 5268 4160
rect 5202 4148 5268 4149
rect 5602 4149 5609 4160
rect 5661 4190 5668 4201
rect 6002 4201 6068 4202
rect 6002 4190 6009 4201
rect 5661 4160 6009 4190
rect 5661 4149 5668 4160
rect 5602 4148 5668 4149
rect 6002 4149 6009 4160
rect 6061 4190 6068 4201
rect 6402 4201 6468 4202
rect 6402 4190 6409 4201
rect 6061 4160 6409 4190
rect 6061 4149 6068 4160
rect 6002 4148 6068 4149
rect 6402 4149 6409 4160
rect 6461 4190 6468 4201
rect 6802 4201 6868 4202
rect 6802 4190 6809 4201
rect 6461 4160 6809 4190
rect 6461 4149 6468 4160
rect 6402 4148 6468 4149
rect 6802 4149 6809 4160
rect 6861 4190 6868 4201
rect 7202 4201 7268 4202
rect 7202 4190 7209 4201
rect 6861 4160 7209 4190
rect 6861 4149 6868 4160
rect 6802 4148 6868 4149
rect 7202 4149 7209 4160
rect 7261 4190 7268 4201
rect 7602 4201 7668 4202
rect 7602 4190 7609 4201
rect 7261 4160 7609 4190
rect 7261 4149 7268 4160
rect 7202 4148 7268 4149
rect 7602 4149 7609 4160
rect 7661 4190 7668 4201
rect 8002 4201 8068 4202
rect 8002 4190 8009 4201
rect 7661 4160 8009 4190
rect 7661 4149 7668 4160
rect 7602 4148 7668 4149
rect 8002 4149 8009 4160
rect 8061 4190 8068 4201
rect 8402 4201 8468 4202
rect 8402 4190 8409 4201
rect 8061 4160 8409 4190
rect 8061 4149 8068 4160
rect 8002 4148 8068 4149
rect 8402 4149 8409 4160
rect 8461 4190 8468 4201
rect 8802 4201 8868 4202
rect 8802 4190 8809 4201
rect 8461 4160 8809 4190
rect 8461 4149 8468 4160
rect 8402 4148 8468 4149
rect 8802 4149 8809 4160
rect 8861 4190 8868 4201
rect 9202 4201 9268 4202
rect 9202 4190 9209 4201
rect 8861 4160 9209 4190
rect 8861 4149 8868 4160
rect 8802 4148 8868 4149
rect 9202 4149 9209 4160
rect 9261 4190 9268 4201
rect 9602 4201 9668 4202
rect 9602 4190 9609 4201
rect 9261 4160 9609 4190
rect 9261 4149 9268 4160
rect 9202 4148 9268 4149
rect 9602 4149 9609 4160
rect 9661 4190 9668 4201
rect 10002 4201 10068 4202
rect 10002 4190 10009 4201
rect 9661 4160 10009 4190
rect 9661 4149 9668 4160
rect 9602 4148 9668 4149
rect 10002 4149 10009 4160
rect 10061 4190 10068 4201
rect 10402 4201 10468 4202
rect 10402 4190 10409 4201
rect 10061 4160 10409 4190
rect 10061 4149 10068 4160
rect 10002 4148 10068 4149
rect 10402 4149 10409 4160
rect 10461 4190 10468 4201
rect 10802 4201 10868 4202
rect 10802 4190 10809 4201
rect 10461 4160 10809 4190
rect 10461 4149 10468 4160
rect 10402 4148 10468 4149
rect 10802 4149 10809 4160
rect 10861 4190 10868 4201
rect 11202 4201 11268 4202
rect 11202 4190 11209 4201
rect 10861 4160 11209 4190
rect 10861 4149 10868 4160
rect 10802 4148 10868 4149
rect 11202 4149 11209 4160
rect 11261 4190 11268 4201
rect 11602 4201 11668 4202
rect 11602 4190 11609 4201
rect 11261 4160 11609 4190
rect 11261 4149 11268 4160
rect 11202 4148 11268 4149
rect 11602 4149 11609 4160
rect 11661 4190 11668 4201
rect 12002 4201 12068 4202
rect 12002 4190 12009 4201
rect 11661 4160 12009 4190
rect 11661 4149 11668 4160
rect 11602 4148 11668 4149
rect 12002 4149 12009 4160
rect 12061 4190 12068 4201
rect 12402 4201 12468 4202
rect 12402 4190 12409 4201
rect 12061 4160 12409 4190
rect 12061 4149 12068 4160
rect 12002 4148 12068 4149
rect 12402 4149 12409 4160
rect 12461 4190 12468 4201
rect 12802 4201 12868 4202
rect 12802 4190 12809 4201
rect 12461 4160 12809 4190
rect 12461 4149 12468 4160
rect 12402 4148 12468 4149
rect 12802 4149 12809 4160
rect 12861 4190 12868 4201
rect 12900 4201 12966 4202
rect 12900 4190 12907 4201
rect 12861 4160 12907 4190
rect 12861 4149 12868 4160
rect 12802 4148 12868 4149
rect 12900 4149 12907 4160
rect 12959 4149 12966 4201
rect 12900 4148 12966 4149
rect 202 4131 268 4132
rect 202 4120 209 4131
rect 0 4090 209 4120
rect 202 4079 209 4090
rect 261 4120 268 4131
rect 602 4131 668 4132
rect 602 4120 609 4131
rect 261 4090 609 4120
rect 261 4079 268 4090
rect 202 4078 268 4079
rect 602 4079 609 4090
rect 661 4120 668 4131
rect 1002 4131 1068 4132
rect 1002 4120 1009 4131
rect 661 4090 1009 4120
rect 661 4079 668 4090
rect 602 4078 668 4079
rect 1002 4079 1009 4090
rect 1061 4120 1068 4131
rect 1402 4131 1468 4132
rect 1402 4120 1409 4131
rect 1061 4090 1409 4120
rect 1061 4079 1068 4090
rect 1002 4078 1068 4079
rect 1402 4079 1409 4090
rect 1461 4120 1468 4131
rect 1802 4131 1868 4132
rect 1802 4120 1809 4131
rect 1461 4090 1809 4120
rect 1461 4079 1468 4090
rect 1402 4078 1468 4079
rect 1802 4079 1809 4090
rect 1861 4120 1868 4131
rect 2202 4131 2268 4132
rect 2202 4120 2209 4131
rect 1861 4090 2209 4120
rect 1861 4079 1868 4090
rect 1802 4078 1868 4079
rect 2202 4079 2209 4090
rect 2261 4120 2268 4131
rect 2602 4131 2668 4132
rect 2602 4120 2609 4131
rect 2261 4090 2609 4120
rect 2261 4079 2268 4090
rect 2202 4078 2268 4079
rect 2602 4079 2609 4090
rect 2661 4120 2668 4131
rect 3002 4131 3068 4132
rect 3002 4120 3009 4131
rect 2661 4090 3009 4120
rect 2661 4079 2668 4090
rect 2602 4078 2668 4079
rect 3002 4079 3009 4090
rect 3061 4120 3068 4131
rect 3402 4131 3468 4132
rect 3402 4120 3409 4131
rect 3061 4090 3409 4120
rect 3061 4079 3068 4090
rect 3002 4078 3068 4079
rect 3402 4079 3409 4090
rect 3461 4120 3468 4131
rect 3802 4131 3868 4132
rect 3802 4120 3809 4131
rect 3461 4090 3809 4120
rect 3461 4079 3468 4090
rect 3402 4078 3468 4079
rect 3802 4079 3809 4090
rect 3861 4120 3868 4131
rect 4202 4131 4268 4132
rect 4202 4120 4209 4131
rect 3861 4090 4209 4120
rect 3861 4079 3868 4090
rect 3802 4078 3868 4079
rect 4202 4079 4209 4090
rect 4261 4120 4268 4131
rect 4602 4131 4668 4132
rect 4602 4120 4609 4131
rect 4261 4090 4609 4120
rect 4261 4079 4268 4090
rect 4202 4078 4268 4079
rect 4602 4079 4609 4090
rect 4661 4120 4668 4131
rect 5002 4131 5068 4132
rect 5002 4120 5009 4131
rect 4661 4090 5009 4120
rect 4661 4079 4668 4090
rect 4602 4078 4668 4079
rect 5002 4079 5009 4090
rect 5061 4120 5068 4131
rect 5402 4131 5468 4132
rect 5402 4120 5409 4131
rect 5061 4090 5409 4120
rect 5061 4079 5068 4090
rect 5002 4078 5068 4079
rect 5402 4079 5409 4090
rect 5461 4120 5468 4131
rect 5802 4131 5868 4132
rect 5802 4120 5809 4131
rect 5461 4090 5809 4120
rect 5461 4079 5468 4090
rect 5402 4078 5468 4079
rect 5802 4079 5809 4090
rect 5861 4120 5868 4131
rect 6202 4131 6268 4132
rect 6202 4120 6209 4131
rect 5861 4090 6209 4120
rect 5861 4079 5868 4090
rect 5802 4078 5868 4079
rect 6202 4079 6209 4090
rect 6261 4120 6268 4131
rect 6602 4131 6668 4132
rect 6602 4120 6609 4131
rect 6261 4090 6609 4120
rect 6261 4079 6268 4090
rect 6202 4078 6268 4079
rect 6602 4079 6609 4090
rect 6661 4120 6668 4131
rect 7002 4131 7068 4132
rect 7002 4120 7009 4131
rect 6661 4090 7009 4120
rect 6661 4079 6668 4090
rect 6602 4078 6668 4079
rect 7002 4079 7009 4090
rect 7061 4120 7068 4131
rect 7402 4131 7468 4132
rect 7402 4120 7409 4131
rect 7061 4090 7409 4120
rect 7061 4079 7068 4090
rect 7002 4078 7068 4079
rect 7402 4079 7409 4090
rect 7461 4120 7468 4131
rect 7802 4131 7868 4132
rect 7802 4120 7809 4131
rect 7461 4090 7809 4120
rect 7461 4079 7468 4090
rect 7402 4078 7468 4079
rect 7802 4079 7809 4090
rect 7861 4120 7868 4131
rect 8202 4131 8268 4132
rect 8202 4120 8209 4131
rect 7861 4090 8209 4120
rect 7861 4079 7868 4090
rect 7802 4078 7868 4079
rect 8202 4079 8209 4090
rect 8261 4120 8268 4131
rect 8602 4131 8668 4132
rect 8602 4120 8609 4131
rect 8261 4090 8609 4120
rect 8261 4079 8268 4090
rect 8202 4078 8268 4079
rect 8602 4079 8609 4090
rect 8661 4120 8668 4131
rect 9002 4131 9068 4132
rect 9002 4120 9009 4131
rect 8661 4090 9009 4120
rect 8661 4079 8668 4090
rect 8602 4078 8668 4079
rect 9002 4079 9009 4090
rect 9061 4120 9068 4131
rect 9402 4131 9468 4132
rect 9402 4120 9409 4131
rect 9061 4090 9409 4120
rect 9061 4079 9068 4090
rect 9002 4078 9068 4079
rect 9402 4079 9409 4090
rect 9461 4120 9468 4131
rect 9802 4131 9868 4132
rect 9802 4120 9809 4131
rect 9461 4090 9809 4120
rect 9461 4079 9468 4090
rect 9402 4078 9468 4079
rect 9802 4079 9809 4090
rect 9861 4120 9868 4131
rect 10202 4131 10268 4132
rect 10202 4120 10209 4131
rect 9861 4090 10209 4120
rect 9861 4079 9868 4090
rect 9802 4078 9868 4079
rect 10202 4079 10209 4090
rect 10261 4120 10268 4131
rect 10602 4131 10668 4132
rect 10602 4120 10609 4131
rect 10261 4090 10609 4120
rect 10261 4079 10268 4090
rect 10202 4078 10268 4079
rect 10602 4079 10609 4090
rect 10661 4120 10668 4131
rect 11002 4131 11068 4132
rect 11002 4120 11009 4131
rect 10661 4090 11009 4120
rect 10661 4079 10668 4090
rect 10602 4078 10668 4079
rect 11002 4079 11009 4090
rect 11061 4120 11068 4131
rect 11402 4131 11468 4132
rect 11402 4120 11409 4131
rect 11061 4090 11409 4120
rect 11061 4079 11068 4090
rect 11002 4078 11068 4079
rect 11402 4079 11409 4090
rect 11461 4120 11468 4131
rect 11802 4131 11868 4132
rect 11802 4120 11809 4131
rect 11461 4090 11809 4120
rect 11461 4079 11468 4090
rect 11402 4078 11468 4079
rect 11802 4079 11809 4090
rect 11861 4120 11868 4131
rect 12202 4131 12268 4132
rect 12202 4120 12209 4131
rect 11861 4090 12209 4120
rect 11861 4079 11868 4090
rect 11802 4078 11868 4079
rect 12202 4079 12209 4090
rect 12261 4120 12268 4131
rect 12602 4131 12668 4132
rect 12602 4120 12609 4131
rect 12261 4090 12609 4120
rect 12261 4079 12268 4090
rect 12202 4078 12268 4079
rect 12602 4079 12609 4090
rect 12661 4120 12668 4131
rect 13104 4131 13170 4132
rect 13104 4120 13111 4131
rect 12661 4090 13111 4120
rect 12661 4079 12668 4090
rect 12602 4078 12668 4079
rect 13104 4079 13111 4090
rect 13163 4079 13170 4131
rect 13104 4078 13170 4079
rect 2 4061 68 4062
rect 2 4050 9 4061
rect 0 4020 9 4050
rect 2 4009 9 4020
rect 61 4050 68 4061
rect 402 4061 468 4062
rect 402 4050 409 4061
rect 61 4020 409 4050
rect 61 4009 68 4020
rect 2 4008 68 4009
rect 402 4009 409 4020
rect 461 4050 468 4061
rect 802 4061 868 4062
rect 802 4050 809 4061
rect 461 4020 809 4050
rect 461 4009 468 4020
rect 402 4008 468 4009
rect 802 4009 809 4020
rect 861 4050 868 4061
rect 1202 4061 1268 4062
rect 1202 4050 1209 4061
rect 861 4020 1209 4050
rect 861 4009 868 4020
rect 802 4008 868 4009
rect 1202 4009 1209 4020
rect 1261 4050 1268 4061
rect 1602 4061 1668 4062
rect 1602 4050 1609 4061
rect 1261 4020 1609 4050
rect 1261 4009 1268 4020
rect 1202 4008 1268 4009
rect 1602 4009 1609 4020
rect 1661 4050 1668 4061
rect 2002 4061 2068 4062
rect 2002 4050 2009 4061
rect 1661 4020 2009 4050
rect 1661 4009 1668 4020
rect 1602 4008 1668 4009
rect 2002 4009 2009 4020
rect 2061 4050 2068 4061
rect 2402 4061 2468 4062
rect 2402 4050 2409 4061
rect 2061 4020 2409 4050
rect 2061 4009 2068 4020
rect 2002 4008 2068 4009
rect 2402 4009 2409 4020
rect 2461 4050 2468 4061
rect 2802 4061 2868 4062
rect 2802 4050 2809 4061
rect 2461 4020 2809 4050
rect 2461 4009 2468 4020
rect 2402 4008 2468 4009
rect 2802 4009 2809 4020
rect 2861 4050 2868 4061
rect 3202 4061 3268 4062
rect 3202 4050 3209 4061
rect 2861 4020 3209 4050
rect 2861 4009 2868 4020
rect 2802 4008 2868 4009
rect 3202 4009 3209 4020
rect 3261 4050 3268 4061
rect 3602 4061 3668 4062
rect 3602 4050 3609 4061
rect 3261 4020 3609 4050
rect 3261 4009 3268 4020
rect 3202 4008 3268 4009
rect 3602 4009 3609 4020
rect 3661 4050 3668 4061
rect 4002 4061 4068 4062
rect 4002 4050 4009 4061
rect 3661 4020 4009 4050
rect 3661 4009 3668 4020
rect 3602 4008 3668 4009
rect 4002 4009 4009 4020
rect 4061 4050 4068 4061
rect 4402 4061 4468 4062
rect 4402 4050 4409 4061
rect 4061 4020 4409 4050
rect 4061 4009 4068 4020
rect 4002 4008 4068 4009
rect 4402 4009 4409 4020
rect 4461 4050 4468 4061
rect 4802 4061 4868 4062
rect 4802 4050 4809 4061
rect 4461 4020 4809 4050
rect 4461 4009 4468 4020
rect 4402 4008 4468 4009
rect 4802 4009 4809 4020
rect 4861 4050 4868 4061
rect 5202 4061 5268 4062
rect 5202 4050 5209 4061
rect 4861 4020 5209 4050
rect 4861 4009 4868 4020
rect 4802 4008 4868 4009
rect 5202 4009 5209 4020
rect 5261 4050 5268 4061
rect 5602 4061 5668 4062
rect 5602 4050 5609 4061
rect 5261 4020 5609 4050
rect 5261 4009 5268 4020
rect 5202 4008 5268 4009
rect 5602 4009 5609 4020
rect 5661 4050 5668 4061
rect 6002 4061 6068 4062
rect 6002 4050 6009 4061
rect 5661 4020 6009 4050
rect 5661 4009 5668 4020
rect 5602 4008 5668 4009
rect 6002 4009 6009 4020
rect 6061 4050 6068 4061
rect 6402 4061 6468 4062
rect 6402 4050 6409 4061
rect 6061 4020 6409 4050
rect 6061 4009 6068 4020
rect 6002 4008 6068 4009
rect 6402 4009 6409 4020
rect 6461 4050 6468 4061
rect 6802 4061 6868 4062
rect 6802 4050 6809 4061
rect 6461 4020 6809 4050
rect 6461 4009 6468 4020
rect 6402 4008 6468 4009
rect 6802 4009 6809 4020
rect 6861 4050 6868 4061
rect 7202 4061 7268 4062
rect 7202 4050 7209 4061
rect 6861 4020 7209 4050
rect 6861 4009 6868 4020
rect 6802 4008 6868 4009
rect 7202 4009 7209 4020
rect 7261 4050 7268 4061
rect 7602 4061 7668 4062
rect 7602 4050 7609 4061
rect 7261 4020 7609 4050
rect 7261 4009 7268 4020
rect 7202 4008 7268 4009
rect 7602 4009 7609 4020
rect 7661 4050 7668 4061
rect 8002 4061 8068 4062
rect 8002 4050 8009 4061
rect 7661 4020 8009 4050
rect 7661 4009 7668 4020
rect 7602 4008 7668 4009
rect 8002 4009 8009 4020
rect 8061 4050 8068 4061
rect 8402 4061 8468 4062
rect 8402 4050 8409 4061
rect 8061 4020 8409 4050
rect 8061 4009 8068 4020
rect 8002 4008 8068 4009
rect 8402 4009 8409 4020
rect 8461 4050 8468 4061
rect 8802 4061 8868 4062
rect 8802 4050 8809 4061
rect 8461 4020 8809 4050
rect 8461 4009 8468 4020
rect 8402 4008 8468 4009
rect 8802 4009 8809 4020
rect 8861 4050 8868 4061
rect 9202 4061 9268 4062
rect 9202 4050 9209 4061
rect 8861 4020 9209 4050
rect 8861 4009 8868 4020
rect 8802 4008 8868 4009
rect 9202 4009 9209 4020
rect 9261 4050 9268 4061
rect 9602 4061 9668 4062
rect 9602 4050 9609 4061
rect 9261 4020 9609 4050
rect 9261 4009 9268 4020
rect 9202 4008 9268 4009
rect 9602 4009 9609 4020
rect 9661 4050 9668 4061
rect 10002 4061 10068 4062
rect 10002 4050 10009 4061
rect 9661 4020 10009 4050
rect 9661 4009 9668 4020
rect 9602 4008 9668 4009
rect 10002 4009 10009 4020
rect 10061 4050 10068 4061
rect 10402 4061 10468 4062
rect 10402 4050 10409 4061
rect 10061 4020 10409 4050
rect 10061 4009 10068 4020
rect 10002 4008 10068 4009
rect 10402 4009 10409 4020
rect 10461 4050 10468 4061
rect 10802 4061 10868 4062
rect 10802 4050 10809 4061
rect 10461 4020 10809 4050
rect 10461 4009 10468 4020
rect 10402 4008 10468 4009
rect 10802 4009 10809 4020
rect 10861 4050 10868 4061
rect 11202 4061 11268 4062
rect 11202 4050 11209 4061
rect 10861 4020 11209 4050
rect 10861 4009 10868 4020
rect 10802 4008 10868 4009
rect 11202 4009 11209 4020
rect 11261 4050 11268 4061
rect 11602 4061 11668 4062
rect 11602 4050 11609 4061
rect 11261 4020 11609 4050
rect 11261 4009 11268 4020
rect 11202 4008 11268 4009
rect 11602 4009 11609 4020
rect 11661 4050 11668 4061
rect 12002 4061 12068 4062
rect 12002 4050 12009 4061
rect 11661 4020 12009 4050
rect 11661 4009 11668 4020
rect 11602 4008 11668 4009
rect 12002 4009 12009 4020
rect 12061 4050 12068 4061
rect 12402 4061 12468 4062
rect 12402 4050 12409 4061
rect 12061 4020 12409 4050
rect 12061 4009 12068 4020
rect 12002 4008 12068 4009
rect 12402 4009 12409 4020
rect 12461 4050 12468 4061
rect 12802 4061 12868 4062
rect 12802 4050 12809 4061
rect 12461 4020 12809 4050
rect 12461 4009 12468 4020
rect 12402 4008 12468 4009
rect 12802 4009 12809 4020
rect 12861 4050 12868 4061
rect 12900 4061 12966 4062
rect 12900 4050 12907 4061
rect 12861 4020 12907 4050
rect 12861 4009 12868 4020
rect 12802 4008 12868 4009
rect 12900 4009 12907 4020
rect 12959 4009 12966 4061
rect 12900 4008 12966 4009
rect 202 3991 268 3992
rect 202 3980 209 3991
rect 0 3950 209 3980
rect 202 3939 209 3950
rect 261 3980 268 3991
rect 602 3991 668 3992
rect 602 3980 609 3991
rect 261 3950 609 3980
rect 261 3939 268 3950
rect 202 3938 268 3939
rect 602 3939 609 3950
rect 661 3980 668 3991
rect 1002 3991 1068 3992
rect 1002 3980 1009 3991
rect 661 3950 1009 3980
rect 661 3939 668 3950
rect 602 3938 668 3939
rect 1002 3939 1009 3950
rect 1061 3980 1068 3991
rect 1402 3991 1468 3992
rect 1402 3980 1409 3991
rect 1061 3950 1409 3980
rect 1061 3939 1068 3950
rect 1002 3938 1068 3939
rect 1402 3939 1409 3950
rect 1461 3980 1468 3991
rect 1802 3991 1868 3992
rect 1802 3980 1809 3991
rect 1461 3950 1809 3980
rect 1461 3939 1468 3950
rect 1402 3938 1468 3939
rect 1802 3939 1809 3950
rect 1861 3980 1868 3991
rect 2202 3991 2268 3992
rect 2202 3980 2209 3991
rect 1861 3950 2209 3980
rect 1861 3939 1868 3950
rect 1802 3938 1868 3939
rect 2202 3939 2209 3950
rect 2261 3980 2268 3991
rect 2602 3991 2668 3992
rect 2602 3980 2609 3991
rect 2261 3950 2609 3980
rect 2261 3939 2268 3950
rect 2202 3938 2268 3939
rect 2602 3939 2609 3950
rect 2661 3980 2668 3991
rect 3002 3991 3068 3992
rect 3002 3980 3009 3991
rect 2661 3950 3009 3980
rect 2661 3939 2668 3950
rect 2602 3938 2668 3939
rect 3002 3939 3009 3950
rect 3061 3980 3068 3991
rect 3402 3991 3468 3992
rect 3402 3980 3409 3991
rect 3061 3950 3409 3980
rect 3061 3939 3068 3950
rect 3002 3938 3068 3939
rect 3402 3939 3409 3950
rect 3461 3980 3468 3991
rect 3802 3991 3868 3992
rect 3802 3980 3809 3991
rect 3461 3950 3809 3980
rect 3461 3939 3468 3950
rect 3402 3938 3468 3939
rect 3802 3939 3809 3950
rect 3861 3980 3868 3991
rect 4202 3991 4268 3992
rect 4202 3980 4209 3991
rect 3861 3950 4209 3980
rect 3861 3939 3868 3950
rect 3802 3938 3868 3939
rect 4202 3939 4209 3950
rect 4261 3980 4268 3991
rect 4602 3991 4668 3992
rect 4602 3980 4609 3991
rect 4261 3950 4609 3980
rect 4261 3939 4268 3950
rect 4202 3938 4268 3939
rect 4602 3939 4609 3950
rect 4661 3980 4668 3991
rect 5002 3991 5068 3992
rect 5002 3980 5009 3991
rect 4661 3950 5009 3980
rect 4661 3939 4668 3950
rect 4602 3938 4668 3939
rect 5002 3939 5009 3950
rect 5061 3980 5068 3991
rect 5402 3991 5468 3992
rect 5402 3980 5409 3991
rect 5061 3950 5409 3980
rect 5061 3939 5068 3950
rect 5002 3938 5068 3939
rect 5402 3939 5409 3950
rect 5461 3980 5468 3991
rect 5802 3991 5868 3992
rect 5802 3980 5809 3991
rect 5461 3950 5809 3980
rect 5461 3939 5468 3950
rect 5402 3938 5468 3939
rect 5802 3939 5809 3950
rect 5861 3980 5868 3991
rect 6202 3991 6268 3992
rect 6202 3980 6209 3991
rect 5861 3950 6209 3980
rect 5861 3939 5868 3950
rect 5802 3938 5868 3939
rect 6202 3939 6209 3950
rect 6261 3980 6268 3991
rect 6602 3991 6668 3992
rect 6602 3980 6609 3991
rect 6261 3950 6609 3980
rect 6261 3939 6268 3950
rect 6202 3938 6268 3939
rect 6602 3939 6609 3950
rect 6661 3980 6668 3991
rect 7002 3991 7068 3992
rect 7002 3980 7009 3991
rect 6661 3950 7009 3980
rect 6661 3939 6668 3950
rect 6602 3938 6668 3939
rect 7002 3939 7009 3950
rect 7061 3980 7068 3991
rect 7402 3991 7468 3992
rect 7402 3980 7409 3991
rect 7061 3950 7409 3980
rect 7061 3939 7068 3950
rect 7002 3938 7068 3939
rect 7402 3939 7409 3950
rect 7461 3980 7468 3991
rect 7802 3991 7868 3992
rect 7802 3980 7809 3991
rect 7461 3950 7809 3980
rect 7461 3939 7468 3950
rect 7402 3938 7468 3939
rect 7802 3939 7809 3950
rect 7861 3980 7868 3991
rect 8202 3991 8268 3992
rect 8202 3980 8209 3991
rect 7861 3950 8209 3980
rect 7861 3939 7868 3950
rect 7802 3938 7868 3939
rect 8202 3939 8209 3950
rect 8261 3980 8268 3991
rect 8602 3991 8668 3992
rect 8602 3980 8609 3991
rect 8261 3950 8609 3980
rect 8261 3939 8268 3950
rect 8202 3938 8268 3939
rect 8602 3939 8609 3950
rect 8661 3980 8668 3991
rect 9002 3991 9068 3992
rect 9002 3980 9009 3991
rect 8661 3950 9009 3980
rect 8661 3939 8668 3950
rect 8602 3938 8668 3939
rect 9002 3939 9009 3950
rect 9061 3980 9068 3991
rect 9402 3991 9468 3992
rect 9402 3980 9409 3991
rect 9061 3950 9409 3980
rect 9061 3939 9068 3950
rect 9002 3938 9068 3939
rect 9402 3939 9409 3950
rect 9461 3980 9468 3991
rect 9802 3991 9868 3992
rect 9802 3980 9809 3991
rect 9461 3950 9809 3980
rect 9461 3939 9468 3950
rect 9402 3938 9468 3939
rect 9802 3939 9809 3950
rect 9861 3980 9868 3991
rect 10202 3991 10268 3992
rect 10202 3980 10209 3991
rect 9861 3950 10209 3980
rect 9861 3939 9868 3950
rect 9802 3938 9868 3939
rect 10202 3939 10209 3950
rect 10261 3980 10268 3991
rect 10602 3991 10668 3992
rect 10602 3980 10609 3991
rect 10261 3950 10609 3980
rect 10261 3939 10268 3950
rect 10202 3938 10268 3939
rect 10602 3939 10609 3950
rect 10661 3980 10668 3991
rect 11002 3991 11068 3992
rect 11002 3980 11009 3991
rect 10661 3950 11009 3980
rect 10661 3939 10668 3950
rect 10602 3938 10668 3939
rect 11002 3939 11009 3950
rect 11061 3980 11068 3991
rect 11402 3991 11468 3992
rect 11402 3980 11409 3991
rect 11061 3950 11409 3980
rect 11061 3939 11068 3950
rect 11002 3938 11068 3939
rect 11402 3939 11409 3950
rect 11461 3980 11468 3991
rect 11802 3991 11868 3992
rect 11802 3980 11809 3991
rect 11461 3950 11809 3980
rect 11461 3939 11468 3950
rect 11402 3938 11468 3939
rect 11802 3939 11809 3950
rect 11861 3980 11868 3991
rect 12202 3991 12268 3992
rect 12202 3980 12209 3991
rect 11861 3950 12209 3980
rect 11861 3939 11868 3950
rect 11802 3938 11868 3939
rect 12202 3939 12209 3950
rect 12261 3980 12268 3991
rect 12602 3991 12668 3992
rect 12602 3980 12609 3991
rect 12261 3950 12609 3980
rect 12261 3939 12268 3950
rect 12202 3938 12268 3939
rect 12602 3939 12609 3950
rect 12661 3980 12668 3991
rect 13104 3991 13170 3992
rect 13104 3980 13111 3991
rect 12661 3950 13111 3980
rect 12661 3939 12668 3950
rect 12602 3938 12668 3939
rect 13104 3939 13111 3950
rect 13163 3939 13170 3991
rect 13104 3938 13170 3939
rect 2 3921 68 3922
rect 2 3910 9 3921
rect 0 3880 9 3910
rect 2 3869 9 3880
rect 61 3910 68 3921
rect 402 3921 468 3922
rect 402 3910 409 3921
rect 61 3880 409 3910
rect 61 3869 68 3880
rect 2 3868 68 3869
rect 402 3869 409 3880
rect 461 3910 468 3921
rect 802 3921 868 3922
rect 802 3910 809 3921
rect 461 3880 809 3910
rect 461 3869 468 3880
rect 402 3868 468 3869
rect 802 3869 809 3880
rect 861 3910 868 3921
rect 1202 3921 1268 3922
rect 1202 3910 1209 3921
rect 861 3880 1209 3910
rect 861 3869 868 3880
rect 802 3868 868 3869
rect 1202 3869 1209 3880
rect 1261 3910 1268 3921
rect 1602 3921 1668 3922
rect 1602 3910 1609 3921
rect 1261 3880 1609 3910
rect 1261 3869 1268 3880
rect 1202 3868 1268 3869
rect 1602 3869 1609 3880
rect 1661 3910 1668 3921
rect 2002 3921 2068 3922
rect 2002 3910 2009 3921
rect 1661 3880 2009 3910
rect 1661 3869 1668 3880
rect 1602 3868 1668 3869
rect 2002 3869 2009 3880
rect 2061 3910 2068 3921
rect 2402 3921 2468 3922
rect 2402 3910 2409 3921
rect 2061 3880 2409 3910
rect 2061 3869 2068 3880
rect 2002 3868 2068 3869
rect 2402 3869 2409 3880
rect 2461 3910 2468 3921
rect 2802 3921 2868 3922
rect 2802 3910 2809 3921
rect 2461 3880 2809 3910
rect 2461 3869 2468 3880
rect 2402 3868 2468 3869
rect 2802 3869 2809 3880
rect 2861 3910 2868 3921
rect 3202 3921 3268 3922
rect 3202 3910 3209 3921
rect 2861 3880 3209 3910
rect 2861 3869 2868 3880
rect 2802 3868 2868 3869
rect 3202 3869 3209 3880
rect 3261 3910 3268 3921
rect 3602 3921 3668 3922
rect 3602 3910 3609 3921
rect 3261 3880 3609 3910
rect 3261 3869 3268 3880
rect 3202 3868 3268 3869
rect 3602 3869 3609 3880
rect 3661 3910 3668 3921
rect 4002 3921 4068 3922
rect 4002 3910 4009 3921
rect 3661 3880 4009 3910
rect 3661 3869 3668 3880
rect 3602 3868 3668 3869
rect 4002 3869 4009 3880
rect 4061 3910 4068 3921
rect 4402 3921 4468 3922
rect 4402 3910 4409 3921
rect 4061 3880 4409 3910
rect 4061 3869 4068 3880
rect 4002 3868 4068 3869
rect 4402 3869 4409 3880
rect 4461 3910 4468 3921
rect 4802 3921 4868 3922
rect 4802 3910 4809 3921
rect 4461 3880 4809 3910
rect 4461 3869 4468 3880
rect 4402 3868 4468 3869
rect 4802 3869 4809 3880
rect 4861 3910 4868 3921
rect 5202 3921 5268 3922
rect 5202 3910 5209 3921
rect 4861 3880 5209 3910
rect 4861 3869 4868 3880
rect 4802 3868 4868 3869
rect 5202 3869 5209 3880
rect 5261 3910 5268 3921
rect 5602 3921 5668 3922
rect 5602 3910 5609 3921
rect 5261 3880 5609 3910
rect 5261 3869 5268 3880
rect 5202 3868 5268 3869
rect 5602 3869 5609 3880
rect 5661 3910 5668 3921
rect 6002 3921 6068 3922
rect 6002 3910 6009 3921
rect 5661 3880 6009 3910
rect 5661 3869 5668 3880
rect 5602 3868 5668 3869
rect 6002 3869 6009 3880
rect 6061 3910 6068 3921
rect 6402 3921 6468 3922
rect 6402 3910 6409 3921
rect 6061 3880 6409 3910
rect 6061 3869 6068 3880
rect 6002 3868 6068 3869
rect 6402 3869 6409 3880
rect 6461 3910 6468 3921
rect 6802 3921 6868 3922
rect 6802 3910 6809 3921
rect 6461 3880 6809 3910
rect 6461 3869 6468 3880
rect 6402 3868 6468 3869
rect 6802 3869 6809 3880
rect 6861 3910 6868 3921
rect 7202 3921 7268 3922
rect 7202 3910 7209 3921
rect 6861 3880 7209 3910
rect 6861 3869 6868 3880
rect 6802 3868 6868 3869
rect 7202 3869 7209 3880
rect 7261 3910 7268 3921
rect 7602 3921 7668 3922
rect 7602 3910 7609 3921
rect 7261 3880 7609 3910
rect 7261 3869 7268 3880
rect 7202 3868 7268 3869
rect 7602 3869 7609 3880
rect 7661 3910 7668 3921
rect 8002 3921 8068 3922
rect 8002 3910 8009 3921
rect 7661 3880 8009 3910
rect 7661 3869 7668 3880
rect 7602 3868 7668 3869
rect 8002 3869 8009 3880
rect 8061 3910 8068 3921
rect 8402 3921 8468 3922
rect 8402 3910 8409 3921
rect 8061 3880 8409 3910
rect 8061 3869 8068 3880
rect 8002 3868 8068 3869
rect 8402 3869 8409 3880
rect 8461 3910 8468 3921
rect 8802 3921 8868 3922
rect 8802 3910 8809 3921
rect 8461 3880 8809 3910
rect 8461 3869 8468 3880
rect 8402 3868 8468 3869
rect 8802 3869 8809 3880
rect 8861 3910 8868 3921
rect 9202 3921 9268 3922
rect 9202 3910 9209 3921
rect 8861 3880 9209 3910
rect 8861 3869 8868 3880
rect 8802 3868 8868 3869
rect 9202 3869 9209 3880
rect 9261 3910 9268 3921
rect 9602 3921 9668 3922
rect 9602 3910 9609 3921
rect 9261 3880 9609 3910
rect 9261 3869 9268 3880
rect 9202 3868 9268 3869
rect 9602 3869 9609 3880
rect 9661 3910 9668 3921
rect 10002 3921 10068 3922
rect 10002 3910 10009 3921
rect 9661 3880 10009 3910
rect 9661 3869 9668 3880
rect 9602 3868 9668 3869
rect 10002 3869 10009 3880
rect 10061 3910 10068 3921
rect 10402 3921 10468 3922
rect 10402 3910 10409 3921
rect 10061 3880 10409 3910
rect 10061 3869 10068 3880
rect 10002 3868 10068 3869
rect 10402 3869 10409 3880
rect 10461 3910 10468 3921
rect 10802 3921 10868 3922
rect 10802 3910 10809 3921
rect 10461 3880 10809 3910
rect 10461 3869 10468 3880
rect 10402 3868 10468 3869
rect 10802 3869 10809 3880
rect 10861 3910 10868 3921
rect 11202 3921 11268 3922
rect 11202 3910 11209 3921
rect 10861 3880 11209 3910
rect 10861 3869 10868 3880
rect 10802 3868 10868 3869
rect 11202 3869 11209 3880
rect 11261 3910 11268 3921
rect 11602 3921 11668 3922
rect 11602 3910 11609 3921
rect 11261 3880 11609 3910
rect 11261 3869 11268 3880
rect 11202 3868 11268 3869
rect 11602 3869 11609 3880
rect 11661 3910 11668 3921
rect 12002 3921 12068 3922
rect 12002 3910 12009 3921
rect 11661 3880 12009 3910
rect 11661 3869 11668 3880
rect 11602 3868 11668 3869
rect 12002 3869 12009 3880
rect 12061 3910 12068 3921
rect 12402 3921 12468 3922
rect 12402 3910 12409 3921
rect 12061 3880 12409 3910
rect 12061 3869 12068 3880
rect 12002 3868 12068 3869
rect 12402 3869 12409 3880
rect 12461 3910 12468 3921
rect 12802 3921 12868 3922
rect 12802 3910 12809 3921
rect 12461 3880 12809 3910
rect 12461 3869 12468 3880
rect 12402 3868 12468 3869
rect 12802 3869 12809 3880
rect 12861 3910 12868 3921
rect 12900 3921 12966 3922
rect 12900 3910 12907 3921
rect 12861 3880 12907 3910
rect 12861 3869 12868 3880
rect 12802 3868 12868 3869
rect 12900 3869 12907 3880
rect 12959 3869 12966 3921
rect 12900 3868 12966 3869
rect 202 3851 268 3852
rect 202 3840 209 3851
rect 0 3810 209 3840
rect 202 3799 209 3810
rect 261 3840 268 3851
rect 602 3851 668 3852
rect 602 3840 609 3851
rect 261 3810 609 3840
rect 261 3799 268 3810
rect 202 3798 268 3799
rect 602 3799 609 3810
rect 661 3840 668 3851
rect 1002 3851 1068 3852
rect 1002 3840 1009 3851
rect 661 3810 1009 3840
rect 661 3799 668 3810
rect 602 3798 668 3799
rect 1002 3799 1009 3810
rect 1061 3840 1068 3851
rect 1402 3851 1468 3852
rect 1402 3840 1409 3851
rect 1061 3810 1409 3840
rect 1061 3799 1068 3810
rect 1002 3798 1068 3799
rect 1402 3799 1409 3810
rect 1461 3840 1468 3851
rect 1802 3851 1868 3852
rect 1802 3840 1809 3851
rect 1461 3810 1809 3840
rect 1461 3799 1468 3810
rect 1402 3798 1468 3799
rect 1802 3799 1809 3810
rect 1861 3840 1868 3851
rect 2202 3851 2268 3852
rect 2202 3840 2209 3851
rect 1861 3810 2209 3840
rect 1861 3799 1868 3810
rect 1802 3798 1868 3799
rect 2202 3799 2209 3810
rect 2261 3840 2268 3851
rect 2602 3851 2668 3852
rect 2602 3840 2609 3851
rect 2261 3810 2609 3840
rect 2261 3799 2268 3810
rect 2202 3798 2268 3799
rect 2602 3799 2609 3810
rect 2661 3840 2668 3851
rect 3002 3851 3068 3852
rect 3002 3840 3009 3851
rect 2661 3810 3009 3840
rect 2661 3799 2668 3810
rect 2602 3798 2668 3799
rect 3002 3799 3009 3810
rect 3061 3840 3068 3851
rect 3402 3851 3468 3852
rect 3402 3840 3409 3851
rect 3061 3810 3409 3840
rect 3061 3799 3068 3810
rect 3002 3798 3068 3799
rect 3402 3799 3409 3810
rect 3461 3840 3468 3851
rect 3802 3851 3868 3852
rect 3802 3840 3809 3851
rect 3461 3810 3809 3840
rect 3461 3799 3468 3810
rect 3402 3798 3468 3799
rect 3802 3799 3809 3810
rect 3861 3840 3868 3851
rect 4202 3851 4268 3852
rect 4202 3840 4209 3851
rect 3861 3810 4209 3840
rect 3861 3799 3868 3810
rect 3802 3798 3868 3799
rect 4202 3799 4209 3810
rect 4261 3840 4268 3851
rect 4602 3851 4668 3852
rect 4602 3840 4609 3851
rect 4261 3810 4609 3840
rect 4261 3799 4268 3810
rect 4202 3798 4268 3799
rect 4602 3799 4609 3810
rect 4661 3840 4668 3851
rect 5002 3851 5068 3852
rect 5002 3840 5009 3851
rect 4661 3810 5009 3840
rect 4661 3799 4668 3810
rect 4602 3798 4668 3799
rect 5002 3799 5009 3810
rect 5061 3840 5068 3851
rect 5402 3851 5468 3852
rect 5402 3840 5409 3851
rect 5061 3810 5409 3840
rect 5061 3799 5068 3810
rect 5002 3798 5068 3799
rect 5402 3799 5409 3810
rect 5461 3840 5468 3851
rect 5802 3851 5868 3852
rect 5802 3840 5809 3851
rect 5461 3810 5809 3840
rect 5461 3799 5468 3810
rect 5402 3798 5468 3799
rect 5802 3799 5809 3810
rect 5861 3840 5868 3851
rect 6202 3851 6268 3852
rect 6202 3840 6209 3851
rect 5861 3810 6209 3840
rect 5861 3799 5868 3810
rect 5802 3798 5868 3799
rect 6202 3799 6209 3810
rect 6261 3840 6268 3851
rect 6602 3851 6668 3852
rect 6602 3840 6609 3851
rect 6261 3810 6609 3840
rect 6261 3799 6268 3810
rect 6202 3798 6268 3799
rect 6602 3799 6609 3810
rect 6661 3840 6668 3851
rect 7002 3851 7068 3852
rect 7002 3840 7009 3851
rect 6661 3810 7009 3840
rect 6661 3799 6668 3810
rect 6602 3798 6668 3799
rect 7002 3799 7009 3810
rect 7061 3840 7068 3851
rect 7402 3851 7468 3852
rect 7402 3840 7409 3851
rect 7061 3810 7409 3840
rect 7061 3799 7068 3810
rect 7002 3798 7068 3799
rect 7402 3799 7409 3810
rect 7461 3840 7468 3851
rect 7802 3851 7868 3852
rect 7802 3840 7809 3851
rect 7461 3810 7809 3840
rect 7461 3799 7468 3810
rect 7402 3798 7468 3799
rect 7802 3799 7809 3810
rect 7861 3840 7868 3851
rect 8202 3851 8268 3852
rect 8202 3840 8209 3851
rect 7861 3810 8209 3840
rect 7861 3799 7868 3810
rect 7802 3798 7868 3799
rect 8202 3799 8209 3810
rect 8261 3840 8268 3851
rect 8602 3851 8668 3852
rect 8602 3840 8609 3851
rect 8261 3810 8609 3840
rect 8261 3799 8268 3810
rect 8202 3798 8268 3799
rect 8602 3799 8609 3810
rect 8661 3840 8668 3851
rect 9002 3851 9068 3852
rect 9002 3840 9009 3851
rect 8661 3810 9009 3840
rect 8661 3799 8668 3810
rect 8602 3798 8668 3799
rect 9002 3799 9009 3810
rect 9061 3840 9068 3851
rect 9402 3851 9468 3852
rect 9402 3840 9409 3851
rect 9061 3810 9409 3840
rect 9061 3799 9068 3810
rect 9002 3798 9068 3799
rect 9402 3799 9409 3810
rect 9461 3840 9468 3851
rect 9802 3851 9868 3852
rect 9802 3840 9809 3851
rect 9461 3810 9809 3840
rect 9461 3799 9468 3810
rect 9402 3798 9468 3799
rect 9802 3799 9809 3810
rect 9861 3840 9868 3851
rect 10202 3851 10268 3852
rect 10202 3840 10209 3851
rect 9861 3810 10209 3840
rect 9861 3799 9868 3810
rect 9802 3798 9868 3799
rect 10202 3799 10209 3810
rect 10261 3840 10268 3851
rect 10602 3851 10668 3852
rect 10602 3840 10609 3851
rect 10261 3810 10609 3840
rect 10261 3799 10268 3810
rect 10202 3798 10268 3799
rect 10602 3799 10609 3810
rect 10661 3840 10668 3851
rect 11002 3851 11068 3852
rect 11002 3840 11009 3851
rect 10661 3810 11009 3840
rect 10661 3799 10668 3810
rect 10602 3798 10668 3799
rect 11002 3799 11009 3810
rect 11061 3840 11068 3851
rect 11402 3851 11468 3852
rect 11402 3840 11409 3851
rect 11061 3810 11409 3840
rect 11061 3799 11068 3810
rect 11002 3798 11068 3799
rect 11402 3799 11409 3810
rect 11461 3840 11468 3851
rect 11802 3851 11868 3852
rect 11802 3840 11809 3851
rect 11461 3810 11809 3840
rect 11461 3799 11468 3810
rect 11402 3798 11468 3799
rect 11802 3799 11809 3810
rect 11861 3840 11868 3851
rect 12202 3851 12268 3852
rect 12202 3840 12209 3851
rect 11861 3810 12209 3840
rect 11861 3799 11868 3810
rect 11802 3798 11868 3799
rect 12202 3799 12209 3810
rect 12261 3840 12268 3851
rect 12602 3851 12668 3852
rect 12602 3840 12609 3851
rect 12261 3810 12609 3840
rect 12261 3799 12268 3810
rect 12202 3798 12268 3799
rect 12602 3799 12609 3810
rect 12661 3840 12668 3851
rect 13104 3851 13170 3852
rect 13104 3840 13111 3851
rect 12661 3810 13111 3840
rect 12661 3799 12668 3810
rect 12602 3798 12668 3799
rect 13104 3799 13111 3810
rect 13163 3799 13170 3851
rect 13104 3798 13170 3799
rect 2 3781 68 3782
rect 2 3770 9 3781
rect 0 3740 9 3770
rect 2 3729 9 3740
rect 61 3770 68 3781
rect 402 3781 468 3782
rect 402 3770 409 3781
rect 61 3740 409 3770
rect 61 3729 68 3740
rect 2 3728 68 3729
rect 402 3729 409 3740
rect 461 3770 468 3781
rect 802 3781 868 3782
rect 802 3770 809 3781
rect 461 3740 809 3770
rect 461 3729 468 3740
rect 402 3728 468 3729
rect 802 3729 809 3740
rect 861 3770 868 3781
rect 1202 3781 1268 3782
rect 1202 3770 1209 3781
rect 861 3740 1209 3770
rect 861 3729 868 3740
rect 802 3728 868 3729
rect 1202 3729 1209 3740
rect 1261 3770 1268 3781
rect 1602 3781 1668 3782
rect 1602 3770 1609 3781
rect 1261 3740 1609 3770
rect 1261 3729 1268 3740
rect 1202 3728 1268 3729
rect 1602 3729 1609 3740
rect 1661 3770 1668 3781
rect 2002 3781 2068 3782
rect 2002 3770 2009 3781
rect 1661 3740 2009 3770
rect 1661 3729 1668 3740
rect 1602 3728 1668 3729
rect 2002 3729 2009 3740
rect 2061 3770 2068 3781
rect 2402 3781 2468 3782
rect 2402 3770 2409 3781
rect 2061 3740 2409 3770
rect 2061 3729 2068 3740
rect 2002 3728 2068 3729
rect 2402 3729 2409 3740
rect 2461 3770 2468 3781
rect 2802 3781 2868 3782
rect 2802 3770 2809 3781
rect 2461 3740 2809 3770
rect 2461 3729 2468 3740
rect 2402 3728 2468 3729
rect 2802 3729 2809 3740
rect 2861 3770 2868 3781
rect 3202 3781 3268 3782
rect 3202 3770 3209 3781
rect 2861 3740 3209 3770
rect 2861 3729 2868 3740
rect 2802 3728 2868 3729
rect 3202 3729 3209 3740
rect 3261 3770 3268 3781
rect 3602 3781 3668 3782
rect 3602 3770 3609 3781
rect 3261 3740 3609 3770
rect 3261 3729 3268 3740
rect 3202 3728 3268 3729
rect 3602 3729 3609 3740
rect 3661 3770 3668 3781
rect 4002 3781 4068 3782
rect 4002 3770 4009 3781
rect 3661 3740 4009 3770
rect 3661 3729 3668 3740
rect 3602 3728 3668 3729
rect 4002 3729 4009 3740
rect 4061 3770 4068 3781
rect 4402 3781 4468 3782
rect 4402 3770 4409 3781
rect 4061 3740 4409 3770
rect 4061 3729 4068 3740
rect 4002 3728 4068 3729
rect 4402 3729 4409 3740
rect 4461 3770 4468 3781
rect 4802 3781 4868 3782
rect 4802 3770 4809 3781
rect 4461 3740 4809 3770
rect 4461 3729 4468 3740
rect 4402 3728 4468 3729
rect 4802 3729 4809 3740
rect 4861 3770 4868 3781
rect 5202 3781 5268 3782
rect 5202 3770 5209 3781
rect 4861 3740 5209 3770
rect 4861 3729 4868 3740
rect 4802 3728 4868 3729
rect 5202 3729 5209 3740
rect 5261 3770 5268 3781
rect 5602 3781 5668 3782
rect 5602 3770 5609 3781
rect 5261 3740 5609 3770
rect 5261 3729 5268 3740
rect 5202 3728 5268 3729
rect 5602 3729 5609 3740
rect 5661 3770 5668 3781
rect 6002 3781 6068 3782
rect 6002 3770 6009 3781
rect 5661 3740 6009 3770
rect 5661 3729 5668 3740
rect 5602 3728 5668 3729
rect 6002 3729 6009 3740
rect 6061 3770 6068 3781
rect 6402 3781 6468 3782
rect 6402 3770 6409 3781
rect 6061 3740 6409 3770
rect 6061 3729 6068 3740
rect 6002 3728 6068 3729
rect 6402 3729 6409 3740
rect 6461 3770 6468 3781
rect 6802 3781 6868 3782
rect 6802 3770 6809 3781
rect 6461 3740 6809 3770
rect 6461 3729 6468 3740
rect 6402 3728 6468 3729
rect 6802 3729 6809 3740
rect 6861 3770 6868 3781
rect 7202 3781 7268 3782
rect 7202 3770 7209 3781
rect 6861 3740 7209 3770
rect 6861 3729 6868 3740
rect 6802 3728 6868 3729
rect 7202 3729 7209 3740
rect 7261 3770 7268 3781
rect 7602 3781 7668 3782
rect 7602 3770 7609 3781
rect 7261 3740 7609 3770
rect 7261 3729 7268 3740
rect 7202 3728 7268 3729
rect 7602 3729 7609 3740
rect 7661 3770 7668 3781
rect 8002 3781 8068 3782
rect 8002 3770 8009 3781
rect 7661 3740 8009 3770
rect 7661 3729 7668 3740
rect 7602 3728 7668 3729
rect 8002 3729 8009 3740
rect 8061 3770 8068 3781
rect 8402 3781 8468 3782
rect 8402 3770 8409 3781
rect 8061 3740 8409 3770
rect 8061 3729 8068 3740
rect 8002 3728 8068 3729
rect 8402 3729 8409 3740
rect 8461 3770 8468 3781
rect 8802 3781 8868 3782
rect 8802 3770 8809 3781
rect 8461 3740 8809 3770
rect 8461 3729 8468 3740
rect 8402 3728 8468 3729
rect 8802 3729 8809 3740
rect 8861 3770 8868 3781
rect 9202 3781 9268 3782
rect 9202 3770 9209 3781
rect 8861 3740 9209 3770
rect 8861 3729 8868 3740
rect 8802 3728 8868 3729
rect 9202 3729 9209 3740
rect 9261 3770 9268 3781
rect 9602 3781 9668 3782
rect 9602 3770 9609 3781
rect 9261 3740 9609 3770
rect 9261 3729 9268 3740
rect 9202 3728 9268 3729
rect 9602 3729 9609 3740
rect 9661 3770 9668 3781
rect 10002 3781 10068 3782
rect 10002 3770 10009 3781
rect 9661 3740 10009 3770
rect 9661 3729 9668 3740
rect 9602 3728 9668 3729
rect 10002 3729 10009 3740
rect 10061 3770 10068 3781
rect 10402 3781 10468 3782
rect 10402 3770 10409 3781
rect 10061 3740 10409 3770
rect 10061 3729 10068 3740
rect 10002 3728 10068 3729
rect 10402 3729 10409 3740
rect 10461 3770 10468 3781
rect 10802 3781 10868 3782
rect 10802 3770 10809 3781
rect 10461 3740 10809 3770
rect 10461 3729 10468 3740
rect 10402 3728 10468 3729
rect 10802 3729 10809 3740
rect 10861 3770 10868 3781
rect 11202 3781 11268 3782
rect 11202 3770 11209 3781
rect 10861 3740 11209 3770
rect 10861 3729 10868 3740
rect 10802 3728 10868 3729
rect 11202 3729 11209 3740
rect 11261 3770 11268 3781
rect 11602 3781 11668 3782
rect 11602 3770 11609 3781
rect 11261 3740 11609 3770
rect 11261 3729 11268 3740
rect 11202 3728 11268 3729
rect 11602 3729 11609 3740
rect 11661 3770 11668 3781
rect 12002 3781 12068 3782
rect 12002 3770 12009 3781
rect 11661 3740 12009 3770
rect 11661 3729 11668 3740
rect 11602 3728 11668 3729
rect 12002 3729 12009 3740
rect 12061 3770 12068 3781
rect 12402 3781 12468 3782
rect 12402 3770 12409 3781
rect 12061 3740 12409 3770
rect 12061 3729 12068 3740
rect 12002 3728 12068 3729
rect 12402 3729 12409 3740
rect 12461 3770 12468 3781
rect 12802 3781 12868 3782
rect 12802 3770 12809 3781
rect 12461 3740 12809 3770
rect 12461 3729 12468 3740
rect 12402 3728 12468 3729
rect 12802 3729 12809 3740
rect 12861 3770 12868 3781
rect 12900 3781 12966 3782
rect 12900 3770 12907 3781
rect 12861 3740 12907 3770
rect 12861 3729 12868 3740
rect 12802 3728 12868 3729
rect 12900 3729 12907 3740
rect 12959 3729 12966 3781
rect 12900 3728 12966 3729
rect 196 3711 274 3712
rect -4 3695 74 3696
rect -4 3639 7 3695
rect 63 3639 74 3695
rect 196 3655 207 3711
rect 263 3655 274 3711
rect 596 3711 674 3712
rect 196 3654 274 3655
rect 396 3695 474 3696
rect -4 3638 74 3639
rect 396 3639 407 3695
rect 463 3639 474 3695
rect 596 3655 607 3711
rect 663 3655 674 3711
rect 996 3711 1074 3712
rect 596 3654 674 3655
rect 796 3695 874 3696
rect 396 3638 474 3639
rect 796 3639 807 3695
rect 863 3639 874 3695
rect 996 3655 1007 3711
rect 1063 3655 1074 3711
rect 1396 3711 1474 3712
rect 996 3654 1074 3655
rect 1196 3695 1274 3696
rect 796 3638 874 3639
rect 1196 3639 1207 3695
rect 1263 3639 1274 3695
rect 1396 3655 1407 3711
rect 1463 3655 1474 3711
rect 1796 3711 1874 3712
rect 1396 3654 1474 3655
rect 1596 3695 1674 3696
rect 1196 3638 1274 3639
rect 1596 3639 1607 3695
rect 1663 3639 1674 3695
rect 1796 3655 1807 3711
rect 1863 3655 1874 3711
rect 2196 3711 2274 3712
rect 1796 3654 1874 3655
rect 1996 3695 2074 3696
rect 1596 3638 1674 3639
rect 1996 3639 2007 3695
rect 2063 3639 2074 3695
rect 2196 3655 2207 3711
rect 2263 3655 2274 3711
rect 2596 3711 2674 3712
rect 2196 3654 2274 3655
rect 2396 3695 2474 3696
rect 1996 3638 2074 3639
rect 2396 3639 2407 3695
rect 2463 3639 2474 3695
rect 2596 3655 2607 3711
rect 2663 3655 2674 3711
rect 2996 3711 3074 3712
rect 2596 3654 2674 3655
rect 2796 3695 2874 3696
rect 2396 3638 2474 3639
rect 2796 3639 2807 3695
rect 2863 3639 2874 3695
rect 2996 3655 3007 3711
rect 3063 3655 3074 3711
rect 3396 3711 3474 3712
rect 2996 3654 3074 3655
rect 3196 3695 3274 3696
rect 2796 3638 2874 3639
rect 3196 3639 3207 3695
rect 3263 3639 3274 3695
rect 3396 3655 3407 3711
rect 3463 3655 3474 3711
rect 3796 3711 3874 3712
rect 3396 3654 3474 3655
rect 3596 3695 3674 3696
rect 3196 3638 3274 3639
rect 3596 3639 3607 3695
rect 3663 3639 3674 3695
rect 3796 3655 3807 3711
rect 3863 3655 3874 3711
rect 4196 3711 4274 3712
rect 3796 3654 3874 3655
rect 3996 3695 4074 3696
rect 3596 3638 3674 3639
rect 3996 3639 4007 3695
rect 4063 3639 4074 3695
rect 4196 3655 4207 3711
rect 4263 3655 4274 3711
rect 4596 3711 4674 3712
rect 4196 3654 4274 3655
rect 4396 3695 4474 3696
rect 3996 3638 4074 3639
rect 4396 3639 4407 3695
rect 4463 3639 4474 3695
rect 4596 3655 4607 3711
rect 4663 3655 4674 3711
rect 4996 3711 5074 3712
rect 4596 3654 4674 3655
rect 4796 3695 4874 3696
rect 4396 3638 4474 3639
rect 4796 3639 4807 3695
rect 4863 3639 4874 3695
rect 4996 3655 5007 3711
rect 5063 3655 5074 3711
rect 5396 3711 5474 3712
rect 4996 3654 5074 3655
rect 5196 3695 5274 3696
rect 4796 3638 4874 3639
rect 5196 3639 5207 3695
rect 5263 3639 5274 3695
rect 5396 3655 5407 3711
rect 5463 3655 5474 3711
rect 5796 3711 5874 3712
rect 5396 3654 5474 3655
rect 5596 3695 5674 3696
rect 5196 3638 5274 3639
rect 5596 3639 5607 3695
rect 5663 3639 5674 3695
rect 5796 3655 5807 3711
rect 5863 3655 5874 3711
rect 6196 3711 6274 3712
rect 5796 3654 5874 3655
rect 5996 3695 6074 3696
rect 5596 3638 5674 3639
rect 5996 3639 6007 3695
rect 6063 3639 6074 3695
rect 6196 3655 6207 3711
rect 6263 3655 6274 3711
rect 6596 3711 6674 3712
rect 6196 3654 6274 3655
rect 6396 3695 6474 3696
rect 5996 3638 6074 3639
rect 6396 3639 6407 3695
rect 6463 3639 6474 3695
rect 6596 3655 6607 3711
rect 6663 3655 6674 3711
rect 6996 3711 7074 3712
rect 6596 3654 6674 3655
rect 6796 3695 6874 3696
rect 6396 3638 6474 3639
rect 6796 3639 6807 3695
rect 6863 3639 6874 3695
rect 6996 3655 7007 3711
rect 7063 3655 7074 3711
rect 7396 3711 7474 3712
rect 6996 3654 7074 3655
rect 7196 3695 7274 3696
rect 6796 3638 6874 3639
rect 7196 3639 7207 3695
rect 7263 3639 7274 3695
rect 7396 3655 7407 3711
rect 7463 3655 7474 3711
rect 7796 3711 7874 3712
rect 7396 3654 7474 3655
rect 7596 3695 7674 3696
rect 7196 3638 7274 3639
rect 7596 3639 7607 3695
rect 7663 3639 7674 3695
rect 7796 3655 7807 3711
rect 7863 3655 7874 3711
rect 8196 3711 8274 3712
rect 7796 3654 7874 3655
rect 7996 3695 8074 3696
rect 7596 3638 7674 3639
rect 7996 3639 8007 3695
rect 8063 3639 8074 3695
rect 8196 3655 8207 3711
rect 8263 3655 8274 3711
rect 8596 3711 8674 3712
rect 8196 3654 8274 3655
rect 8396 3695 8474 3696
rect 7996 3638 8074 3639
rect 8396 3639 8407 3695
rect 8463 3639 8474 3695
rect 8596 3655 8607 3711
rect 8663 3655 8674 3711
rect 8996 3711 9074 3712
rect 8596 3654 8674 3655
rect 8796 3695 8874 3696
rect 8396 3638 8474 3639
rect 8796 3639 8807 3695
rect 8863 3639 8874 3695
rect 8996 3655 9007 3711
rect 9063 3655 9074 3711
rect 9396 3711 9474 3712
rect 8996 3654 9074 3655
rect 9196 3695 9274 3696
rect 8796 3638 8874 3639
rect 9196 3639 9207 3695
rect 9263 3639 9274 3695
rect 9396 3655 9407 3711
rect 9463 3655 9474 3711
rect 9796 3711 9874 3712
rect 9396 3654 9474 3655
rect 9596 3695 9674 3696
rect 9196 3638 9274 3639
rect 9596 3639 9607 3695
rect 9663 3639 9674 3695
rect 9796 3655 9807 3711
rect 9863 3655 9874 3711
rect 10196 3711 10274 3712
rect 9796 3654 9874 3655
rect 9996 3695 10074 3696
rect 9596 3638 9674 3639
rect 9996 3639 10007 3695
rect 10063 3639 10074 3695
rect 10196 3655 10207 3711
rect 10263 3655 10274 3711
rect 10596 3711 10674 3712
rect 10196 3654 10274 3655
rect 10396 3695 10474 3696
rect 9996 3638 10074 3639
rect 10396 3639 10407 3695
rect 10463 3639 10474 3695
rect 10596 3655 10607 3711
rect 10663 3655 10674 3711
rect 10996 3711 11074 3712
rect 10596 3654 10674 3655
rect 10796 3695 10874 3696
rect 10396 3638 10474 3639
rect 10796 3639 10807 3695
rect 10863 3639 10874 3695
rect 10996 3655 11007 3711
rect 11063 3655 11074 3711
rect 11396 3711 11474 3712
rect 10996 3654 11074 3655
rect 11196 3695 11274 3696
rect 10796 3638 10874 3639
rect 11196 3639 11207 3695
rect 11263 3639 11274 3695
rect 11396 3655 11407 3711
rect 11463 3655 11474 3711
rect 11796 3711 11874 3712
rect 11396 3654 11474 3655
rect 11596 3695 11674 3696
rect 11196 3638 11274 3639
rect 11596 3639 11607 3695
rect 11663 3639 11674 3695
rect 11796 3655 11807 3711
rect 11863 3655 11874 3711
rect 12196 3711 12274 3712
rect 11796 3654 11874 3655
rect 11996 3695 12074 3696
rect 11596 3638 11674 3639
rect 11996 3639 12007 3695
rect 12063 3639 12074 3695
rect 12196 3655 12207 3711
rect 12263 3655 12274 3711
rect 12596 3711 12674 3712
rect 12196 3654 12274 3655
rect 12396 3695 12474 3696
rect 11996 3638 12074 3639
rect 12396 3639 12407 3695
rect 12463 3639 12474 3695
rect 12596 3655 12607 3711
rect 12663 3655 12674 3711
rect 12596 3654 12674 3655
rect 12396 3638 12474 3639
rect 202 3621 268 3622
rect 202 3610 209 3621
rect 0 3580 209 3610
rect 202 3569 209 3580
rect 261 3610 268 3621
rect 602 3621 668 3622
rect 602 3610 609 3621
rect 261 3580 609 3610
rect 261 3569 268 3580
rect 202 3568 268 3569
rect 602 3569 609 3580
rect 661 3610 668 3621
rect 1002 3621 1068 3622
rect 1002 3610 1009 3621
rect 661 3580 1009 3610
rect 661 3569 668 3580
rect 602 3568 668 3569
rect 1002 3569 1009 3580
rect 1061 3610 1068 3621
rect 1402 3621 1468 3622
rect 1402 3610 1409 3621
rect 1061 3580 1409 3610
rect 1061 3569 1068 3580
rect 1002 3568 1068 3569
rect 1402 3569 1409 3580
rect 1461 3610 1468 3621
rect 1802 3621 1868 3622
rect 1802 3610 1809 3621
rect 1461 3580 1809 3610
rect 1461 3569 1468 3580
rect 1402 3568 1468 3569
rect 1802 3569 1809 3580
rect 1861 3610 1868 3621
rect 2202 3621 2268 3622
rect 2202 3610 2209 3621
rect 1861 3580 2209 3610
rect 1861 3569 1868 3580
rect 1802 3568 1868 3569
rect 2202 3569 2209 3580
rect 2261 3610 2268 3621
rect 2602 3621 2668 3622
rect 2602 3610 2609 3621
rect 2261 3580 2609 3610
rect 2261 3569 2268 3580
rect 2202 3568 2268 3569
rect 2602 3569 2609 3580
rect 2661 3610 2668 3621
rect 3002 3621 3068 3622
rect 3002 3610 3009 3621
rect 2661 3580 3009 3610
rect 2661 3569 2668 3580
rect 2602 3568 2668 3569
rect 3002 3569 3009 3580
rect 3061 3610 3068 3621
rect 3402 3621 3468 3622
rect 3402 3610 3409 3621
rect 3061 3580 3409 3610
rect 3061 3569 3068 3580
rect 3002 3568 3068 3569
rect 3402 3569 3409 3580
rect 3461 3610 3468 3621
rect 3802 3621 3868 3622
rect 3802 3610 3809 3621
rect 3461 3580 3809 3610
rect 3461 3569 3468 3580
rect 3402 3568 3468 3569
rect 3802 3569 3809 3580
rect 3861 3610 3868 3621
rect 4202 3621 4268 3622
rect 4202 3610 4209 3621
rect 3861 3580 4209 3610
rect 3861 3569 3868 3580
rect 3802 3568 3868 3569
rect 4202 3569 4209 3580
rect 4261 3610 4268 3621
rect 4602 3621 4668 3622
rect 4602 3610 4609 3621
rect 4261 3580 4609 3610
rect 4261 3569 4268 3580
rect 4202 3568 4268 3569
rect 4602 3569 4609 3580
rect 4661 3610 4668 3621
rect 5002 3621 5068 3622
rect 5002 3610 5009 3621
rect 4661 3580 5009 3610
rect 4661 3569 4668 3580
rect 4602 3568 4668 3569
rect 5002 3569 5009 3580
rect 5061 3610 5068 3621
rect 5402 3621 5468 3622
rect 5402 3610 5409 3621
rect 5061 3580 5409 3610
rect 5061 3569 5068 3580
rect 5002 3568 5068 3569
rect 5402 3569 5409 3580
rect 5461 3610 5468 3621
rect 5802 3621 5868 3622
rect 5802 3610 5809 3621
rect 5461 3580 5809 3610
rect 5461 3569 5468 3580
rect 5402 3568 5468 3569
rect 5802 3569 5809 3580
rect 5861 3610 5868 3621
rect 6202 3621 6268 3622
rect 6202 3610 6209 3621
rect 5861 3580 6209 3610
rect 5861 3569 5868 3580
rect 5802 3568 5868 3569
rect 6202 3569 6209 3580
rect 6261 3610 6268 3621
rect 6602 3621 6668 3622
rect 6602 3610 6609 3621
rect 6261 3580 6609 3610
rect 6261 3569 6268 3580
rect 6202 3568 6268 3569
rect 6602 3569 6609 3580
rect 6661 3610 6668 3621
rect 7002 3621 7068 3622
rect 7002 3610 7009 3621
rect 6661 3580 7009 3610
rect 6661 3569 6668 3580
rect 6602 3568 6668 3569
rect 7002 3569 7009 3580
rect 7061 3610 7068 3621
rect 7402 3621 7468 3622
rect 7402 3610 7409 3621
rect 7061 3580 7409 3610
rect 7061 3569 7068 3580
rect 7002 3568 7068 3569
rect 7402 3569 7409 3580
rect 7461 3610 7468 3621
rect 7802 3621 7868 3622
rect 7802 3610 7809 3621
rect 7461 3580 7809 3610
rect 7461 3569 7468 3580
rect 7402 3568 7468 3569
rect 7802 3569 7809 3580
rect 7861 3610 7868 3621
rect 8202 3621 8268 3622
rect 8202 3610 8209 3621
rect 7861 3580 8209 3610
rect 7861 3569 7868 3580
rect 7802 3568 7868 3569
rect 8202 3569 8209 3580
rect 8261 3610 8268 3621
rect 8602 3621 8668 3622
rect 8602 3610 8609 3621
rect 8261 3580 8609 3610
rect 8261 3569 8268 3580
rect 8202 3568 8268 3569
rect 8602 3569 8609 3580
rect 8661 3610 8668 3621
rect 9002 3621 9068 3622
rect 9002 3610 9009 3621
rect 8661 3580 9009 3610
rect 8661 3569 8668 3580
rect 8602 3568 8668 3569
rect 9002 3569 9009 3580
rect 9061 3610 9068 3621
rect 9402 3621 9468 3622
rect 9402 3610 9409 3621
rect 9061 3580 9409 3610
rect 9061 3569 9068 3580
rect 9002 3568 9068 3569
rect 9402 3569 9409 3580
rect 9461 3610 9468 3621
rect 9802 3621 9868 3622
rect 9802 3610 9809 3621
rect 9461 3580 9809 3610
rect 9461 3569 9468 3580
rect 9402 3568 9468 3569
rect 9802 3569 9809 3580
rect 9861 3610 9868 3621
rect 10202 3621 10268 3622
rect 10202 3610 10209 3621
rect 9861 3580 10209 3610
rect 9861 3569 9868 3580
rect 9802 3568 9868 3569
rect 10202 3569 10209 3580
rect 10261 3610 10268 3621
rect 10602 3621 10668 3622
rect 10602 3610 10609 3621
rect 10261 3580 10609 3610
rect 10261 3569 10268 3580
rect 10202 3568 10268 3569
rect 10602 3569 10609 3580
rect 10661 3610 10668 3621
rect 11002 3621 11068 3622
rect 11002 3610 11009 3621
rect 10661 3580 11009 3610
rect 10661 3569 10668 3580
rect 10602 3568 10668 3569
rect 11002 3569 11009 3580
rect 11061 3610 11068 3621
rect 11402 3621 11468 3622
rect 11402 3610 11409 3621
rect 11061 3580 11409 3610
rect 11061 3569 11068 3580
rect 11002 3568 11068 3569
rect 11402 3569 11409 3580
rect 11461 3610 11468 3621
rect 11802 3621 11868 3622
rect 11802 3610 11809 3621
rect 11461 3580 11809 3610
rect 11461 3569 11468 3580
rect 11402 3568 11468 3569
rect 11802 3569 11809 3580
rect 11861 3610 11868 3621
rect 12202 3621 12268 3622
rect 12202 3610 12209 3621
rect 11861 3580 12209 3610
rect 11861 3569 11868 3580
rect 11802 3568 11868 3569
rect 12202 3569 12209 3580
rect 12261 3610 12268 3621
rect 12602 3621 12668 3622
rect 12602 3610 12609 3621
rect 12261 3580 12609 3610
rect 12261 3569 12268 3580
rect 12202 3568 12268 3569
rect 12602 3569 12609 3580
rect 12661 3610 12668 3621
rect 13104 3621 13170 3622
rect 13104 3610 13111 3621
rect 12661 3580 13111 3610
rect 12661 3569 12668 3580
rect 12602 3568 12668 3569
rect 13104 3569 13111 3580
rect 13163 3569 13170 3621
rect 13104 3568 13170 3569
rect 2 3551 68 3552
rect 2 3540 9 3551
rect 0 3510 9 3540
rect 2 3499 9 3510
rect 61 3540 68 3551
rect 402 3551 468 3552
rect 402 3540 409 3551
rect 61 3510 409 3540
rect 61 3499 68 3510
rect 2 3498 68 3499
rect 402 3499 409 3510
rect 461 3540 468 3551
rect 802 3551 868 3552
rect 802 3540 809 3551
rect 461 3510 809 3540
rect 461 3499 468 3510
rect 402 3498 468 3499
rect 802 3499 809 3510
rect 861 3540 868 3551
rect 1202 3551 1268 3552
rect 1202 3540 1209 3551
rect 861 3510 1209 3540
rect 861 3499 868 3510
rect 802 3498 868 3499
rect 1202 3499 1209 3510
rect 1261 3540 1268 3551
rect 1602 3551 1668 3552
rect 1602 3540 1609 3551
rect 1261 3510 1609 3540
rect 1261 3499 1268 3510
rect 1202 3498 1268 3499
rect 1602 3499 1609 3510
rect 1661 3540 1668 3551
rect 2002 3551 2068 3552
rect 2002 3540 2009 3551
rect 1661 3510 2009 3540
rect 1661 3499 1668 3510
rect 1602 3498 1668 3499
rect 2002 3499 2009 3510
rect 2061 3540 2068 3551
rect 2402 3551 2468 3552
rect 2402 3540 2409 3551
rect 2061 3510 2409 3540
rect 2061 3499 2068 3510
rect 2002 3498 2068 3499
rect 2402 3499 2409 3510
rect 2461 3540 2468 3551
rect 2802 3551 2868 3552
rect 2802 3540 2809 3551
rect 2461 3510 2809 3540
rect 2461 3499 2468 3510
rect 2402 3498 2468 3499
rect 2802 3499 2809 3510
rect 2861 3540 2868 3551
rect 3202 3551 3268 3552
rect 3202 3540 3209 3551
rect 2861 3510 3209 3540
rect 2861 3499 2868 3510
rect 2802 3498 2868 3499
rect 3202 3499 3209 3510
rect 3261 3540 3268 3551
rect 3602 3551 3668 3552
rect 3602 3540 3609 3551
rect 3261 3510 3609 3540
rect 3261 3499 3268 3510
rect 3202 3498 3268 3499
rect 3602 3499 3609 3510
rect 3661 3540 3668 3551
rect 4002 3551 4068 3552
rect 4002 3540 4009 3551
rect 3661 3510 4009 3540
rect 3661 3499 3668 3510
rect 3602 3498 3668 3499
rect 4002 3499 4009 3510
rect 4061 3540 4068 3551
rect 4402 3551 4468 3552
rect 4402 3540 4409 3551
rect 4061 3510 4409 3540
rect 4061 3499 4068 3510
rect 4002 3498 4068 3499
rect 4402 3499 4409 3510
rect 4461 3540 4468 3551
rect 4802 3551 4868 3552
rect 4802 3540 4809 3551
rect 4461 3510 4809 3540
rect 4461 3499 4468 3510
rect 4402 3498 4468 3499
rect 4802 3499 4809 3510
rect 4861 3540 4868 3551
rect 5202 3551 5268 3552
rect 5202 3540 5209 3551
rect 4861 3510 5209 3540
rect 4861 3499 4868 3510
rect 4802 3498 4868 3499
rect 5202 3499 5209 3510
rect 5261 3540 5268 3551
rect 5602 3551 5668 3552
rect 5602 3540 5609 3551
rect 5261 3510 5609 3540
rect 5261 3499 5268 3510
rect 5202 3498 5268 3499
rect 5602 3499 5609 3510
rect 5661 3540 5668 3551
rect 6002 3551 6068 3552
rect 6002 3540 6009 3551
rect 5661 3510 6009 3540
rect 5661 3499 5668 3510
rect 5602 3498 5668 3499
rect 6002 3499 6009 3510
rect 6061 3540 6068 3551
rect 6402 3551 6468 3552
rect 6402 3540 6409 3551
rect 6061 3510 6409 3540
rect 6061 3499 6068 3510
rect 6002 3498 6068 3499
rect 6402 3499 6409 3510
rect 6461 3540 6468 3551
rect 6802 3551 6868 3552
rect 6802 3540 6809 3551
rect 6461 3510 6809 3540
rect 6461 3499 6468 3510
rect 6402 3498 6468 3499
rect 6802 3499 6809 3510
rect 6861 3540 6868 3551
rect 7202 3551 7268 3552
rect 7202 3540 7209 3551
rect 6861 3510 7209 3540
rect 6861 3499 6868 3510
rect 6802 3498 6868 3499
rect 7202 3499 7209 3510
rect 7261 3540 7268 3551
rect 7602 3551 7668 3552
rect 7602 3540 7609 3551
rect 7261 3510 7609 3540
rect 7261 3499 7268 3510
rect 7202 3498 7268 3499
rect 7602 3499 7609 3510
rect 7661 3540 7668 3551
rect 8002 3551 8068 3552
rect 8002 3540 8009 3551
rect 7661 3510 8009 3540
rect 7661 3499 7668 3510
rect 7602 3498 7668 3499
rect 8002 3499 8009 3510
rect 8061 3540 8068 3551
rect 8402 3551 8468 3552
rect 8402 3540 8409 3551
rect 8061 3510 8409 3540
rect 8061 3499 8068 3510
rect 8002 3498 8068 3499
rect 8402 3499 8409 3510
rect 8461 3540 8468 3551
rect 8802 3551 8868 3552
rect 8802 3540 8809 3551
rect 8461 3510 8809 3540
rect 8461 3499 8468 3510
rect 8402 3498 8468 3499
rect 8802 3499 8809 3510
rect 8861 3540 8868 3551
rect 9202 3551 9268 3552
rect 9202 3540 9209 3551
rect 8861 3510 9209 3540
rect 8861 3499 8868 3510
rect 8802 3498 8868 3499
rect 9202 3499 9209 3510
rect 9261 3540 9268 3551
rect 9602 3551 9668 3552
rect 9602 3540 9609 3551
rect 9261 3510 9609 3540
rect 9261 3499 9268 3510
rect 9202 3498 9268 3499
rect 9602 3499 9609 3510
rect 9661 3540 9668 3551
rect 10002 3551 10068 3552
rect 10002 3540 10009 3551
rect 9661 3510 10009 3540
rect 9661 3499 9668 3510
rect 9602 3498 9668 3499
rect 10002 3499 10009 3510
rect 10061 3540 10068 3551
rect 10402 3551 10468 3552
rect 10402 3540 10409 3551
rect 10061 3510 10409 3540
rect 10061 3499 10068 3510
rect 10002 3498 10068 3499
rect 10402 3499 10409 3510
rect 10461 3540 10468 3551
rect 10802 3551 10868 3552
rect 10802 3540 10809 3551
rect 10461 3510 10809 3540
rect 10461 3499 10468 3510
rect 10402 3498 10468 3499
rect 10802 3499 10809 3510
rect 10861 3540 10868 3551
rect 11202 3551 11268 3552
rect 11202 3540 11209 3551
rect 10861 3510 11209 3540
rect 10861 3499 10868 3510
rect 10802 3498 10868 3499
rect 11202 3499 11209 3510
rect 11261 3540 11268 3551
rect 11602 3551 11668 3552
rect 11602 3540 11609 3551
rect 11261 3510 11609 3540
rect 11261 3499 11268 3510
rect 11202 3498 11268 3499
rect 11602 3499 11609 3510
rect 11661 3540 11668 3551
rect 12002 3551 12068 3552
rect 12002 3540 12009 3551
rect 11661 3510 12009 3540
rect 11661 3499 11668 3510
rect 11602 3498 11668 3499
rect 12002 3499 12009 3510
rect 12061 3540 12068 3551
rect 12402 3551 12468 3552
rect 12402 3540 12409 3551
rect 12061 3510 12409 3540
rect 12061 3499 12068 3510
rect 12002 3498 12068 3499
rect 12402 3499 12409 3510
rect 12461 3540 12468 3551
rect 12802 3551 12868 3552
rect 12802 3540 12809 3551
rect 12461 3510 12809 3540
rect 12461 3499 12468 3510
rect 12402 3498 12468 3499
rect 12802 3499 12809 3510
rect 12861 3540 12868 3551
rect 12900 3551 12966 3552
rect 12900 3540 12907 3551
rect 12861 3510 12907 3540
rect 12861 3499 12868 3510
rect 12802 3498 12868 3499
rect 12900 3499 12907 3510
rect 12959 3499 12966 3551
rect 12900 3498 12966 3499
rect 202 3481 268 3482
rect 202 3470 209 3481
rect 0 3440 209 3470
rect 202 3429 209 3440
rect 261 3470 268 3481
rect 602 3481 668 3482
rect 602 3470 609 3481
rect 261 3440 609 3470
rect 261 3429 268 3440
rect 202 3428 268 3429
rect 602 3429 609 3440
rect 661 3470 668 3481
rect 1002 3481 1068 3482
rect 1002 3470 1009 3481
rect 661 3440 1009 3470
rect 661 3429 668 3440
rect 602 3428 668 3429
rect 1002 3429 1009 3440
rect 1061 3470 1068 3481
rect 1402 3481 1468 3482
rect 1402 3470 1409 3481
rect 1061 3440 1409 3470
rect 1061 3429 1068 3440
rect 1002 3428 1068 3429
rect 1402 3429 1409 3440
rect 1461 3470 1468 3481
rect 1802 3481 1868 3482
rect 1802 3470 1809 3481
rect 1461 3440 1809 3470
rect 1461 3429 1468 3440
rect 1402 3428 1468 3429
rect 1802 3429 1809 3440
rect 1861 3470 1868 3481
rect 2202 3481 2268 3482
rect 2202 3470 2209 3481
rect 1861 3440 2209 3470
rect 1861 3429 1868 3440
rect 1802 3428 1868 3429
rect 2202 3429 2209 3440
rect 2261 3470 2268 3481
rect 2602 3481 2668 3482
rect 2602 3470 2609 3481
rect 2261 3440 2609 3470
rect 2261 3429 2268 3440
rect 2202 3428 2268 3429
rect 2602 3429 2609 3440
rect 2661 3470 2668 3481
rect 3002 3481 3068 3482
rect 3002 3470 3009 3481
rect 2661 3440 3009 3470
rect 2661 3429 2668 3440
rect 2602 3428 2668 3429
rect 3002 3429 3009 3440
rect 3061 3470 3068 3481
rect 3402 3481 3468 3482
rect 3402 3470 3409 3481
rect 3061 3440 3409 3470
rect 3061 3429 3068 3440
rect 3002 3428 3068 3429
rect 3402 3429 3409 3440
rect 3461 3470 3468 3481
rect 3802 3481 3868 3482
rect 3802 3470 3809 3481
rect 3461 3440 3809 3470
rect 3461 3429 3468 3440
rect 3402 3428 3468 3429
rect 3802 3429 3809 3440
rect 3861 3470 3868 3481
rect 4202 3481 4268 3482
rect 4202 3470 4209 3481
rect 3861 3440 4209 3470
rect 3861 3429 3868 3440
rect 3802 3428 3868 3429
rect 4202 3429 4209 3440
rect 4261 3470 4268 3481
rect 4602 3481 4668 3482
rect 4602 3470 4609 3481
rect 4261 3440 4609 3470
rect 4261 3429 4268 3440
rect 4202 3428 4268 3429
rect 4602 3429 4609 3440
rect 4661 3470 4668 3481
rect 5002 3481 5068 3482
rect 5002 3470 5009 3481
rect 4661 3440 5009 3470
rect 4661 3429 4668 3440
rect 4602 3428 4668 3429
rect 5002 3429 5009 3440
rect 5061 3470 5068 3481
rect 5402 3481 5468 3482
rect 5402 3470 5409 3481
rect 5061 3440 5409 3470
rect 5061 3429 5068 3440
rect 5002 3428 5068 3429
rect 5402 3429 5409 3440
rect 5461 3470 5468 3481
rect 5802 3481 5868 3482
rect 5802 3470 5809 3481
rect 5461 3440 5809 3470
rect 5461 3429 5468 3440
rect 5402 3428 5468 3429
rect 5802 3429 5809 3440
rect 5861 3470 5868 3481
rect 6202 3481 6268 3482
rect 6202 3470 6209 3481
rect 5861 3440 6209 3470
rect 5861 3429 5868 3440
rect 5802 3428 5868 3429
rect 6202 3429 6209 3440
rect 6261 3470 6268 3481
rect 6602 3481 6668 3482
rect 6602 3470 6609 3481
rect 6261 3440 6609 3470
rect 6261 3429 6268 3440
rect 6202 3428 6268 3429
rect 6602 3429 6609 3440
rect 6661 3470 6668 3481
rect 7002 3481 7068 3482
rect 7002 3470 7009 3481
rect 6661 3440 7009 3470
rect 6661 3429 6668 3440
rect 6602 3428 6668 3429
rect 7002 3429 7009 3440
rect 7061 3470 7068 3481
rect 7402 3481 7468 3482
rect 7402 3470 7409 3481
rect 7061 3440 7409 3470
rect 7061 3429 7068 3440
rect 7002 3428 7068 3429
rect 7402 3429 7409 3440
rect 7461 3470 7468 3481
rect 7802 3481 7868 3482
rect 7802 3470 7809 3481
rect 7461 3440 7809 3470
rect 7461 3429 7468 3440
rect 7402 3428 7468 3429
rect 7802 3429 7809 3440
rect 7861 3470 7868 3481
rect 8202 3481 8268 3482
rect 8202 3470 8209 3481
rect 7861 3440 8209 3470
rect 7861 3429 7868 3440
rect 7802 3428 7868 3429
rect 8202 3429 8209 3440
rect 8261 3470 8268 3481
rect 8602 3481 8668 3482
rect 8602 3470 8609 3481
rect 8261 3440 8609 3470
rect 8261 3429 8268 3440
rect 8202 3428 8268 3429
rect 8602 3429 8609 3440
rect 8661 3470 8668 3481
rect 9002 3481 9068 3482
rect 9002 3470 9009 3481
rect 8661 3440 9009 3470
rect 8661 3429 8668 3440
rect 8602 3428 8668 3429
rect 9002 3429 9009 3440
rect 9061 3470 9068 3481
rect 9402 3481 9468 3482
rect 9402 3470 9409 3481
rect 9061 3440 9409 3470
rect 9061 3429 9068 3440
rect 9002 3428 9068 3429
rect 9402 3429 9409 3440
rect 9461 3470 9468 3481
rect 9802 3481 9868 3482
rect 9802 3470 9809 3481
rect 9461 3440 9809 3470
rect 9461 3429 9468 3440
rect 9402 3428 9468 3429
rect 9802 3429 9809 3440
rect 9861 3470 9868 3481
rect 10202 3481 10268 3482
rect 10202 3470 10209 3481
rect 9861 3440 10209 3470
rect 9861 3429 9868 3440
rect 9802 3428 9868 3429
rect 10202 3429 10209 3440
rect 10261 3470 10268 3481
rect 10602 3481 10668 3482
rect 10602 3470 10609 3481
rect 10261 3440 10609 3470
rect 10261 3429 10268 3440
rect 10202 3428 10268 3429
rect 10602 3429 10609 3440
rect 10661 3470 10668 3481
rect 11002 3481 11068 3482
rect 11002 3470 11009 3481
rect 10661 3440 11009 3470
rect 10661 3429 10668 3440
rect 10602 3428 10668 3429
rect 11002 3429 11009 3440
rect 11061 3470 11068 3481
rect 11402 3481 11468 3482
rect 11402 3470 11409 3481
rect 11061 3440 11409 3470
rect 11061 3429 11068 3440
rect 11002 3428 11068 3429
rect 11402 3429 11409 3440
rect 11461 3470 11468 3481
rect 11802 3481 11868 3482
rect 11802 3470 11809 3481
rect 11461 3440 11809 3470
rect 11461 3429 11468 3440
rect 11402 3428 11468 3429
rect 11802 3429 11809 3440
rect 11861 3470 11868 3481
rect 12202 3481 12268 3482
rect 12202 3470 12209 3481
rect 11861 3440 12209 3470
rect 11861 3429 11868 3440
rect 11802 3428 11868 3429
rect 12202 3429 12209 3440
rect 12261 3470 12268 3481
rect 12602 3481 12668 3482
rect 12602 3470 12609 3481
rect 12261 3440 12609 3470
rect 12261 3429 12268 3440
rect 12202 3428 12268 3429
rect 12602 3429 12609 3440
rect 12661 3470 12668 3481
rect 13104 3481 13170 3482
rect 13104 3470 13111 3481
rect 12661 3440 13111 3470
rect 12661 3429 12668 3440
rect 12602 3428 12668 3429
rect 13104 3429 13111 3440
rect 13163 3429 13170 3481
rect 13104 3428 13170 3429
rect 2 3411 68 3412
rect 2 3400 9 3411
rect 0 3370 9 3400
rect 2 3359 9 3370
rect 61 3400 68 3411
rect 402 3411 468 3412
rect 402 3400 409 3411
rect 61 3370 409 3400
rect 61 3359 68 3370
rect 2 3358 68 3359
rect 402 3359 409 3370
rect 461 3400 468 3411
rect 802 3411 868 3412
rect 802 3400 809 3411
rect 461 3370 809 3400
rect 461 3359 468 3370
rect 402 3358 468 3359
rect 802 3359 809 3370
rect 861 3400 868 3411
rect 1202 3411 1268 3412
rect 1202 3400 1209 3411
rect 861 3370 1209 3400
rect 861 3359 868 3370
rect 802 3358 868 3359
rect 1202 3359 1209 3370
rect 1261 3400 1268 3411
rect 1602 3411 1668 3412
rect 1602 3400 1609 3411
rect 1261 3370 1609 3400
rect 1261 3359 1268 3370
rect 1202 3358 1268 3359
rect 1602 3359 1609 3370
rect 1661 3400 1668 3411
rect 2002 3411 2068 3412
rect 2002 3400 2009 3411
rect 1661 3370 2009 3400
rect 1661 3359 1668 3370
rect 1602 3358 1668 3359
rect 2002 3359 2009 3370
rect 2061 3400 2068 3411
rect 2402 3411 2468 3412
rect 2402 3400 2409 3411
rect 2061 3370 2409 3400
rect 2061 3359 2068 3370
rect 2002 3358 2068 3359
rect 2402 3359 2409 3370
rect 2461 3400 2468 3411
rect 2802 3411 2868 3412
rect 2802 3400 2809 3411
rect 2461 3370 2809 3400
rect 2461 3359 2468 3370
rect 2402 3358 2468 3359
rect 2802 3359 2809 3370
rect 2861 3400 2868 3411
rect 3202 3411 3268 3412
rect 3202 3400 3209 3411
rect 2861 3370 3209 3400
rect 2861 3359 2868 3370
rect 2802 3358 2868 3359
rect 3202 3359 3209 3370
rect 3261 3400 3268 3411
rect 3602 3411 3668 3412
rect 3602 3400 3609 3411
rect 3261 3370 3609 3400
rect 3261 3359 3268 3370
rect 3202 3358 3268 3359
rect 3602 3359 3609 3370
rect 3661 3400 3668 3411
rect 4002 3411 4068 3412
rect 4002 3400 4009 3411
rect 3661 3370 4009 3400
rect 3661 3359 3668 3370
rect 3602 3358 3668 3359
rect 4002 3359 4009 3370
rect 4061 3400 4068 3411
rect 4402 3411 4468 3412
rect 4402 3400 4409 3411
rect 4061 3370 4409 3400
rect 4061 3359 4068 3370
rect 4002 3358 4068 3359
rect 4402 3359 4409 3370
rect 4461 3400 4468 3411
rect 4802 3411 4868 3412
rect 4802 3400 4809 3411
rect 4461 3370 4809 3400
rect 4461 3359 4468 3370
rect 4402 3358 4468 3359
rect 4802 3359 4809 3370
rect 4861 3400 4868 3411
rect 5202 3411 5268 3412
rect 5202 3400 5209 3411
rect 4861 3370 5209 3400
rect 4861 3359 4868 3370
rect 4802 3358 4868 3359
rect 5202 3359 5209 3370
rect 5261 3400 5268 3411
rect 5602 3411 5668 3412
rect 5602 3400 5609 3411
rect 5261 3370 5609 3400
rect 5261 3359 5268 3370
rect 5202 3358 5268 3359
rect 5602 3359 5609 3370
rect 5661 3400 5668 3411
rect 6002 3411 6068 3412
rect 6002 3400 6009 3411
rect 5661 3370 6009 3400
rect 5661 3359 5668 3370
rect 5602 3358 5668 3359
rect 6002 3359 6009 3370
rect 6061 3400 6068 3411
rect 6402 3411 6468 3412
rect 6402 3400 6409 3411
rect 6061 3370 6409 3400
rect 6061 3359 6068 3370
rect 6002 3358 6068 3359
rect 6402 3359 6409 3370
rect 6461 3400 6468 3411
rect 6802 3411 6868 3412
rect 6802 3400 6809 3411
rect 6461 3370 6809 3400
rect 6461 3359 6468 3370
rect 6402 3358 6468 3359
rect 6802 3359 6809 3370
rect 6861 3400 6868 3411
rect 7202 3411 7268 3412
rect 7202 3400 7209 3411
rect 6861 3370 7209 3400
rect 6861 3359 6868 3370
rect 6802 3358 6868 3359
rect 7202 3359 7209 3370
rect 7261 3400 7268 3411
rect 7602 3411 7668 3412
rect 7602 3400 7609 3411
rect 7261 3370 7609 3400
rect 7261 3359 7268 3370
rect 7202 3358 7268 3359
rect 7602 3359 7609 3370
rect 7661 3400 7668 3411
rect 8002 3411 8068 3412
rect 8002 3400 8009 3411
rect 7661 3370 8009 3400
rect 7661 3359 7668 3370
rect 7602 3358 7668 3359
rect 8002 3359 8009 3370
rect 8061 3400 8068 3411
rect 8402 3411 8468 3412
rect 8402 3400 8409 3411
rect 8061 3370 8409 3400
rect 8061 3359 8068 3370
rect 8002 3358 8068 3359
rect 8402 3359 8409 3370
rect 8461 3400 8468 3411
rect 8802 3411 8868 3412
rect 8802 3400 8809 3411
rect 8461 3370 8809 3400
rect 8461 3359 8468 3370
rect 8402 3358 8468 3359
rect 8802 3359 8809 3370
rect 8861 3400 8868 3411
rect 9202 3411 9268 3412
rect 9202 3400 9209 3411
rect 8861 3370 9209 3400
rect 8861 3359 8868 3370
rect 8802 3358 8868 3359
rect 9202 3359 9209 3370
rect 9261 3400 9268 3411
rect 9602 3411 9668 3412
rect 9602 3400 9609 3411
rect 9261 3370 9609 3400
rect 9261 3359 9268 3370
rect 9202 3358 9268 3359
rect 9602 3359 9609 3370
rect 9661 3400 9668 3411
rect 10002 3411 10068 3412
rect 10002 3400 10009 3411
rect 9661 3370 10009 3400
rect 9661 3359 9668 3370
rect 9602 3358 9668 3359
rect 10002 3359 10009 3370
rect 10061 3400 10068 3411
rect 10402 3411 10468 3412
rect 10402 3400 10409 3411
rect 10061 3370 10409 3400
rect 10061 3359 10068 3370
rect 10002 3358 10068 3359
rect 10402 3359 10409 3370
rect 10461 3400 10468 3411
rect 10802 3411 10868 3412
rect 10802 3400 10809 3411
rect 10461 3370 10809 3400
rect 10461 3359 10468 3370
rect 10402 3358 10468 3359
rect 10802 3359 10809 3370
rect 10861 3400 10868 3411
rect 11202 3411 11268 3412
rect 11202 3400 11209 3411
rect 10861 3370 11209 3400
rect 10861 3359 10868 3370
rect 10802 3358 10868 3359
rect 11202 3359 11209 3370
rect 11261 3400 11268 3411
rect 11602 3411 11668 3412
rect 11602 3400 11609 3411
rect 11261 3370 11609 3400
rect 11261 3359 11268 3370
rect 11202 3358 11268 3359
rect 11602 3359 11609 3370
rect 11661 3400 11668 3411
rect 12002 3411 12068 3412
rect 12002 3400 12009 3411
rect 11661 3370 12009 3400
rect 11661 3359 11668 3370
rect 11602 3358 11668 3359
rect 12002 3359 12009 3370
rect 12061 3400 12068 3411
rect 12402 3411 12468 3412
rect 12402 3400 12409 3411
rect 12061 3370 12409 3400
rect 12061 3359 12068 3370
rect 12002 3358 12068 3359
rect 12402 3359 12409 3370
rect 12461 3400 12468 3411
rect 12802 3411 12868 3412
rect 12802 3400 12809 3411
rect 12461 3370 12809 3400
rect 12461 3359 12468 3370
rect 12402 3358 12468 3359
rect 12802 3359 12809 3370
rect 12861 3400 12868 3411
rect 12900 3411 12966 3412
rect 12900 3400 12907 3411
rect 12861 3370 12907 3400
rect 12861 3359 12868 3370
rect 12802 3358 12868 3359
rect 12900 3359 12907 3370
rect 12959 3359 12966 3411
rect 12900 3358 12966 3359
rect 202 3341 268 3342
rect 202 3330 209 3341
rect 0 3300 209 3330
rect 202 3289 209 3300
rect 261 3330 268 3341
rect 602 3341 668 3342
rect 602 3330 609 3341
rect 261 3300 609 3330
rect 261 3289 268 3300
rect 202 3288 268 3289
rect 602 3289 609 3300
rect 661 3330 668 3341
rect 1002 3341 1068 3342
rect 1002 3330 1009 3341
rect 661 3300 1009 3330
rect 661 3289 668 3300
rect 602 3288 668 3289
rect 1002 3289 1009 3300
rect 1061 3330 1068 3341
rect 1402 3341 1468 3342
rect 1402 3330 1409 3341
rect 1061 3300 1409 3330
rect 1061 3289 1068 3300
rect 1002 3288 1068 3289
rect 1402 3289 1409 3300
rect 1461 3330 1468 3341
rect 1802 3341 1868 3342
rect 1802 3330 1809 3341
rect 1461 3300 1809 3330
rect 1461 3289 1468 3300
rect 1402 3288 1468 3289
rect 1802 3289 1809 3300
rect 1861 3330 1868 3341
rect 2202 3341 2268 3342
rect 2202 3330 2209 3341
rect 1861 3300 2209 3330
rect 1861 3289 1868 3300
rect 1802 3288 1868 3289
rect 2202 3289 2209 3300
rect 2261 3330 2268 3341
rect 2602 3341 2668 3342
rect 2602 3330 2609 3341
rect 2261 3300 2609 3330
rect 2261 3289 2268 3300
rect 2202 3288 2268 3289
rect 2602 3289 2609 3300
rect 2661 3330 2668 3341
rect 3002 3341 3068 3342
rect 3002 3330 3009 3341
rect 2661 3300 3009 3330
rect 2661 3289 2668 3300
rect 2602 3288 2668 3289
rect 3002 3289 3009 3300
rect 3061 3330 3068 3341
rect 3402 3341 3468 3342
rect 3402 3330 3409 3341
rect 3061 3300 3409 3330
rect 3061 3289 3068 3300
rect 3002 3288 3068 3289
rect 3402 3289 3409 3300
rect 3461 3330 3468 3341
rect 3802 3341 3868 3342
rect 3802 3330 3809 3341
rect 3461 3300 3809 3330
rect 3461 3289 3468 3300
rect 3402 3288 3468 3289
rect 3802 3289 3809 3300
rect 3861 3330 3868 3341
rect 4202 3341 4268 3342
rect 4202 3330 4209 3341
rect 3861 3300 4209 3330
rect 3861 3289 3868 3300
rect 3802 3288 3868 3289
rect 4202 3289 4209 3300
rect 4261 3330 4268 3341
rect 4602 3341 4668 3342
rect 4602 3330 4609 3341
rect 4261 3300 4609 3330
rect 4261 3289 4268 3300
rect 4202 3288 4268 3289
rect 4602 3289 4609 3300
rect 4661 3330 4668 3341
rect 5002 3341 5068 3342
rect 5002 3330 5009 3341
rect 4661 3300 5009 3330
rect 4661 3289 4668 3300
rect 4602 3288 4668 3289
rect 5002 3289 5009 3300
rect 5061 3330 5068 3341
rect 5402 3341 5468 3342
rect 5402 3330 5409 3341
rect 5061 3300 5409 3330
rect 5061 3289 5068 3300
rect 5002 3288 5068 3289
rect 5402 3289 5409 3300
rect 5461 3330 5468 3341
rect 5802 3341 5868 3342
rect 5802 3330 5809 3341
rect 5461 3300 5809 3330
rect 5461 3289 5468 3300
rect 5402 3288 5468 3289
rect 5802 3289 5809 3300
rect 5861 3330 5868 3341
rect 6202 3341 6268 3342
rect 6202 3330 6209 3341
rect 5861 3300 6209 3330
rect 5861 3289 5868 3300
rect 5802 3288 5868 3289
rect 6202 3289 6209 3300
rect 6261 3330 6268 3341
rect 6602 3341 6668 3342
rect 6602 3330 6609 3341
rect 6261 3300 6609 3330
rect 6261 3289 6268 3300
rect 6202 3288 6268 3289
rect 6602 3289 6609 3300
rect 6661 3330 6668 3341
rect 7002 3341 7068 3342
rect 7002 3330 7009 3341
rect 6661 3300 7009 3330
rect 6661 3289 6668 3300
rect 6602 3288 6668 3289
rect 7002 3289 7009 3300
rect 7061 3330 7068 3341
rect 7402 3341 7468 3342
rect 7402 3330 7409 3341
rect 7061 3300 7409 3330
rect 7061 3289 7068 3300
rect 7002 3288 7068 3289
rect 7402 3289 7409 3300
rect 7461 3330 7468 3341
rect 7802 3341 7868 3342
rect 7802 3330 7809 3341
rect 7461 3300 7809 3330
rect 7461 3289 7468 3300
rect 7402 3288 7468 3289
rect 7802 3289 7809 3300
rect 7861 3330 7868 3341
rect 8202 3341 8268 3342
rect 8202 3330 8209 3341
rect 7861 3300 8209 3330
rect 7861 3289 7868 3300
rect 7802 3288 7868 3289
rect 8202 3289 8209 3300
rect 8261 3330 8268 3341
rect 8602 3341 8668 3342
rect 8602 3330 8609 3341
rect 8261 3300 8609 3330
rect 8261 3289 8268 3300
rect 8202 3288 8268 3289
rect 8602 3289 8609 3300
rect 8661 3330 8668 3341
rect 9002 3341 9068 3342
rect 9002 3330 9009 3341
rect 8661 3300 9009 3330
rect 8661 3289 8668 3300
rect 8602 3288 8668 3289
rect 9002 3289 9009 3300
rect 9061 3330 9068 3341
rect 9402 3341 9468 3342
rect 9402 3330 9409 3341
rect 9061 3300 9409 3330
rect 9061 3289 9068 3300
rect 9002 3288 9068 3289
rect 9402 3289 9409 3300
rect 9461 3330 9468 3341
rect 9802 3341 9868 3342
rect 9802 3330 9809 3341
rect 9461 3300 9809 3330
rect 9461 3289 9468 3300
rect 9402 3288 9468 3289
rect 9802 3289 9809 3300
rect 9861 3330 9868 3341
rect 10202 3341 10268 3342
rect 10202 3330 10209 3341
rect 9861 3300 10209 3330
rect 9861 3289 9868 3300
rect 9802 3288 9868 3289
rect 10202 3289 10209 3300
rect 10261 3330 10268 3341
rect 10602 3341 10668 3342
rect 10602 3330 10609 3341
rect 10261 3300 10609 3330
rect 10261 3289 10268 3300
rect 10202 3288 10268 3289
rect 10602 3289 10609 3300
rect 10661 3330 10668 3341
rect 11002 3341 11068 3342
rect 11002 3330 11009 3341
rect 10661 3300 11009 3330
rect 10661 3289 10668 3300
rect 10602 3288 10668 3289
rect 11002 3289 11009 3300
rect 11061 3330 11068 3341
rect 11402 3341 11468 3342
rect 11402 3330 11409 3341
rect 11061 3300 11409 3330
rect 11061 3289 11068 3300
rect 11002 3288 11068 3289
rect 11402 3289 11409 3300
rect 11461 3330 11468 3341
rect 11802 3341 11868 3342
rect 11802 3330 11809 3341
rect 11461 3300 11809 3330
rect 11461 3289 11468 3300
rect 11402 3288 11468 3289
rect 11802 3289 11809 3300
rect 11861 3330 11868 3341
rect 12202 3341 12268 3342
rect 12202 3330 12209 3341
rect 11861 3300 12209 3330
rect 11861 3289 11868 3300
rect 11802 3288 11868 3289
rect 12202 3289 12209 3300
rect 12261 3330 12268 3341
rect 12602 3341 12668 3342
rect 12602 3330 12609 3341
rect 12261 3300 12609 3330
rect 12261 3289 12268 3300
rect 12202 3288 12268 3289
rect 12602 3289 12609 3300
rect 12661 3330 12668 3341
rect 13104 3341 13170 3342
rect 13104 3330 13111 3341
rect 12661 3300 13111 3330
rect 12661 3289 12668 3300
rect 12602 3288 12668 3289
rect 13104 3289 13111 3300
rect 13163 3289 13170 3341
rect 13104 3288 13170 3289
rect 2 3271 68 3272
rect 2 3260 9 3271
rect 0 3230 9 3260
rect 2 3219 9 3230
rect 61 3260 68 3271
rect 402 3271 468 3272
rect 402 3260 409 3271
rect 61 3230 409 3260
rect 61 3219 68 3230
rect 2 3218 68 3219
rect 402 3219 409 3230
rect 461 3260 468 3271
rect 802 3271 868 3272
rect 802 3260 809 3271
rect 461 3230 809 3260
rect 461 3219 468 3230
rect 402 3218 468 3219
rect 802 3219 809 3230
rect 861 3260 868 3271
rect 1202 3271 1268 3272
rect 1202 3260 1209 3271
rect 861 3230 1209 3260
rect 861 3219 868 3230
rect 802 3218 868 3219
rect 1202 3219 1209 3230
rect 1261 3260 1268 3271
rect 1602 3271 1668 3272
rect 1602 3260 1609 3271
rect 1261 3230 1609 3260
rect 1261 3219 1268 3230
rect 1202 3218 1268 3219
rect 1602 3219 1609 3230
rect 1661 3260 1668 3271
rect 2002 3271 2068 3272
rect 2002 3260 2009 3271
rect 1661 3230 2009 3260
rect 1661 3219 1668 3230
rect 1602 3218 1668 3219
rect 2002 3219 2009 3230
rect 2061 3260 2068 3271
rect 2402 3271 2468 3272
rect 2402 3260 2409 3271
rect 2061 3230 2409 3260
rect 2061 3219 2068 3230
rect 2002 3218 2068 3219
rect 2402 3219 2409 3230
rect 2461 3260 2468 3271
rect 2802 3271 2868 3272
rect 2802 3260 2809 3271
rect 2461 3230 2809 3260
rect 2461 3219 2468 3230
rect 2402 3218 2468 3219
rect 2802 3219 2809 3230
rect 2861 3260 2868 3271
rect 3202 3271 3268 3272
rect 3202 3260 3209 3271
rect 2861 3230 3209 3260
rect 2861 3219 2868 3230
rect 2802 3218 2868 3219
rect 3202 3219 3209 3230
rect 3261 3260 3268 3271
rect 3602 3271 3668 3272
rect 3602 3260 3609 3271
rect 3261 3230 3609 3260
rect 3261 3219 3268 3230
rect 3202 3218 3268 3219
rect 3602 3219 3609 3230
rect 3661 3260 3668 3271
rect 4002 3271 4068 3272
rect 4002 3260 4009 3271
rect 3661 3230 4009 3260
rect 3661 3219 3668 3230
rect 3602 3218 3668 3219
rect 4002 3219 4009 3230
rect 4061 3260 4068 3271
rect 4402 3271 4468 3272
rect 4402 3260 4409 3271
rect 4061 3230 4409 3260
rect 4061 3219 4068 3230
rect 4002 3218 4068 3219
rect 4402 3219 4409 3230
rect 4461 3260 4468 3271
rect 4802 3271 4868 3272
rect 4802 3260 4809 3271
rect 4461 3230 4809 3260
rect 4461 3219 4468 3230
rect 4402 3218 4468 3219
rect 4802 3219 4809 3230
rect 4861 3260 4868 3271
rect 5202 3271 5268 3272
rect 5202 3260 5209 3271
rect 4861 3230 5209 3260
rect 4861 3219 4868 3230
rect 4802 3218 4868 3219
rect 5202 3219 5209 3230
rect 5261 3260 5268 3271
rect 5602 3271 5668 3272
rect 5602 3260 5609 3271
rect 5261 3230 5609 3260
rect 5261 3219 5268 3230
rect 5202 3218 5268 3219
rect 5602 3219 5609 3230
rect 5661 3260 5668 3271
rect 6002 3271 6068 3272
rect 6002 3260 6009 3271
rect 5661 3230 6009 3260
rect 5661 3219 5668 3230
rect 5602 3218 5668 3219
rect 6002 3219 6009 3230
rect 6061 3260 6068 3271
rect 6402 3271 6468 3272
rect 6402 3260 6409 3271
rect 6061 3230 6409 3260
rect 6061 3219 6068 3230
rect 6002 3218 6068 3219
rect 6402 3219 6409 3230
rect 6461 3260 6468 3271
rect 6802 3271 6868 3272
rect 6802 3260 6809 3271
rect 6461 3230 6809 3260
rect 6461 3219 6468 3230
rect 6402 3218 6468 3219
rect 6802 3219 6809 3230
rect 6861 3260 6868 3271
rect 7202 3271 7268 3272
rect 7202 3260 7209 3271
rect 6861 3230 7209 3260
rect 6861 3219 6868 3230
rect 6802 3218 6868 3219
rect 7202 3219 7209 3230
rect 7261 3260 7268 3271
rect 7602 3271 7668 3272
rect 7602 3260 7609 3271
rect 7261 3230 7609 3260
rect 7261 3219 7268 3230
rect 7202 3218 7268 3219
rect 7602 3219 7609 3230
rect 7661 3260 7668 3271
rect 8002 3271 8068 3272
rect 8002 3260 8009 3271
rect 7661 3230 8009 3260
rect 7661 3219 7668 3230
rect 7602 3218 7668 3219
rect 8002 3219 8009 3230
rect 8061 3260 8068 3271
rect 8402 3271 8468 3272
rect 8402 3260 8409 3271
rect 8061 3230 8409 3260
rect 8061 3219 8068 3230
rect 8002 3218 8068 3219
rect 8402 3219 8409 3230
rect 8461 3260 8468 3271
rect 8802 3271 8868 3272
rect 8802 3260 8809 3271
rect 8461 3230 8809 3260
rect 8461 3219 8468 3230
rect 8402 3218 8468 3219
rect 8802 3219 8809 3230
rect 8861 3260 8868 3271
rect 9202 3271 9268 3272
rect 9202 3260 9209 3271
rect 8861 3230 9209 3260
rect 8861 3219 8868 3230
rect 8802 3218 8868 3219
rect 9202 3219 9209 3230
rect 9261 3260 9268 3271
rect 9602 3271 9668 3272
rect 9602 3260 9609 3271
rect 9261 3230 9609 3260
rect 9261 3219 9268 3230
rect 9202 3218 9268 3219
rect 9602 3219 9609 3230
rect 9661 3260 9668 3271
rect 10002 3271 10068 3272
rect 10002 3260 10009 3271
rect 9661 3230 10009 3260
rect 9661 3219 9668 3230
rect 9602 3218 9668 3219
rect 10002 3219 10009 3230
rect 10061 3260 10068 3271
rect 10402 3271 10468 3272
rect 10402 3260 10409 3271
rect 10061 3230 10409 3260
rect 10061 3219 10068 3230
rect 10002 3218 10068 3219
rect 10402 3219 10409 3230
rect 10461 3260 10468 3271
rect 10802 3271 10868 3272
rect 10802 3260 10809 3271
rect 10461 3230 10809 3260
rect 10461 3219 10468 3230
rect 10402 3218 10468 3219
rect 10802 3219 10809 3230
rect 10861 3260 10868 3271
rect 11202 3271 11268 3272
rect 11202 3260 11209 3271
rect 10861 3230 11209 3260
rect 10861 3219 10868 3230
rect 10802 3218 10868 3219
rect 11202 3219 11209 3230
rect 11261 3260 11268 3271
rect 11602 3271 11668 3272
rect 11602 3260 11609 3271
rect 11261 3230 11609 3260
rect 11261 3219 11268 3230
rect 11202 3218 11268 3219
rect 11602 3219 11609 3230
rect 11661 3260 11668 3271
rect 12002 3271 12068 3272
rect 12002 3260 12009 3271
rect 11661 3230 12009 3260
rect 11661 3219 11668 3230
rect 11602 3218 11668 3219
rect 12002 3219 12009 3230
rect 12061 3260 12068 3271
rect 12402 3271 12468 3272
rect 12402 3260 12409 3271
rect 12061 3230 12409 3260
rect 12061 3219 12068 3230
rect 12002 3218 12068 3219
rect 12402 3219 12409 3230
rect 12461 3260 12468 3271
rect 12802 3271 12868 3272
rect 12802 3260 12809 3271
rect 12461 3230 12809 3260
rect 12461 3219 12468 3230
rect 12402 3218 12468 3219
rect 12802 3219 12809 3230
rect 12861 3260 12868 3271
rect 12900 3271 12966 3272
rect 12900 3260 12907 3271
rect 12861 3230 12907 3260
rect 12861 3219 12868 3230
rect 12802 3218 12868 3219
rect 12900 3219 12907 3230
rect 12959 3219 12966 3271
rect 12900 3218 12966 3219
rect 202 3201 268 3202
rect 202 3190 209 3201
rect 0 3160 209 3190
rect 202 3149 209 3160
rect 261 3190 268 3201
rect 602 3201 668 3202
rect 602 3190 609 3201
rect 261 3160 609 3190
rect 261 3149 268 3160
rect 202 3148 268 3149
rect 602 3149 609 3160
rect 661 3190 668 3201
rect 1002 3201 1068 3202
rect 1002 3190 1009 3201
rect 661 3160 1009 3190
rect 661 3149 668 3160
rect 602 3148 668 3149
rect 1002 3149 1009 3160
rect 1061 3190 1068 3201
rect 1402 3201 1468 3202
rect 1402 3190 1409 3201
rect 1061 3160 1409 3190
rect 1061 3149 1068 3160
rect 1002 3148 1068 3149
rect 1402 3149 1409 3160
rect 1461 3190 1468 3201
rect 1802 3201 1868 3202
rect 1802 3190 1809 3201
rect 1461 3160 1809 3190
rect 1461 3149 1468 3160
rect 1402 3148 1468 3149
rect 1802 3149 1809 3160
rect 1861 3190 1868 3201
rect 2202 3201 2268 3202
rect 2202 3190 2209 3201
rect 1861 3160 2209 3190
rect 1861 3149 1868 3160
rect 1802 3148 1868 3149
rect 2202 3149 2209 3160
rect 2261 3190 2268 3201
rect 2602 3201 2668 3202
rect 2602 3190 2609 3201
rect 2261 3160 2609 3190
rect 2261 3149 2268 3160
rect 2202 3148 2268 3149
rect 2602 3149 2609 3160
rect 2661 3190 2668 3201
rect 3002 3201 3068 3202
rect 3002 3190 3009 3201
rect 2661 3160 3009 3190
rect 2661 3149 2668 3160
rect 2602 3148 2668 3149
rect 3002 3149 3009 3160
rect 3061 3190 3068 3201
rect 3402 3201 3468 3202
rect 3402 3190 3409 3201
rect 3061 3160 3409 3190
rect 3061 3149 3068 3160
rect 3002 3148 3068 3149
rect 3402 3149 3409 3160
rect 3461 3190 3468 3201
rect 3802 3201 3868 3202
rect 3802 3190 3809 3201
rect 3461 3160 3809 3190
rect 3461 3149 3468 3160
rect 3402 3148 3468 3149
rect 3802 3149 3809 3160
rect 3861 3190 3868 3201
rect 4202 3201 4268 3202
rect 4202 3190 4209 3201
rect 3861 3160 4209 3190
rect 3861 3149 3868 3160
rect 3802 3148 3868 3149
rect 4202 3149 4209 3160
rect 4261 3190 4268 3201
rect 4602 3201 4668 3202
rect 4602 3190 4609 3201
rect 4261 3160 4609 3190
rect 4261 3149 4268 3160
rect 4202 3148 4268 3149
rect 4602 3149 4609 3160
rect 4661 3190 4668 3201
rect 5002 3201 5068 3202
rect 5002 3190 5009 3201
rect 4661 3160 5009 3190
rect 4661 3149 4668 3160
rect 4602 3148 4668 3149
rect 5002 3149 5009 3160
rect 5061 3190 5068 3201
rect 5402 3201 5468 3202
rect 5402 3190 5409 3201
rect 5061 3160 5409 3190
rect 5061 3149 5068 3160
rect 5002 3148 5068 3149
rect 5402 3149 5409 3160
rect 5461 3190 5468 3201
rect 5802 3201 5868 3202
rect 5802 3190 5809 3201
rect 5461 3160 5809 3190
rect 5461 3149 5468 3160
rect 5402 3148 5468 3149
rect 5802 3149 5809 3160
rect 5861 3190 5868 3201
rect 6202 3201 6268 3202
rect 6202 3190 6209 3201
rect 5861 3160 6209 3190
rect 5861 3149 5868 3160
rect 5802 3148 5868 3149
rect 6202 3149 6209 3160
rect 6261 3190 6268 3201
rect 6602 3201 6668 3202
rect 6602 3190 6609 3201
rect 6261 3160 6609 3190
rect 6261 3149 6268 3160
rect 6202 3148 6268 3149
rect 6602 3149 6609 3160
rect 6661 3190 6668 3201
rect 7002 3201 7068 3202
rect 7002 3190 7009 3201
rect 6661 3160 7009 3190
rect 6661 3149 6668 3160
rect 6602 3148 6668 3149
rect 7002 3149 7009 3160
rect 7061 3190 7068 3201
rect 7402 3201 7468 3202
rect 7402 3190 7409 3201
rect 7061 3160 7409 3190
rect 7061 3149 7068 3160
rect 7002 3148 7068 3149
rect 7402 3149 7409 3160
rect 7461 3190 7468 3201
rect 7802 3201 7868 3202
rect 7802 3190 7809 3201
rect 7461 3160 7809 3190
rect 7461 3149 7468 3160
rect 7402 3148 7468 3149
rect 7802 3149 7809 3160
rect 7861 3190 7868 3201
rect 8202 3201 8268 3202
rect 8202 3190 8209 3201
rect 7861 3160 8209 3190
rect 7861 3149 7868 3160
rect 7802 3148 7868 3149
rect 8202 3149 8209 3160
rect 8261 3190 8268 3201
rect 8602 3201 8668 3202
rect 8602 3190 8609 3201
rect 8261 3160 8609 3190
rect 8261 3149 8268 3160
rect 8202 3148 8268 3149
rect 8602 3149 8609 3160
rect 8661 3190 8668 3201
rect 9002 3201 9068 3202
rect 9002 3190 9009 3201
rect 8661 3160 9009 3190
rect 8661 3149 8668 3160
rect 8602 3148 8668 3149
rect 9002 3149 9009 3160
rect 9061 3190 9068 3201
rect 9402 3201 9468 3202
rect 9402 3190 9409 3201
rect 9061 3160 9409 3190
rect 9061 3149 9068 3160
rect 9002 3148 9068 3149
rect 9402 3149 9409 3160
rect 9461 3190 9468 3201
rect 9802 3201 9868 3202
rect 9802 3190 9809 3201
rect 9461 3160 9809 3190
rect 9461 3149 9468 3160
rect 9402 3148 9468 3149
rect 9802 3149 9809 3160
rect 9861 3190 9868 3201
rect 10202 3201 10268 3202
rect 10202 3190 10209 3201
rect 9861 3160 10209 3190
rect 9861 3149 9868 3160
rect 9802 3148 9868 3149
rect 10202 3149 10209 3160
rect 10261 3190 10268 3201
rect 10602 3201 10668 3202
rect 10602 3190 10609 3201
rect 10261 3160 10609 3190
rect 10261 3149 10268 3160
rect 10202 3148 10268 3149
rect 10602 3149 10609 3160
rect 10661 3190 10668 3201
rect 11002 3201 11068 3202
rect 11002 3190 11009 3201
rect 10661 3160 11009 3190
rect 10661 3149 10668 3160
rect 10602 3148 10668 3149
rect 11002 3149 11009 3160
rect 11061 3190 11068 3201
rect 11402 3201 11468 3202
rect 11402 3190 11409 3201
rect 11061 3160 11409 3190
rect 11061 3149 11068 3160
rect 11002 3148 11068 3149
rect 11402 3149 11409 3160
rect 11461 3190 11468 3201
rect 11802 3201 11868 3202
rect 11802 3190 11809 3201
rect 11461 3160 11809 3190
rect 11461 3149 11468 3160
rect 11402 3148 11468 3149
rect 11802 3149 11809 3160
rect 11861 3190 11868 3201
rect 12202 3201 12268 3202
rect 12202 3190 12209 3201
rect 11861 3160 12209 3190
rect 11861 3149 11868 3160
rect 11802 3148 11868 3149
rect 12202 3149 12209 3160
rect 12261 3190 12268 3201
rect 12602 3201 12668 3202
rect 12602 3190 12609 3201
rect 12261 3160 12609 3190
rect 12261 3149 12268 3160
rect 12202 3148 12268 3149
rect 12602 3149 12609 3160
rect 12661 3190 12668 3201
rect 13104 3201 13170 3202
rect 13104 3190 13111 3201
rect 12661 3160 13111 3190
rect 12661 3149 12668 3160
rect 12602 3148 12668 3149
rect 13104 3149 13111 3160
rect 13163 3149 13170 3201
rect 13104 3148 13170 3149
rect 2 3131 68 3132
rect 2 3120 9 3131
rect 0 3090 9 3120
rect 2 3079 9 3090
rect 61 3120 68 3131
rect 402 3131 468 3132
rect 402 3120 409 3131
rect 61 3090 409 3120
rect 61 3079 68 3090
rect 2 3078 68 3079
rect 402 3079 409 3090
rect 461 3120 468 3131
rect 802 3131 868 3132
rect 802 3120 809 3131
rect 461 3090 809 3120
rect 461 3079 468 3090
rect 402 3078 468 3079
rect 802 3079 809 3090
rect 861 3120 868 3131
rect 1202 3131 1268 3132
rect 1202 3120 1209 3131
rect 861 3090 1209 3120
rect 861 3079 868 3090
rect 802 3078 868 3079
rect 1202 3079 1209 3090
rect 1261 3120 1268 3131
rect 1602 3131 1668 3132
rect 1602 3120 1609 3131
rect 1261 3090 1609 3120
rect 1261 3079 1268 3090
rect 1202 3078 1268 3079
rect 1602 3079 1609 3090
rect 1661 3120 1668 3131
rect 2002 3131 2068 3132
rect 2002 3120 2009 3131
rect 1661 3090 2009 3120
rect 1661 3079 1668 3090
rect 1602 3078 1668 3079
rect 2002 3079 2009 3090
rect 2061 3120 2068 3131
rect 2402 3131 2468 3132
rect 2402 3120 2409 3131
rect 2061 3090 2409 3120
rect 2061 3079 2068 3090
rect 2002 3078 2068 3079
rect 2402 3079 2409 3090
rect 2461 3120 2468 3131
rect 2802 3131 2868 3132
rect 2802 3120 2809 3131
rect 2461 3090 2809 3120
rect 2461 3079 2468 3090
rect 2402 3078 2468 3079
rect 2802 3079 2809 3090
rect 2861 3120 2868 3131
rect 3202 3131 3268 3132
rect 3202 3120 3209 3131
rect 2861 3090 3209 3120
rect 2861 3079 2868 3090
rect 2802 3078 2868 3079
rect 3202 3079 3209 3090
rect 3261 3120 3268 3131
rect 3602 3131 3668 3132
rect 3602 3120 3609 3131
rect 3261 3090 3609 3120
rect 3261 3079 3268 3090
rect 3202 3078 3268 3079
rect 3602 3079 3609 3090
rect 3661 3120 3668 3131
rect 4002 3131 4068 3132
rect 4002 3120 4009 3131
rect 3661 3090 4009 3120
rect 3661 3079 3668 3090
rect 3602 3078 3668 3079
rect 4002 3079 4009 3090
rect 4061 3120 4068 3131
rect 4402 3131 4468 3132
rect 4402 3120 4409 3131
rect 4061 3090 4409 3120
rect 4061 3079 4068 3090
rect 4002 3078 4068 3079
rect 4402 3079 4409 3090
rect 4461 3120 4468 3131
rect 4802 3131 4868 3132
rect 4802 3120 4809 3131
rect 4461 3090 4809 3120
rect 4461 3079 4468 3090
rect 4402 3078 4468 3079
rect 4802 3079 4809 3090
rect 4861 3120 4868 3131
rect 5202 3131 5268 3132
rect 5202 3120 5209 3131
rect 4861 3090 5209 3120
rect 4861 3079 4868 3090
rect 4802 3078 4868 3079
rect 5202 3079 5209 3090
rect 5261 3120 5268 3131
rect 5602 3131 5668 3132
rect 5602 3120 5609 3131
rect 5261 3090 5609 3120
rect 5261 3079 5268 3090
rect 5202 3078 5268 3079
rect 5602 3079 5609 3090
rect 5661 3120 5668 3131
rect 6002 3131 6068 3132
rect 6002 3120 6009 3131
rect 5661 3090 6009 3120
rect 5661 3079 5668 3090
rect 5602 3078 5668 3079
rect 6002 3079 6009 3090
rect 6061 3120 6068 3131
rect 6402 3131 6468 3132
rect 6402 3120 6409 3131
rect 6061 3090 6409 3120
rect 6061 3079 6068 3090
rect 6002 3078 6068 3079
rect 6402 3079 6409 3090
rect 6461 3120 6468 3131
rect 6802 3131 6868 3132
rect 6802 3120 6809 3131
rect 6461 3090 6809 3120
rect 6461 3079 6468 3090
rect 6402 3078 6468 3079
rect 6802 3079 6809 3090
rect 6861 3120 6868 3131
rect 7202 3131 7268 3132
rect 7202 3120 7209 3131
rect 6861 3090 7209 3120
rect 6861 3079 6868 3090
rect 6802 3078 6868 3079
rect 7202 3079 7209 3090
rect 7261 3120 7268 3131
rect 7602 3131 7668 3132
rect 7602 3120 7609 3131
rect 7261 3090 7609 3120
rect 7261 3079 7268 3090
rect 7202 3078 7268 3079
rect 7602 3079 7609 3090
rect 7661 3120 7668 3131
rect 8002 3131 8068 3132
rect 8002 3120 8009 3131
rect 7661 3090 8009 3120
rect 7661 3079 7668 3090
rect 7602 3078 7668 3079
rect 8002 3079 8009 3090
rect 8061 3120 8068 3131
rect 8402 3131 8468 3132
rect 8402 3120 8409 3131
rect 8061 3090 8409 3120
rect 8061 3079 8068 3090
rect 8002 3078 8068 3079
rect 8402 3079 8409 3090
rect 8461 3120 8468 3131
rect 8802 3131 8868 3132
rect 8802 3120 8809 3131
rect 8461 3090 8809 3120
rect 8461 3079 8468 3090
rect 8402 3078 8468 3079
rect 8802 3079 8809 3090
rect 8861 3120 8868 3131
rect 9202 3131 9268 3132
rect 9202 3120 9209 3131
rect 8861 3090 9209 3120
rect 8861 3079 8868 3090
rect 8802 3078 8868 3079
rect 9202 3079 9209 3090
rect 9261 3120 9268 3131
rect 9602 3131 9668 3132
rect 9602 3120 9609 3131
rect 9261 3090 9609 3120
rect 9261 3079 9268 3090
rect 9202 3078 9268 3079
rect 9602 3079 9609 3090
rect 9661 3120 9668 3131
rect 10002 3131 10068 3132
rect 10002 3120 10009 3131
rect 9661 3090 10009 3120
rect 9661 3079 9668 3090
rect 9602 3078 9668 3079
rect 10002 3079 10009 3090
rect 10061 3120 10068 3131
rect 10402 3131 10468 3132
rect 10402 3120 10409 3131
rect 10061 3090 10409 3120
rect 10061 3079 10068 3090
rect 10002 3078 10068 3079
rect 10402 3079 10409 3090
rect 10461 3120 10468 3131
rect 10802 3131 10868 3132
rect 10802 3120 10809 3131
rect 10461 3090 10809 3120
rect 10461 3079 10468 3090
rect 10402 3078 10468 3079
rect 10802 3079 10809 3090
rect 10861 3120 10868 3131
rect 11202 3131 11268 3132
rect 11202 3120 11209 3131
rect 10861 3090 11209 3120
rect 10861 3079 10868 3090
rect 10802 3078 10868 3079
rect 11202 3079 11209 3090
rect 11261 3120 11268 3131
rect 11602 3131 11668 3132
rect 11602 3120 11609 3131
rect 11261 3090 11609 3120
rect 11261 3079 11268 3090
rect 11202 3078 11268 3079
rect 11602 3079 11609 3090
rect 11661 3120 11668 3131
rect 12002 3131 12068 3132
rect 12002 3120 12009 3131
rect 11661 3090 12009 3120
rect 11661 3079 11668 3090
rect 11602 3078 11668 3079
rect 12002 3079 12009 3090
rect 12061 3120 12068 3131
rect 12402 3131 12468 3132
rect 12402 3120 12409 3131
rect 12061 3090 12409 3120
rect 12061 3079 12068 3090
rect 12002 3078 12068 3079
rect 12402 3079 12409 3090
rect 12461 3120 12468 3131
rect 12802 3131 12868 3132
rect 12802 3120 12809 3131
rect 12461 3090 12809 3120
rect 12461 3079 12468 3090
rect 12402 3078 12468 3079
rect 12802 3079 12809 3090
rect 12861 3120 12868 3131
rect 12900 3131 12966 3132
rect 12900 3120 12907 3131
rect 12861 3090 12907 3120
rect 12861 3079 12868 3090
rect 12802 3078 12868 3079
rect 12900 3079 12907 3090
rect 12959 3079 12966 3131
rect 12900 3078 12966 3079
rect 202 3061 268 3062
rect 202 3050 209 3061
rect 0 3020 209 3050
rect 202 3009 209 3020
rect 261 3050 268 3061
rect 602 3061 668 3062
rect 602 3050 609 3061
rect 261 3020 609 3050
rect 261 3009 268 3020
rect 202 3008 268 3009
rect 602 3009 609 3020
rect 661 3050 668 3061
rect 1002 3061 1068 3062
rect 1002 3050 1009 3061
rect 661 3020 1009 3050
rect 661 3009 668 3020
rect 602 3008 668 3009
rect 1002 3009 1009 3020
rect 1061 3050 1068 3061
rect 1402 3061 1468 3062
rect 1402 3050 1409 3061
rect 1061 3020 1409 3050
rect 1061 3009 1068 3020
rect 1002 3008 1068 3009
rect 1402 3009 1409 3020
rect 1461 3050 1468 3061
rect 1802 3061 1868 3062
rect 1802 3050 1809 3061
rect 1461 3020 1809 3050
rect 1461 3009 1468 3020
rect 1402 3008 1468 3009
rect 1802 3009 1809 3020
rect 1861 3050 1868 3061
rect 2202 3061 2268 3062
rect 2202 3050 2209 3061
rect 1861 3020 2209 3050
rect 1861 3009 1868 3020
rect 1802 3008 1868 3009
rect 2202 3009 2209 3020
rect 2261 3050 2268 3061
rect 2602 3061 2668 3062
rect 2602 3050 2609 3061
rect 2261 3020 2609 3050
rect 2261 3009 2268 3020
rect 2202 3008 2268 3009
rect 2602 3009 2609 3020
rect 2661 3050 2668 3061
rect 3002 3061 3068 3062
rect 3002 3050 3009 3061
rect 2661 3020 3009 3050
rect 2661 3009 2668 3020
rect 2602 3008 2668 3009
rect 3002 3009 3009 3020
rect 3061 3050 3068 3061
rect 3402 3061 3468 3062
rect 3402 3050 3409 3061
rect 3061 3020 3409 3050
rect 3061 3009 3068 3020
rect 3002 3008 3068 3009
rect 3402 3009 3409 3020
rect 3461 3050 3468 3061
rect 3802 3061 3868 3062
rect 3802 3050 3809 3061
rect 3461 3020 3809 3050
rect 3461 3009 3468 3020
rect 3402 3008 3468 3009
rect 3802 3009 3809 3020
rect 3861 3050 3868 3061
rect 4202 3061 4268 3062
rect 4202 3050 4209 3061
rect 3861 3020 4209 3050
rect 3861 3009 3868 3020
rect 3802 3008 3868 3009
rect 4202 3009 4209 3020
rect 4261 3050 4268 3061
rect 4602 3061 4668 3062
rect 4602 3050 4609 3061
rect 4261 3020 4609 3050
rect 4261 3009 4268 3020
rect 4202 3008 4268 3009
rect 4602 3009 4609 3020
rect 4661 3050 4668 3061
rect 5002 3061 5068 3062
rect 5002 3050 5009 3061
rect 4661 3020 5009 3050
rect 4661 3009 4668 3020
rect 4602 3008 4668 3009
rect 5002 3009 5009 3020
rect 5061 3050 5068 3061
rect 5402 3061 5468 3062
rect 5402 3050 5409 3061
rect 5061 3020 5409 3050
rect 5061 3009 5068 3020
rect 5002 3008 5068 3009
rect 5402 3009 5409 3020
rect 5461 3050 5468 3061
rect 5802 3061 5868 3062
rect 5802 3050 5809 3061
rect 5461 3020 5809 3050
rect 5461 3009 5468 3020
rect 5402 3008 5468 3009
rect 5802 3009 5809 3020
rect 5861 3050 5868 3061
rect 6202 3061 6268 3062
rect 6202 3050 6209 3061
rect 5861 3020 6209 3050
rect 5861 3009 5868 3020
rect 5802 3008 5868 3009
rect 6202 3009 6209 3020
rect 6261 3050 6268 3061
rect 6602 3061 6668 3062
rect 6602 3050 6609 3061
rect 6261 3020 6609 3050
rect 6261 3009 6268 3020
rect 6202 3008 6268 3009
rect 6602 3009 6609 3020
rect 6661 3050 6668 3061
rect 7002 3061 7068 3062
rect 7002 3050 7009 3061
rect 6661 3020 7009 3050
rect 6661 3009 6668 3020
rect 6602 3008 6668 3009
rect 7002 3009 7009 3020
rect 7061 3050 7068 3061
rect 7402 3061 7468 3062
rect 7402 3050 7409 3061
rect 7061 3020 7409 3050
rect 7061 3009 7068 3020
rect 7002 3008 7068 3009
rect 7402 3009 7409 3020
rect 7461 3050 7468 3061
rect 7802 3061 7868 3062
rect 7802 3050 7809 3061
rect 7461 3020 7809 3050
rect 7461 3009 7468 3020
rect 7402 3008 7468 3009
rect 7802 3009 7809 3020
rect 7861 3050 7868 3061
rect 8202 3061 8268 3062
rect 8202 3050 8209 3061
rect 7861 3020 8209 3050
rect 7861 3009 7868 3020
rect 7802 3008 7868 3009
rect 8202 3009 8209 3020
rect 8261 3050 8268 3061
rect 8602 3061 8668 3062
rect 8602 3050 8609 3061
rect 8261 3020 8609 3050
rect 8261 3009 8268 3020
rect 8202 3008 8268 3009
rect 8602 3009 8609 3020
rect 8661 3050 8668 3061
rect 9002 3061 9068 3062
rect 9002 3050 9009 3061
rect 8661 3020 9009 3050
rect 8661 3009 8668 3020
rect 8602 3008 8668 3009
rect 9002 3009 9009 3020
rect 9061 3050 9068 3061
rect 9402 3061 9468 3062
rect 9402 3050 9409 3061
rect 9061 3020 9409 3050
rect 9061 3009 9068 3020
rect 9002 3008 9068 3009
rect 9402 3009 9409 3020
rect 9461 3050 9468 3061
rect 9802 3061 9868 3062
rect 9802 3050 9809 3061
rect 9461 3020 9809 3050
rect 9461 3009 9468 3020
rect 9402 3008 9468 3009
rect 9802 3009 9809 3020
rect 9861 3050 9868 3061
rect 10202 3061 10268 3062
rect 10202 3050 10209 3061
rect 9861 3020 10209 3050
rect 9861 3009 9868 3020
rect 9802 3008 9868 3009
rect 10202 3009 10209 3020
rect 10261 3050 10268 3061
rect 10602 3061 10668 3062
rect 10602 3050 10609 3061
rect 10261 3020 10609 3050
rect 10261 3009 10268 3020
rect 10202 3008 10268 3009
rect 10602 3009 10609 3020
rect 10661 3050 10668 3061
rect 11002 3061 11068 3062
rect 11002 3050 11009 3061
rect 10661 3020 11009 3050
rect 10661 3009 10668 3020
rect 10602 3008 10668 3009
rect 11002 3009 11009 3020
rect 11061 3050 11068 3061
rect 11402 3061 11468 3062
rect 11402 3050 11409 3061
rect 11061 3020 11409 3050
rect 11061 3009 11068 3020
rect 11002 3008 11068 3009
rect 11402 3009 11409 3020
rect 11461 3050 11468 3061
rect 11802 3061 11868 3062
rect 11802 3050 11809 3061
rect 11461 3020 11809 3050
rect 11461 3009 11468 3020
rect 11402 3008 11468 3009
rect 11802 3009 11809 3020
rect 11861 3050 11868 3061
rect 12202 3061 12268 3062
rect 12202 3050 12209 3061
rect 11861 3020 12209 3050
rect 11861 3009 11868 3020
rect 11802 3008 11868 3009
rect 12202 3009 12209 3020
rect 12261 3050 12268 3061
rect 12602 3061 12668 3062
rect 12602 3050 12609 3061
rect 12261 3020 12609 3050
rect 12261 3009 12268 3020
rect 12202 3008 12268 3009
rect 12602 3009 12609 3020
rect 12661 3050 12668 3061
rect 13104 3061 13170 3062
rect 13104 3050 13111 3061
rect 12661 3020 13111 3050
rect 12661 3009 12668 3020
rect 12602 3008 12668 3009
rect 13104 3009 13111 3020
rect 13163 3009 13170 3061
rect 13104 3008 13170 3009
rect 2 2991 68 2992
rect 2 2980 9 2991
rect 0 2950 9 2980
rect 2 2939 9 2950
rect 61 2980 68 2991
rect 402 2991 468 2992
rect 402 2980 409 2991
rect 61 2950 409 2980
rect 61 2939 68 2950
rect 2 2938 68 2939
rect 402 2939 409 2950
rect 461 2980 468 2991
rect 802 2991 868 2992
rect 802 2980 809 2991
rect 461 2950 809 2980
rect 461 2939 468 2950
rect 402 2938 468 2939
rect 802 2939 809 2950
rect 861 2980 868 2991
rect 1202 2991 1268 2992
rect 1202 2980 1209 2991
rect 861 2950 1209 2980
rect 861 2939 868 2950
rect 802 2938 868 2939
rect 1202 2939 1209 2950
rect 1261 2980 1268 2991
rect 1602 2991 1668 2992
rect 1602 2980 1609 2991
rect 1261 2950 1609 2980
rect 1261 2939 1268 2950
rect 1202 2938 1268 2939
rect 1602 2939 1609 2950
rect 1661 2980 1668 2991
rect 2002 2991 2068 2992
rect 2002 2980 2009 2991
rect 1661 2950 2009 2980
rect 1661 2939 1668 2950
rect 1602 2938 1668 2939
rect 2002 2939 2009 2950
rect 2061 2980 2068 2991
rect 2402 2991 2468 2992
rect 2402 2980 2409 2991
rect 2061 2950 2409 2980
rect 2061 2939 2068 2950
rect 2002 2938 2068 2939
rect 2402 2939 2409 2950
rect 2461 2980 2468 2991
rect 2802 2991 2868 2992
rect 2802 2980 2809 2991
rect 2461 2950 2809 2980
rect 2461 2939 2468 2950
rect 2402 2938 2468 2939
rect 2802 2939 2809 2950
rect 2861 2980 2868 2991
rect 3202 2991 3268 2992
rect 3202 2980 3209 2991
rect 2861 2950 3209 2980
rect 2861 2939 2868 2950
rect 2802 2938 2868 2939
rect 3202 2939 3209 2950
rect 3261 2980 3268 2991
rect 3602 2991 3668 2992
rect 3602 2980 3609 2991
rect 3261 2950 3609 2980
rect 3261 2939 3268 2950
rect 3202 2938 3268 2939
rect 3602 2939 3609 2950
rect 3661 2980 3668 2991
rect 4002 2991 4068 2992
rect 4002 2980 4009 2991
rect 3661 2950 4009 2980
rect 3661 2939 3668 2950
rect 3602 2938 3668 2939
rect 4002 2939 4009 2950
rect 4061 2980 4068 2991
rect 4402 2991 4468 2992
rect 4402 2980 4409 2991
rect 4061 2950 4409 2980
rect 4061 2939 4068 2950
rect 4002 2938 4068 2939
rect 4402 2939 4409 2950
rect 4461 2980 4468 2991
rect 4802 2991 4868 2992
rect 4802 2980 4809 2991
rect 4461 2950 4809 2980
rect 4461 2939 4468 2950
rect 4402 2938 4468 2939
rect 4802 2939 4809 2950
rect 4861 2980 4868 2991
rect 5202 2991 5268 2992
rect 5202 2980 5209 2991
rect 4861 2950 5209 2980
rect 4861 2939 4868 2950
rect 4802 2938 4868 2939
rect 5202 2939 5209 2950
rect 5261 2980 5268 2991
rect 5602 2991 5668 2992
rect 5602 2980 5609 2991
rect 5261 2950 5609 2980
rect 5261 2939 5268 2950
rect 5202 2938 5268 2939
rect 5602 2939 5609 2950
rect 5661 2980 5668 2991
rect 6002 2991 6068 2992
rect 6002 2980 6009 2991
rect 5661 2950 6009 2980
rect 5661 2939 5668 2950
rect 5602 2938 5668 2939
rect 6002 2939 6009 2950
rect 6061 2980 6068 2991
rect 6402 2991 6468 2992
rect 6402 2980 6409 2991
rect 6061 2950 6409 2980
rect 6061 2939 6068 2950
rect 6002 2938 6068 2939
rect 6402 2939 6409 2950
rect 6461 2980 6468 2991
rect 6802 2991 6868 2992
rect 6802 2980 6809 2991
rect 6461 2950 6809 2980
rect 6461 2939 6468 2950
rect 6402 2938 6468 2939
rect 6802 2939 6809 2950
rect 6861 2980 6868 2991
rect 7202 2991 7268 2992
rect 7202 2980 7209 2991
rect 6861 2950 7209 2980
rect 6861 2939 6868 2950
rect 6802 2938 6868 2939
rect 7202 2939 7209 2950
rect 7261 2980 7268 2991
rect 7602 2991 7668 2992
rect 7602 2980 7609 2991
rect 7261 2950 7609 2980
rect 7261 2939 7268 2950
rect 7202 2938 7268 2939
rect 7602 2939 7609 2950
rect 7661 2980 7668 2991
rect 8002 2991 8068 2992
rect 8002 2980 8009 2991
rect 7661 2950 8009 2980
rect 7661 2939 7668 2950
rect 7602 2938 7668 2939
rect 8002 2939 8009 2950
rect 8061 2980 8068 2991
rect 8402 2991 8468 2992
rect 8402 2980 8409 2991
rect 8061 2950 8409 2980
rect 8061 2939 8068 2950
rect 8002 2938 8068 2939
rect 8402 2939 8409 2950
rect 8461 2980 8468 2991
rect 8802 2991 8868 2992
rect 8802 2980 8809 2991
rect 8461 2950 8809 2980
rect 8461 2939 8468 2950
rect 8402 2938 8468 2939
rect 8802 2939 8809 2950
rect 8861 2980 8868 2991
rect 9202 2991 9268 2992
rect 9202 2980 9209 2991
rect 8861 2950 9209 2980
rect 8861 2939 8868 2950
rect 8802 2938 8868 2939
rect 9202 2939 9209 2950
rect 9261 2980 9268 2991
rect 9602 2991 9668 2992
rect 9602 2980 9609 2991
rect 9261 2950 9609 2980
rect 9261 2939 9268 2950
rect 9202 2938 9268 2939
rect 9602 2939 9609 2950
rect 9661 2980 9668 2991
rect 10002 2991 10068 2992
rect 10002 2980 10009 2991
rect 9661 2950 10009 2980
rect 9661 2939 9668 2950
rect 9602 2938 9668 2939
rect 10002 2939 10009 2950
rect 10061 2980 10068 2991
rect 10402 2991 10468 2992
rect 10402 2980 10409 2991
rect 10061 2950 10409 2980
rect 10061 2939 10068 2950
rect 10002 2938 10068 2939
rect 10402 2939 10409 2950
rect 10461 2980 10468 2991
rect 10802 2991 10868 2992
rect 10802 2980 10809 2991
rect 10461 2950 10809 2980
rect 10461 2939 10468 2950
rect 10402 2938 10468 2939
rect 10802 2939 10809 2950
rect 10861 2980 10868 2991
rect 11202 2991 11268 2992
rect 11202 2980 11209 2991
rect 10861 2950 11209 2980
rect 10861 2939 10868 2950
rect 10802 2938 10868 2939
rect 11202 2939 11209 2950
rect 11261 2980 11268 2991
rect 11602 2991 11668 2992
rect 11602 2980 11609 2991
rect 11261 2950 11609 2980
rect 11261 2939 11268 2950
rect 11202 2938 11268 2939
rect 11602 2939 11609 2950
rect 11661 2980 11668 2991
rect 12002 2991 12068 2992
rect 12002 2980 12009 2991
rect 11661 2950 12009 2980
rect 11661 2939 11668 2950
rect 11602 2938 11668 2939
rect 12002 2939 12009 2950
rect 12061 2980 12068 2991
rect 12402 2991 12468 2992
rect 12402 2980 12409 2991
rect 12061 2950 12409 2980
rect 12061 2939 12068 2950
rect 12002 2938 12068 2939
rect 12402 2939 12409 2950
rect 12461 2980 12468 2991
rect 12802 2991 12868 2992
rect 12802 2980 12809 2991
rect 12461 2950 12809 2980
rect 12461 2939 12468 2950
rect 12402 2938 12468 2939
rect 12802 2939 12809 2950
rect 12861 2980 12868 2991
rect 12900 2991 12966 2992
rect 12900 2980 12907 2991
rect 12861 2950 12907 2980
rect 12861 2939 12868 2950
rect 12802 2938 12868 2939
rect 12900 2939 12907 2950
rect 12959 2939 12966 2991
rect 12900 2938 12966 2939
rect 202 2921 268 2922
rect 202 2910 209 2921
rect 0 2880 209 2910
rect 202 2869 209 2880
rect 261 2910 268 2921
rect 602 2921 668 2922
rect 602 2910 609 2921
rect 261 2880 609 2910
rect 261 2869 268 2880
rect 202 2868 268 2869
rect 602 2869 609 2880
rect 661 2910 668 2921
rect 1002 2921 1068 2922
rect 1002 2910 1009 2921
rect 661 2880 1009 2910
rect 661 2869 668 2880
rect 602 2868 668 2869
rect 1002 2869 1009 2880
rect 1061 2910 1068 2921
rect 1402 2921 1468 2922
rect 1402 2910 1409 2921
rect 1061 2880 1409 2910
rect 1061 2869 1068 2880
rect 1002 2868 1068 2869
rect 1402 2869 1409 2880
rect 1461 2910 1468 2921
rect 1802 2921 1868 2922
rect 1802 2910 1809 2921
rect 1461 2880 1809 2910
rect 1461 2869 1468 2880
rect 1402 2868 1468 2869
rect 1802 2869 1809 2880
rect 1861 2910 1868 2921
rect 2202 2921 2268 2922
rect 2202 2910 2209 2921
rect 1861 2880 2209 2910
rect 1861 2869 1868 2880
rect 1802 2868 1868 2869
rect 2202 2869 2209 2880
rect 2261 2910 2268 2921
rect 2602 2921 2668 2922
rect 2602 2910 2609 2921
rect 2261 2880 2609 2910
rect 2261 2869 2268 2880
rect 2202 2868 2268 2869
rect 2602 2869 2609 2880
rect 2661 2910 2668 2921
rect 3002 2921 3068 2922
rect 3002 2910 3009 2921
rect 2661 2880 3009 2910
rect 2661 2869 2668 2880
rect 2602 2868 2668 2869
rect 3002 2869 3009 2880
rect 3061 2910 3068 2921
rect 3402 2921 3468 2922
rect 3402 2910 3409 2921
rect 3061 2880 3409 2910
rect 3061 2869 3068 2880
rect 3002 2868 3068 2869
rect 3402 2869 3409 2880
rect 3461 2910 3468 2921
rect 3802 2921 3868 2922
rect 3802 2910 3809 2921
rect 3461 2880 3809 2910
rect 3461 2869 3468 2880
rect 3402 2868 3468 2869
rect 3802 2869 3809 2880
rect 3861 2910 3868 2921
rect 4202 2921 4268 2922
rect 4202 2910 4209 2921
rect 3861 2880 4209 2910
rect 3861 2869 3868 2880
rect 3802 2868 3868 2869
rect 4202 2869 4209 2880
rect 4261 2910 4268 2921
rect 4602 2921 4668 2922
rect 4602 2910 4609 2921
rect 4261 2880 4609 2910
rect 4261 2869 4268 2880
rect 4202 2868 4268 2869
rect 4602 2869 4609 2880
rect 4661 2910 4668 2921
rect 5002 2921 5068 2922
rect 5002 2910 5009 2921
rect 4661 2880 5009 2910
rect 4661 2869 4668 2880
rect 4602 2868 4668 2869
rect 5002 2869 5009 2880
rect 5061 2910 5068 2921
rect 5402 2921 5468 2922
rect 5402 2910 5409 2921
rect 5061 2880 5409 2910
rect 5061 2869 5068 2880
rect 5002 2868 5068 2869
rect 5402 2869 5409 2880
rect 5461 2910 5468 2921
rect 5802 2921 5868 2922
rect 5802 2910 5809 2921
rect 5461 2880 5809 2910
rect 5461 2869 5468 2880
rect 5402 2868 5468 2869
rect 5802 2869 5809 2880
rect 5861 2910 5868 2921
rect 6202 2921 6268 2922
rect 6202 2910 6209 2921
rect 5861 2880 6209 2910
rect 5861 2869 5868 2880
rect 5802 2868 5868 2869
rect 6202 2869 6209 2880
rect 6261 2910 6268 2921
rect 6602 2921 6668 2922
rect 6602 2910 6609 2921
rect 6261 2880 6609 2910
rect 6261 2869 6268 2880
rect 6202 2868 6268 2869
rect 6602 2869 6609 2880
rect 6661 2910 6668 2921
rect 7002 2921 7068 2922
rect 7002 2910 7009 2921
rect 6661 2880 7009 2910
rect 6661 2869 6668 2880
rect 6602 2868 6668 2869
rect 7002 2869 7009 2880
rect 7061 2910 7068 2921
rect 7402 2921 7468 2922
rect 7402 2910 7409 2921
rect 7061 2880 7409 2910
rect 7061 2869 7068 2880
rect 7002 2868 7068 2869
rect 7402 2869 7409 2880
rect 7461 2910 7468 2921
rect 7802 2921 7868 2922
rect 7802 2910 7809 2921
rect 7461 2880 7809 2910
rect 7461 2869 7468 2880
rect 7402 2868 7468 2869
rect 7802 2869 7809 2880
rect 7861 2910 7868 2921
rect 8202 2921 8268 2922
rect 8202 2910 8209 2921
rect 7861 2880 8209 2910
rect 7861 2869 7868 2880
rect 7802 2868 7868 2869
rect 8202 2869 8209 2880
rect 8261 2910 8268 2921
rect 8602 2921 8668 2922
rect 8602 2910 8609 2921
rect 8261 2880 8609 2910
rect 8261 2869 8268 2880
rect 8202 2868 8268 2869
rect 8602 2869 8609 2880
rect 8661 2910 8668 2921
rect 9002 2921 9068 2922
rect 9002 2910 9009 2921
rect 8661 2880 9009 2910
rect 8661 2869 8668 2880
rect 8602 2868 8668 2869
rect 9002 2869 9009 2880
rect 9061 2910 9068 2921
rect 9402 2921 9468 2922
rect 9402 2910 9409 2921
rect 9061 2880 9409 2910
rect 9061 2869 9068 2880
rect 9002 2868 9068 2869
rect 9402 2869 9409 2880
rect 9461 2910 9468 2921
rect 9802 2921 9868 2922
rect 9802 2910 9809 2921
rect 9461 2880 9809 2910
rect 9461 2869 9468 2880
rect 9402 2868 9468 2869
rect 9802 2869 9809 2880
rect 9861 2910 9868 2921
rect 10202 2921 10268 2922
rect 10202 2910 10209 2921
rect 9861 2880 10209 2910
rect 9861 2869 9868 2880
rect 9802 2868 9868 2869
rect 10202 2869 10209 2880
rect 10261 2910 10268 2921
rect 10602 2921 10668 2922
rect 10602 2910 10609 2921
rect 10261 2880 10609 2910
rect 10261 2869 10268 2880
rect 10202 2868 10268 2869
rect 10602 2869 10609 2880
rect 10661 2910 10668 2921
rect 11002 2921 11068 2922
rect 11002 2910 11009 2921
rect 10661 2880 11009 2910
rect 10661 2869 10668 2880
rect 10602 2868 10668 2869
rect 11002 2869 11009 2880
rect 11061 2910 11068 2921
rect 11402 2921 11468 2922
rect 11402 2910 11409 2921
rect 11061 2880 11409 2910
rect 11061 2869 11068 2880
rect 11002 2868 11068 2869
rect 11402 2869 11409 2880
rect 11461 2910 11468 2921
rect 11802 2921 11868 2922
rect 11802 2910 11809 2921
rect 11461 2880 11809 2910
rect 11461 2869 11468 2880
rect 11402 2868 11468 2869
rect 11802 2869 11809 2880
rect 11861 2910 11868 2921
rect 12202 2921 12268 2922
rect 12202 2910 12209 2921
rect 11861 2880 12209 2910
rect 11861 2869 11868 2880
rect 11802 2868 11868 2869
rect 12202 2869 12209 2880
rect 12261 2910 12268 2921
rect 12602 2921 12668 2922
rect 12602 2910 12609 2921
rect 12261 2880 12609 2910
rect 12261 2869 12268 2880
rect 12202 2868 12268 2869
rect 12602 2869 12609 2880
rect 12661 2910 12668 2921
rect 13104 2921 13170 2922
rect 13104 2910 13111 2921
rect 12661 2880 13111 2910
rect 12661 2869 12668 2880
rect 12602 2868 12668 2869
rect 13104 2869 13111 2880
rect 13163 2869 13170 2921
rect 13104 2868 13170 2869
rect 2 2851 68 2852
rect 2 2840 9 2851
rect 0 2810 9 2840
rect 2 2799 9 2810
rect 61 2840 68 2851
rect 402 2851 468 2852
rect 402 2840 409 2851
rect 61 2810 409 2840
rect 61 2799 68 2810
rect 2 2798 68 2799
rect 402 2799 409 2810
rect 461 2840 468 2851
rect 802 2851 868 2852
rect 802 2840 809 2851
rect 461 2810 809 2840
rect 461 2799 468 2810
rect 402 2798 468 2799
rect 802 2799 809 2810
rect 861 2840 868 2851
rect 1202 2851 1268 2852
rect 1202 2840 1209 2851
rect 861 2810 1209 2840
rect 861 2799 868 2810
rect 802 2798 868 2799
rect 1202 2799 1209 2810
rect 1261 2840 1268 2851
rect 1602 2851 1668 2852
rect 1602 2840 1609 2851
rect 1261 2810 1609 2840
rect 1261 2799 1268 2810
rect 1202 2798 1268 2799
rect 1602 2799 1609 2810
rect 1661 2840 1668 2851
rect 2002 2851 2068 2852
rect 2002 2840 2009 2851
rect 1661 2810 2009 2840
rect 1661 2799 1668 2810
rect 1602 2798 1668 2799
rect 2002 2799 2009 2810
rect 2061 2840 2068 2851
rect 2402 2851 2468 2852
rect 2402 2840 2409 2851
rect 2061 2810 2409 2840
rect 2061 2799 2068 2810
rect 2002 2798 2068 2799
rect 2402 2799 2409 2810
rect 2461 2840 2468 2851
rect 2802 2851 2868 2852
rect 2802 2840 2809 2851
rect 2461 2810 2809 2840
rect 2461 2799 2468 2810
rect 2402 2798 2468 2799
rect 2802 2799 2809 2810
rect 2861 2840 2868 2851
rect 3202 2851 3268 2852
rect 3202 2840 3209 2851
rect 2861 2810 3209 2840
rect 2861 2799 2868 2810
rect 2802 2798 2868 2799
rect 3202 2799 3209 2810
rect 3261 2840 3268 2851
rect 3602 2851 3668 2852
rect 3602 2840 3609 2851
rect 3261 2810 3609 2840
rect 3261 2799 3268 2810
rect 3202 2798 3268 2799
rect 3602 2799 3609 2810
rect 3661 2840 3668 2851
rect 4002 2851 4068 2852
rect 4002 2840 4009 2851
rect 3661 2810 4009 2840
rect 3661 2799 3668 2810
rect 3602 2798 3668 2799
rect 4002 2799 4009 2810
rect 4061 2840 4068 2851
rect 4402 2851 4468 2852
rect 4402 2840 4409 2851
rect 4061 2810 4409 2840
rect 4061 2799 4068 2810
rect 4002 2798 4068 2799
rect 4402 2799 4409 2810
rect 4461 2840 4468 2851
rect 4802 2851 4868 2852
rect 4802 2840 4809 2851
rect 4461 2810 4809 2840
rect 4461 2799 4468 2810
rect 4402 2798 4468 2799
rect 4802 2799 4809 2810
rect 4861 2840 4868 2851
rect 5202 2851 5268 2852
rect 5202 2840 5209 2851
rect 4861 2810 5209 2840
rect 4861 2799 4868 2810
rect 4802 2798 4868 2799
rect 5202 2799 5209 2810
rect 5261 2840 5268 2851
rect 5602 2851 5668 2852
rect 5602 2840 5609 2851
rect 5261 2810 5609 2840
rect 5261 2799 5268 2810
rect 5202 2798 5268 2799
rect 5602 2799 5609 2810
rect 5661 2840 5668 2851
rect 6002 2851 6068 2852
rect 6002 2840 6009 2851
rect 5661 2810 6009 2840
rect 5661 2799 5668 2810
rect 5602 2798 5668 2799
rect 6002 2799 6009 2810
rect 6061 2840 6068 2851
rect 6402 2851 6468 2852
rect 6402 2840 6409 2851
rect 6061 2810 6409 2840
rect 6061 2799 6068 2810
rect 6002 2798 6068 2799
rect 6402 2799 6409 2810
rect 6461 2840 6468 2851
rect 6802 2851 6868 2852
rect 6802 2840 6809 2851
rect 6461 2810 6809 2840
rect 6461 2799 6468 2810
rect 6402 2798 6468 2799
rect 6802 2799 6809 2810
rect 6861 2840 6868 2851
rect 7202 2851 7268 2852
rect 7202 2840 7209 2851
rect 6861 2810 7209 2840
rect 6861 2799 6868 2810
rect 6802 2798 6868 2799
rect 7202 2799 7209 2810
rect 7261 2840 7268 2851
rect 7602 2851 7668 2852
rect 7602 2840 7609 2851
rect 7261 2810 7609 2840
rect 7261 2799 7268 2810
rect 7202 2798 7268 2799
rect 7602 2799 7609 2810
rect 7661 2840 7668 2851
rect 8002 2851 8068 2852
rect 8002 2840 8009 2851
rect 7661 2810 8009 2840
rect 7661 2799 7668 2810
rect 7602 2798 7668 2799
rect 8002 2799 8009 2810
rect 8061 2840 8068 2851
rect 8402 2851 8468 2852
rect 8402 2840 8409 2851
rect 8061 2810 8409 2840
rect 8061 2799 8068 2810
rect 8002 2798 8068 2799
rect 8402 2799 8409 2810
rect 8461 2840 8468 2851
rect 8802 2851 8868 2852
rect 8802 2840 8809 2851
rect 8461 2810 8809 2840
rect 8461 2799 8468 2810
rect 8402 2798 8468 2799
rect 8802 2799 8809 2810
rect 8861 2840 8868 2851
rect 9202 2851 9268 2852
rect 9202 2840 9209 2851
rect 8861 2810 9209 2840
rect 8861 2799 8868 2810
rect 8802 2798 8868 2799
rect 9202 2799 9209 2810
rect 9261 2840 9268 2851
rect 9602 2851 9668 2852
rect 9602 2840 9609 2851
rect 9261 2810 9609 2840
rect 9261 2799 9268 2810
rect 9202 2798 9268 2799
rect 9602 2799 9609 2810
rect 9661 2840 9668 2851
rect 10002 2851 10068 2852
rect 10002 2840 10009 2851
rect 9661 2810 10009 2840
rect 9661 2799 9668 2810
rect 9602 2798 9668 2799
rect 10002 2799 10009 2810
rect 10061 2840 10068 2851
rect 10402 2851 10468 2852
rect 10402 2840 10409 2851
rect 10061 2810 10409 2840
rect 10061 2799 10068 2810
rect 10002 2798 10068 2799
rect 10402 2799 10409 2810
rect 10461 2840 10468 2851
rect 10802 2851 10868 2852
rect 10802 2840 10809 2851
rect 10461 2810 10809 2840
rect 10461 2799 10468 2810
rect 10402 2798 10468 2799
rect 10802 2799 10809 2810
rect 10861 2840 10868 2851
rect 11202 2851 11268 2852
rect 11202 2840 11209 2851
rect 10861 2810 11209 2840
rect 10861 2799 10868 2810
rect 10802 2798 10868 2799
rect 11202 2799 11209 2810
rect 11261 2840 11268 2851
rect 11602 2851 11668 2852
rect 11602 2840 11609 2851
rect 11261 2810 11609 2840
rect 11261 2799 11268 2810
rect 11202 2798 11268 2799
rect 11602 2799 11609 2810
rect 11661 2840 11668 2851
rect 12002 2851 12068 2852
rect 12002 2840 12009 2851
rect 11661 2810 12009 2840
rect 11661 2799 11668 2810
rect 11602 2798 11668 2799
rect 12002 2799 12009 2810
rect 12061 2840 12068 2851
rect 12402 2851 12468 2852
rect 12402 2840 12409 2851
rect 12061 2810 12409 2840
rect 12061 2799 12068 2810
rect 12002 2798 12068 2799
rect 12402 2799 12409 2810
rect 12461 2840 12468 2851
rect 12802 2851 12868 2852
rect 12802 2840 12809 2851
rect 12461 2810 12809 2840
rect 12461 2799 12468 2810
rect 12402 2798 12468 2799
rect 12802 2799 12809 2810
rect 12861 2840 12868 2851
rect 12900 2851 12966 2852
rect 12900 2840 12907 2851
rect 12861 2810 12907 2840
rect 12861 2799 12868 2810
rect 12802 2798 12868 2799
rect 12900 2799 12907 2810
rect 12959 2799 12966 2851
rect 12900 2798 12966 2799
rect 202 2781 268 2782
rect 202 2770 209 2781
rect 0 2740 209 2770
rect 202 2729 209 2740
rect 261 2770 268 2781
rect 602 2781 668 2782
rect 602 2770 609 2781
rect 261 2740 609 2770
rect 261 2729 268 2740
rect 202 2728 268 2729
rect 602 2729 609 2740
rect 661 2770 668 2781
rect 1002 2781 1068 2782
rect 1002 2770 1009 2781
rect 661 2740 1009 2770
rect 661 2729 668 2740
rect 602 2728 668 2729
rect 1002 2729 1009 2740
rect 1061 2770 1068 2781
rect 1402 2781 1468 2782
rect 1402 2770 1409 2781
rect 1061 2740 1409 2770
rect 1061 2729 1068 2740
rect 1002 2728 1068 2729
rect 1402 2729 1409 2740
rect 1461 2770 1468 2781
rect 1802 2781 1868 2782
rect 1802 2770 1809 2781
rect 1461 2740 1809 2770
rect 1461 2729 1468 2740
rect 1402 2728 1468 2729
rect 1802 2729 1809 2740
rect 1861 2770 1868 2781
rect 2202 2781 2268 2782
rect 2202 2770 2209 2781
rect 1861 2740 2209 2770
rect 1861 2729 1868 2740
rect 1802 2728 1868 2729
rect 2202 2729 2209 2740
rect 2261 2770 2268 2781
rect 2602 2781 2668 2782
rect 2602 2770 2609 2781
rect 2261 2740 2609 2770
rect 2261 2729 2268 2740
rect 2202 2728 2268 2729
rect 2602 2729 2609 2740
rect 2661 2770 2668 2781
rect 3002 2781 3068 2782
rect 3002 2770 3009 2781
rect 2661 2740 3009 2770
rect 2661 2729 2668 2740
rect 2602 2728 2668 2729
rect 3002 2729 3009 2740
rect 3061 2770 3068 2781
rect 3402 2781 3468 2782
rect 3402 2770 3409 2781
rect 3061 2740 3409 2770
rect 3061 2729 3068 2740
rect 3002 2728 3068 2729
rect 3402 2729 3409 2740
rect 3461 2770 3468 2781
rect 3802 2781 3868 2782
rect 3802 2770 3809 2781
rect 3461 2740 3809 2770
rect 3461 2729 3468 2740
rect 3402 2728 3468 2729
rect 3802 2729 3809 2740
rect 3861 2770 3868 2781
rect 4202 2781 4268 2782
rect 4202 2770 4209 2781
rect 3861 2740 4209 2770
rect 3861 2729 3868 2740
rect 3802 2728 3868 2729
rect 4202 2729 4209 2740
rect 4261 2770 4268 2781
rect 4602 2781 4668 2782
rect 4602 2770 4609 2781
rect 4261 2740 4609 2770
rect 4261 2729 4268 2740
rect 4202 2728 4268 2729
rect 4602 2729 4609 2740
rect 4661 2770 4668 2781
rect 5002 2781 5068 2782
rect 5002 2770 5009 2781
rect 4661 2740 5009 2770
rect 4661 2729 4668 2740
rect 4602 2728 4668 2729
rect 5002 2729 5009 2740
rect 5061 2770 5068 2781
rect 5402 2781 5468 2782
rect 5402 2770 5409 2781
rect 5061 2740 5409 2770
rect 5061 2729 5068 2740
rect 5002 2728 5068 2729
rect 5402 2729 5409 2740
rect 5461 2770 5468 2781
rect 5802 2781 5868 2782
rect 5802 2770 5809 2781
rect 5461 2740 5809 2770
rect 5461 2729 5468 2740
rect 5402 2728 5468 2729
rect 5802 2729 5809 2740
rect 5861 2770 5868 2781
rect 6202 2781 6268 2782
rect 6202 2770 6209 2781
rect 5861 2740 6209 2770
rect 5861 2729 5868 2740
rect 5802 2728 5868 2729
rect 6202 2729 6209 2740
rect 6261 2770 6268 2781
rect 6602 2781 6668 2782
rect 6602 2770 6609 2781
rect 6261 2740 6609 2770
rect 6261 2729 6268 2740
rect 6202 2728 6268 2729
rect 6602 2729 6609 2740
rect 6661 2770 6668 2781
rect 7002 2781 7068 2782
rect 7002 2770 7009 2781
rect 6661 2740 7009 2770
rect 6661 2729 6668 2740
rect 6602 2728 6668 2729
rect 7002 2729 7009 2740
rect 7061 2770 7068 2781
rect 7402 2781 7468 2782
rect 7402 2770 7409 2781
rect 7061 2740 7409 2770
rect 7061 2729 7068 2740
rect 7002 2728 7068 2729
rect 7402 2729 7409 2740
rect 7461 2770 7468 2781
rect 7802 2781 7868 2782
rect 7802 2770 7809 2781
rect 7461 2740 7809 2770
rect 7461 2729 7468 2740
rect 7402 2728 7468 2729
rect 7802 2729 7809 2740
rect 7861 2770 7868 2781
rect 8202 2781 8268 2782
rect 8202 2770 8209 2781
rect 7861 2740 8209 2770
rect 7861 2729 7868 2740
rect 7802 2728 7868 2729
rect 8202 2729 8209 2740
rect 8261 2770 8268 2781
rect 8602 2781 8668 2782
rect 8602 2770 8609 2781
rect 8261 2740 8609 2770
rect 8261 2729 8268 2740
rect 8202 2728 8268 2729
rect 8602 2729 8609 2740
rect 8661 2770 8668 2781
rect 9002 2781 9068 2782
rect 9002 2770 9009 2781
rect 8661 2740 9009 2770
rect 8661 2729 8668 2740
rect 8602 2728 8668 2729
rect 9002 2729 9009 2740
rect 9061 2770 9068 2781
rect 9402 2781 9468 2782
rect 9402 2770 9409 2781
rect 9061 2740 9409 2770
rect 9061 2729 9068 2740
rect 9002 2728 9068 2729
rect 9402 2729 9409 2740
rect 9461 2770 9468 2781
rect 9802 2781 9868 2782
rect 9802 2770 9809 2781
rect 9461 2740 9809 2770
rect 9461 2729 9468 2740
rect 9402 2728 9468 2729
rect 9802 2729 9809 2740
rect 9861 2770 9868 2781
rect 10202 2781 10268 2782
rect 10202 2770 10209 2781
rect 9861 2740 10209 2770
rect 9861 2729 9868 2740
rect 9802 2728 9868 2729
rect 10202 2729 10209 2740
rect 10261 2770 10268 2781
rect 10602 2781 10668 2782
rect 10602 2770 10609 2781
rect 10261 2740 10609 2770
rect 10261 2729 10268 2740
rect 10202 2728 10268 2729
rect 10602 2729 10609 2740
rect 10661 2770 10668 2781
rect 11002 2781 11068 2782
rect 11002 2770 11009 2781
rect 10661 2740 11009 2770
rect 10661 2729 10668 2740
rect 10602 2728 10668 2729
rect 11002 2729 11009 2740
rect 11061 2770 11068 2781
rect 11402 2781 11468 2782
rect 11402 2770 11409 2781
rect 11061 2740 11409 2770
rect 11061 2729 11068 2740
rect 11002 2728 11068 2729
rect 11402 2729 11409 2740
rect 11461 2770 11468 2781
rect 11802 2781 11868 2782
rect 11802 2770 11809 2781
rect 11461 2740 11809 2770
rect 11461 2729 11468 2740
rect 11402 2728 11468 2729
rect 11802 2729 11809 2740
rect 11861 2770 11868 2781
rect 12202 2781 12268 2782
rect 12202 2770 12209 2781
rect 11861 2740 12209 2770
rect 11861 2729 11868 2740
rect 11802 2728 11868 2729
rect 12202 2729 12209 2740
rect 12261 2770 12268 2781
rect 12602 2781 12668 2782
rect 12602 2770 12609 2781
rect 12261 2740 12609 2770
rect 12261 2729 12268 2740
rect 12202 2728 12268 2729
rect 12602 2729 12609 2740
rect 12661 2770 12668 2781
rect 13104 2781 13170 2782
rect 13104 2770 13111 2781
rect 12661 2740 13111 2770
rect 12661 2729 12668 2740
rect 12602 2728 12668 2729
rect 13104 2729 13111 2740
rect 13163 2729 13170 2781
rect 13104 2728 13170 2729
rect 2 2711 68 2712
rect 2 2700 9 2711
rect 0 2670 9 2700
rect 2 2659 9 2670
rect 61 2700 68 2711
rect 402 2711 468 2712
rect 402 2700 409 2711
rect 61 2670 409 2700
rect 61 2659 68 2670
rect 2 2658 68 2659
rect 402 2659 409 2670
rect 461 2700 468 2711
rect 802 2711 868 2712
rect 802 2700 809 2711
rect 461 2670 809 2700
rect 461 2659 468 2670
rect 402 2658 468 2659
rect 802 2659 809 2670
rect 861 2700 868 2711
rect 1202 2711 1268 2712
rect 1202 2700 1209 2711
rect 861 2670 1209 2700
rect 861 2659 868 2670
rect 802 2658 868 2659
rect 1202 2659 1209 2670
rect 1261 2700 1268 2711
rect 1602 2711 1668 2712
rect 1602 2700 1609 2711
rect 1261 2670 1609 2700
rect 1261 2659 1268 2670
rect 1202 2658 1268 2659
rect 1602 2659 1609 2670
rect 1661 2700 1668 2711
rect 2002 2711 2068 2712
rect 2002 2700 2009 2711
rect 1661 2670 2009 2700
rect 1661 2659 1668 2670
rect 1602 2658 1668 2659
rect 2002 2659 2009 2670
rect 2061 2700 2068 2711
rect 2402 2711 2468 2712
rect 2402 2700 2409 2711
rect 2061 2670 2409 2700
rect 2061 2659 2068 2670
rect 2002 2658 2068 2659
rect 2402 2659 2409 2670
rect 2461 2700 2468 2711
rect 2802 2711 2868 2712
rect 2802 2700 2809 2711
rect 2461 2670 2809 2700
rect 2461 2659 2468 2670
rect 2402 2658 2468 2659
rect 2802 2659 2809 2670
rect 2861 2700 2868 2711
rect 3202 2711 3268 2712
rect 3202 2700 3209 2711
rect 2861 2670 3209 2700
rect 2861 2659 2868 2670
rect 2802 2658 2868 2659
rect 3202 2659 3209 2670
rect 3261 2700 3268 2711
rect 3602 2711 3668 2712
rect 3602 2700 3609 2711
rect 3261 2670 3609 2700
rect 3261 2659 3268 2670
rect 3202 2658 3268 2659
rect 3602 2659 3609 2670
rect 3661 2700 3668 2711
rect 4002 2711 4068 2712
rect 4002 2700 4009 2711
rect 3661 2670 4009 2700
rect 3661 2659 3668 2670
rect 3602 2658 3668 2659
rect 4002 2659 4009 2670
rect 4061 2700 4068 2711
rect 4402 2711 4468 2712
rect 4402 2700 4409 2711
rect 4061 2670 4409 2700
rect 4061 2659 4068 2670
rect 4002 2658 4068 2659
rect 4402 2659 4409 2670
rect 4461 2700 4468 2711
rect 4802 2711 4868 2712
rect 4802 2700 4809 2711
rect 4461 2670 4809 2700
rect 4461 2659 4468 2670
rect 4402 2658 4468 2659
rect 4802 2659 4809 2670
rect 4861 2700 4868 2711
rect 5202 2711 5268 2712
rect 5202 2700 5209 2711
rect 4861 2670 5209 2700
rect 4861 2659 4868 2670
rect 4802 2658 4868 2659
rect 5202 2659 5209 2670
rect 5261 2700 5268 2711
rect 5602 2711 5668 2712
rect 5602 2700 5609 2711
rect 5261 2670 5609 2700
rect 5261 2659 5268 2670
rect 5202 2658 5268 2659
rect 5602 2659 5609 2670
rect 5661 2700 5668 2711
rect 6002 2711 6068 2712
rect 6002 2700 6009 2711
rect 5661 2670 6009 2700
rect 5661 2659 5668 2670
rect 5602 2658 5668 2659
rect 6002 2659 6009 2670
rect 6061 2700 6068 2711
rect 6402 2711 6468 2712
rect 6402 2700 6409 2711
rect 6061 2670 6409 2700
rect 6061 2659 6068 2670
rect 6002 2658 6068 2659
rect 6402 2659 6409 2670
rect 6461 2700 6468 2711
rect 6802 2711 6868 2712
rect 6802 2700 6809 2711
rect 6461 2670 6809 2700
rect 6461 2659 6468 2670
rect 6402 2658 6468 2659
rect 6802 2659 6809 2670
rect 6861 2700 6868 2711
rect 7202 2711 7268 2712
rect 7202 2700 7209 2711
rect 6861 2670 7209 2700
rect 6861 2659 6868 2670
rect 6802 2658 6868 2659
rect 7202 2659 7209 2670
rect 7261 2700 7268 2711
rect 7602 2711 7668 2712
rect 7602 2700 7609 2711
rect 7261 2670 7609 2700
rect 7261 2659 7268 2670
rect 7202 2658 7268 2659
rect 7602 2659 7609 2670
rect 7661 2700 7668 2711
rect 8002 2711 8068 2712
rect 8002 2700 8009 2711
rect 7661 2670 8009 2700
rect 7661 2659 7668 2670
rect 7602 2658 7668 2659
rect 8002 2659 8009 2670
rect 8061 2700 8068 2711
rect 8402 2711 8468 2712
rect 8402 2700 8409 2711
rect 8061 2670 8409 2700
rect 8061 2659 8068 2670
rect 8002 2658 8068 2659
rect 8402 2659 8409 2670
rect 8461 2700 8468 2711
rect 8802 2711 8868 2712
rect 8802 2700 8809 2711
rect 8461 2670 8809 2700
rect 8461 2659 8468 2670
rect 8402 2658 8468 2659
rect 8802 2659 8809 2670
rect 8861 2700 8868 2711
rect 9202 2711 9268 2712
rect 9202 2700 9209 2711
rect 8861 2670 9209 2700
rect 8861 2659 8868 2670
rect 8802 2658 8868 2659
rect 9202 2659 9209 2670
rect 9261 2700 9268 2711
rect 9602 2711 9668 2712
rect 9602 2700 9609 2711
rect 9261 2670 9609 2700
rect 9261 2659 9268 2670
rect 9202 2658 9268 2659
rect 9602 2659 9609 2670
rect 9661 2700 9668 2711
rect 10002 2711 10068 2712
rect 10002 2700 10009 2711
rect 9661 2670 10009 2700
rect 9661 2659 9668 2670
rect 9602 2658 9668 2659
rect 10002 2659 10009 2670
rect 10061 2700 10068 2711
rect 10402 2711 10468 2712
rect 10402 2700 10409 2711
rect 10061 2670 10409 2700
rect 10061 2659 10068 2670
rect 10002 2658 10068 2659
rect 10402 2659 10409 2670
rect 10461 2700 10468 2711
rect 10802 2711 10868 2712
rect 10802 2700 10809 2711
rect 10461 2670 10809 2700
rect 10461 2659 10468 2670
rect 10402 2658 10468 2659
rect 10802 2659 10809 2670
rect 10861 2700 10868 2711
rect 11202 2711 11268 2712
rect 11202 2700 11209 2711
rect 10861 2670 11209 2700
rect 10861 2659 10868 2670
rect 10802 2658 10868 2659
rect 11202 2659 11209 2670
rect 11261 2700 11268 2711
rect 11602 2711 11668 2712
rect 11602 2700 11609 2711
rect 11261 2670 11609 2700
rect 11261 2659 11268 2670
rect 11202 2658 11268 2659
rect 11602 2659 11609 2670
rect 11661 2700 11668 2711
rect 12002 2711 12068 2712
rect 12002 2700 12009 2711
rect 11661 2670 12009 2700
rect 11661 2659 11668 2670
rect 11602 2658 11668 2659
rect 12002 2659 12009 2670
rect 12061 2700 12068 2711
rect 12402 2711 12468 2712
rect 12402 2700 12409 2711
rect 12061 2670 12409 2700
rect 12061 2659 12068 2670
rect 12002 2658 12068 2659
rect 12402 2659 12409 2670
rect 12461 2700 12468 2711
rect 12802 2711 12868 2712
rect 12802 2700 12809 2711
rect 12461 2670 12809 2700
rect 12461 2659 12468 2670
rect 12402 2658 12468 2659
rect 12802 2659 12809 2670
rect 12861 2700 12868 2711
rect 12900 2711 12966 2712
rect 12900 2700 12907 2711
rect 12861 2670 12907 2700
rect 12861 2659 12868 2670
rect 12802 2658 12868 2659
rect 12900 2659 12907 2670
rect 12959 2659 12966 2711
rect 12900 2658 12966 2659
rect 202 2641 268 2642
rect 202 2630 209 2641
rect 0 2600 209 2630
rect 202 2589 209 2600
rect 261 2630 268 2641
rect 602 2641 668 2642
rect 602 2630 609 2641
rect 261 2600 609 2630
rect 261 2589 268 2600
rect 202 2588 268 2589
rect 602 2589 609 2600
rect 661 2630 668 2641
rect 1002 2641 1068 2642
rect 1002 2630 1009 2641
rect 661 2600 1009 2630
rect 661 2589 668 2600
rect 602 2588 668 2589
rect 1002 2589 1009 2600
rect 1061 2630 1068 2641
rect 1402 2641 1468 2642
rect 1402 2630 1409 2641
rect 1061 2600 1409 2630
rect 1061 2589 1068 2600
rect 1002 2588 1068 2589
rect 1402 2589 1409 2600
rect 1461 2630 1468 2641
rect 1802 2641 1868 2642
rect 1802 2630 1809 2641
rect 1461 2600 1809 2630
rect 1461 2589 1468 2600
rect 1402 2588 1468 2589
rect 1802 2589 1809 2600
rect 1861 2630 1868 2641
rect 2202 2641 2268 2642
rect 2202 2630 2209 2641
rect 1861 2600 2209 2630
rect 1861 2589 1868 2600
rect 1802 2588 1868 2589
rect 2202 2589 2209 2600
rect 2261 2630 2268 2641
rect 2602 2641 2668 2642
rect 2602 2630 2609 2641
rect 2261 2600 2609 2630
rect 2261 2589 2268 2600
rect 2202 2588 2268 2589
rect 2602 2589 2609 2600
rect 2661 2630 2668 2641
rect 3002 2641 3068 2642
rect 3002 2630 3009 2641
rect 2661 2600 3009 2630
rect 2661 2589 2668 2600
rect 2602 2588 2668 2589
rect 3002 2589 3009 2600
rect 3061 2630 3068 2641
rect 3402 2641 3468 2642
rect 3402 2630 3409 2641
rect 3061 2600 3409 2630
rect 3061 2589 3068 2600
rect 3002 2588 3068 2589
rect 3402 2589 3409 2600
rect 3461 2630 3468 2641
rect 3802 2641 3868 2642
rect 3802 2630 3809 2641
rect 3461 2600 3809 2630
rect 3461 2589 3468 2600
rect 3402 2588 3468 2589
rect 3802 2589 3809 2600
rect 3861 2630 3868 2641
rect 4202 2641 4268 2642
rect 4202 2630 4209 2641
rect 3861 2600 4209 2630
rect 3861 2589 3868 2600
rect 3802 2588 3868 2589
rect 4202 2589 4209 2600
rect 4261 2630 4268 2641
rect 4602 2641 4668 2642
rect 4602 2630 4609 2641
rect 4261 2600 4609 2630
rect 4261 2589 4268 2600
rect 4202 2588 4268 2589
rect 4602 2589 4609 2600
rect 4661 2630 4668 2641
rect 5002 2641 5068 2642
rect 5002 2630 5009 2641
rect 4661 2600 5009 2630
rect 4661 2589 4668 2600
rect 4602 2588 4668 2589
rect 5002 2589 5009 2600
rect 5061 2630 5068 2641
rect 5402 2641 5468 2642
rect 5402 2630 5409 2641
rect 5061 2600 5409 2630
rect 5061 2589 5068 2600
rect 5002 2588 5068 2589
rect 5402 2589 5409 2600
rect 5461 2630 5468 2641
rect 5802 2641 5868 2642
rect 5802 2630 5809 2641
rect 5461 2600 5809 2630
rect 5461 2589 5468 2600
rect 5402 2588 5468 2589
rect 5802 2589 5809 2600
rect 5861 2630 5868 2641
rect 6202 2641 6268 2642
rect 6202 2630 6209 2641
rect 5861 2600 6209 2630
rect 5861 2589 5868 2600
rect 5802 2588 5868 2589
rect 6202 2589 6209 2600
rect 6261 2630 6268 2641
rect 6602 2641 6668 2642
rect 6602 2630 6609 2641
rect 6261 2600 6609 2630
rect 6261 2589 6268 2600
rect 6202 2588 6268 2589
rect 6602 2589 6609 2600
rect 6661 2630 6668 2641
rect 7002 2641 7068 2642
rect 7002 2630 7009 2641
rect 6661 2600 7009 2630
rect 6661 2589 6668 2600
rect 6602 2588 6668 2589
rect 7002 2589 7009 2600
rect 7061 2630 7068 2641
rect 7402 2641 7468 2642
rect 7402 2630 7409 2641
rect 7061 2600 7409 2630
rect 7061 2589 7068 2600
rect 7002 2588 7068 2589
rect 7402 2589 7409 2600
rect 7461 2630 7468 2641
rect 7802 2641 7868 2642
rect 7802 2630 7809 2641
rect 7461 2600 7809 2630
rect 7461 2589 7468 2600
rect 7402 2588 7468 2589
rect 7802 2589 7809 2600
rect 7861 2630 7868 2641
rect 8202 2641 8268 2642
rect 8202 2630 8209 2641
rect 7861 2600 8209 2630
rect 7861 2589 7868 2600
rect 7802 2588 7868 2589
rect 8202 2589 8209 2600
rect 8261 2630 8268 2641
rect 8602 2641 8668 2642
rect 8602 2630 8609 2641
rect 8261 2600 8609 2630
rect 8261 2589 8268 2600
rect 8202 2588 8268 2589
rect 8602 2589 8609 2600
rect 8661 2630 8668 2641
rect 9002 2641 9068 2642
rect 9002 2630 9009 2641
rect 8661 2600 9009 2630
rect 8661 2589 8668 2600
rect 8602 2588 8668 2589
rect 9002 2589 9009 2600
rect 9061 2630 9068 2641
rect 9402 2641 9468 2642
rect 9402 2630 9409 2641
rect 9061 2600 9409 2630
rect 9061 2589 9068 2600
rect 9002 2588 9068 2589
rect 9402 2589 9409 2600
rect 9461 2630 9468 2641
rect 9802 2641 9868 2642
rect 9802 2630 9809 2641
rect 9461 2600 9809 2630
rect 9461 2589 9468 2600
rect 9402 2588 9468 2589
rect 9802 2589 9809 2600
rect 9861 2630 9868 2641
rect 10202 2641 10268 2642
rect 10202 2630 10209 2641
rect 9861 2600 10209 2630
rect 9861 2589 9868 2600
rect 9802 2588 9868 2589
rect 10202 2589 10209 2600
rect 10261 2630 10268 2641
rect 10602 2641 10668 2642
rect 10602 2630 10609 2641
rect 10261 2600 10609 2630
rect 10261 2589 10268 2600
rect 10202 2588 10268 2589
rect 10602 2589 10609 2600
rect 10661 2630 10668 2641
rect 11002 2641 11068 2642
rect 11002 2630 11009 2641
rect 10661 2600 11009 2630
rect 10661 2589 10668 2600
rect 10602 2588 10668 2589
rect 11002 2589 11009 2600
rect 11061 2630 11068 2641
rect 11402 2641 11468 2642
rect 11402 2630 11409 2641
rect 11061 2600 11409 2630
rect 11061 2589 11068 2600
rect 11002 2588 11068 2589
rect 11402 2589 11409 2600
rect 11461 2630 11468 2641
rect 11802 2641 11868 2642
rect 11802 2630 11809 2641
rect 11461 2600 11809 2630
rect 11461 2589 11468 2600
rect 11402 2588 11468 2589
rect 11802 2589 11809 2600
rect 11861 2630 11868 2641
rect 12202 2641 12268 2642
rect 12202 2630 12209 2641
rect 11861 2600 12209 2630
rect 11861 2589 11868 2600
rect 11802 2588 11868 2589
rect 12202 2589 12209 2600
rect 12261 2630 12268 2641
rect 12602 2641 12668 2642
rect 12602 2630 12609 2641
rect 12261 2600 12609 2630
rect 12261 2589 12268 2600
rect 12202 2588 12268 2589
rect 12602 2589 12609 2600
rect 12661 2630 12668 2641
rect 13104 2641 13170 2642
rect 13104 2630 13111 2641
rect 12661 2600 13111 2630
rect 12661 2589 12668 2600
rect 12602 2588 12668 2589
rect 13104 2589 13111 2600
rect 13163 2589 13170 2641
rect 13104 2588 13170 2589
rect 2 2571 68 2572
rect 2 2560 9 2571
rect 0 2530 9 2560
rect 2 2519 9 2530
rect 61 2560 68 2571
rect 402 2571 468 2572
rect 402 2560 409 2571
rect 61 2530 409 2560
rect 61 2519 68 2530
rect 2 2518 68 2519
rect 402 2519 409 2530
rect 461 2560 468 2571
rect 802 2571 868 2572
rect 802 2560 809 2571
rect 461 2530 809 2560
rect 461 2519 468 2530
rect 402 2518 468 2519
rect 802 2519 809 2530
rect 861 2560 868 2571
rect 1202 2571 1268 2572
rect 1202 2560 1209 2571
rect 861 2530 1209 2560
rect 861 2519 868 2530
rect 802 2518 868 2519
rect 1202 2519 1209 2530
rect 1261 2560 1268 2571
rect 1602 2571 1668 2572
rect 1602 2560 1609 2571
rect 1261 2530 1609 2560
rect 1261 2519 1268 2530
rect 1202 2518 1268 2519
rect 1602 2519 1609 2530
rect 1661 2560 1668 2571
rect 2002 2571 2068 2572
rect 2002 2560 2009 2571
rect 1661 2530 2009 2560
rect 1661 2519 1668 2530
rect 1602 2518 1668 2519
rect 2002 2519 2009 2530
rect 2061 2560 2068 2571
rect 2402 2571 2468 2572
rect 2402 2560 2409 2571
rect 2061 2530 2409 2560
rect 2061 2519 2068 2530
rect 2002 2518 2068 2519
rect 2402 2519 2409 2530
rect 2461 2560 2468 2571
rect 2802 2571 2868 2572
rect 2802 2560 2809 2571
rect 2461 2530 2809 2560
rect 2461 2519 2468 2530
rect 2402 2518 2468 2519
rect 2802 2519 2809 2530
rect 2861 2560 2868 2571
rect 3202 2571 3268 2572
rect 3202 2560 3209 2571
rect 2861 2530 3209 2560
rect 2861 2519 2868 2530
rect 2802 2518 2868 2519
rect 3202 2519 3209 2530
rect 3261 2560 3268 2571
rect 3602 2571 3668 2572
rect 3602 2560 3609 2571
rect 3261 2530 3609 2560
rect 3261 2519 3268 2530
rect 3202 2518 3268 2519
rect 3602 2519 3609 2530
rect 3661 2560 3668 2571
rect 4002 2571 4068 2572
rect 4002 2560 4009 2571
rect 3661 2530 4009 2560
rect 3661 2519 3668 2530
rect 3602 2518 3668 2519
rect 4002 2519 4009 2530
rect 4061 2560 4068 2571
rect 4402 2571 4468 2572
rect 4402 2560 4409 2571
rect 4061 2530 4409 2560
rect 4061 2519 4068 2530
rect 4002 2518 4068 2519
rect 4402 2519 4409 2530
rect 4461 2560 4468 2571
rect 4802 2571 4868 2572
rect 4802 2560 4809 2571
rect 4461 2530 4809 2560
rect 4461 2519 4468 2530
rect 4402 2518 4468 2519
rect 4802 2519 4809 2530
rect 4861 2560 4868 2571
rect 5202 2571 5268 2572
rect 5202 2560 5209 2571
rect 4861 2530 5209 2560
rect 4861 2519 4868 2530
rect 4802 2518 4868 2519
rect 5202 2519 5209 2530
rect 5261 2560 5268 2571
rect 5602 2571 5668 2572
rect 5602 2560 5609 2571
rect 5261 2530 5609 2560
rect 5261 2519 5268 2530
rect 5202 2518 5268 2519
rect 5602 2519 5609 2530
rect 5661 2560 5668 2571
rect 6002 2571 6068 2572
rect 6002 2560 6009 2571
rect 5661 2530 6009 2560
rect 5661 2519 5668 2530
rect 5602 2518 5668 2519
rect 6002 2519 6009 2530
rect 6061 2560 6068 2571
rect 6402 2571 6468 2572
rect 6402 2560 6409 2571
rect 6061 2530 6409 2560
rect 6061 2519 6068 2530
rect 6002 2518 6068 2519
rect 6402 2519 6409 2530
rect 6461 2560 6468 2571
rect 6802 2571 6868 2572
rect 6802 2560 6809 2571
rect 6461 2530 6809 2560
rect 6461 2519 6468 2530
rect 6402 2518 6468 2519
rect 6802 2519 6809 2530
rect 6861 2560 6868 2571
rect 7202 2571 7268 2572
rect 7202 2560 7209 2571
rect 6861 2530 7209 2560
rect 6861 2519 6868 2530
rect 6802 2518 6868 2519
rect 7202 2519 7209 2530
rect 7261 2560 7268 2571
rect 7602 2571 7668 2572
rect 7602 2560 7609 2571
rect 7261 2530 7609 2560
rect 7261 2519 7268 2530
rect 7202 2518 7268 2519
rect 7602 2519 7609 2530
rect 7661 2560 7668 2571
rect 8002 2571 8068 2572
rect 8002 2560 8009 2571
rect 7661 2530 8009 2560
rect 7661 2519 7668 2530
rect 7602 2518 7668 2519
rect 8002 2519 8009 2530
rect 8061 2560 8068 2571
rect 8402 2571 8468 2572
rect 8402 2560 8409 2571
rect 8061 2530 8409 2560
rect 8061 2519 8068 2530
rect 8002 2518 8068 2519
rect 8402 2519 8409 2530
rect 8461 2560 8468 2571
rect 8802 2571 8868 2572
rect 8802 2560 8809 2571
rect 8461 2530 8809 2560
rect 8461 2519 8468 2530
rect 8402 2518 8468 2519
rect 8802 2519 8809 2530
rect 8861 2560 8868 2571
rect 9202 2571 9268 2572
rect 9202 2560 9209 2571
rect 8861 2530 9209 2560
rect 8861 2519 8868 2530
rect 8802 2518 8868 2519
rect 9202 2519 9209 2530
rect 9261 2560 9268 2571
rect 9602 2571 9668 2572
rect 9602 2560 9609 2571
rect 9261 2530 9609 2560
rect 9261 2519 9268 2530
rect 9202 2518 9268 2519
rect 9602 2519 9609 2530
rect 9661 2560 9668 2571
rect 10002 2571 10068 2572
rect 10002 2560 10009 2571
rect 9661 2530 10009 2560
rect 9661 2519 9668 2530
rect 9602 2518 9668 2519
rect 10002 2519 10009 2530
rect 10061 2560 10068 2571
rect 10402 2571 10468 2572
rect 10402 2560 10409 2571
rect 10061 2530 10409 2560
rect 10061 2519 10068 2530
rect 10002 2518 10068 2519
rect 10402 2519 10409 2530
rect 10461 2560 10468 2571
rect 10802 2571 10868 2572
rect 10802 2560 10809 2571
rect 10461 2530 10809 2560
rect 10461 2519 10468 2530
rect 10402 2518 10468 2519
rect 10802 2519 10809 2530
rect 10861 2560 10868 2571
rect 11202 2571 11268 2572
rect 11202 2560 11209 2571
rect 10861 2530 11209 2560
rect 10861 2519 10868 2530
rect 10802 2518 10868 2519
rect 11202 2519 11209 2530
rect 11261 2560 11268 2571
rect 11602 2571 11668 2572
rect 11602 2560 11609 2571
rect 11261 2530 11609 2560
rect 11261 2519 11268 2530
rect 11202 2518 11268 2519
rect 11602 2519 11609 2530
rect 11661 2560 11668 2571
rect 12002 2571 12068 2572
rect 12002 2560 12009 2571
rect 11661 2530 12009 2560
rect 11661 2519 11668 2530
rect 11602 2518 11668 2519
rect 12002 2519 12009 2530
rect 12061 2560 12068 2571
rect 12402 2571 12468 2572
rect 12402 2560 12409 2571
rect 12061 2530 12409 2560
rect 12061 2519 12068 2530
rect 12002 2518 12068 2519
rect 12402 2519 12409 2530
rect 12461 2560 12468 2571
rect 12802 2571 12868 2572
rect 12802 2560 12809 2571
rect 12461 2530 12809 2560
rect 12461 2519 12468 2530
rect 12402 2518 12468 2519
rect 12802 2519 12809 2530
rect 12861 2560 12868 2571
rect 12900 2571 12966 2572
rect 12900 2560 12907 2571
rect 12861 2530 12907 2560
rect 12861 2519 12868 2530
rect 12802 2518 12868 2519
rect 12900 2519 12907 2530
rect 12959 2519 12966 2571
rect 12900 2518 12966 2519
rect 196 2501 274 2502
rect -4 2485 74 2486
rect -4 2429 7 2485
rect 63 2429 74 2485
rect 196 2445 207 2501
rect 263 2445 274 2501
rect 596 2501 674 2502
rect 196 2444 274 2445
rect 396 2485 474 2486
rect -4 2428 74 2429
rect 396 2429 407 2485
rect 463 2429 474 2485
rect 596 2445 607 2501
rect 663 2445 674 2501
rect 996 2501 1074 2502
rect 596 2444 674 2445
rect 796 2485 874 2486
rect 396 2428 474 2429
rect 796 2429 807 2485
rect 863 2429 874 2485
rect 996 2445 1007 2501
rect 1063 2445 1074 2501
rect 1396 2501 1474 2502
rect 996 2444 1074 2445
rect 1196 2485 1274 2486
rect 796 2428 874 2429
rect 1196 2429 1207 2485
rect 1263 2429 1274 2485
rect 1396 2445 1407 2501
rect 1463 2445 1474 2501
rect 1796 2501 1874 2502
rect 1396 2444 1474 2445
rect 1596 2485 1674 2486
rect 1196 2428 1274 2429
rect 1596 2429 1607 2485
rect 1663 2429 1674 2485
rect 1796 2445 1807 2501
rect 1863 2445 1874 2501
rect 2196 2501 2274 2502
rect 1796 2444 1874 2445
rect 1996 2485 2074 2486
rect 1596 2428 1674 2429
rect 1996 2429 2007 2485
rect 2063 2429 2074 2485
rect 2196 2445 2207 2501
rect 2263 2445 2274 2501
rect 2596 2501 2674 2502
rect 2196 2444 2274 2445
rect 2396 2485 2474 2486
rect 1996 2428 2074 2429
rect 2396 2429 2407 2485
rect 2463 2429 2474 2485
rect 2596 2445 2607 2501
rect 2663 2445 2674 2501
rect 2996 2501 3074 2502
rect 2596 2444 2674 2445
rect 2796 2485 2874 2486
rect 2396 2428 2474 2429
rect 2796 2429 2807 2485
rect 2863 2429 2874 2485
rect 2996 2445 3007 2501
rect 3063 2445 3074 2501
rect 3396 2501 3474 2502
rect 2996 2444 3074 2445
rect 3196 2485 3274 2486
rect 2796 2428 2874 2429
rect 3196 2429 3207 2485
rect 3263 2429 3274 2485
rect 3396 2445 3407 2501
rect 3463 2445 3474 2501
rect 3796 2501 3874 2502
rect 3396 2444 3474 2445
rect 3596 2485 3674 2486
rect 3196 2428 3274 2429
rect 3596 2429 3607 2485
rect 3663 2429 3674 2485
rect 3796 2445 3807 2501
rect 3863 2445 3874 2501
rect 4196 2501 4274 2502
rect 3796 2444 3874 2445
rect 3996 2485 4074 2486
rect 3596 2428 3674 2429
rect 3996 2429 4007 2485
rect 4063 2429 4074 2485
rect 4196 2445 4207 2501
rect 4263 2445 4274 2501
rect 4596 2501 4674 2502
rect 4196 2444 4274 2445
rect 4396 2485 4474 2486
rect 3996 2428 4074 2429
rect 4396 2429 4407 2485
rect 4463 2429 4474 2485
rect 4596 2445 4607 2501
rect 4663 2445 4674 2501
rect 4996 2501 5074 2502
rect 4596 2444 4674 2445
rect 4796 2485 4874 2486
rect 4396 2428 4474 2429
rect 4796 2429 4807 2485
rect 4863 2429 4874 2485
rect 4996 2445 5007 2501
rect 5063 2445 5074 2501
rect 5396 2501 5474 2502
rect 4996 2444 5074 2445
rect 5196 2485 5274 2486
rect 4796 2428 4874 2429
rect 5196 2429 5207 2485
rect 5263 2429 5274 2485
rect 5396 2445 5407 2501
rect 5463 2445 5474 2501
rect 5796 2501 5874 2502
rect 5396 2444 5474 2445
rect 5596 2485 5674 2486
rect 5196 2428 5274 2429
rect 5596 2429 5607 2485
rect 5663 2429 5674 2485
rect 5796 2445 5807 2501
rect 5863 2445 5874 2501
rect 6196 2501 6274 2502
rect 5796 2444 5874 2445
rect 5996 2485 6074 2486
rect 5596 2428 5674 2429
rect 5996 2429 6007 2485
rect 6063 2429 6074 2485
rect 6196 2445 6207 2501
rect 6263 2445 6274 2501
rect 6596 2501 6674 2502
rect 6196 2444 6274 2445
rect 6396 2485 6474 2486
rect 5996 2428 6074 2429
rect 6396 2429 6407 2485
rect 6463 2429 6474 2485
rect 6596 2445 6607 2501
rect 6663 2445 6674 2501
rect 6996 2501 7074 2502
rect 6596 2444 6674 2445
rect 6796 2485 6874 2486
rect 6396 2428 6474 2429
rect 6796 2429 6807 2485
rect 6863 2429 6874 2485
rect 6996 2445 7007 2501
rect 7063 2445 7074 2501
rect 7396 2501 7474 2502
rect 6996 2444 7074 2445
rect 7196 2485 7274 2486
rect 6796 2428 6874 2429
rect 7196 2429 7207 2485
rect 7263 2429 7274 2485
rect 7396 2445 7407 2501
rect 7463 2445 7474 2501
rect 7796 2501 7874 2502
rect 7396 2444 7474 2445
rect 7596 2485 7674 2486
rect 7196 2428 7274 2429
rect 7596 2429 7607 2485
rect 7663 2429 7674 2485
rect 7796 2445 7807 2501
rect 7863 2445 7874 2501
rect 8196 2501 8274 2502
rect 7796 2444 7874 2445
rect 7996 2485 8074 2486
rect 7596 2428 7674 2429
rect 7996 2429 8007 2485
rect 8063 2429 8074 2485
rect 8196 2445 8207 2501
rect 8263 2445 8274 2501
rect 8596 2501 8674 2502
rect 8196 2444 8274 2445
rect 8396 2485 8474 2486
rect 7996 2428 8074 2429
rect 8396 2429 8407 2485
rect 8463 2429 8474 2485
rect 8596 2445 8607 2501
rect 8663 2445 8674 2501
rect 8996 2501 9074 2502
rect 8596 2444 8674 2445
rect 8796 2485 8874 2486
rect 8396 2428 8474 2429
rect 8796 2429 8807 2485
rect 8863 2429 8874 2485
rect 8996 2445 9007 2501
rect 9063 2445 9074 2501
rect 9396 2501 9474 2502
rect 8996 2444 9074 2445
rect 9196 2485 9274 2486
rect 8796 2428 8874 2429
rect 9196 2429 9207 2485
rect 9263 2429 9274 2485
rect 9396 2445 9407 2501
rect 9463 2445 9474 2501
rect 9796 2501 9874 2502
rect 9396 2444 9474 2445
rect 9596 2485 9674 2486
rect 9196 2428 9274 2429
rect 9596 2429 9607 2485
rect 9663 2429 9674 2485
rect 9796 2445 9807 2501
rect 9863 2445 9874 2501
rect 10196 2501 10274 2502
rect 9796 2444 9874 2445
rect 9996 2485 10074 2486
rect 9596 2428 9674 2429
rect 9996 2429 10007 2485
rect 10063 2429 10074 2485
rect 10196 2445 10207 2501
rect 10263 2445 10274 2501
rect 10596 2501 10674 2502
rect 10196 2444 10274 2445
rect 10396 2485 10474 2486
rect 9996 2428 10074 2429
rect 10396 2429 10407 2485
rect 10463 2429 10474 2485
rect 10596 2445 10607 2501
rect 10663 2445 10674 2501
rect 10996 2501 11074 2502
rect 10596 2444 10674 2445
rect 10796 2485 10874 2486
rect 10396 2428 10474 2429
rect 10796 2429 10807 2485
rect 10863 2429 10874 2485
rect 10996 2445 11007 2501
rect 11063 2445 11074 2501
rect 11396 2501 11474 2502
rect 10996 2444 11074 2445
rect 11196 2485 11274 2486
rect 10796 2428 10874 2429
rect 11196 2429 11207 2485
rect 11263 2429 11274 2485
rect 11396 2445 11407 2501
rect 11463 2445 11474 2501
rect 11796 2501 11874 2502
rect 11396 2444 11474 2445
rect 11596 2485 11674 2486
rect 11196 2428 11274 2429
rect 11596 2429 11607 2485
rect 11663 2429 11674 2485
rect 11796 2445 11807 2501
rect 11863 2445 11874 2501
rect 12196 2501 12274 2502
rect 11796 2444 11874 2445
rect 11996 2485 12074 2486
rect 11596 2428 11674 2429
rect 11996 2429 12007 2485
rect 12063 2429 12074 2485
rect 12196 2445 12207 2501
rect 12263 2445 12274 2501
rect 12596 2501 12674 2502
rect 12196 2444 12274 2445
rect 12396 2485 12474 2486
rect 11996 2428 12074 2429
rect 12396 2429 12407 2485
rect 12463 2429 12474 2485
rect 12596 2445 12607 2501
rect 12663 2445 12674 2501
rect 12596 2444 12674 2445
rect 12396 2428 12474 2429
rect 202 2411 268 2412
rect 202 2400 209 2411
rect 0 2370 209 2400
rect 202 2359 209 2370
rect 261 2400 268 2411
rect 602 2411 668 2412
rect 602 2400 609 2411
rect 261 2370 609 2400
rect 261 2359 268 2370
rect 202 2358 268 2359
rect 602 2359 609 2370
rect 661 2400 668 2411
rect 1002 2411 1068 2412
rect 1002 2400 1009 2411
rect 661 2370 1009 2400
rect 661 2359 668 2370
rect 602 2358 668 2359
rect 1002 2359 1009 2370
rect 1061 2400 1068 2411
rect 1402 2411 1468 2412
rect 1402 2400 1409 2411
rect 1061 2370 1409 2400
rect 1061 2359 1068 2370
rect 1002 2358 1068 2359
rect 1402 2359 1409 2370
rect 1461 2400 1468 2411
rect 1802 2411 1868 2412
rect 1802 2400 1809 2411
rect 1461 2370 1809 2400
rect 1461 2359 1468 2370
rect 1402 2358 1468 2359
rect 1802 2359 1809 2370
rect 1861 2400 1868 2411
rect 2202 2411 2268 2412
rect 2202 2400 2209 2411
rect 1861 2370 2209 2400
rect 1861 2359 1868 2370
rect 1802 2358 1868 2359
rect 2202 2359 2209 2370
rect 2261 2400 2268 2411
rect 2602 2411 2668 2412
rect 2602 2400 2609 2411
rect 2261 2370 2609 2400
rect 2261 2359 2268 2370
rect 2202 2358 2268 2359
rect 2602 2359 2609 2370
rect 2661 2400 2668 2411
rect 3002 2411 3068 2412
rect 3002 2400 3009 2411
rect 2661 2370 3009 2400
rect 2661 2359 2668 2370
rect 2602 2358 2668 2359
rect 3002 2359 3009 2370
rect 3061 2400 3068 2411
rect 3402 2411 3468 2412
rect 3402 2400 3409 2411
rect 3061 2370 3409 2400
rect 3061 2359 3068 2370
rect 3002 2358 3068 2359
rect 3402 2359 3409 2370
rect 3461 2400 3468 2411
rect 3802 2411 3868 2412
rect 3802 2400 3809 2411
rect 3461 2370 3809 2400
rect 3461 2359 3468 2370
rect 3402 2358 3468 2359
rect 3802 2359 3809 2370
rect 3861 2400 3868 2411
rect 4202 2411 4268 2412
rect 4202 2400 4209 2411
rect 3861 2370 4209 2400
rect 3861 2359 3868 2370
rect 3802 2358 3868 2359
rect 4202 2359 4209 2370
rect 4261 2400 4268 2411
rect 4602 2411 4668 2412
rect 4602 2400 4609 2411
rect 4261 2370 4609 2400
rect 4261 2359 4268 2370
rect 4202 2358 4268 2359
rect 4602 2359 4609 2370
rect 4661 2400 4668 2411
rect 5002 2411 5068 2412
rect 5002 2400 5009 2411
rect 4661 2370 5009 2400
rect 4661 2359 4668 2370
rect 4602 2358 4668 2359
rect 5002 2359 5009 2370
rect 5061 2400 5068 2411
rect 5402 2411 5468 2412
rect 5402 2400 5409 2411
rect 5061 2370 5409 2400
rect 5061 2359 5068 2370
rect 5002 2358 5068 2359
rect 5402 2359 5409 2370
rect 5461 2400 5468 2411
rect 5802 2411 5868 2412
rect 5802 2400 5809 2411
rect 5461 2370 5809 2400
rect 5461 2359 5468 2370
rect 5402 2358 5468 2359
rect 5802 2359 5809 2370
rect 5861 2400 5868 2411
rect 6202 2411 6268 2412
rect 6202 2400 6209 2411
rect 5861 2370 6209 2400
rect 5861 2359 5868 2370
rect 5802 2358 5868 2359
rect 6202 2359 6209 2370
rect 6261 2400 6268 2411
rect 6602 2411 6668 2412
rect 6602 2400 6609 2411
rect 6261 2370 6609 2400
rect 6261 2359 6268 2370
rect 6202 2358 6268 2359
rect 6602 2359 6609 2370
rect 6661 2400 6668 2411
rect 7002 2411 7068 2412
rect 7002 2400 7009 2411
rect 6661 2370 7009 2400
rect 6661 2359 6668 2370
rect 6602 2358 6668 2359
rect 7002 2359 7009 2370
rect 7061 2400 7068 2411
rect 7402 2411 7468 2412
rect 7402 2400 7409 2411
rect 7061 2370 7409 2400
rect 7061 2359 7068 2370
rect 7002 2358 7068 2359
rect 7402 2359 7409 2370
rect 7461 2400 7468 2411
rect 7802 2411 7868 2412
rect 7802 2400 7809 2411
rect 7461 2370 7809 2400
rect 7461 2359 7468 2370
rect 7402 2358 7468 2359
rect 7802 2359 7809 2370
rect 7861 2400 7868 2411
rect 8202 2411 8268 2412
rect 8202 2400 8209 2411
rect 7861 2370 8209 2400
rect 7861 2359 7868 2370
rect 7802 2358 7868 2359
rect 8202 2359 8209 2370
rect 8261 2400 8268 2411
rect 8602 2411 8668 2412
rect 8602 2400 8609 2411
rect 8261 2370 8609 2400
rect 8261 2359 8268 2370
rect 8202 2358 8268 2359
rect 8602 2359 8609 2370
rect 8661 2400 8668 2411
rect 9002 2411 9068 2412
rect 9002 2400 9009 2411
rect 8661 2370 9009 2400
rect 8661 2359 8668 2370
rect 8602 2358 8668 2359
rect 9002 2359 9009 2370
rect 9061 2400 9068 2411
rect 9402 2411 9468 2412
rect 9402 2400 9409 2411
rect 9061 2370 9409 2400
rect 9061 2359 9068 2370
rect 9002 2358 9068 2359
rect 9402 2359 9409 2370
rect 9461 2400 9468 2411
rect 9802 2411 9868 2412
rect 9802 2400 9809 2411
rect 9461 2370 9809 2400
rect 9461 2359 9468 2370
rect 9402 2358 9468 2359
rect 9802 2359 9809 2370
rect 9861 2400 9868 2411
rect 10202 2411 10268 2412
rect 10202 2400 10209 2411
rect 9861 2370 10209 2400
rect 9861 2359 9868 2370
rect 9802 2358 9868 2359
rect 10202 2359 10209 2370
rect 10261 2400 10268 2411
rect 10602 2411 10668 2412
rect 10602 2400 10609 2411
rect 10261 2370 10609 2400
rect 10261 2359 10268 2370
rect 10202 2358 10268 2359
rect 10602 2359 10609 2370
rect 10661 2400 10668 2411
rect 11002 2411 11068 2412
rect 11002 2400 11009 2411
rect 10661 2370 11009 2400
rect 10661 2359 10668 2370
rect 10602 2358 10668 2359
rect 11002 2359 11009 2370
rect 11061 2400 11068 2411
rect 11402 2411 11468 2412
rect 11402 2400 11409 2411
rect 11061 2370 11409 2400
rect 11061 2359 11068 2370
rect 11002 2358 11068 2359
rect 11402 2359 11409 2370
rect 11461 2400 11468 2411
rect 11802 2411 11868 2412
rect 11802 2400 11809 2411
rect 11461 2370 11809 2400
rect 11461 2359 11468 2370
rect 11402 2358 11468 2359
rect 11802 2359 11809 2370
rect 11861 2400 11868 2411
rect 12202 2411 12268 2412
rect 12202 2400 12209 2411
rect 11861 2370 12209 2400
rect 11861 2359 11868 2370
rect 11802 2358 11868 2359
rect 12202 2359 12209 2370
rect 12261 2400 12268 2411
rect 12602 2411 12668 2412
rect 12602 2400 12609 2411
rect 12261 2370 12609 2400
rect 12261 2359 12268 2370
rect 12202 2358 12268 2359
rect 12602 2359 12609 2370
rect 12661 2400 12668 2411
rect 13104 2411 13170 2412
rect 13104 2400 13111 2411
rect 12661 2370 13111 2400
rect 12661 2359 12668 2370
rect 12602 2358 12668 2359
rect 13104 2359 13111 2370
rect 13163 2359 13170 2411
rect 13104 2358 13170 2359
rect 2 2341 68 2342
rect 2 2330 9 2341
rect 0 2300 9 2330
rect 2 2289 9 2300
rect 61 2330 68 2341
rect 402 2341 468 2342
rect 402 2330 409 2341
rect 61 2300 409 2330
rect 61 2289 68 2300
rect 2 2288 68 2289
rect 402 2289 409 2300
rect 461 2330 468 2341
rect 802 2341 868 2342
rect 802 2330 809 2341
rect 461 2300 809 2330
rect 461 2289 468 2300
rect 402 2288 468 2289
rect 802 2289 809 2300
rect 861 2330 868 2341
rect 1202 2341 1268 2342
rect 1202 2330 1209 2341
rect 861 2300 1209 2330
rect 861 2289 868 2300
rect 802 2288 868 2289
rect 1202 2289 1209 2300
rect 1261 2330 1268 2341
rect 1602 2341 1668 2342
rect 1602 2330 1609 2341
rect 1261 2300 1609 2330
rect 1261 2289 1268 2300
rect 1202 2288 1268 2289
rect 1602 2289 1609 2300
rect 1661 2330 1668 2341
rect 2002 2341 2068 2342
rect 2002 2330 2009 2341
rect 1661 2300 2009 2330
rect 1661 2289 1668 2300
rect 1602 2288 1668 2289
rect 2002 2289 2009 2300
rect 2061 2330 2068 2341
rect 2402 2341 2468 2342
rect 2402 2330 2409 2341
rect 2061 2300 2409 2330
rect 2061 2289 2068 2300
rect 2002 2288 2068 2289
rect 2402 2289 2409 2300
rect 2461 2330 2468 2341
rect 2802 2341 2868 2342
rect 2802 2330 2809 2341
rect 2461 2300 2809 2330
rect 2461 2289 2468 2300
rect 2402 2288 2468 2289
rect 2802 2289 2809 2300
rect 2861 2330 2868 2341
rect 3202 2341 3268 2342
rect 3202 2330 3209 2341
rect 2861 2300 3209 2330
rect 2861 2289 2868 2300
rect 2802 2288 2868 2289
rect 3202 2289 3209 2300
rect 3261 2330 3268 2341
rect 3602 2341 3668 2342
rect 3602 2330 3609 2341
rect 3261 2300 3609 2330
rect 3261 2289 3268 2300
rect 3202 2288 3268 2289
rect 3602 2289 3609 2300
rect 3661 2330 3668 2341
rect 4002 2341 4068 2342
rect 4002 2330 4009 2341
rect 3661 2300 4009 2330
rect 3661 2289 3668 2300
rect 3602 2288 3668 2289
rect 4002 2289 4009 2300
rect 4061 2330 4068 2341
rect 4402 2341 4468 2342
rect 4402 2330 4409 2341
rect 4061 2300 4409 2330
rect 4061 2289 4068 2300
rect 4002 2288 4068 2289
rect 4402 2289 4409 2300
rect 4461 2330 4468 2341
rect 4802 2341 4868 2342
rect 4802 2330 4809 2341
rect 4461 2300 4809 2330
rect 4461 2289 4468 2300
rect 4402 2288 4468 2289
rect 4802 2289 4809 2300
rect 4861 2330 4868 2341
rect 5202 2341 5268 2342
rect 5202 2330 5209 2341
rect 4861 2300 5209 2330
rect 4861 2289 4868 2300
rect 4802 2288 4868 2289
rect 5202 2289 5209 2300
rect 5261 2330 5268 2341
rect 5602 2341 5668 2342
rect 5602 2330 5609 2341
rect 5261 2300 5609 2330
rect 5261 2289 5268 2300
rect 5202 2288 5268 2289
rect 5602 2289 5609 2300
rect 5661 2330 5668 2341
rect 6002 2341 6068 2342
rect 6002 2330 6009 2341
rect 5661 2300 6009 2330
rect 5661 2289 5668 2300
rect 5602 2288 5668 2289
rect 6002 2289 6009 2300
rect 6061 2330 6068 2341
rect 6402 2341 6468 2342
rect 6402 2330 6409 2341
rect 6061 2300 6409 2330
rect 6061 2289 6068 2300
rect 6002 2288 6068 2289
rect 6402 2289 6409 2300
rect 6461 2330 6468 2341
rect 6802 2341 6868 2342
rect 6802 2330 6809 2341
rect 6461 2300 6809 2330
rect 6461 2289 6468 2300
rect 6402 2288 6468 2289
rect 6802 2289 6809 2300
rect 6861 2330 6868 2341
rect 7202 2341 7268 2342
rect 7202 2330 7209 2341
rect 6861 2300 7209 2330
rect 6861 2289 6868 2300
rect 6802 2288 6868 2289
rect 7202 2289 7209 2300
rect 7261 2330 7268 2341
rect 7602 2341 7668 2342
rect 7602 2330 7609 2341
rect 7261 2300 7609 2330
rect 7261 2289 7268 2300
rect 7202 2288 7268 2289
rect 7602 2289 7609 2300
rect 7661 2330 7668 2341
rect 8002 2341 8068 2342
rect 8002 2330 8009 2341
rect 7661 2300 8009 2330
rect 7661 2289 7668 2300
rect 7602 2288 7668 2289
rect 8002 2289 8009 2300
rect 8061 2330 8068 2341
rect 8402 2341 8468 2342
rect 8402 2330 8409 2341
rect 8061 2300 8409 2330
rect 8061 2289 8068 2300
rect 8002 2288 8068 2289
rect 8402 2289 8409 2300
rect 8461 2330 8468 2341
rect 8802 2341 8868 2342
rect 8802 2330 8809 2341
rect 8461 2300 8809 2330
rect 8461 2289 8468 2300
rect 8402 2288 8468 2289
rect 8802 2289 8809 2300
rect 8861 2330 8868 2341
rect 9202 2341 9268 2342
rect 9202 2330 9209 2341
rect 8861 2300 9209 2330
rect 8861 2289 8868 2300
rect 8802 2288 8868 2289
rect 9202 2289 9209 2300
rect 9261 2330 9268 2341
rect 9602 2341 9668 2342
rect 9602 2330 9609 2341
rect 9261 2300 9609 2330
rect 9261 2289 9268 2300
rect 9202 2288 9268 2289
rect 9602 2289 9609 2300
rect 9661 2330 9668 2341
rect 10002 2341 10068 2342
rect 10002 2330 10009 2341
rect 9661 2300 10009 2330
rect 9661 2289 9668 2300
rect 9602 2288 9668 2289
rect 10002 2289 10009 2300
rect 10061 2330 10068 2341
rect 10402 2341 10468 2342
rect 10402 2330 10409 2341
rect 10061 2300 10409 2330
rect 10061 2289 10068 2300
rect 10002 2288 10068 2289
rect 10402 2289 10409 2300
rect 10461 2330 10468 2341
rect 10802 2341 10868 2342
rect 10802 2330 10809 2341
rect 10461 2300 10809 2330
rect 10461 2289 10468 2300
rect 10402 2288 10468 2289
rect 10802 2289 10809 2300
rect 10861 2330 10868 2341
rect 11202 2341 11268 2342
rect 11202 2330 11209 2341
rect 10861 2300 11209 2330
rect 10861 2289 10868 2300
rect 10802 2288 10868 2289
rect 11202 2289 11209 2300
rect 11261 2330 11268 2341
rect 11602 2341 11668 2342
rect 11602 2330 11609 2341
rect 11261 2300 11609 2330
rect 11261 2289 11268 2300
rect 11202 2288 11268 2289
rect 11602 2289 11609 2300
rect 11661 2330 11668 2341
rect 12002 2341 12068 2342
rect 12002 2330 12009 2341
rect 11661 2300 12009 2330
rect 11661 2289 11668 2300
rect 11602 2288 11668 2289
rect 12002 2289 12009 2300
rect 12061 2330 12068 2341
rect 12402 2341 12468 2342
rect 12402 2330 12409 2341
rect 12061 2300 12409 2330
rect 12061 2289 12068 2300
rect 12002 2288 12068 2289
rect 12402 2289 12409 2300
rect 12461 2330 12468 2341
rect 12802 2341 12868 2342
rect 12802 2330 12809 2341
rect 12461 2300 12809 2330
rect 12461 2289 12468 2300
rect 12402 2288 12468 2289
rect 12802 2289 12809 2300
rect 12861 2330 12868 2341
rect 12900 2341 12966 2342
rect 12900 2330 12907 2341
rect 12861 2300 12907 2330
rect 12861 2289 12868 2300
rect 12802 2288 12868 2289
rect 12900 2289 12907 2300
rect 12959 2289 12966 2341
rect 12900 2288 12966 2289
rect 202 2271 268 2272
rect 202 2260 209 2271
rect 0 2230 209 2260
rect 202 2219 209 2230
rect 261 2260 268 2271
rect 602 2271 668 2272
rect 602 2260 609 2271
rect 261 2230 609 2260
rect 261 2219 268 2230
rect 202 2218 268 2219
rect 602 2219 609 2230
rect 661 2260 668 2271
rect 1002 2271 1068 2272
rect 1002 2260 1009 2271
rect 661 2230 1009 2260
rect 661 2219 668 2230
rect 602 2218 668 2219
rect 1002 2219 1009 2230
rect 1061 2260 1068 2271
rect 1402 2271 1468 2272
rect 1402 2260 1409 2271
rect 1061 2230 1409 2260
rect 1061 2219 1068 2230
rect 1002 2218 1068 2219
rect 1402 2219 1409 2230
rect 1461 2260 1468 2271
rect 1802 2271 1868 2272
rect 1802 2260 1809 2271
rect 1461 2230 1809 2260
rect 1461 2219 1468 2230
rect 1402 2218 1468 2219
rect 1802 2219 1809 2230
rect 1861 2260 1868 2271
rect 2202 2271 2268 2272
rect 2202 2260 2209 2271
rect 1861 2230 2209 2260
rect 1861 2219 1868 2230
rect 1802 2218 1868 2219
rect 2202 2219 2209 2230
rect 2261 2260 2268 2271
rect 2602 2271 2668 2272
rect 2602 2260 2609 2271
rect 2261 2230 2609 2260
rect 2261 2219 2268 2230
rect 2202 2218 2268 2219
rect 2602 2219 2609 2230
rect 2661 2260 2668 2271
rect 3002 2271 3068 2272
rect 3002 2260 3009 2271
rect 2661 2230 3009 2260
rect 2661 2219 2668 2230
rect 2602 2218 2668 2219
rect 3002 2219 3009 2230
rect 3061 2260 3068 2271
rect 3402 2271 3468 2272
rect 3402 2260 3409 2271
rect 3061 2230 3409 2260
rect 3061 2219 3068 2230
rect 3002 2218 3068 2219
rect 3402 2219 3409 2230
rect 3461 2260 3468 2271
rect 3802 2271 3868 2272
rect 3802 2260 3809 2271
rect 3461 2230 3809 2260
rect 3461 2219 3468 2230
rect 3402 2218 3468 2219
rect 3802 2219 3809 2230
rect 3861 2260 3868 2271
rect 4202 2271 4268 2272
rect 4202 2260 4209 2271
rect 3861 2230 4209 2260
rect 3861 2219 3868 2230
rect 3802 2218 3868 2219
rect 4202 2219 4209 2230
rect 4261 2260 4268 2271
rect 4602 2271 4668 2272
rect 4602 2260 4609 2271
rect 4261 2230 4609 2260
rect 4261 2219 4268 2230
rect 4202 2218 4268 2219
rect 4602 2219 4609 2230
rect 4661 2260 4668 2271
rect 5002 2271 5068 2272
rect 5002 2260 5009 2271
rect 4661 2230 5009 2260
rect 4661 2219 4668 2230
rect 4602 2218 4668 2219
rect 5002 2219 5009 2230
rect 5061 2260 5068 2271
rect 5402 2271 5468 2272
rect 5402 2260 5409 2271
rect 5061 2230 5409 2260
rect 5061 2219 5068 2230
rect 5002 2218 5068 2219
rect 5402 2219 5409 2230
rect 5461 2260 5468 2271
rect 5802 2271 5868 2272
rect 5802 2260 5809 2271
rect 5461 2230 5809 2260
rect 5461 2219 5468 2230
rect 5402 2218 5468 2219
rect 5802 2219 5809 2230
rect 5861 2260 5868 2271
rect 6202 2271 6268 2272
rect 6202 2260 6209 2271
rect 5861 2230 6209 2260
rect 5861 2219 5868 2230
rect 5802 2218 5868 2219
rect 6202 2219 6209 2230
rect 6261 2260 6268 2271
rect 6602 2271 6668 2272
rect 6602 2260 6609 2271
rect 6261 2230 6609 2260
rect 6261 2219 6268 2230
rect 6202 2218 6268 2219
rect 6602 2219 6609 2230
rect 6661 2260 6668 2271
rect 7002 2271 7068 2272
rect 7002 2260 7009 2271
rect 6661 2230 7009 2260
rect 6661 2219 6668 2230
rect 6602 2218 6668 2219
rect 7002 2219 7009 2230
rect 7061 2260 7068 2271
rect 7402 2271 7468 2272
rect 7402 2260 7409 2271
rect 7061 2230 7409 2260
rect 7061 2219 7068 2230
rect 7002 2218 7068 2219
rect 7402 2219 7409 2230
rect 7461 2260 7468 2271
rect 7802 2271 7868 2272
rect 7802 2260 7809 2271
rect 7461 2230 7809 2260
rect 7461 2219 7468 2230
rect 7402 2218 7468 2219
rect 7802 2219 7809 2230
rect 7861 2260 7868 2271
rect 8202 2271 8268 2272
rect 8202 2260 8209 2271
rect 7861 2230 8209 2260
rect 7861 2219 7868 2230
rect 7802 2218 7868 2219
rect 8202 2219 8209 2230
rect 8261 2260 8268 2271
rect 8602 2271 8668 2272
rect 8602 2260 8609 2271
rect 8261 2230 8609 2260
rect 8261 2219 8268 2230
rect 8202 2218 8268 2219
rect 8602 2219 8609 2230
rect 8661 2260 8668 2271
rect 9002 2271 9068 2272
rect 9002 2260 9009 2271
rect 8661 2230 9009 2260
rect 8661 2219 8668 2230
rect 8602 2218 8668 2219
rect 9002 2219 9009 2230
rect 9061 2260 9068 2271
rect 9402 2271 9468 2272
rect 9402 2260 9409 2271
rect 9061 2230 9409 2260
rect 9061 2219 9068 2230
rect 9002 2218 9068 2219
rect 9402 2219 9409 2230
rect 9461 2260 9468 2271
rect 9802 2271 9868 2272
rect 9802 2260 9809 2271
rect 9461 2230 9809 2260
rect 9461 2219 9468 2230
rect 9402 2218 9468 2219
rect 9802 2219 9809 2230
rect 9861 2260 9868 2271
rect 10202 2271 10268 2272
rect 10202 2260 10209 2271
rect 9861 2230 10209 2260
rect 9861 2219 9868 2230
rect 9802 2218 9868 2219
rect 10202 2219 10209 2230
rect 10261 2260 10268 2271
rect 10602 2271 10668 2272
rect 10602 2260 10609 2271
rect 10261 2230 10609 2260
rect 10261 2219 10268 2230
rect 10202 2218 10268 2219
rect 10602 2219 10609 2230
rect 10661 2260 10668 2271
rect 11002 2271 11068 2272
rect 11002 2260 11009 2271
rect 10661 2230 11009 2260
rect 10661 2219 10668 2230
rect 10602 2218 10668 2219
rect 11002 2219 11009 2230
rect 11061 2260 11068 2271
rect 11402 2271 11468 2272
rect 11402 2260 11409 2271
rect 11061 2230 11409 2260
rect 11061 2219 11068 2230
rect 11002 2218 11068 2219
rect 11402 2219 11409 2230
rect 11461 2260 11468 2271
rect 11802 2271 11868 2272
rect 11802 2260 11809 2271
rect 11461 2230 11809 2260
rect 11461 2219 11468 2230
rect 11402 2218 11468 2219
rect 11802 2219 11809 2230
rect 11861 2260 11868 2271
rect 12202 2271 12268 2272
rect 12202 2260 12209 2271
rect 11861 2230 12209 2260
rect 11861 2219 11868 2230
rect 11802 2218 11868 2219
rect 12202 2219 12209 2230
rect 12261 2260 12268 2271
rect 12602 2271 12668 2272
rect 12602 2260 12609 2271
rect 12261 2230 12609 2260
rect 12261 2219 12268 2230
rect 12202 2218 12268 2219
rect 12602 2219 12609 2230
rect 12661 2260 12668 2271
rect 13104 2271 13170 2272
rect 13104 2260 13111 2271
rect 12661 2230 13111 2260
rect 12661 2219 12668 2230
rect 12602 2218 12668 2219
rect 13104 2219 13111 2230
rect 13163 2219 13170 2271
rect 13104 2218 13170 2219
rect 2 2201 68 2202
rect 2 2190 9 2201
rect 0 2160 9 2190
rect 2 2149 9 2160
rect 61 2190 68 2201
rect 402 2201 468 2202
rect 402 2190 409 2201
rect 61 2160 409 2190
rect 61 2149 68 2160
rect 2 2148 68 2149
rect 402 2149 409 2160
rect 461 2190 468 2201
rect 802 2201 868 2202
rect 802 2190 809 2201
rect 461 2160 809 2190
rect 461 2149 468 2160
rect 402 2148 468 2149
rect 802 2149 809 2160
rect 861 2190 868 2201
rect 1202 2201 1268 2202
rect 1202 2190 1209 2201
rect 861 2160 1209 2190
rect 861 2149 868 2160
rect 802 2148 868 2149
rect 1202 2149 1209 2160
rect 1261 2190 1268 2201
rect 1602 2201 1668 2202
rect 1602 2190 1609 2201
rect 1261 2160 1609 2190
rect 1261 2149 1268 2160
rect 1202 2148 1268 2149
rect 1602 2149 1609 2160
rect 1661 2190 1668 2201
rect 2002 2201 2068 2202
rect 2002 2190 2009 2201
rect 1661 2160 2009 2190
rect 1661 2149 1668 2160
rect 1602 2148 1668 2149
rect 2002 2149 2009 2160
rect 2061 2190 2068 2201
rect 2402 2201 2468 2202
rect 2402 2190 2409 2201
rect 2061 2160 2409 2190
rect 2061 2149 2068 2160
rect 2002 2148 2068 2149
rect 2402 2149 2409 2160
rect 2461 2190 2468 2201
rect 2802 2201 2868 2202
rect 2802 2190 2809 2201
rect 2461 2160 2809 2190
rect 2461 2149 2468 2160
rect 2402 2148 2468 2149
rect 2802 2149 2809 2160
rect 2861 2190 2868 2201
rect 3202 2201 3268 2202
rect 3202 2190 3209 2201
rect 2861 2160 3209 2190
rect 2861 2149 2868 2160
rect 2802 2148 2868 2149
rect 3202 2149 3209 2160
rect 3261 2190 3268 2201
rect 3602 2201 3668 2202
rect 3602 2190 3609 2201
rect 3261 2160 3609 2190
rect 3261 2149 3268 2160
rect 3202 2148 3268 2149
rect 3602 2149 3609 2160
rect 3661 2190 3668 2201
rect 4002 2201 4068 2202
rect 4002 2190 4009 2201
rect 3661 2160 4009 2190
rect 3661 2149 3668 2160
rect 3602 2148 3668 2149
rect 4002 2149 4009 2160
rect 4061 2190 4068 2201
rect 4402 2201 4468 2202
rect 4402 2190 4409 2201
rect 4061 2160 4409 2190
rect 4061 2149 4068 2160
rect 4002 2148 4068 2149
rect 4402 2149 4409 2160
rect 4461 2190 4468 2201
rect 4802 2201 4868 2202
rect 4802 2190 4809 2201
rect 4461 2160 4809 2190
rect 4461 2149 4468 2160
rect 4402 2148 4468 2149
rect 4802 2149 4809 2160
rect 4861 2190 4868 2201
rect 5202 2201 5268 2202
rect 5202 2190 5209 2201
rect 4861 2160 5209 2190
rect 4861 2149 4868 2160
rect 4802 2148 4868 2149
rect 5202 2149 5209 2160
rect 5261 2190 5268 2201
rect 5602 2201 5668 2202
rect 5602 2190 5609 2201
rect 5261 2160 5609 2190
rect 5261 2149 5268 2160
rect 5202 2148 5268 2149
rect 5602 2149 5609 2160
rect 5661 2190 5668 2201
rect 6002 2201 6068 2202
rect 6002 2190 6009 2201
rect 5661 2160 6009 2190
rect 5661 2149 5668 2160
rect 5602 2148 5668 2149
rect 6002 2149 6009 2160
rect 6061 2190 6068 2201
rect 6402 2201 6468 2202
rect 6402 2190 6409 2201
rect 6061 2160 6409 2190
rect 6061 2149 6068 2160
rect 6002 2148 6068 2149
rect 6402 2149 6409 2160
rect 6461 2190 6468 2201
rect 6802 2201 6868 2202
rect 6802 2190 6809 2201
rect 6461 2160 6809 2190
rect 6461 2149 6468 2160
rect 6402 2148 6468 2149
rect 6802 2149 6809 2160
rect 6861 2190 6868 2201
rect 7202 2201 7268 2202
rect 7202 2190 7209 2201
rect 6861 2160 7209 2190
rect 6861 2149 6868 2160
rect 6802 2148 6868 2149
rect 7202 2149 7209 2160
rect 7261 2190 7268 2201
rect 7602 2201 7668 2202
rect 7602 2190 7609 2201
rect 7261 2160 7609 2190
rect 7261 2149 7268 2160
rect 7202 2148 7268 2149
rect 7602 2149 7609 2160
rect 7661 2190 7668 2201
rect 8002 2201 8068 2202
rect 8002 2190 8009 2201
rect 7661 2160 8009 2190
rect 7661 2149 7668 2160
rect 7602 2148 7668 2149
rect 8002 2149 8009 2160
rect 8061 2190 8068 2201
rect 8402 2201 8468 2202
rect 8402 2190 8409 2201
rect 8061 2160 8409 2190
rect 8061 2149 8068 2160
rect 8002 2148 8068 2149
rect 8402 2149 8409 2160
rect 8461 2190 8468 2201
rect 8802 2201 8868 2202
rect 8802 2190 8809 2201
rect 8461 2160 8809 2190
rect 8461 2149 8468 2160
rect 8402 2148 8468 2149
rect 8802 2149 8809 2160
rect 8861 2190 8868 2201
rect 9202 2201 9268 2202
rect 9202 2190 9209 2201
rect 8861 2160 9209 2190
rect 8861 2149 8868 2160
rect 8802 2148 8868 2149
rect 9202 2149 9209 2160
rect 9261 2190 9268 2201
rect 9602 2201 9668 2202
rect 9602 2190 9609 2201
rect 9261 2160 9609 2190
rect 9261 2149 9268 2160
rect 9202 2148 9268 2149
rect 9602 2149 9609 2160
rect 9661 2190 9668 2201
rect 10002 2201 10068 2202
rect 10002 2190 10009 2201
rect 9661 2160 10009 2190
rect 9661 2149 9668 2160
rect 9602 2148 9668 2149
rect 10002 2149 10009 2160
rect 10061 2190 10068 2201
rect 10402 2201 10468 2202
rect 10402 2190 10409 2201
rect 10061 2160 10409 2190
rect 10061 2149 10068 2160
rect 10002 2148 10068 2149
rect 10402 2149 10409 2160
rect 10461 2190 10468 2201
rect 10802 2201 10868 2202
rect 10802 2190 10809 2201
rect 10461 2160 10809 2190
rect 10461 2149 10468 2160
rect 10402 2148 10468 2149
rect 10802 2149 10809 2160
rect 10861 2190 10868 2201
rect 11202 2201 11268 2202
rect 11202 2190 11209 2201
rect 10861 2160 11209 2190
rect 10861 2149 10868 2160
rect 10802 2148 10868 2149
rect 11202 2149 11209 2160
rect 11261 2190 11268 2201
rect 11602 2201 11668 2202
rect 11602 2190 11609 2201
rect 11261 2160 11609 2190
rect 11261 2149 11268 2160
rect 11202 2148 11268 2149
rect 11602 2149 11609 2160
rect 11661 2190 11668 2201
rect 12002 2201 12068 2202
rect 12002 2190 12009 2201
rect 11661 2160 12009 2190
rect 11661 2149 11668 2160
rect 11602 2148 11668 2149
rect 12002 2149 12009 2160
rect 12061 2190 12068 2201
rect 12402 2201 12468 2202
rect 12402 2190 12409 2201
rect 12061 2160 12409 2190
rect 12061 2149 12068 2160
rect 12002 2148 12068 2149
rect 12402 2149 12409 2160
rect 12461 2190 12468 2201
rect 12802 2201 12868 2202
rect 12802 2190 12809 2201
rect 12461 2160 12809 2190
rect 12461 2149 12468 2160
rect 12402 2148 12468 2149
rect 12802 2149 12809 2160
rect 12861 2190 12868 2201
rect 12900 2201 12966 2202
rect 12900 2190 12907 2201
rect 12861 2160 12907 2190
rect 12861 2149 12868 2160
rect 12802 2148 12868 2149
rect 12900 2149 12907 2160
rect 12959 2149 12966 2201
rect 12900 2148 12966 2149
rect 202 2131 268 2132
rect 202 2120 209 2131
rect 0 2090 209 2120
rect 202 2079 209 2090
rect 261 2120 268 2131
rect 602 2131 668 2132
rect 602 2120 609 2131
rect 261 2090 609 2120
rect 261 2079 268 2090
rect 202 2078 268 2079
rect 602 2079 609 2090
rect 661 2120 668 2131
rect 1002 2131 1068 2132
rect 1002 2120 1009 2131
rect 661 2090 1009 2120
rect 661 2079 668 2090
rect 602 2078 668 2079
rect 1002 2079 1009 2090
rect 1061 2120 1068 2131
rect 1402 2131 1468 2132
rect 1402 2120 1409 2131
rect 1061 2090 1409 2120
rect 1061 2079 1068 2090
rect 1002 2078 1068 2079
rect 1402 2079 1409 2090
rect 1461 2120 1468 2131
rect 1802 2131 1868 2132
rect 1802 2120 1809 2131
rect 1461 2090 1809 2120
rect 1461 2079 1468 2090
rect 1402 2078 1468 2079
rect 1802 2079 1809 2090
rect 1861 2120 1868 2131
rect 2202 2131 2268 2132
rect 2202 2120 2209 2131
rect 1861 2090 2209 2120
rect 1861 2079 1868 2090
rect 1802 2078 1868 2079
rect 2202 2079 2209 2090
rect 2261 2120 2268 2131
rect 2602 2131 2668 2132
rect 2602 2120 2609 2131
rect 2261 2090 2609 2120
rect 2261 2079 2268 2090
rect 2202 2078 2268 2079
rect 2602 2079 2609 2090
rect 2661 2120 2668 2131
rect 3002 2131 3068 2132
rect 3002 2120 3009 2131
rect 2661 2090 3009 2120
rect 2661 2079 2668 2090
rect 2602 2078 2668 2079
rect 3002 2079 3009 2090
rect 3061 2120 3068 2131
rect 3402 2131 3468 2132
rect 3402 2120 3409 2131
rect 3061 2090 3409 2120
rect 3061 2079 3068 2090
rect 3002 2078 3068 2079
rect 3402 2079 3409 2090
rect 3461 2120 3468 2131
rect 3802 2131 3868 2132
rect 3802 2120 3809 2131
rect 3461 2090 3809 2120
rect 3461 2079 3468 2090
rect 3402 2078 3468 2079
rect 3802 2079 3809 2090
rect 3861 2120 3868 2131
rect 4202 2131 4268 2132
rect 4202 2120 4209 2131
rect 3861 2090 4209 2120
rect 3861 2079 3868 2090
rect 3802 2078 3868 2079
rect 4202 2079 4209 2090
rect 4261 2120 4268 2131
rect 4602 2131 4668 2132
rect 4602 2120 4609 2131
rect 4261 2090 4609 2120
rect 4261 2079 4268 2090
rect 4202 2078 4268 2079
rect 4602 2079 4609 2090
rect 4661 2120 4668 2131
rect 5002 2131 5068 2132
rect 5002 2120 5009 2131
rect 4661 2090 5009 2120
rect 4661 2079 4668 2090
rect 4602 2078 4668 2079
rect 5002 2079 5009 2090
rect 5061 2120 5068 2131
rect 5402 2131 5468 2132
rect 5402 2120 5409 2131
rect 5061 2090 5409 2120
rect 5061 2079 5068 2090
rect 5002 2078 5068 2079
rect 5402 2079 5409 2090
rect 5461 2120 5468 2131
rect 5802 2131 5868 2132
rect 5802 2120 5809 2131
rect 5461 2090 5809 2120
rect 5461 2079 5468 2090
rect 5402 2078 5468 2079
rect 5802 2079 5809 2090
rect 5861 2120 5868 2131
rect 6202 2131 6268 2132
rect 6202 2120 6209 2131
rect 5861 2090 6209 2120
rect 5861 2079 5868 2090
rect 5802 2078 5868 2079
rect 6202 2079 6209 2090
rect 6261 2120 6268 2131
rect 6602 2131 6668 2132
rect 6602 2120 6609 2131
rect 6261 2090 6609 2120
rect 6261 2079 6268 2090
rect 6202 2078 6268 2079
rect 6602 2079 6609 2090
rect 6661 2120 6668 2131
rect 7002 2131 7068 2132
rect 7002 2120 7009 2131
rect 6661 2090 7009 2120
rect 6661 2079 6668 2090
rect 6602 2078 6668 2079
rect 7002 2079 7009 2090
rect 7061 2120 7068 2131
rect 7402 2131 7468 2132
rect 7402 2120 7409 2131
rect 7061 2090 7409 2120
rect 7061 2079 7068 2090
rect 7002 2078 7068 2079
rect 7402 2079 7409 2090
rect 7461 2120 7468 2131
rect 7802 2131 7868 2132
rect 7802 2120 7809 2131
rect 7461 2090 7809 2120
rect 7461 2079 7468 2090
rect 7402 2078 7468 2079
rect 7802 2079 7809 2090
rect 7861 2120 7868 2131
rect 8202 2131 8268 2132
rect 8202 2120 8209 2131
rect 7861 2090 8209 2120
rect 7861 2079 7868 2090
rect 7802 2078 7868 2079
rect 8202 2079 8209 2090
rect 8261 2120 8268 2131
rect 8602 2131 8668 2132
rect 8602 2120 8609 2131
rect 8261 2090 8609 2120
rect 8261 2079 8268 2090
rect 8202 2078 8268 2079
rect 8602 2079 8609 2090
rect 8661 2120 8668 2131
rect 9002 2131 9068 2132
rect 9002 2120 9009 2131
rect 8661 2090 9009 2120
rect 8661 2079 8668 2090
rect 8602 2078 8668 2079
rect 9002 2079 9009 2090
rect 9061 2120 9068 2131
rect 9402 2131 9468 2132
rect 9402 2120 9409 2131
rect 9061 2090 9409 2120
rect 9061 2079 9068 2090
rect 9002 2078 9068 2079
rect 9402 2079 9409 2090
rect 9461 2120 9468 2131
rect 9802 2131 9868 2132
rect 9802 2120 9809 2131
rect 9461 2090 9809 2120
rect 9461 2079 9468 2090
rect 9402 2078 9468 2079
rect 9802 2079 9809 2090
rect 9861 2120 9868 2131
rect 10202 2131 10268 2132
rect 10202 2120 10209 2131
rect 9861 2090 10209 2120
rect 9861 2079 9868 2090
rect 9802 2078 9868 2079
rect 10202 2079 10209 2090
rect 10261 2120 10268 2131
rect 10602 2131 10668 2132
rect 10602 2120 10609 2131
rect 10261 2090 10609 2120
rect 10261 2079 10268 2090
rect 10202 2078 10268 2079
rect 10602 2079 10609 2090
rect 10661 2120 10668 2131
rect 11002 2131 11068 2132
rect 11002 2120 11009 2131
rect 10661 2090 11009 2120
rect 10661 2079 10668 2090
rect 10602 2078 10668 2079
rect 11002 2079 11009 2090
rect 11061 2120 11068 2131
rect 11402 2131 11468 2132
rect 11402 2120 11409 2131
rect 11061 2090 11409 2120
rect 11061 2079 11068 2090
rect 11002 2078 11068 2079
rect 11402 2079 11409 2090
rect 11461 2120 11468 2131
rect 11802 2131 11868 2132
rect 11802 2120 11809 2131
rect 11461 2090 11809 2120
rect 11461 2079 11468 2090
rect 11402 2078 11468 2079
rect 11802 2079 11809 2090
rect 11861 2120 11868 2131
rect 12202 2131 12268 2132
rect 12202 2120 12209 2131
rect 11861 2090 12209 2120
rect 11861 2079 11868 2090
rect 11802 2078 11868 2079
rect 12202 2079 12209 2090
rect 12261 2120 12268 2131
rect 12602 2131 12668 2132
rect 12602 2120 12609 2131
rect 12261 2090 12609 2120
rect 12261 2079 12268 2090
rect 12202 2078 12268 2079
rect 12602 2079 12609 2090
rect 12661 2120 12668 2131
rect 13104 2131 13170 2132
rect 13104 2120 13111 2131
rect 12661 2090 13111 2120
rect 12661 2079 12668 2090
rect 12602 2078 12668 2079
rect 13104 2079 13111 2090
rect 13163 2079 13170 2131
rect 13104 2078 13170 2079
rect 2 2061 68 2062
rect 2 2050 9 2061
rect 0 2020 9 2050
rect 2 2009 9 2020
rect 61 2050 68 2061
rect 402 2061 468 2062
rect 402 2050 409 2061
rect 61 2020 409 2050
rect 61 2009 68 2020
rect 2 2008 68 2009
rect 402 2009 409 2020
rect 461 2050 468 2061
rect 802 2061 868 2062
rect 802 2050 809 2061
rect 461 2020 809 2050
rect 461 2009 468 2020
rect 402 2008 468 2009
rect 802 2009 809 2020
rect 861 2050 868 2061
rect 1202 2061 1268 2062
rect 1202 2050 1209 2061
rect 861 2020 1209 2050
rect 861 2009 868 2020
rect 802 2008 868 2009
rect 1202 2009 1209 2020
rect 1261 2050 1268 2061
rect 1602 2061 1668 2062
rect 1602 2050 1609 2061
rect 1261 2020 1609 2050
rect 1261 2009 1268 2020
rect 1202 2008 1268 2009
rect 1602 2009 1609 2020
rect 1661 2050 1668 2061
rect 2002 2061 2068 2062
rect 2002 2050 2009 2061
rect 1661 2020 2009 2050
rect 1661 2009 1668 2020
rect 1602 2008 1668 2009
rect 2002 2009 2009 2020
rect 2061 2050 2068 2061
rect 2402 2061 2468 2062
rect 2402 2050 2409 2061
rect 2061 2020 2409 2050
rect 2061 2009 2068 2020
rect 2002 2008 2068 2009
rect 2402 2009 2409 2020
rect 2461 2050 2468 2061
rect 2802 2061 2868 2062
rect 2802 2050 2809 2061
rect 2461 2020 2809 2050
rect 2461 2009 2468 2020
rect 2402 2008 2468 2009
rect 2802 2009 2809 2020
rect 2861 2050 2868 2061
rect 3202 2061 3268 2062
rect 3202 2050 3209 2061
rect 2861 2020 3209 2050
rect 2861 2009 2868 2020
rect 2802 2008 2868 2009
rect 3202 2009 3209 2020
rect 3261 2050 3268 2061
rect 3602 2061 3668 2062
rect 3602 2050 3609 2061
rect 3261 2020 3609 2050
rect 3261 2009 3268 2020
rect 3202 2008 3268 2009
rect 3602 2009 3609 2020
rect 3661 2050 3668 2061
rect 4002 2061 4068 2062
rect 4002 2050 4009 2061
rect 3661 2020 4009 2050
rect 3661 2009 3668 2020
rect 3602 2008 3668 2009
rect 4002 2009 4009 2020
rect 4061 2050 4068 2061
rect 4402 2061 4468 2062
rect 4402 2050 4409 2061
rect 4061 2020 4409 2050
rect 4061 2009 4068 2020
rect 4002 2008 4068 2009
rect 4402 2009 4409 2020
rect 4461 2050 4468 2061
rect 4802 2061 4868 2062
rect 4802 2050 4809 2061
rect 4461 2020 4809 2050
rect 4461 2009 4468 2020
rect 4402 2008 4468 2009
rect 4802 2009 4809 2020
rect 4861 2050 4868 2061
rect 5202 2061 5268 2062
rect 5202 2050 5209 2061
rect 4861 2020 5209 2050
rect 4861 2009 4868 2020
rect 4802 2008 4868 2009
rect 5202 2009 5209 2020
rect 5261 2050 5268 2061
rect 5602 2061 5668 2062
rect 5602 2050 5609 2061
rect 5261 2020 5609 2050
rect 5261 2009 5268 2020
rect 5202 2008 5268 2009
rect 5602 2009 5609 2020
rect 5661 2050 5668 2061
rect 6002 2061 6068 2062
rect 6002 2050 6009 2061
rect 5661 2020 6009 2050
rect 5661 2009 5668 2020
rect 5602 2008 5668 2009
rect 6002 2009 6009 2020
rect 6061 2050 6068 2061
rect 6402 2061 6468 2062
rect 6402 2050 6409 2061
rect 6061 2020 6409 2050
rect 6061 2009 6068 2020
rect 6002 2008 6068 2009
rect 6402 2009 6409 2020
rect 6461 2050 6468 2061
rect 6802 2061 6868 2062
rect 6802 2050 6809 2061
rect 6461 2020 6809 2050
rect 6461 2009 6468 2020
rect 6402 2008 6468 2009
rect 6802 2009 6809 2020
rect 6861 2050 6868 2061
rect 7202 2061 7268 2062
rect 7202 2050 7209 2061
rect 6861 2020 7209 2050
rect 6861 2009 6868 2020
rect 6802 2008 6868 2009
rect 7202 2009 7209 2020
rect 7261 2050 7268 2061
rect 7602 2061 7668 2062
rect 7602 2050 7609 2061
rect 7261 2020 7609 2050
rect 7261 2009 7268 2020
rect 7202 2008 7268 2009
rect 7602 2009 7609 2020
rect 7661 2050 7668 2061
rect 8002 2061 8068 2062
rect 8002 2050 8009 2061
rect 7661 2020 8009 2050
rect 7661 2009 7668 2020
rect 7602 2008 7668 2009
rect 8002 2009 8009 2020
rect 8061 2050 8068 2061
rect 8402 2061 8468 2062
rect 8402 2050 8409 2061
rect 8061 2020 8409 2050
rect 8061 2009 8068 2020
rect 8002 2008 8068 2009
rect 8402 2009 8409 2020
rect 8461 2050 8468 2061
rect 8802 2061 8868 2062
rect 8802 2050 8809 2061
rect 8461 2020 8809 2050
rect 8461 2009 8468 2020
rect 8402 2008 8468 2009
rect 8802 2009 8809 2020
rect 8861 2050 8868 2061
rect 9202 2061 9268 2062
rect 9202 2050 9209 2061
rect 8861 2020 9209 2050
rect 8861 2009 8868 2020
rect 8802 2008 8868 2009
rect 9202 2009 9209 2020
rect 9261 2050 9268 2061
rect 9602 2061 9668 2062
rect 9602 2050 9609 2061
rect 9261 2020 9609 2050
rect 9261 2009 9268 2020
rect 9202 2008 9268 2009
rect 9602 2009 9609 2020
rect 9661 2050 9668 2061
rect 10002 2061 10068 2062
rect 10002 2050 10009 2061
rect 9661 2020 10009 2050
rect 9661 2009 9668 2020
rect 9602 2008 9668 2009
rect 10002 2009 10009 2020
rect 10061 2050 10068 2061
rect 10402 2061 10468 2062
rect 10402 2050 10409 2061
rect 10061 2020 10409 2050
rect 10061 2009 10068 2020
rect 10002 2008 10068 2009
rect 10402 2009 10409 2020
rect 10461 2050 10468 2061
rect 10802 2061 10868 2062
rect 10802 2050 10809 2061
rect 10461 2020 10809 2050
rect 10461 2009 10468 2020
rect 10402 2008 10468 2009
rect 10802 2009 10809 2020
rect 10861 2050 10868 2061
rect 11202 2061 11268 2062
rect 11202 2050 11209 2061
rect 10861 2020 11209 2050
rect 10861 2009 10868 2020
rect 10802 2008 10868 2009
rect 11202 2009 11209 2020
rect 11261 2050 11268 2061
rect 11602 2061 11668 2062
rect 11602 2050 11609 2061
rect 11261 2020 11609 2050
rect 11261 2009 11268 2020
rect 11202 2008 11268 2009
rect 11602 2009 11609 2020
rect 11661 2050 11668 2061
rect 12002 2061 12068 2062
rect 12002 2050 12009 2061
rect 11661 2020 12009 2050
rect 11661 2009 11668 2020
rect 11602 2008 11668 2009
rect 12002 2009 12009 2020
rect 12061 2050 12068 2061
rect 12402 2061 12468 2062
rect 12402 2050 12409 2061
rect 12061 2020 12409 2050
rect 12061 2009 12068 2020
rect 12002 2008 12068 2009
rect 12402 2009 12409 2020
rect 12461 2050 12468 2061
rect 12802 2061 12868 2062
rect 12802 2050 12809 2061
rect 12461 2020 12809 2050
rect 12461 2009 12468 2020
rect 12402 2008 12468 2009
rect 12802 2009 12809 2020
rect 12861 2050 12868 2061
rect 12900 2061 12966 2062
rect 12900 2050 12907 2061
rect 12861 2020 12907 2050
rect 12861 2009 12868 2020
rect 12802 2008 12868 2009
rect 12900 2009 12907 2020
rect 12959 2009 12966 2061
rect 12900 2008 12966 2009
rect 202 1991 268 1992
rect 202 1980 209 1991
rect 0 1950 209 1980
rect 202 1939 209 1950
rect 261 1980 268 1991
rect 602 1991 668 1992
rect 602 1980 609 1991
rect 261 1950 609 1980
rect 261 1939 268 1950
rect 202 1938 268 1939
rect 602 1939 609 1950
rect 661 1980 668 1991
rect 1002 1991 1068 1992
rect 1002 1980 1009 1991
rect 661 1950 1009 1980
rect 661 1939 668 1950
rect 602 1938 668 1939
rect 1002 1939 1009 1950
rect 1061 1980 1068 1991
rect 1402 1991 1468 1992
rect 1402 1980 1409 1991
rect 1061 1950 1409 1980
rect 1061 1939 1068 1950
rect 1002 1938 1068 1939
rect 1402 1939 1409 1950
rect 1461 1980 1468 1991
rect 1802 1991 1868 1992
rect 1802 1980 1809 1991
rect 1461 1950 1809 1980
rect 1461 1939 1468 1950
rect 1402 1938 1468 1939
rect 1802 1939 1809 1950
rect 1861 1980 1868 1991
rect 2202 1991 2268 1992
rect 2202 1980 2209 1991
rect 1861 1950 2209 1980
rect 1861 1939 1868 1950
rect 1802 1938 1868 1939
rect 2202 1939 2209 1950
rect 2261 1980 2268 1991
rect 2602 1991 2668 1992
rect 2602 1980 2609 1991
rect 2261 1950 2609 1980
rect 2261 1939 2268 1950
rect 2202 1938 2268 1939
rect 2602 1939 2609 1950
rect 2661 1980 2668 1991
rect 3002 1991 3068 1992
rect 3002 1980 3009 1991
rect 2661 1950 3009 1980
rect 2661 1939 2668 1950
rect 2602 1938 2668 1939
rect 3002 1939 3009 1950
rect 3061 1980 3068 1991
rect 3402 1991 3468 1992
rect 3402 1980 3409 1991
rect 3061 1950 3409 1980
rect 3061 1939 3068 1950
rect 3002 1938 3068 1939
rect 3402 1939 3409 1950
rect 3461 1980 3468 1991
rect 3802 1991 3868 1992
rect 3802 1980 3809 1991
rect 3461 1950 3809 1980
rect 3461 1939 3468 1950
rect 3402 1938 3468 1939
rect 3802 1939 3809 1950
rect 3861 1980 3868 1991
rect 4202 1991 4268 1992
rect 4202 1980 4209 1991
rect 3861 1950 4209 1980
rect 3861 1939 3868 1950
rect 3802 1938 3868 1939
rect 4202 1939 4209 1950
rect 4261 1980 4268 1991
rect 4602 1991 4668 1992
rect 4602 1980 4609 1991
rect 4261 1950 4609 1980
rect 4261 1939 4268 1950
rect 4202 1938 4268 1939
rect 4602 1939 4609 1950
rect 4661 1980 4668 1991
rect 5002 1991 5068 1992
rect 5002 1980 5009 1991
rect 4661 1950 5009 1980
rect 4661 1939 4668 1950
rect 4602 1938 4668 1939
rect 5002 1939 5009 1950
rect 5061 1980 5068 1991
rect 5402 1991 5468 1992
rect 5402 1980 5409 1991
rect 5061 1950 5409 1980
rect 5061 1939 5068 1950
rect 5002 1938 5068 1939
rect 5402 1939 5409 1950
rect 5461 1980 5468 1991
rect 5802 1991 5868 1992
rect 5802 1980 5809 1991
rect 5461 1950 5809 1980
rect 5461 1939 5468 1950
rect 5402 1938 5468 1939
rect 5802 1939 5809 1950
rect 5861 1980 5868 1991
rect 6202 1991 6268 1992
rect 6202 1980 6209 1991
rect 5861 1950 6209 1980
rect 5861 1939 5868 1950
rect 5802 1938 5868 1939
rect 6202 1939 6209 1950
rect 6261 1980 6268 1991
rect 6602 1991 6668 1992
rect 6602 1980 6609 1991
rect 6261 1950 6609 1980
rect 6261 1939 6268 1950
rect 6202 1938 6268 1939
rect 6602 1939 6609 1950
rect 6661 1980 6668 1991
rect 7002 1991 7068 1992
rect 7002 1980 7009 1991
rect 6661 1950 7009 1980
rect 6661 1939 6668 1950
rect 6602 1938 6668 1939
rect 7002 1939 7009 1950
rect 7061 1980 7068 1991
rect 7402 1991 7468 1992
rect 7402 1980 7409 1991
rect 7061 1950 7409 1980
rect 7061 1939 7068 1950
rect 7002 1938 7068 1939
rect 7402 1939 7409 1950
rect 7461 1980 7468 1991
rect 7802 1991 7868 1992
rect 7802 1980 7809 1991
rect 7461 1950 7809 1980
rect 7461 1939 7468 1950
rect 7402 1938 7468 1939
rect 7802 1939 7809 1950
rect 7861 1980 7868 1991
rect 8202 1991 8268 1992
rect 8202 1980 8209 1991
rect 7861 1950 8209 1980
rect 7861 1939 7868 1950
rect 7802 1938 7868 1939
rect 8202 1939 8209 1950
rect 8261 1980 8268 1991
rect 8602 1991 8668 1992
rect 8602 1980 8609 1991
rect 8261 1950 8609 1980
rect 8261 1939 8268 1950
rect 8202 1938 8268 1939
rect 8602 1939 8609 1950
rect 8661 1980 8668 1991
rect 9002 1991 9068 1992
rect 9002 1980 9009 1991
rect 8661 1950 9009 1980
rect 8661 1939 8668 1950
rect 8602 1938 8668 1939
rect 9002 1939 9009 1950
rect 9061 1980 9068 1991
rect 9402 1991 9468 1992
rect 9402 1980 9409 1991
rect 9061 1950 9409 1980
rect 9061 1939 9068 1950
rect 9002 1938 9068 1939
rect 9402 1939 9409 1950
rect 9461 1980 9468 1991
rect 9802 1991 9868 1992
rect 9802 1980 9809 1991
rect 9461 1950 9809 1980
rect 9461 1939 9468 1950
rect 9402 1938 9468 1939
rect 9802 1939 9809 1950
rect 9861 1980 9868 1991
rect 10202 1991 10268 1992
rect 10202 1980 10209 1991
rect 9861 1950 10209 1980
rect 9861 1939 9868 1950
rect 9802 1938 9868 1939
rect 10202 1939 10209 1950
rect 10261 1980 10268 1991
rect 10602 1991 10668 1992
rect 10602 1980 10609 1991
rect 10261 1950 10609 1980
rect 10261 1939 10268 1950
rect 10202 1938 10268 1939
rect 10602 1939 10609 1950
rect 10661 1980 10668 1991
rect 11002 1991 11068 1992
rect 11002 1980 11009 1991
rect 10661 1950 11009 1980
rect 10661 1939 10668 1950
rect 10602 1938 10668 1939
rect 11002 1939 11009 1950
rect 11061 1980 11068 1991
rect 11402 1991 11468 1992
rect 11402 1980 11409 1991
rect 11061 1950 11409 1980
rect 11061 1939 11068 1950
rect 11002 1938 11068 1939
rect 11402 1939 11409 1950
rect 11461 1980 11468 1991
rect 11802 1991 11868 1992
rect 11802 1980 11809 1991
rect 11461 1950 11809 1980
rect 11461 1939 11468 1950
rect 11402 1938 11468 1939
rect 11802 1939 11809 1950
rect 11861 1980 11868 1991
rect 12202 1991 12268 1992
rect 12202 1980 12209 1991
rect 11861 1950 12209 1980
rect 11861 1939 11868 1950
rect 11802 1938 11868 1939
rect 12202 1939 12209 1950
rect 12261 1980 12268 1991
rect 12602 1991 12668 1992
rect 12602 1980 12609 1991
rect 12261 1950 12609 1980
rect 12261 1939 12268 1950
rect 12202 1938 12268 1939
rect 12602 1939 12609 1950
rect 12661 1980 12668 1991
rect 13104 1991 13170 1992
rect 13104 1980 13111 1991
rect 12661 1950 13111 1980
rect 12661 1939 12668 1950
rect 12602 1938 12668 1939
rect 13104 1939 13111 1950
rect 13163 1939 13170 1991
rect 13104 1938 13170 1939
rect 2 1921 68 1922
rect 2 1910 9 1921
rect 0 1880 9 1910
rect 2 1869 9 1880
rect 61 1910 68 1921
rect 402 1921 468 1922
rect 402 1910 409 1921
rect 61 1880 409 1910
rect 61 1869 68 1880
rect 2 1868 68 1869
rect 402 1869 409 1880
rect 461 1910 468 1921
rect 802 1921 868 1922
rect 802 1910 809 1921
rect 461 1880 809 1910
rect 461 1869 468 1880
rect 402 1868 468 1869
rect 802 1869 809 1880
rect 861 1910 868 1921
rect 1202 1921 1268 1922
rect 1202 1910 1209 1921
rect 861 1880 1209 1910
rect 861 1869 868 1880
rect 802 1868 868 1869
rect 1202 1869 1209 1880
rect 1261 1910 1268 1921
rect 1602 1921 1668 1922
rect 1602 1910 1609 1921
rect 1261 1880 1609 1910
rect 1261 1869 1268 1880
rect 1202 1868 1268 1869
rect 1602 1869 1609 1880
rect 1661 1910 1668 1921
rect 2002 1921 2068 1922
rect 2002 1910 2009 1921
rect 1661 1880 2009 1910
rect 1661 1869 1668 1880
rect 1602 1868 1668 1869
rect 2002 1869 2009 1880
rect 2061 1910 2068 1921
rect 2402 1921 2468 1922
rect 2402 1910 2409 1921
rect 2061 1880 2409 1910
rect 2061 1869 2068 1880
rect 2002 1868 2068 1869
rect 2402 1869 2409 1880
rect 2461 1910 2468 1921
rect 2802 1921 2868 1922
rect 2802 1910 2809 1921
rect 2461 1880 2809 1910
rect 2461 1869 2468 1880
rect 2402 1868 2468 1869
rect 2802 1869 2809 1880
rect 2861 1910 2868 1921
rect 3202 1921 3268 1922
rect 3202 1910 3209 1921
rect 2861 1880 3209 1910
rect 2861 1869 2868 1880
rect 2802 1868 2868 1869
rect 3202 1869 3209 1880
rect 3261 1910 3268 1921
rect 3602 1921 3668 1922
rect 3602 1910 3609 1921
rect 3261 1880 3609 1910
rect 3261 1869 3268 1880
rect 3202 1868 3268 1869
rect 3602 1869 3609 1880
rect 3661 1910 3668 1921
rect 4002 1921 4068 1922
rect 4002 1910 4009 1921
rect 3661 1880 4009 1910
rect 3661 1869 3668 1880
rect 3602 1868 3668 1869
rect 4002 1869 4009 1880
rect 4061 1910 4068 1921
rect 4402 1921 4468 1922
rect 4402 1910 4409 1921
rect 4061 1880 4409 1910
rect 4061 1869 4068 1880
rect 4002 1868 4068 1869
rect 4402 1869 4409 1880
rect 4461 1910 4468 1921
rect 4802 1921 4868 1922
rect 4802 1910 4809 1921
rect 4461 1880 4809 1910
rect 4461 1869 4468 1880
rect 4402 1868 4468 1869
rect 4802 1869 4809 1880
rect 4861 1910 4868 1921
rect 5202 1921 5268 1922
rect 5202 1910 5209 1921
rect 4861 1880 5209 1910
rect 4861 1869 4868 1880
rect 4802 1868 4868 1869
rect 5202 1869 5209 1880
rect 5261 1910 5268 1921
rect 5602 1921 5668 1922
rect 5602 1910 5609 1921
rect 5261 1880 5609 1910
rect 5261 1869 5268 1880
rect 5202 1868 5268 1869
rect 5602 1869 5609 1880
rect 5661 1910 5668 1921
rect 6002 1921 6068 1922
rect 6002 1910 6009 1921
rect 5661 1880 6009 1910
rect 5661 1869 5668 1880
rect 5602 1868 5668 1869
rect 6002 1869 6009 1880
rect 6061 1910 6068 1921
rect 6402 1921 6468 1922
rect 6402 1910 6409 1921
rect 6061 1880 6409 1910
rect 6061 1869 6068 1880
rect 6002 1868 6068 1869
rect 6402 1869 6409 1880
rect 6461 1910 6468 1921
rect 6802 1921 6868 1922
rect 6802 1910 6809 1921
rect 6461 1880 6809 1910
rect 6461 1869 6468 1880
rect 6402 1868 6468 1869
rect 6802 1869 6809 1880
rect 6861 1910 6868 1921
rect 7202 1921 7268 1922
rect 7202 1910 7209 1921
rect 6861 1880 7209 1910
rect 6861 1869 6868 1880
rect 6802 1868 6868 1869
rect 7202 1869 7209 1880
rect 7261 1910 7268 1921
rect 7602 1921 7668 1922
rect 7602 1910 7609 1921
rect 7261 1880 7609 1910
rect 7261 1869 7268 1880
rect 7202 1868 7268 1869
rect 7602 1869 7609 1880
rect 7661 1910 7668 1921
rect 8002 1921 8068 1922
rect 8002 1910 8009 1921
rect 7661 1880 8009 1910
rect 7661 1869 7668 1880
rect 7602 1868 7668 1869
rect 8002 1869 8009 1880
rect 8061 1910 8068 1921
rect 8402 1921 8468 1922
rect 8402 1910 8409 1921
rect 8061 1880 8409 1910
rect 8061 1869 8068 1880
rect 8002 1868 8068 1869
rect 8402 1869 8409 1880
rect 8461 1910 8468 1921
rect 8802 1921 8868 1922
rect 8802 1910 8809 1921
rect 8461 1880 8809 1910
rect 8461 1869 8468 1880
rect 8402 1868 8468 1869
rect 8802 1869 8809 1880
rect 8861 1910 8868 1921
rect 9202 1921 9268 1922
rect 9202 1910 9209 1921
rect 8861 1880 9209 1910
rect 8861 1869 8868 1880
rect 8802 1868 8868 1869
rect 9202 1869 9209 1880
rect 9261 1910 9268 1921
rect 9602 1921 9668 1922
rect 9602 1910 9609 1921
rect 9261 1880 9609 1910
rect 9261 1869 9268 1880
rect 9202 1868 9268 1869
rect 9602 1869 9609 1880
rect 9661 1910 9668 1921
rect 10002 1921 10068 1922
rect 10002 1910 10009 1921
rect 9661 1880 10009 1910
rect 9661 1869 9668 1880
rect 9602 1868 9668 1869
rect 10002 1869 10009 1880
rect 10061 1910 10068 1921
rect 10402 1921 10468 1922
rect 10402 1910 10409 1921
rect 10061 1880 10409 1910
rect 10061 1869 10068 1880
rect 10002 1868 10068 1869
rect 10402 1869 10409 1880
rect 10461 1910 10468 1921
rect 10802 1921 10868 1922
rect 10802 1910 10809 1921
rect 10461 1880 10809 1910
rect 10461 1869 10468 1880
rect 10402 1868 10468 1869
rect 10802 1869 10809 1880
rect 10861 1910 10868 1921
rect 11202 1921 11268 1922
rect 11202 1910 11209 1921
rect 10861 1880 11209 1910
rect 10861 1869 10868 1880
rect 10802 1868 10868 1869
rect 11202 1869 11209 1880
rect 11261 1910 11268 1921
rect 11602 1921 11668 1922
rect 11602 1910 11609 1921
rect 11261 1880 11609 1910
rect 11261 1869 11268 1880
rect 11202 1868 11268 1869
rect 11602 1869 11609 1880
rect 11661 1910 11668 1921
rect 12002 1921 12068 1922
rect 12002 1910 12009 1921
rect 11661 1880 12009 1910
rect 11661 1869 11668 1880
rect 11602 1868 11668 1869
rect 12002 1869 12009 1880
rect 12061 1910 12068 1921
rect 12402 1921 12468 1922
rect 12402 1910 12409 1921
rect 12061 1880 12409 1910
rect 12061 1869 12068 1880
rect 12002 1868 12068 1869
rect 12402 1869 12409 1880
rect 12461 1910 12468 1921
rect 12802 1921 12868 1922
rect 12802 1910 12809 1921
rect 12461 1880 12809 1910
rect 12461 1869 12468 1880
rect 12402 1868 12468 1869
rect 12802 1869 12809 1880
rect 12861 1910 12868 1921
rect 12900 1921 12966 1922
rect 12900 1910 12907 1921
rect 12861 1880 12907 1910
rect 12861 1869 12868 1880
rect 12802 1868 12868 1869
rect 12900 1869 12907 1880
rect 12959 1869 12966 1921
rect 12900 1868 12966 1869
rect 202 1851 268 1852
rect 202 1840 209 1851
rect 0 1810 209 1840
rect 202 1799 209 1810
rect 261 1840 268 1851
rect 602 1851 668 1852
rect 602 1840 609 1851
rect 261 1810 609 1840
rect 261 1799 268 1810
rect 202 1798 268 1799
rect 602 1799 609 1810
rect 661 1840 668 1851
rect 1002 1851 1068 1852
rect 1002 1840 1009 1851
rect 661 1810 1009 1840
rect 661 1799 668 1810
rect 602 1798 668 1799
rect 1002 1799 1009 1810
rect 1061 1840 1068 1851
rect 1402 1851 1468 1852
rect 1402 1840 1409 1851
rect 1061 1810 1409 1840
rect 1061 1799 1068 1810
rect 1002 1798 1068 1799
rect 1402 1799 1409 1810
rect 1461 1840 1468 1851
rect 1802 1851 1868 1852
rect 1802 1840 1809 1851
rect 1461 1810 1809 1840
rect 1461 1799 1468 1810
rect 1402 1798 1468 1799
rect 1802 1799 1809 1810
rect 1861 1840 1868 1851
rect 2202 1851 2268 1852
rect 2202 1840 2209 1851
rect 1861 1810 2209 1840
rect 1861 1799 1868 1810
rect 1802 1798 1868 1799
rect 2202 1799 2209 1810
rect 2261 1840 2268 1851
rect 2602 1851 2668 1852
rect 2602 1840 2609 1851
rect 2261 1810 2609 1840
rect 2261 1799 2268 1810
rect 2202 1798 2268 1799
rect 2602 1799 2609 1810
rect 2661 1840 2668 1851
rect 3002 1851 3068 1852
rect 3002 1840 3009 1851
rect 2661 1810 3009 1840
rect 2661 1799 2668 1810
rect 2602 1798 2668 1799
rect 3002 1799 3009 1810
rect 3061 1840 3068 1851
rect 3402 1851 3468 1852
rect 3402 1840 3409 1851
rect 3061 1810 3409 1840
rect 3061 1799 3068 1810
rect 3002 1798 3068 1799
rect 3402 1799 3409 1810
rect 3461 1840 3468 1851
rect 3802 1851 3868 1852
rect 3802 1840 3809 1851
rect 3461 1810 3809 1840
rect 3461 1799 3468 1810
rect 3402 1798 3468 1799
rect 3802 1799 3809 1810
rect 3861 1840 3868 1851
rect 4202 1851 4268 1852
rect 4202 1840 4209 1851
rect 3861 1810 4209 1840
rect 3861 1799 3868 1810
rect 3802 1798 3868 1799
rect 4202 1799 4209 1810
rect 4261 1840 4268 1851
rect 4602 1851 4668 1852
rect 4602 1840 4609 1851
rect 4261 1810 4609 1840
rect 4261 1799 4268 1810
rect 4202 1798 4268 1799
rect 4602 1799 4609 1810
rect 4661 1840 4668 1851
rect 5002 1851 5068 1852
rect 5002 1840 5009 1851
rect 4661 1810 5009 1840
rect 4661 1799 4668 1810
rect 4602 1798 4668 1799
rect 5002 1799 5009 1810
rect 5061 1840 5068 1851
rect 5402 1851 5468 1852
rect 5402 1840 5409 1851
rect 5061 1810 5409 1840
rect 5061 1799 5068 1810
rect 5002 1798 5068 1799
rect 5402 1799 5409 1810
rect 5461 1840 5468 1851
rect 5802 1851 5868 1852
rect 5802 1840 5809 1851
rect 5461 1810 5809 1840
rect 5461 1799 5468 1810
rect 5402 1798 5468 1799
rect 5802 1799 5809 1810
rect 5861 1840 5868 1851
rect 6202 1851 6268 1852
rect 6202 1840 6209 1851
rect 5861 1810 6209 1840
rect 5861 1799 5868 1810
rect 5802 1798 5868 1799
rect 6202 1799 6209 1810
rect 6261 1840 6268 1851
rect 6602 1851 6668 1852
rect 6602 1840 6609 1851
rect 6261 1810 6609 1840
rect 6261 1799 6268 1810
rect 6202 1798 6268 1799
rect 6602 1799 6609 1810
rect 6661 1840 6668 1851
rect 7002 1851 7068 1852
rect 7002 1840 7009 1851
rect 6661 1810 7009 1840
rect 6661 1799 6668 1810
rect 6602 1798 6668 1799
rect 7002 1799 7009 1810
rect 7061 1840 7068 1851
rect 7402 1851 7468 1852
rect 7402 1840 7409 1851
rect 7061 1810 7409 1840
rect 7061 1799 7068 1810
rect 7002 1798 7068 1799
rect 7402 1799 7409 1810
rect 7461 1840 7468 1851
rect 7802 1851 7868 1852
rect 7802 1840 7809 1851
rect 7461 1810 7809 1840
rect 7461 1799 7468 1810
rect 7402 1798 7468 1799
rect 7802 1799 7809 1810
rect 7861 1840 7868 1851
rect 8202 1851 8268 1852
rect 8202 1840 8209 1851
rect 7861 1810 8209 1840
rect 7861 1799 7868 1810
rect 7802 1798 7868 1799
rect 8202 1799 8209 1810
rect 8261 1840 8268 1851
rect 8602 1851 8668 1852
rect 8602 1840 8609 1851
rect 8261 1810 8609 1840
rect 8261 1799 8268 1810
rect 8202 1798 8268 1799
rect 8602 1799 8609 1810
rect 8661 1840 8668 1851
rect 9002 1851 9068 1852
rect 9002 1840 9009 1851
rect 8661 1810 9009 1840
rect 8661 1799 8668 1810
rect 8602 1798 8668 1799
rect 9002 1799 9009 1810
rect 9061 1840 9068 1851
rect 9402 1851 9468 1852
rect 9402 1840 9409 1851
rect 9061 1810 9409 1840
rect 9061 1799 9068 1810
rect 9002 1798 9068 1799
rect 9402 1799 9409 1810
rect 9461 1840 9468 1851
rect 9802 1851 9868 1852
rect 9802 1840 9809 1851
rect 9461 1810 9809 1840
rect 9461 1799 9468 1810
rect 9402 1798 9468 1799
rect 9802 1799 9809 1810
rect 9861 1840 9868 1851
rect 10202 1851 10268 1852
rect 10202 1840 10209 1851
rect 9861 1810 10209 1840
rect 9861 1799 9868 1810
rect 9802 1798 9868 1799
rect 10202 1799 10209 1810
rect 10261 1840 10268 1851
rect 10602 1851 10668 1852
rect 10602 1840 10609 1851
rect 10261 1810 10609 1840
rect 10261 1799 10268 1810
rect 10202 1798 10268 1799
rect 10602 1799 10609 1810
rect 10661 1840 10668 1851
rect 11002 1851 11068 1852
rect 11002 1840 11009 1851
rect 10661 1810 11009 1840
rect 10661 1799 10668 1810
rect 10602 1798 10668 1799
rect 11002 1799 11009 1810
rect 11061 1840 11068 1851
rect 11402 1851 11468 1852
rect 11402 1840 11409 1851
rect 11061 1810 11409 1840
rect 11061 1799 11068 1810
rect 11002 1798 11068 1799
rect 11402 1799 11409 1810
rect 11461 1840 11468 1851
rect 11802 1851 11868 1852
rect 11802 1840 11809 1851
rect 11461 1810 11809 1840
rect 11461 1799 11468 1810
rect 11402 1798 11468 1799
rect 11802 1799 11809 1810
rect 11861 1840 11868 1851
rect 12202 1851 12268 1852
rect 12202 1840 12209 1851
rect 11861 1810 12209 1840
rect 11861 1799 11868 1810
rect 11802 1798 11868 1799
rect 12202 1799 12209 1810
rect 12261 1840 12268 1851
rect 12602 1851 12668 1852
rect 12602 1840 12609 1851
rect 12261 1810 12609 1840
rect 12261 1799 12268 1810
rect 12202 1798 12268 1799
rect 12602 1799 12609 1810
rect 12661 1840 12668 1851
rect 13104 1851 13170 1852
rect 13104 1840 13111 1851
rect 12661 1810 13111 1840
rect 12661 1799 12668 1810
rect 12602 1798 12668 1799
rect 13104 1799 13111 1810
rect 13163 1799 13170 1851
rect 13104 1798 13170 1799
rect 2 1781 68 1782
rect 2 1770 9 1781
rect 0 1740 9 1770
rect 2 1729 9 1740
rect 61 1770 68 1781
rect 402 1781 468 1782
rect 402 1770 409 1781
rect 61 1740 409 1770
rect 61 1729 68 1740
rect 2 1728 68 1729
rect 402 1729 409 1740
rect 461 1770 468 1781
rect 802 1781 868 1782
rect 802 1770 809 1781
rect 461 1740 809 1770
rect 461 1729 468 1740
rect 402 1728 468 1729
rect 802 1729 809 1740
rect 861 1770 868 1781
rect 1202 1781 1268 1782
rect 1202 1770 1209 1781
rect 861 1740 1209 1770
rect 861 1729 868 1740
rect 802 1728 868 1729
rect 1202 1729 1209 1740
rect 1261 1770 1268 1781
rect 1602 1781 1668 1782
rect 1602 1770 1609 1781
rect 1261 1740 1609 1770
rect 1261 1729 1268 1740
rect 1202 1728 1268 1729
rect 1602 1729 1609 1740
rect 1661 1770 1668 1781
rect 2002 1781 2068 1782
rect 2002 1770 2009 1781
rect 1661 1740 2009 1770
rect 1661 1729 1668 1740
rect 1602 1728 1668 1729
rect 2002 1729 2009 1740
rect 2061 1770 2068 1781
rect 2402 1781 2468 1782
rect 2402 1770 2409 1781
rect 2061 1740 2409 1770
rect 2061 1729 2068 1740
rect 2002 1728 2068 1729
rect 2402 1729 2409 1740
rect 2461 1770 2468 1781
rect 2802 1781 2868 1782
rect 2802 1770 2809 1781
rect 2461 1740 2809 1770
rect 2461 1729 2468 1740
rect 2402 1728 2468 1729
rect 2802 1729 2809 1740
rect 2861 1770 2868 1781
rect 3202 1781 3268 1782
rect 3202 1770 3209 1781
rect 2861 1740 3209 1770
rect 2861 1729 2868 1740
rect 2802 1728 2868 1729
rect 3202 1729 3209 1740
rect 3261 1770 3268 1781
rect 3602 1781 3668 1782
rect 3602 1770 3609 1781
rect 3261 1740 3609 1770
rect 3261 1729 3268 1740
rect 3202 1728 3268 1729
rect 3602 1729 3609 1740
rect 3661 1770 3668 1781
rect 4002 1781 4068 1782
rect 4002 1770 4009 1781
rect 3661 1740 4009 1770
rect 3661 1729 3668 1740
rect 3602 1728 3668 1729
rect 4002 1729 4009 1740
rect 4061 1770 4068 1781
rect 4402 1781 4468 1782
rect 4402 1770 4409 1781
rect 4061 1740 4409 1770
rect 4061 1729 4068 1740
rect 4002 1728 4068 1729
rect 4402 1729 4409 1740
rect 4461 1770 4468 1781
rect 4802 1781 4868 1782
rect 4802 1770 4809 1781
rect 4461 1740 4809 1770
rect 4461 1729 4468 1740
rect 4402 1728 4468 1729
rect 4802 1729 4809 1740
rect 4861 1770 4868 1781
rect 5202 1781 5268 1782
rect 5202 1770 5209 1781
rect 4861 1740 5209 1770
rect 4861 1729 4868 1740
rect 4802 1728 4868 1729
rect 5202 1729 5209 1740
rect 5261 1770 5268 1781
rect 5602 1781 5668 1782
rect 5602 1770 5609 1781
rect 5261 1740 5609 1770
rect 5261 1729 5268 1740
rect 5202 1728 5268 1729
rect 5602 1729 5609 1740
rect 5661 1770 5668 1781
rect 6002 1781 6068 1782
rect 6002 1770 6009 1781
rect 5661 1740 6009 1770
rect 5661 1729 5668 1740
rect 5602 1728 5668 1729
rect 6002 1729 6009 1740
rect 6061 1770 6068 1781
rect 6402 1781 6468 1782
rect 6402 1770 6409 1781
rect 6061 1740 6409 1770
rect 6061 1729 6068 1740
rect 6002 1728 6068 1729
rect 6402 1729 6409 1740
rect 6461 1770 6468 1781
rect 6802 1781 6868 1782
rect 6802 1770 6809 1781
rect 6461 1740 6809 1770
rect 6461 1729 6468 1740
rect 6402 1728 6468 1729
rect 6802 1729 6809 1740
rect 6861 1770 6868 1781
rect 7202 1781 7268 1782
rect 7202 1770 7209 1781
rect 6861 1740 7209 1770
rect 6861 1729 6868 1740
rect 6802 1728 6868 1729
rect 7202 1729 7209 1740
rect 7261 1770 7268 1781
rect 7602 1781 7668 1782
rect 7602 1770 7609 1781
rect 7261 1740 7609 1770
rect 7261 1729 7268 1740
rect 7202 1728 7268 1729
rect 7602 1729 7609 1740
rect 7661 1770 7668 1781
rect 8002 1781 8068 1782
rect 8002 1770 8009 1781
rect 7661 1740 8009 1770
rect 7661 1729 7668 1740
rect 7602 1728 7668 1729
rect 8002 1729 8009 1740
rect 8061 1770 8068 1781
rect 8402 1781 8468 1782
rect 8402 1770 8409 1781
rect 8061 1740 8409 1770
rect 8061 1729 8068 1740
rect 8002 1728 8068 1729
rect 8402 1729 8409 1740
rect 8461 1770 8468 1781
rect 8802 1781 8868 1782
rect 8802 1770 8809 1781
rect 8461 1740 8809 1770
rect 8461 1729 8468 1740
rect 8402 1728 8468 1729
rect 8802 1729 8809 1740
rect 8861 1770 8868 1781
rect 9202 1781 9268 1782
rect 9202 1770 9209 1781
rect 8861 1740 9209 1770
rect 8861 1729 8868 1740
rect 8802 1728 8868 1729
rect 9202 1729 9209 1740
rect 9261 1770 9268 1781
rect 9602 1781 9668 1782
rect 9602 1770 9609 1781
rect 9261 1740 9609 1770
rect 9261 1729 9268 1740
rect 9202 1728 9268 1729
rect 9602 1729 9609 1740
rect 9661 1770 9668 1781
rect 10002 1781 10068 1782
rect 10002 1770 10009 1781
rect 9661 1740 10009 1770
rect 9661 1729 9668 1740
rect 9602 1728 9668 1729
rect 10002 1729 10009 1740
rect 10061 1770 10068 1781
rect 10402 1781 10468 1782
rect 10402 1770 10409 1781
rect 10061 1740 10409 1770
rect 10061 1729 10068 1740
rect 10002 1728 10068 1729
rect 10402 1729 10409 1740
rect 10461 1770 10468 1781
rect 10802 1781 10868 1782
rect 10802 1770 10809 1781
rect 10461 1740 10809 1770
rect 10461 1729 10468 1740
rect 10402 1728 10468 1729
rect 10802 1729 10809 1740
rect 10861 1770 10868 1781
rect 11202 1781 11268 1782
rect 11202 1770 11209 1781
rect 10861 1740 11209 1770
rect 10861 1729 10868 1740
rect 10802 1728 10868 1729
rect 11202 1729 11209 1740
rect 11261 1770 11268 1781
rect 11602 1781 11668 1782
rect 11602 1770 11609 1781
rect 11261 1740 11609 1770
rect 11261 1729 11268 1740
rect 11202 1728 11268 1729
rect 11602 1729 11609 1740
rect 11661 1770 11668 1781
rect 12002 1781 12068 1782
rect 12002 1770 12009 1781
rect 11661 1740 12009 1770
rect 11661 1729 11668 1740
rect 11602 1728 11668 1729
rect 12002 1729 12009 1740
rect 12061 1770 12068 1781
rect 12402 1781 12468 1782
rect 12402 1770 12409 1781
rect 12061 1740 12409 1770
rect 12061 1729 12068 1740
rect 12002 1728 12068 1729
rect 12402 1729 12409 1740
rect 12461 1770 12468 1781
rect 12802 1781 12868 1782
rect 12802 1770 12809 1781
rect 12461 1740 12809 1770
rect 12461 1729 12468 1740
rect 12402 1728 12468 1729
rect 12802 1729 12809 1740
rect 12861 1770 12868 1781
rect 12900 1781 12966 1782
rect 12900 1770 12907 1781
rect 12861 1740 12907 1770
rect 12861 1729 12868 1740
rect 12802 1728 12868 1729
rect 12900 1729 12907 1740
rect 12959 1729 12966 1781
rect 12900 1728 12966 1729
rect 202 1711 268 1712
rect 202 1700 209 1711
rect 0 1670 209 1700
rect 202 1659 209 1670
rect 261 1700 268 1711
rect 602 1711 668 1712
rect 602 1700 609 1711
rect 261 1670 609 1700
rect 261 1659 268 1670
rect 202 1658 268 1659
rect 602 1659 609 1670
rect 661 1700 668 1711
rect 1002 1711 1068 1712
rect 1002 1700 1009 1711
rect 661 1670 1009 1700
rect 661 1659 668 1670
rect 602 1658 668 1659
rect 1002 1659 1009 1670
rect 1061 1700 1068 1711
rect 1402 1711 1468 1712
rect 1402 1700 1409 1711
rect 1061 1670 1409 1700
rect 1061 1659 1068 1670
rect 1002 1658 1068 1659
rect 1402 1659 1409 1670
rect 1461 1700 1468 1711
rect 1802 1711 1868 1712
rect 1802 1700 1809 1711
rect 1461 1670 1809 1700
rect 1461 1659 1468 1670
rect 1402 1658 1468 1659
rect 1802 1659 1809 1670
rect 1861 1700 1868 1711
rect 2202 1711 2268 1712
rect 2202 1700 2209 1711
rect 1861 1670 2209 1700
rect 1861 1659 1868 1670
rect 1802 1658 1868 1659
rect 2202 1659 2209 1670
rect 2261 1700 2268 1711
rect 2602 1711 2668 1712
rect 2602 1700 2609 1711
rect 2261 1670 2609 1700
rect 2261 1659 2268 1670
rect 2202 1658 2268 1659
rect 2602 1659 2609 1670
rect 2661 1700 2668 1711
rect 3002 1711 3068 1712
rect 3002 1700 3009 1711
rect 2661 1670 3009 1700
rect 2661 1659 2668 1670
rect 2602 1658 2668 1659
rect 3002 1659 3009 1670
rect 3061 1700 3068 1711
rect 3402 1711 3468 1712
rect 3402 1700 3409 1711
rect 3061 1670 3409 1700
rect 3061 1659 3068 1670
rect 3002 1658 3068 1659
rect 3402 1659 3409 1670
rect 3461 1700 3468 1711
rect 3802 1711 3868 1712
rect 3802 1700 3809 1711
rect 3461 1670 3809 1700
rect 3461 1659 3468 1670
rect 3402 1658 3468 1659
rect 3802 1659 3809 1670
rect 3861 1700 3868 1711
rect 4202 1711 4268 1712
rect 4202 1700 4209 1711
rect 3861 1670 4209 1700
rect 3861 1659 3868 1670
rect 3802 1658 3868 1659
rect 4202 1659 4209 1670
rect 4261 1700 4268 1711
rect 4602 1711 4668 1712
rect 4602 1700 4609 1711
rect 4261 1670 4609 1700
rect 4261 1659 4268 1670
rect 4202 1658 4268 1659
rect 4602 1659 4609 1670
rect 4661 1700 4668 1711
rect 5002 1711 5068 1712
rect 5002 1700 5009 1711
rect 4661 1670 5009 1700
rect 4661 1659 4668 1670
rect 4602 1658 4668 1659
rect 5002 1659 5009 1670
rect 5061 1700 5068 1711
rect 5402 1711 5468 1712
rect 5402 1700 5409 1711
rect 5061 1670 5409 1700
rect 5061 1659 5068 1670
rect 5002 1658 5068 1659
rect 5402 1659 5409 1670
rect 5461 1700 5468 1711
rect 5802 1711 5868 1712
rect 5802 1700 5809 1711
rect 5461 1670 5809 1700
rect 5461 1659 5468 1670
rect 5402 1658 5468 1659
rect 5802 1659 5809 1670
rect 5861 1700 5868 1711
rect 6202 1711 6268 1712
rect 6202 1700 6209 1711
rect 5861 1670 6209 1700
rect 5861 1659 5868 1670
rect 5802 1658 5868 1659
rect 6202 1659 6209 1670
rect 6261 1700 6268 1711
rect 6602 1711 6668 1712
rect 6602 1700 6609 1711
rect 6261 1670 6609 1700
rect 6261 1659 6268 1670
rect 6202 1658 6268 1659
rect 6602 1659 6609 1670
rect 6661 1700 6668 1711
rect 7002 1711 7068 1712
rect 7002 1700 7009 1711
rect 6661 1670 7009 1700
rect 6661 1659 6668 1670
rect 6602 1658 6668 1659
rect 7002 1659 7009 1670
rect 7061 1700 7068 1711
rect 7402 1711 7468 1712
rect 7402 1700 7409 1711
rect 7061 1670 7409 1700
rect 7061 1659 7068 1670
rect 7002 1658 7068 1659
rect 7402 1659 7409 1670
rect 7461 1700 7468 1711
rect 7802 1711 7868 1712
rect 7802 1700 7809 1711
rect 7461 1670 7809 1700
rect 7461 1659 7468 1670
rect 7402 1658 7468 1659
rect 7802 1659 7809 1670
rect 7861 1700 7868 1711
rect 8202 1711 8268 1712
rect 8202 1700 8209 1711
rect 7861 1670 8209 1700
rect 7861 1659 7868 1670
rect 7802 1658 7868 1659
rect 8202 1659 8209 1670
rect 8261 1700 8268 1711
rect 8602 1711 8668 1712
rect 8602 1700 8609 1711
rect 8261 1670 8609 1700
rect 8261 1659 8268 1670
rect 8202 1658 8268 1659
rect 8602 1659 8609 1670
rect 8661 1700 8668 1711
rect 9002 1711 9068 1712
rect 9002 1700 9009 1711
rect 8661 1670 9009 1700
rect 8661 1659 8668 1670
rect 8602 1658 8668 1659
rect 9002 1659 9009 1670
rect 9061 1700 9068 1711
rect 9402 1711 9468 1712
rect 9402 1700 9409 1711
rect 9061 1670 9409 1700
rect 9061 1659 9068 1670
rect 9002 1658 9068 1659
rect 9402 1659 9409 1670
rect 9461 1700 9468 1711
rect 9802 1711 9868 1712
rect 9802 1700 9809 1711
rect 9461 1670 9809 1700
rect 9461 1659 9468 1670
rect 9402 1658 9468 1659
rect 9802 1659 9809 1670
rect 9861 1700 9868 1711
rect 10202 1711 10268 1712
rect 10202 1700 10209 1711
rect 9861 1670 10209 1700
rect 9861 1659 9868 1670
rect 9802 1658 9868 1659
rect 10202 1659 10209 1670
rect 10261 1700 10268 1711
rect 10602 1711 10668 1712
rect 10602 1700 10609 1711
rect 10261 1670 10609 1700
rect 10261 1659 10268 1670
rect 10202 1658 10268 1659
rect 10602 1659 10609 1670
rect 10661 1700 10668 1711
rect 11002 1711 11068 1712
rect 11002 1700 11009 1711
rect 10661 1670 11009 1700
rect 10661 1659 10668 1670
rect 10602 1658 10668 1659
rect 11002 1659 11009 1670
rect 11061 1700 11068 1711
rect 11402 1711 11468 1712
rect 11402 1700 11409 1711
rect 11061 1670 11409 1700
rect 11061 1659 11068 1670
rect 11002 1658 11068 1659
rect 11402 1659 11409 1670
rect 11461 1700 11468 1711
rect 11802 1711 11868 1712
rect 11802 1700 11809 1711
rect 11461 1670 11809 1700
rect 11461 1659 11468 1670
rect 11402 1658 11468 1659
rect 11802 1659 11809 1670
rect 11861 1700 11868 1711
rect 12202 1711 12268 1712
rect 12202 1700 12209 1711
rect 11861 1670 12209 1700
rect 11861 1659 11868 1670
rect 11802 1658 11868 1659
rect 12202 1659 12209 1670
rect 12261 1700 12268 1711
rect 12602 1711 12668 1712
rect 12602 1700 12609 1711
rect 12261 1670 12609 1700
rect 12261 1659 12268 1670
rect 12202 1658 12268 1659
rect 12602 1659 12609 1670
rect 12661 1700 12668 1711
rect 13104 1711 13170 1712
rect 13104 1700 13111 1711
rect 12661 1670 13111 1700
rect 12661 1659 12668 1670
rect 12602 1658 12668 1659
rect 13104 1659 13111 1670
rect 13163 1659 13170 1711
rect 13104 1658 13170 1659
rect 2 1641 68 1642
rect 2 1630 9 1641
rect 0 1600 9 1630
rect 2 1589 9 1600
rect 61 1630 68 1641
rect 402 1641 468 1642
rect 402 1630 409 1641
rect 61 1600 409 1630
rect 61 1589 68 1600
rect 2 1588 68 1589
rect 402 1589 409 1600
rect 461 1630 468 1641
rect 802 1641 868 1642
rect 802 1630 809 1641
rect 461 1600 809 1630
rect 461 1589 468 1600
rect 402 1588 468 1589
rect 802 1589 809 1600
rect 861 1630 868 1641
rect 1202 1641 1268 1642
rect 1202 1630 1209 1641
rect 861 1600 1209 1630
rect 861 1589 868 1600
rect 802 1588 868 1589
rect 1202 1589 1209 1600
rect 1261 1630 1268 1641
rect 1602 1641 1668 1642
rect 1602 1630 1609 1641
rect 1261 1600 1609 1630
rect 1261 1589 1268 1600
rect 1202 1588 1268 1589
rect 1602 1589 1609 1600
rect 1661 1630 1668 1641
rect 2002 1641 2068 1642
rect 2002 1630 2009 1641
rect 1661 1600 2009 1630
rect 1661 1589 1668 1600
rect 1602 1588 1668 1589
rect 2002 1589 2009 1600
rect 2061 1630 2068 1641
rect 2402 1641 2468 1642
rect 2402 1630 2409 1641
rect 2061 1600 2409 1630
rect 2061 1589 2068 1600
rect 2002 1588 2068 1589
rect 2402 1589 2409 1600
rect 2461 1630 2468 1641
rect 2802 1641 2868 1642
rect 2802 1630 2809 1641
rect 2461 1600 2809 1630
rect 2461 1589 2468 1600
rect 2402 1588 2468 1589
rect 2802 1589 2809 1600
rect 2861 1630 2868 1641
rect 3202 1641 3268 1642
rect 3202 1630 3209 1641
rect 2861 1600 3209 1630
rect 2861 1589 2868 1600
rect 2802 1588 2868 1589
rect 3202 1589 3209 1600
rect 3261 1630 3268 1641
rect 3602 1641 3668 1642
rect 3602 1630 3609 1641
rect 3261 1600 3609 1630
rect 3261 1589 3268 1600
rect 3202 1588 3268 1589
rect 3602 1589 3609 1600
rect 3661 1630 3668 1641
rect 4002 1641 4068 1642
rect 4002 1630 4009 1641
rect 3661 1600 4009 1630
rect 3661 1589 3668 1600
rect 3602 1588 3668 1589
rect 4002 1589 4009 1600
rect 4061 1630 4068 1641
rect 4402 1641 4468 1642
rect 4402 1630 4409 1641
rect 4061 1600 4409 1630
rect 4061 1589 4068 1600
rect 4002 1588 4068 1589
rect 4402 1589 4409 1600
rect 4461 1630 4468 1641
rect 4802 1641 4868 1642
rect 4802 1630 4809 1641
rect 4461 1600 4809 1630
rect 4461 1589 4468 1600
rect 4402 1588 4468 1589
rect 4802 1589 4809 1600
rect 4861 1630 4868 1641
rect 5202 1641 5268 1642
rect 5202 1630 5209 1641
rect 4861 1600 5209 1630
rect 4861 1589 4868 1600
rect 4802 1588 4868 1589
rect 5202 1589 5209 1600
rect 5261 1630 5268 1641
rect 5602 1641 5668 1642
rect 5602 1630 5609 1641
rect 5261 1600 5609 1630
rect 5261 1589 5268 1600
rect 5202 1588 5268 1589
rect 5602 1589 5609 1600
rect 5661 1630 5668 1641
rect 6002 1641 6068 1642
rect 6002 1630 6009 1641
rect 5661 1600 6009 1630
rect 5661 1589 5668 1600
rect 5602 1588 5668 1589
rect 6002 1589 6009 1600
rect 6061 1630 6068 1641
rect 6402 1641 6468 1642
rect 6402 1630 6409 1641
rect 6061 1600 6409 1630
rect 6061 1589 6068 1600
rect 6002 1588 6068 1589
rect 6402 1589 6409 1600
rect 6461 1630 6468 1641
rect 6802 1641 6868 1642
rect 6802 1630 6809 1641
rect 6461 1600 6809 1630
rect 6461 1589 6468 1600
rect 6402 1588 6468 1589
rect 6802 1589 6809 1600
rect 6861 1630 6868 1641
rect 7202 1641 7268 1642
rect 7202 1630 7209 1641
rect 6861 1600 7209 1630
rect 6861 1589 6868 1600
rect 6802 1588 6868 1589
rect 7202 1589 7209 1600
rect 7261 1630 7268 1641
rect 7602 1641 7668 1642
rect 7602 1630 7609 1641
rect 7261 1600 7609 1630
rect 7261 1589 7268 1600
rect 7202 1588 7268 1589
rect 7602 1589 7609 1600
rect 7661 1630 7668 1641
rect 8002 1641 8068 1642
rect 8002 1630 8009 1641
rect 7661 1600 8009 1630
rect 7661 1589 7668 1600
rect 7602 1588 7668 1589
rect 8002 1589 8009 1600
rect 8061 1630 8068 1641
rect 8402 1641 8468 1642
rect 8402 1630 8409 1641
rect 8061 1600 8409 1630
rect 8061 1589 8068 1600
rect 8002 1588 8068 1589
rect 8402 1589 8409 1600
rect 8461 1630 8468 1641
rect 8802 1641 8868 1642
rect 8802 1630 8809 1641
rect 8461 1600 8809 1630
rect 8461 1589 8468 1600
rect 8402 1588 8468 1589
rect 8802 1589 8809 1600
rect 8861 1630 8868 1641
rect 9202 1641 9268 1642
rect 9202 1630 9209 1641
rect 8861 1600 9209 1630
rect 8861 1589 8868 1600
rect 8802 1588 8868 1589
rect 9202 1589 9209 1600
rect 9261 1630 9268 1641
rect 9602 1641 9668 1642
rect 9602 1630 9609 1641
rect 9261 1600 9609 1630
rect 9261 1589 9268 1600
rect 9202 1588 9268 1589
rect 9602 1589 9609 1600
rect 9661 1630 9668 1641
rect 10002 1641 10068 1642
rect 10002 1630 10009 1641
rect 9661 1600 10009 1630
rect 9661 1589 9668 1600
rect 9602 1588 9668 1589
rect 10002 1589 10009 1600
rect 10061 1630 10068 1641
rect 10402 1641 10468 1642
rect 10402 1630 10409 1641
rect 10061 1600 10409 1630
rect 10061 1589 10068 1600
rect 10002 1588 10068 1589
rect 10402 1589 10409 1600
rect 10461 1630 10468 1641
rect 10802 1641 10868 1642
rect 10802 1630 10809 1641
rect 10461 1600 10809 1630
rect 10461 1589 10468 1600
rect 10402 1588 10468 1589
rect 10802 1589 10809 1600
rect 10861 1630 10868 1641
rect 11202 1641 11268 1642
rect 11202 1630 11209 1641
rect 10861 1600 11209 1630
rect 10861 1589 10868 1600
rect 10802 1588 10868 1589
rect 11202 1589 11209 1600
rect 11261 1630 11268 1641
rect 11602 1641 11668 1642
rect 11602 1630 11609 1641
rect 11261 1600 11609 1630
rect 11261 1589 11268 1600
rect 11202 1588 11268 1589
rect 11602 1589 11609 1600
rect 11661 1630 11668 1641
rect 12002 1641 12068 1642
rect 12002 1630 12009 1641
rect 11661 1600 12009 1630
rect 11661 1589 11668 1600
rect 11602 1588 11668 1589
rect 12002 1589 12009 1600
rect 12061 1630 12068 1641
rect 12402 1641 12468 1642
rect 12402 1630 12409 1641
rect 12061 1600 12409 1630
rect 12061 1589 12068 1600
rect 12002 1588 12068 1589
rect 12402 1589 12409 1600
rect 12461 1630 12468 1641
rect 12802 1641 12868 1642
rect 12802 1630 12809 1641
rect 12461 1600 12809 1630
rect 12461 1589 12468 1600
rect 12402 1588 12468 1589
rect 12802 1589 12809 1600
rect 12861 1630 12868 1641
rect 12900 1641 12966 1642
rect 12900 1630 12907 1641
rect 12861 1600 12907 1630
rect 12861 1589 12868 1600
rect 12802 1588 12868 1589
rect 12900 1589 12907 1600
rect 12959 1589 12966 1641
rect 12900 1588 12966 1589
rect 202 1571 268 1572
rect 202 1560 209 1571
rect 0 1530 209 1560
rect 202 1519 209 1530
rect 261 1560 268 1571
rect 602 1571 668 1572
rect 602 1560 609 1571
rect 261 1530 609 1560
rect 261 1519 268 1530
rect 202 1518 268 1519
rect 602 1519 609 1530
rect 661 1560 668 1571
rect 1002 1571 1068 1572
rect 1002 1560 1009 1571
rect 661 1530 1009 1560
rect 661 1519 668 1530
rect 602 1518 668 1519
rect 1002 1519 1009 1530
rect 1061 1560 1068 1571
rect 1402 1571 1468 1572
rect 1402 1560 1409 1571
rect 1061 1530 1409 1560
rect 1061 1519 1068 1530
rect 1002 1518 1068 1519
rect 1402 1519 1409 1530
rect 1461 1560 1468 1571
rect 1802 1571 1868 1572
rect 1802 1560 1809 1571
rect 1461 1530 1809 1560
rect 1461 1519 1468 1530
rect 1402 1518 1468 1519
rect 1802 1519 1809 1530
rect 1861 1560 1868 1571
rect 2202 1571 2268 1572
rect 2202 1560 2209 1571
rect 1861 1530 2209 1560
rect 1861 1519 1868 1530
rect 1802 1518 1868 1519
rect 2202 1519 2209 1530
rect 2261 1560 2268 1571
rect 2602 1571 2668 1572
rect 2602 1560 2609 1571
rect 2261 1530 2609 1560
rect 2261 1519 2268 1530
rect 2202 1518 2268 1519
rect 2602 1519 2609 1530
rect 2661 1560 2668 1571
rect 3002 1571 3068 1572
rect 3002 1560 3009 1571
rect 2661 1530 3009 1560
rect 2661 1519 2668 1530
rect 2602 1518 2668 1519
rect 3002 1519 3009 1530
rect 3061 1560 3068 1571
rect 3402 1571 3468 1572
rect 3402 1560 3409 1571
rect 3061 1530 3409 1560
rect 3061 1519 3068 1530
rect 3002 1518 3068 1519
rect 3402 1519 3409 1530
rect 3461 1560 3468 1571
rect 3802 1571 3868 1572
rect 3802 1560 3809 1571
rect 3461 1530 3809 1560
rect 3461 1519 3468 1530
rect 3402 1518 3468 1519
rect 3802 1519 3809 1530
rect 3861 1560 3868 1571
rect 4202 1571 4268 1572
rect 4202 1560 4209 1571
rect 3861 1530 4209 1560
rect 3861 1519 3868 1530
rect 3802 1518 3868 1519
rect 4202 1519 4209 1530
rect 4261 1560 4268 1571
rect 4602 1571 4668 1572
rect 4602 1560 4609 1571
rect 4261 1530 4609 1560
rect 4261 1519 4268 1530
rect 4202 1518 4268 1519
rect 4602 1519 4609 1530
rect 4661 1560 4668 1571
rect 5002 1571 5068 1572
rect 5002 1560 5009 1571
rect 4661 1530 5009 1560
rect 4661 1519 4668 1530
rect 4602 1518 4668 1519
rect 5002 1519 5009 1530
rect 5061 1560 5068 1571
rect 5402 1571 5468 1572
rect 5402 1560 5409 1571
rect 5061 1530 5409 1560
rect 5061 1519 5068 1530
rect 5002 1518 5068 1519
rect 5402 1519 5409 1530
rect 5461 1560 5468 1571
rect 5802 1571 5868 1572
rect 5802 1560 5809 1571
rect 5461 1530 5809 1560
rect 5461 1519 5468 1530
rect 5402 1518 5468 1519
rect 5802 1519 5809 1530
rect 5861 1560 5868 1571
rect 6202 1571 6268 1572
rect 6202 1560 6209 1571
rect 5861 1530 6209 1560
rect 5861 1519 5868 1530
rect 5802 1518 5868 1519
rect 6202 1519 6209 1530
rect 6261 1560 6268 1571
rect 6602 1571 6668 1572
rect 6602 1560 6609 1571
rect 6261 1530 6609 1560
rect 6261 1519 6268 1530
rect 6202 1518 6268 1519
rect 6602 1519 6609 1530
rect 6661 1560 6668 1571
rect 7002 1571 7068 1572
rect 7002 1560 7009 1571
rect 6661 1530 7009 1560
rect 6661 1519 6668 1530
rect 6602 1518 6668 1519
rect 7002 1519 7009 1530
rect 7061 1560 7068 1571
rect 7402 1571 7468 1572
rect 7402 1560 7409 1571
rect 7061 1530 7409 1560
rect 7061 1519 7068 1530
rect 7002 1518 7068 1519
rect 7402 1519 7409 1530
rect 7461 1560 7468 1571
rect 7802 1571 7868 1572
rect 7802 1560 7809 1571
rect 7461 1530 7809 1560
rect 7461 1519 7468 1530
rect 7402 1518 7468 1519
rect 7802 1519 7809 1530
rect 7861 1560 7868 1571
rect 8202 1571 8268 1572
rect 8202 1560 8209 1571
rect 7861 1530 8209 1560
rect 7861 1519 7868 1530
rect 7802 1518 7868 1519
rect 8202 1519 8209 1530
rect 8261 1560 8268 1571
rect 8602 1571 8668 1572
rect 8602 1560 8609 1571
rect 8261 1530 8609 1560
rect 8261 1519 8268 1530
rect 8202 1518 8268 1519
rect 8602 1519 8609 1530
rect 8661 1560 8668 1571
rect 9002 1571 9068 1572
rect 9002 1560 9009 1571
rect 8661 1530 9009 1560
rect 8661 1519 8668 1530
rect 8602 1518 8668 1519
rect 9002 1519 9009 1530
rect 9061 1560 9068 1571
rect 9402 1571 9468 1572
rect 9402 1560 9409 1571
rect 9061 1530 9409 1560
rect 9061 1519 9068 1530
rect 9002 1518 9068 1519
rect 9402 1519 9409 1530
rect 9461 1560 9468 1571
rect 9802 1571 9868 1572
rect 9802 1560 9809 1571
rect 9461 1530 9809 1560
rect 9461 1519 9468 1530
rect 9402 1518 9468 1519
rect 9802 1519 9809 1530
rect 9861 1560 9868 1571
rect 10202 1571 10268 1572
rect 10202 1560 10209 1571
rect 9861 1530 10209 1560
rect 9861 1519 9868 1530
rect 9802 1518 9868 1519
rect 10202 1519 10209 1530
rect 10261 1560 10268 1571
rect 10602 1571 10668 1572
rect 10602 1560 10609 1571
rect 10261 1530 10609 1560
rect 10261 1519 10268 1530
rect 10202 1518 10268 1519
rect 10602 1519 10609 1530
rect 10661 1560 10668 1571
rect 11002 1571 11068 1572
rect 11002 1560 11009 1571
rect 10661 1530 11009 1560
rect 10661 1519 10668 1530
rect 10602 1518 10668 1519
rect 11002 1519 11009 1530
rect 11061 1560 11068 1571
rect 11402 1571 11468 1572
rect 11402 1560 11409 1571
rect 11061 1530 11409 1560
rect 11061 1519 11068 1530
rect 11002 1518 11068 1519
rect 11402 1519 11409 1530
rect 11461 1560 11468 1571
rect 11802 1571 11868 1572
rect 11802 1560 11809 1571
rect 11461 1530 11809 1560
rect 11461 1519 11468 1530
rect 11402 1518 11468 1519
rect 11802 1519 11809 1530
rect 11861 1560 11868 1571
rect 12202 1571 12268 1572
rect 12202 1560 12209 1571
rect 11861 1530 12209 1560
rect 11861 1519 11868 1530
rect 11802 1518 11868 1519
rect 12202 1519 12209 1530
rect 12261 1560 12268 1571
rect 12602 1571 12668 1572
rect 12602 1560 12609 1571
rect 12261 1530 12609 1560
rect 12261 1519 12268 1530
rect 12202 1518 12268 1519
rect 12602 1519 12609 1530
rect 12661 1560 12668 1571
rect 13104 1571 13170 1572
rect 13104 1560 13111 1571
rect 12661 1530 13111 1560
rect 12661 1519 12668 1530
rect 12602 1518 12668 1519
rect 13104 1519 13111 1530
rect 13163 1519 13170 1571
rect 13104 1518 13170 1519
rect 2 1501 68 1502
rect 2 1490 9 1501
rect 0 1460 9 1490
rect 2 1449 9 1460
rect 61 1490 68 1501
rect 402 1501 468 1502
rect 402 1490 409 1501
rect 61 1460 409 1490
rect 61 1449 68 1460
rect 2 1448 68 1449
rect 402 1449 409 1460
rect 461 1490 468 1501
rect 802 1501 868 1502
rect 802 1490 809 1501
rect 461 1460 809 1490
rect 461 1449 468 1460
rect 402 1448 468 1449
rect 802 1449 809 1460
rect 861 1490 868 1501
rect 1202 1501 1268 1502
rect 1202 1490 1209 1501
rect 861 1460 1209 1490
rect 861 1449 868 1460
rect 802 1448 868 1449
rect 1202 1449 1209 1460
rect 1261 1490 1268 1501
rect 1602 1501 1668 1502
rect 1602 1490 1609 1501
rect 1261 1460 1609 1490
rect 1261 1449 1268 1460
rect 1202 1448 1268 1449
rect 1602 1449 1609 1460
rect 1661 1490 1668 1501
rect 2002 1501 2068 1502
rect 2002 1490 2009 1501
rect 1661 1460 2009 1490
rect 1661 1449 1668 1460
rect 1602 1448 1668 1449
rect 2002 1449 2009 1460
rect 2061 1490 2068 1501
rect 2402 1501 2468 1502
rect 2402 1490 2409 1501
rect 2061 1460 2409 1490
rect 2061 1449 2068 1460
rect 2002 1448 2068 1449
rect 2402 1449 2409 1460
rect 2461 1490 2468 1501
rect 2802 1501 2868 1502
rect 2802 1490 2809 1501
rect 2461 1460 2809 1490
rect 2461 1449 2468 1460
rect 2402 1448 2468 1449
rect 2802 1449 2809 1460
rect 2861 1490 2868 1501
rect 3202 1501 3268 1502
rect 3202 1490 3209 1501
rect 2861 1460 3209 1490
rect 2861 1449 2868 1460
rect 2802 1448 2868 1449
rect 3202 1449 3209 1460
rect 3261 1490 3268 1501
rect 3602 1501 3668 1502
rect 3602 1490 3609 1501
rect 3261 1460 3609 1490
rect 3261 1449 3268 1460
rect 3202 1448 3268 1449
rect 3602 1449 3609 1460
rect 3661 1490 3668 1501
rect 4002 1501 4068 1502
rect 4002 1490 4009 1501
rect 3661 1460 4009 1490
rect 3661 1449 3668 1460
rect 3602 1448 3668 1449
rect 4002 1449 4009 1460
rect 4061 1490 4068 1501
rect 4402 1501 4468 1502
rect 4402 1490 4409 1501
rect 4061 1460 4409 1490
rect 4061 1449 4068 1460
rect 4002 1448 4068 1449
rect 4402 1449 4409 1460
rect 4461 1490 4468 1501
rect 4802 1501 4868 1502
rect 4802 1490 4809 1501
rect 4461 1460 4809 1490
rect 4461 1449 4468 1460
rect 4402 1448 4468 1449
rect 4802 1449 4809 1460
rect 4861 1490 4868 1501
rect 5202 1501 5268 1502
rect 5202 1490 5209 1501
rect 4861 1460 5209 1490
rect 4861 1449 4868 1460
rect 4802 1448 4868 1449
rect 5202 1449 5209 1460
rect 5261 1490 5268 1501
rect 5602 1501 5668 1502
rect 5602 1490 5609 1501
rect 5261 1460 5609 1490
rect 5261 1449 5268 1460
rect 5202 1448 5268 1449
rect 5602 1449 5609 1460
rect 5661 1490 5668 1501
rect 6002 1501 6068 1502
rect 6002 1490 6009 1501
rect 5661 1460 6009 1490
rect 5661 1449 5668 1460
rect 5602 1448 5668 1449
rect 6002 1449 6009 1460
rect 6061 1490 6068 1501
rect 6402 1501 6468 1502
rect 6402 1490 6409 1501
rect 6061 1460 6409 1490
rect 6061 1449 6068 1460
rect 6002 1448 6068 1449
rect 6402 1449 6409 1460
rect 6461 1490 6468 1501
rect 6802 1501 6868 1502
rect 6802 1490 6809 1501
rect 6461 1460 6809 1490
rect 6461 1449 6468 1460
rect 6402 1448 6468 1449
rect 6802 1449 6809 1460
rect 6861 1490 6868 1501
rect 7202 1501 7268 1502
rect 7202 1490 7209 1501
rect 6861 1460 7209 1490
rect 6861 1449 6868 1460
rect 6802 1448 6868 1449
rect 7202 1449 7209 1460
rect 7261 1490 7268 1501
rect 7602 1501 7668 1502
rect 7602 1490 7609 1501
rect 7261 1460 7609 1490
rect 7261 1449 7268 1460
rect 7202 1448 7268 1449
rect 7602 1449 7609 1460
rect 7661 1490 7668 1501
rect 8002 1501 8068 1502
rect 8002 1490 8009 1501
rect 7661 1460 8009 1490
rect 7661 1449 7668 1460
rect 7602 1448 7668 1449
rect 8002 1449 8009 1460
rect 8061 1490 8068 1501
rect 8402 1501 8468 1502
rect 8402 1490 8409 1501
rect 8061 1460 8409 1490
rect 8061 1449 8068 1460
rect 8002 1448 8068 1449
rect 8402 1449 8409 1460
rect 8461 1490 8468 1501
rect 8802 1501 8868 1502
rect 8802 1490 8809 1501
rect 8461 1460 8809 1490
rect 8461 1449 8468 1460
rect 8402 1448 8468 1449
rect 8802 1449 8809 1460
rect 8861 1490 8868 1501
rect 9202 1501 9268 1502
rect 9202 1490 9209 1501
rect 8861 1460 9209 1490
rect 8861 1449 8868 1460
rect 8802 1448 8868 1449
rect 9202 1449 9209 1460
rect 9261 1490 9268 1501
rect 9602 1501 9668 1502
rect 9602 1490 9609 1501
rect 9261 1460 9609 1490
rect 9261 1449 9268 1460
rect 9202 1448 9268 1449
rect 9602 1449 9609 1460
rect 9661 1490 9668 1501
rect 10002 1501 10068 1502
rect 10002 1490 10009 1501
rect 9661 1460 10009 1490
rect 9661 1449 9668 1460
rect 9602 1448 9668 1449
rect 10002 1449 10009 1460
rect 10061 1490 10068 1501
rect 10402 1501 10468 1502
rect 10402 1490 10409 1501
rect 10061 1460 10409 1490
rect 10061 1449 10068 1460
rect 10002 1448 10068 1449
rect 10402 1449 10409 1460
rect 10461 1490 10468 1501
rect 10802 1501 10868 1502
rect 10802 1490 10809 1501
rect 10461 1460 10809 1490
rect 10461 1449 10468 1460
rect 10402 1448 10468 1449
rect 10802 1449 10809 1460
rect 10861 1490 10868 1501
rect 11202 1501 11268 1502
rect 11202 1490 11209 1501
rect 10861 1460 11209 1490
rect 10861 1449 10868 1460
rect 10802 1448 10868 1449
rect 11202 1449 11209 1460
rect 11261 1490 11268 1501
rect 11602 1501 11668 1502
rect 11602 1490 11609 1501
rect 11261 1460 11609 1490
rect 11261 1449 11268 1460
rect 11202 1448 11268 1449
rect 11602 1449 11609 1460
rect 11661 1490 11668 1501
rect 12002 1501 12068 1502
rect 12002 1490 12009 1501
rect 11661 1460 12009 1490
rect 11661 1449 11668 1460
rect 11602 1448 11668 1449
rect 12002 1449 12009 1460
rect 12061 1490 12068 1501
rect 12402 1501 12468 1502
rect 12402 1490 12409 1501
rect 12061 1460 12409 1490
rect 12061 1449 12068 1460
rect 12002 1448 12068 1449
rect 12402 1449 12409 1460
rect 12461 1490 12468 1501
rect 12802 1501 12868 1502
rect 12802 1490 12809 1501
rect 12461 1460 12809 1490
rect 12461 1449 12468 1460
rect 12402 1448 12468 1449
rect 12802 1449 12809 1460
rect 12861 1490 12868 1501
rect 12900 1501 12966 1502
rect 12900 1490 12907 1501
rect 12861 1460 12907 1490
rect 12861 1449 12868 1460
rect 12802 1448 12868 1449
rect 12900 1449 12907 1460
rect 12959 1449 12966 1501
rect 12900 1448 12966 1449
rect 202 1431 268 1432
rect 202 1420 209 1431
rect 0 1390 209 1420
rect 202 1379 209 1390
rect 261 1420 268 1431
rect 602 1431 668 1432
rect 602 1420 609 1431
rect 261 1390 609 1420
rect 261 1379 268 1390
rect 202 1378 268 1379
rect 602 1379 609 1390
rect 661 1420 668 1431
rect 1002 1431 1068 1432
rect 1002 1420 1009 1431
rect 661 1390 1009 1420
rect 661 1379 668 1390
rect 602 1378 668 1379
rect 1002 1379 1009 1390
rect 1061 1420 1068 1431
rect 1402 1431 1468 1432
rect 1402 1420 1409 1431
rect 1061 1390 1409 1420
rect 1061 1379 1068 1390
rect 1002 1378 1068 1379
rect 1402 1379 1409 1390
rect 1461 1420 1468 1431
rect 1802 1431 1868 1432
rect 1802 1420 1809 1431
rect 1461 1390 1809 1420
rect 1461 1379 1468 1390
rect 1402 1378 1468 1379
rect 1802 1379 1809 1390
rect 1861 1420 1868 1431
rect 2202 1431 2268 1432
rect 2202 1420 2209 1431
rect 1861 1390 2209 1420
rect 1861 1379 1868 1390
rect 1802 1378 1868 1379
rect 2202 1379 2209 1390
rect 2261 1420 2268 1431
rect 2602 1431 2668 1432
rect 2602 1420 2609 1431
rect 2261 1390 2609 1420
rect 2261 1379 2268 1390
rect 2202 1378 2268 1379
rect 2602 1379 2609 1390
rect 2661 1420 2668 1431
rect 3002 1431 3068 1432
rect 3002 1420 3009 1431
rect 2661 1390 3009 1420
rect 2661 1379 2668 1390
rect 2602 1378 2668 1379
rect 3002 1379 3009 1390
rect 3061 1420 3068 1431
rect 3402 1431 3468 1432
rect 3402 1420 3409 1431
rect 3061 1390 3409 1420
rect 3061 1379 3068 1390
rect 3002 1378 3068 1379
rect 3402 1379 3409 1390
rect 3461 1420 3468 1431
rect 3802 1431 3868 1432
rect 3802 1420 3809 1431
rect 3461 1390 3809 1420
rect 3461 1379 3468 1390
rect 3402 1378 3468 1379
rect 3802 1379 3809 1390
rect 3861 1420 3868 1431
rect 4202 1431 4268 1432
rect 4202 1420 4209 1431
rect 3861 1390 4209 1420
rect 3861 1379 3868 1390
rect 3802 1378 3868 1379
rect 4202 1379 4209 1390
rect 4261 1420 4268 1431
rect 4602 1431 4668 1432
rect 4602 1420 4609 1431
rect 4261 1390 4609 1420
rect 4261 1379 4268 1390
rect 4202 1378 4268 1379
rect 4602 1379 4609 1390
rect 4661 1420 4668 1431
rect 5002 1431 5068 1432
rect 5002 1420 5009 1431
rect 4661 1390 5009 1420
rect 4661 1379 4668 1390
rect 4602 1378 4668 1379
rect 5002 1379 5009 1390
rect 5061 1420 5068 1431
rect 5402 1431 5468 1432
rect 5402 1420 5409 1431
rect 5061 1390 5409 1420
rect 5061 1379 5068 1390
rect 5002 1378 5068 1379
rect 5402 1379 5409 1390
rect 5461 1420 5468 1431
rect 5802 1431 5868 1432
rect 5802 1420 5809 1431
rect 5461 1390 5809 1420
rect 5461 1379 5468 1390
rect 5402 1378 5468 1379
rect 5802 1379 5809 1390
rect 5861 1420 5868 1431
rect 6202 1431 6268 1432
rect 6202 1420 6209 1431
rect 5861 1390 6209 1420
rect 5861 1379 5868 1390
rect 5802 1378 5868 1379
rect 6202 1379 6209 1390
rect 6261 1420 6268 1431
rect 6602 1431 6668 1432
rect 6602 1420 6609 1431
rect 6261 1390 6609 1420
rect 6261 1379 6268 1390
rect 6202 1378 6268 1379
rect 6602 1379 6609 1390
rect 6661 1420 6668 1431
rect 7002 1431 7068 1432
rect 7002 1420 7009 1431
rect 6661 1390 7009 1420
rect 6661 1379 6668 1390
rect 6602 1378 6668 1379
rect 7002 1379 7009 1390
rect 7061 1420 7068 1431
rect 7402 1431 7468 1432
rect 7402 1420 7409 1431
rect 7061 1390 7409 1420
rect 7061 1379 7068 1390
rect 7002 1378 7068 1379
rect 7402 1379 7409 1390
rect 7461 1420 7468 1431
rect 7802 1431 7868 1432
rect 7802 1420 7809 1431
rect 7461 1390 7809 1420
rect 7461 1379 7468 1390
rect 7402 1378 7468 1379
rect 7802 1379 7809 1390
rect 7861 1420 7868 1431
rect 8202 1431 8268 1432
rect 8202 1420 8209 1431
rect 7861 1390 8209 1420
rect 7861 1379 7868 1390
rect 7802 1378 7868 1379
rect 8202 1379 8209 1390
rect 8261 1420 8268 1431
rect 8602 1431 8668 1432
rect 8602 1420 8609 1431
rect 8261 1390 8609 1420
rect 8261 1379 8268 1390
rect 8202 1378 8268 1379
rect 8602 1379 8609 1390
rect 8661 1420 8668 1431
rect 9002 1431 9068 1432
rect 9002 1420 9009 1431
rect 8661 1390 9009 1420
rect 8661 1379 8668 1390
rect 8602 1378 8668 1379
rect 9002 1379 9009 1390
rect 9061 1420 9068 1431
rect 9402 1431 9468 1432
rect 9402 1420 9409 1431
rect 9061 1390 9409 1420
rect 9061 1379 9068 1390
rect 9002 1378 9068 1379
rect 9402 1379 9409 1390
rect 9461 1420 9468 1431
rect 9802 1431 9868 1432
rect 9802 1420 9809 1431
rect 9461 1390 9809 1420
rect 9461 1379 9468 1390
rect 9402 1378 9468 1379
rect 9802 1379 9809 1390
rect 9861 1420 9868 1431
rect 10202 1431 10268 1432
rect 10202 1420 10209 1431
rect 9861 1390 10209 1420
rect 9861 1379 9868 1390
rect 9802 1378 9868 1379
rect 10202 1379 10209 1390
rect 10261 1420 10268 1431
rect 10602 1431 10668 1432
rect 10602 1420 10609 1431
rect 10261 1390 10609 1420
rect 10261 1379 10268 1390
rect 10202 1378 10268 1379
rect 10602 1379 10609 1390
rect 10661 1420 10668 1431
rect 11002 1431 11068 1432
rect 11002 1420 11009 1431
rect 10661 1390 11009 1420
rect 10661 1379 10668 1390
rect 10602 1378 10668 1379
rect 11002 1379 11009 1390
rect 11061 1420 11068 1431
rect 11402 1431 11468 1432
rect 11402 1420 11409 1431
rect 11061 1390 11409 1420
rect 11061 1379 11068 1390
rect 11002 1378 11068 1379
rect 11402 1379 11409 1390
rect 11461 1420 11468 1431
rect 11802 1431 11868 1432
rect 11802 1420 11809 1431
rect 11461 1390 11809 1420
rect 11461 1379 11468 1390
rect 11402 1378 11468 1379
rect 11802 1379 11809 1390
rect 11861 1420 11868 1431
rect 12202 1431 12268 1432
rect 12202 1420 12209 1431
rect 11861 1390 12209 1420
rect 11861 1379 11868 1390
rect 11802 1378 11868 1379
rect 12202 1379 12209 1390
rect 12261 1420 12268 1431
rect 12602 1431 12668 1432
rect 12602 1420 12609 1431
rect 12261 1390 12609 1420
rect 12261 1379 12268 1390
rect 12202 1378 12268 1379
rect 12602 1379 12609 1390
rect 12661 1420 12668 1431
rect 13104 1431 13170 1432
rect 13104 1420 13111 1431
rect 12661 1390 13111 1420
rect 12661 1379 12668 1390
rect 12602 1378 12668 1379
rect 13104 1379 13111 1390
rect 13163 1379 13170 1431
rect 13104 1378 13170 1379
rect 2 1361 68 1362
rect 2 1350 9 1361
rect 0 1320 9 1350
rect 2 1309 9 1320
rect 61 1350 68 1361
rect 402 1361 468 1362
rect 402 1350 409 1361
rect 61 1320 409 1350
rect 61 1309 68 1320
rect 2 1308 68 1309
rect 402 1309 409 1320
rect 461 1350 468 1361
rect 802 1361 868 1362
rect 802 1350 809 1361
rect 461 1320 809 1350
rect 461 1309 468 1320
rect 402 1308 468 1309
rect 802 1309 809 1320
rect 861 1350 868 1361
rect 1202 1361 1268 1362
rect 1202 1350 1209 1361
rect 861 1320 1209 1350
rect 861 1309 868 1320
rect 802 1308 868 1309
rect 1202 1309 1209 1320
rect 1261 1350 1268 1361
rect 1602 1361 1668 1362
rect 1602 1350 1609 1361
rect 1261 1320 1609 1350
rect 1261 1309 1268 1320
rect 1202 1308 1268 1309
rect 1602 1309 1609 1320
rect 1661 1350 1668 1361
rect 2002 1361 2068 1362
rect 2002 1350 2009 1361
rect 1661 1320 2009 1350
rect 1661 1309 1668 1320
rect 1602 1308 1668 1309
rect 2002 1309 2009 1320
rect 2061 1350 2068 1361
rect 2402 1361 2468 1362
rect 2402 1350 2409 1361
rect 2061 1320 2409 1350
rect 2061 1309 2068 1320
rect 2002 1308 2068 1309
rect 2402 1309 2409 1320
rect 2461 1350 2468 1361
rect 2802 1361 2868 1362
rect 2802 1350 2809 1361
rect 2461 1320 2809 1350
rect 2461 1309 2468 1320
rect 2402 1308 2468 1309
rect 2802 1309 2809 1320
rect 2861 1350 2868 1361
rect 3202 1361 3268 1362
rect 3202 1350 3209 1361
rect 2861 1320 3209 1350
rect 2861 1309 2868 1320
rect 2802 1308 2868 1309
rect 3202 1309 3209 1320
rect 3261 1350 3268 1361
rect 3602 1361 3668 1362
rect 3602 1350 3609 1361
rect 3261 1320 3609 1350
rect 3261 1309 3268 1320
rect 3202 1308 3268 1309
rect 3602 1309 3609 1320
rect 3661 1350 3668 1361
rect 4002 1361 4068 1362
rect 4002 1350 4009 1361
rect 3661 1320 4009 1350
rect 3661 1309 3668 1320
rect 3602 1308 3668 1309
rect 4002 1309 4009 1320
rect 4061 1350 4068 1361
rect 4402 1361 4468 1362
rect 4402 1350 4409 1361
rect 4061 1320 4409 1350
rect 4061 1309 4068 1320
rect 4002 1308 4068 1309
rect 4402 1309 4409 1320
rect 4461 1350 4468 1361
rect 4802 1361 4868 1362
rect 4802 1350 4809 1361
rect 4461 1320 4809 1350
rect 4461 1309 4468 1320
rect 4402 1308 4468 1309
rect 4802 1309 4809 1320
rect 4861 1350 4868 1361
rect 5202 1361 5268 1362
rect 5202 1350 5209 1361
rect 4861 1320 5209 1350
rect 4861 1309 4868 1320
rect 4802 1308 4868 1309
rect 5202 1309 5209 1320
rect 5261 1350 5268 1361
rect 5602 1361 5668 1362
rect 5602 1350 5609 1361
rect 5261 1320 5609 1350
rect 5261 1309 5268 1320
rect 5202 1308 5268 1309
rect 5602 1309 5609 1320
rect 5661 1350 5668 1361
rect 6002 1361 6068 1362
rect 6002 1350 6009 1361
rect 5661 1320 6009 1350
rect 5661 1309 5668 1320
rect 5602 1308 5668 1309
rect 6002 1309 6009 1320
rect 6061 1350 6068 1361
rect 6402 1361 6468 1362
rect 6402 1350 6409 1361
rect 6061 1320 6409 1350
rect 6061 1309 6068 1320
rect 6002 1308 6068 1309
rect 6402 1309 6409 1320
rect 6461 1350 6468 1361
rect 6802 1361 6868 1362
rect 6802 1350 6809 1361
rect 6461 1320 6809 1350
rect 6461 1309 6468 1320
rect 6402 1308 6468 1309
rect 6802 1309 6809 1320
rect 6861 1350 6868 1361
rect 7202 1361 7268 1362
rect 7202 1350 7209 1361
rect 6861 1320 7209 1350
rect 6861 1309 6868 1320
rect 6802 1308 6868 1309
rect 7202 1309 7209 1320
rect 7261 1350 7268 1361
rect 7602 1361 7668 1362
rect 7602 1350 7609 1361
rect 7261 1320 7609 1350
rect 7261 1309 7268 1320
rect 7202 1308 7268 1309
rect 7602 1309 7609 1320
rect 7661 1350 7668 1361
rect 8002 1361 8068 1362
rect 8002 1350 8009 1361
rect 7661 1320 8009 1350
rect 7661 1309 7668 1320
rect 7602 1308 7668 1309
rect 8002 1309 8009 1320
rect 8061 1350 8068 1361
rect 8402 1361 8468 1362
rect 8402 1350 8409 1361
rect 8061 1320 8409 1350
rect 8061 1309 8068 1320
rect 8002 1308 8068 1309
rect 8402 1309 8409 1320
rect 8461 1350 8468 1361
rect 8802 1361 8868 1362
rect 8802 1350 8809 1361
rect 8461 1320 8809 1350
rect 8461 1309 8468 1320
rect 8402 1308 8468 1309
rect 8802 1309 8809 1320
rect 8861 1350 8868 1361
rect 9202 1361 9268 1362
rect 9202 1350 9209 1361
rect 8861 1320 9209 1350
rect 8861 1309 8868 1320
rect 8802 1308 8868 1309
rect 9202 1309 9209 1320
rect 9261 1350 9268 1361
rect 9602 1361 9668 1362
rect 9602 1350 9609 1361
rect 9261 1320 9609 1350
rect 9261 1309 9268 1320
rect 9202 1308 9268 1309
rect 9602 1309 9609 1320
rect 9661 1350 9668 1361
rect 10002 1361 10068 1362
rect 10002 1350 10009 1361
rect 9661 1320 10009 1350
rect 9661 1309 9668 1320
rect 9602 1308 9668 1309
rect 10002 1309 10009 1320
rect 10061 1350 10068 1361
rect 10402 1361 10468 1362
rect 10402 1350 10409 1361
rect 10061 1320 10409 1350
rect 10061 1309 10068 1320
rect 10002 1308 10068 1309
rect 10402 1309 10409 1320
rect 10461 1350 10468 1361
rect 10802 1361 10868 1362
rect 10802 1350 10809 1361
rect 10461 1320 10809 1350
rect 10461 1309 10468 1320
rect 10402 1308 10468 1309
rect 10802 1309 10809 1320
rect 10861 1350 10868 1361
rect 11202 1361 11268 1362
rect 11202 1350 11209 1361
rect 10861 1320 11209 1350
rect 10861 1309 10868 1320
rect 10802 1308 10868 1309
rect 11202 1309 11209 1320
rect 11261 1350 11268 1361
rect 11602 1361 11668 1362
rect 11602 1350 11609 1361
rect 11261 1320 11609 1350
rect 11261 1309 11268 1320
rect 11202 1308 11268 1309
rect 11602 1309 11609 1320
rect 11661 1350 11668 1361
rect 12002 1361 12068 1362
rect 12002 1350 12009 1361
rect 11661 1320 12009 1350
rect 11661 1309 11668 1320
rect 11602 1308 11668 1309
rect 12002 1309 12009 1320
rect 12061 1350 12068 1361
rect 12402 1361 12468 1362
rect 12402 1350 12409 1361
rect 12061 1320 12409 1350
rect 12061 1309 12068 1320
rect 12002 1308 12068 1309
rect 12402 1309 12409 1320
rect 12461 1350 12468 1361
rect 12802 1361 12868 1362
rect 12802 1350 12809 1361
rect 12461 1320 12809 1350
rect 12461 1309 12468 1320
rect 12402 1308 12468 1309
rect 12802 1309 12809 1320
rect 12861 1350 12868 1361
rect 12900 1361 12966 1362
rect 12900 1350 12907 1361
rect 12861 1320 12907 1350
rect 12861 1309 12868 1320
rect 12802 1308 12868 1309
rect 12900 1309 12907 1320
rect 12959 1309 12966 1361
rect 12900 1308 12966 1309
rect 196 1291 274 1292
rect -4 1275 74 1276
rect -4 1219 7 1275
rect 63 1219 74 1275
rect 196 1235 207 1291
rect 263 1235 274 1291
rect 596 1291 674 1292
rect 196 1234 274 1235
rect 396 1275 474 1276
rect -4 1218 74 1219
rect 396 1219 407 1275
rect 463 1219 474 1275
rect 596 1235 607 1291
rect 663 1235 674 1291
rect 996 1291 1074 1292
rect 596 1234 674 1235
rect 796 1275 874 1276
rect 396 1218 474 1219
rect 796 1219 807 1275
rect 863 1219 874 1275
rect 996 1235 1007 1291
rect 1063 1235 1074 1291
rect 1396 1291 1474 1292
rect 996 1234 1074 1235
rect 1196 1275 1274 1276
rect 796 1218 874 1219
rect 1196 1219 1207 1275
rect 1263 1219 1274 1275
rect 1396 1235 1407 1291
rect 1463 1235 1474 1291
rect 1796 1291 1874 1292
rect 1396 1234 1474 1235
rect 1596 1275 1674 1276
rect 1196 1218 1274 1219
rect 1596 1219 1607 1275
rect 1663 1219 1674 1275
rect 1796 1235 1807 1291
rect 1863 1235 1874 1291
rect 2196 1291 2274 1292
rect 1796 1234 1874 1235
rect 1996 1275 2074 1276
rect 1596 1218 1674 1219
rect 1996 1219 2007 1275
rect 2063 1219 2074 1275
rect 2196 1235 2207 1291
rect 2263 1235 2274 1291
rect 2596 1291 2674 1292
rect 2196 1234 2274 1235
rect 2396 1275 2474 1276
rect 1996 1218 2074 1219
rect 2396 1219 2407 1275
rect 2463 1219 2474 1275
rect 2596 1235 2607 1291
rect 2663 1235 2674 1291
rect 2996 1291 3074 1292
rect 2596 1234 2674 1235
rect 2796 1275 2874 1276
rect 2396 1218 2474 1219
rect 2796 1219 2807 1275
rect 2863 1219 2874 1275
rect 2996 1235 3007 1291
rect 3063 1235 3074 1291
rect 3396 1291 3474 1292
rect 2996 1234 3074 1235
rect 3196 1275 3274 1276
rect 2796 1218 2874 1219
rect 3196 1219 3207 1275
rect 3263 1219 3274 1275
rect 3396 1235 3407 1291
rect 3463 1235 3474 1291
rect 3796 1291 3874 1292
rect 3396 1234 3474 1235
rect 3596 1275 3674 1276
rect 3196 1218 3274 1219
rect 3596 1219 3607 1275
rect 3663 1219 3674 1275
rect 3796 1235 3807 1291
rect 3863 1235 3874 1291
rect 4196 1291 4274 1292
rect 3796 1234 3874 1235
rect 3996 1275 4074 1276
rect 3596 1218 3674 1219
rect 3996 1219 4007 1275
rect 4063 1219 4074 1275
rect 4196 1235 4207 1291
rect 4263 1235 4274 1291
rect 4596 1291 4674 1292
rect 4196 1234 4274 1235
rect 4396 1275 4474 1276
rect 3996 1218 4074 1219
rect 4396 1219 4407 1275
rect 4463 1219 4474 1275
rect 4596 1235 4607 1291
rect 4663 1235 4674 1291
rect 4996 1291 5074 1292
rect 4596 1234 4674 1235
rect 4796 1275 4874 1276
rect 4396 1218 4474 1219
rect 4796 1219 4807 1275
rect 4863 1219 4874 1275
rect 4996 1235 5007 1291
rect 5063 1235 5074 1291
rect 5396 1291 5474 1292
rect 4996 1234 5074 1235
rect 5196 1275 5274 1276
rect 4796 1218 4874 1219
rect 5196 1219 5207 1275
rect 5263 1219 5274 1275
rect 5396 1235 5407 1291
rect 5463 1235 5474 1291
rect 5796 1291 5874 1292
rect 5396 1234 5474 1235
rect 5596 1275 5674 1276
rect 5196 1218 5274 1219
rect 5596 1219 5607 1275
rect 5663 1219 5674 1275
rect 5796 1235 5807 1291
rect 5863 1235 5874 1291
rect 6196 1291 6274 1292
rect 5796 1234 5874 1235
rect 5996 1275 6074 1276
rect 5596 1218 5674 1219
rect 5996 1219 6007 1275
rect 6063 1219 6074 1275
rect 6196 1235 6207 1291
rect 6263 1235 6274 1291
rect 6596 1291 6674 1292
rect 6196 1234 6274 1235
rect 6396 1275 6474 1276
rect 5996 1218 6074 1219
rect 6396 1219 6407 1275
rect 6463 1219 6474 1275
rect 6596 1235 6607 1291
rect 6663 1235 6674 1291
rect 6996 1291 7074 1292
rect 6596 1234 6674 1235
rect 6796 1275 6874 1276
rect 6396 1218 6474 1219
rect 6796 1219 6807 1275
rect 6863 1219 6874 1275
rect 6996 1235 7007 1291
rect 7063 1235 7074 1291
rect 7396 1291 7474 1292
rect 6996 1234 7074 1235
rect 7196 1275 7274 1276
rect 6796 1218 6874 1219
rect 7196 1219 7207 1275
rect 7263 1219 7274 1275
rect 7396 1235 7407 1291
rect 7463 1235 7474 1291
rect 7796 1291 7874 1292
rect 7396 1234 7474 1235
rect 7596 1275 7674 1276
rect 7196 1218 7274 1219
rect 7596 1219 7607 1275
rect 7663 1219 7674 1275
rect 7796 1235 7807 1291
rect 7863 1235 7874 1291
rect 8196 1291 8274 1292
rect 7796 1234 7874 1235
rect 7996 1275 8074 1276
rect 7596 1218 7674 1219
rect 7996 1219 8007 1275
rect 8063 1219 8074 1275
rect 8196 1235 8207 1291
rect 8263 1235 8274 1291
rect 8596 1291 8674 1292
rect 8196 1234 8274 1235
rect 8396 1275 8474 1276
rect 7996 1218 8074 1219
rect 8396 1219 8407 1275
rect 8463 1219 8474 1275
rect 8596 1235 8607 1291
rect 8663 1235 8674 1291
rect 8996 1291 9074 1292
rect 8596 1234 8674 1235
rect 8796 1275 8874 1276
rect 8396 1218 8474 1219
rect 8796 1219 8807 1275
rect 8863 1219 8874 1275
rect 8996 1235 9007 1291
rect 9063 1235 9074 1291
rect 9396 1291 9474 1292
rect 8996 1234 9074 1235
rect 9196 1275 9274 1276
rect 8796 1218 8874 1219
rect 9196 1219 9207 1275
rect 9263 1219 9274 1275
rect 9396 1235 9407 1291
rect 9463 1235 9474 1291
rect 9796 1291 9874 1292
rect 9396 1234 9474 1235
rect 9596 1275 9674 1276
rect 9196 1218 9274 1219
rect 9596 1219 9607 1275
rect 9663 1219 9674 1275
rect 9796 1235 9807 1291
rect 9863 1235 9874 1291
rect 10196 1291 10274 1292
rect 9796 1234 9874 1235
rect 9996 1275 10074 1276
rect 9596 1218 9674 1219
rect 9996 1219 10007 1275
rect 10063 1219 10074 1275
rect 10196 1235 10207 1291
rect 10263 1235 10274 1291
rect 10596 1291 10674 1292
rect 10196 1234 10274 1235
rect 10396 1275 10474 1276
rect 9996 1218 10074 1219
rect 10396 1219 10407 1275
rect 10463 1219 10474 1275
rect 10596 1235 10607 1291
rect 10663 1235 10674 1291
rect 10996 1291 11074 1292
rect 10596 1234 10674 1235
rect 10796 1275 10874 1276
rect 10396 1218 10474 1219
rect 10796 1219 10807 1275
rect 10863 1219 10874 1275
rect 10996 1235 11007 1291
rect 11063 1235 11074 1291
rect 11396 1291 11474 1292
rect 10996 1234 11074 1235
rect 11196 1275 11274 1276
rect 10796 1218 10874 1219
rect 11196 1219 11207 1275
rect 11263 1219 11274 1275
rect 11396 1235 11407 1291
rect 11463 1235 11474 1291
rect 11796 1291 11874 1292
rect 11396 1234 11474 1235
rect 11596 1275 11674 1276
rect 11196 1218 11274 1219
rect 11596 1219 11607 1275
rect 11663 1219 11674 1275
rect 11796 1235 11807 1291
rect 11863 1235 11874 1291
rect 12196 1291 12274 1292
rect 11796 1234 11874 1235
rect 11996 1275 12074 1276
rect 11596 1218 11674 1219
rect 11996 1219 12007 1275
rect 12063 1219 12074 1275
rect 12196 1235 12207 1291
rect 12263 1235 12274 1291
rect 12596 1291 12674 1292
rect 12196 1234 12274 1235
rect 12396 1275 12474 1276
rect 11996 1218 12074 1219
rect 12396 1219 12407 1275
rect 12463 1219 12474 1275
rect 12596 1235 12607 1291
rect 12663 1235 12674 1291
rect 12596 1234 12674 1235
rect 12396 1218 12474 1219
rect 202 1201 268 1202
rect 202 1190 209 1201
rect 0 1160 209 1190
rect 202 1149 209 1160
rect 261 1190 268 1201
rect 602 1201 668 1202
rect 602 1190 609 1201
rect 261 1160 609 1190
rect 261 1149 268 1160
rect 202 1148 268 1149
rect 602 1149 609 1160
rect 661 1190 668 1201
rect 1002 1201 1068 1202
rect 1002 1190 1009 1201
rect 661 1160 1009 1190
rect 661 1149 668 1160
rect 602 1148 668 1149
rect 1002 1149 1009 1160
rect 1061 1190 1068 1201
rect 1402 1201 1468 1202
rect 1402 1190 1409 1201
rect 1061 1160 1409 1190
rect 1061 1149 1068 1160
rect 1002 1148 1068 1149
rect 1402 1149 1409 1160
rect 1461 1190 1468 1201
rect 1802 1201 1868 1202
rect 1802 1190 1809 1201
rect 1461 1160 1809 1190
rect 1461 1149 1468 1160
rect 1402 1148 1468 1149
rect 1802 1149 1809 1160
rect 1861 1190 1868 1201
rect 2202 1201 2268 1202
rect 2202 1190 2209 1201
rect 1861 1160 2209 1190
rect 1861 1149 1868 1160
rect 1802 1148 1868 1149
rect 2202 1149 2209 1160
rect 2261 1190 2268 1201
rect 2602 1201 2668 1202
rect 2602 1190 2609 1201
rect 2261 1160 2609 1190
rect 2261 1149 2268 1160
rect 2202 1148 2268 1149
rect 2602 1149 2609 1160
rect 2661 1190 2668 1201
rect 3002 1201 3068 1202
rect 3002 1190 3009 1201
rect 2661 1160 3009 1190
rect 2661 1149 2668 1160
rect 2602 1148 2668 1149
rect 3002 1149 3009 1160
rect 3061 1190 3068 1201
rect 3402 1201 3468 1202
rect 3402 1190 3409 1201
rect 3061 1160 3409 1190
rect 3061 1149 3068 1160
rect 3002 1148 3068 1149
rect 3402 1149 3409 1160
rect 3461 1190 3468 1201
rect 3802 1201 3868 1202
rect 3802 1190 3809 1201
rect 3461 1160 3809 1190
rect 3461 1149 3468 1160
rect 3402 1148 3468 1149
rect 3802 1149 3809 1160
rect 3861 1190 3868 1201
rect 4202 1201 4268 1202
rect 4202 1190 4209 1201
rect 3861 1160 4209 1190
rect 3861 1149 3868 1160
rect 3802 1148 3868 1149
rect 4202 1149 4209 1160
rect 4261 1190 4268 1201
rect 4602 1201 4668 1202
rect 4602 1190 4609 1201
rect 4261 1160 4609 1190
rect 4261 1149 4268 1160
rect 4202 1148 4268 1149
rect 4602 1149 4609 1160
rect 4661 1190 4668 1201
rect 5002 1201 5068 1202
rect 5002 1190 5009 1201
rect 4661 1160 5009 1190
rect 4661 1149 4668 1160
rect 4602 1148 4668 1149
rect 5002 1149 5009 1160
rect 5061 1190 5068 1201
rect 5402 1201 5468 1202
rect 5402 1190 5409 1201
rect 5061 1160 5409 1190
rect 5061 1149 5068 1160
rect 5002 1148 5068 1149
rect 5402 1149 5409 1160
rect 5461 1190 5468 1201
rect 5802 1201 5868 1202
rect 5802 1190 5809 1201
rect 5461 1160 5809 1190
rect 5461 1149 5468 1160
rect 5402 1148 5468 1149
rect 5802 1149 5809 1160
rect 5861 1190 5868 1201
rect 6202 1201 6268 1202
rect 6202 1190 6209 1201
rect 5861 1160 6209 1190
rect 5861 1149 5868 1160
rect 5802 1148 5868 1149
rect 6202 1149 6209 1160
rect 6261 1190 6268 1201
rect 6602 1201 6668 1202
rect 6602 1190 6609 1201
rect 6261 1160 6609 1190
rect 6261 1149 6268 1160
rect 6202 1148 6268 1149
rect 6602 1149 6609 1160
rect 6661 1190 6668 1201
rect 7002 1201 7068 1202
rect 7002 1190 7009 1201
rect 6661 1160 7009 1190
rect 6661 1149 6668 1160
rect 6602 1148 6668 1149
rect 7002 1149 7009 1160
rect 7061 1190 7068 1201
rect 7402 1201 7468 1202
rect 7402 1190 7409 1201
rect 7061 1160 7409 1190
rect 7061 1149 7068 1160
rect 7002 1148 7068 1149
rect 7402 1149 7409 1160
rect 7461 1190 7468 1201
rect 7802 1201 7868 1202
rect 7802 1190 7809 1201
rect 7461 1160 7809 1190
rect 7461 1149 7468 1160
rect 7402 1148 7468 1149
rect 7802 1149 7809 1160
rect 7861 1190 7868 1201
rect 8202 1201 8268 1202
rect 8202 1190 8209 1201
rect 7861 1160 8209 1190
rect 7861 1149 7868 1160
rect 7802 1148 7868 1149
rect 8202 1149 8209 1160
rect 8261 1190 8268 1201
rect 8602 1201 8668 1202
rect 8602 1190 8609 1201
rect 8261 1160 8609 1190
rect 8261 1149 8268 1160
rect 8202 1148 8268 1149
rect 8602 1149 8609 1160
rect 8661 1190 8668 1201
rect 9002 1201 9068 1202
rect 9002 1190 9009 1201
rect 8661 1160 9009 1190
rect 8661 1149 8668 1160
rect 8602 1148 8668 1149
rect 9002 1149 9009 1160
rect 9061 1190 9068 1201
rect 9402 1201 9468 1202
rect 9402 1190 9409 1201
rect 9061 1160 9409 1190
rect 9061 1149 9068 1160
rect 9002 1148 9068 1149
rect 9402 1149 9409 1160
rect 9461 1190 9468 1201
rect 9802 1201 9868 1202
rect 9802 1190 9809 1201
rect 9461 1160 9809 1190
rect 9461 1149 9468 1160
rect 9402 1148 9468 1149
rect 9802 1149 9809 1160
rect 9861 1190 9868 1201
rect 10202 1201 10268 1202
rect 10202 1190 10209 1201
rect 9861 1160 10209 1190
rect 9861 1149 9868 1160
rect 9802 1148 9868 1149
rect 10202 1149 10209 1160
rect 10261 1190 10268 1201
rect 10602 1201 10668 1202
rect 10602 1190 10609 1201
rect 10261 1160 10609 1190
rect 10261 1149 10268 1160
rect 10202 1148 10268 1149
rect 10602 1149 10609 1160
rect 10661 1190 10668 1201
rect 11002 1201 11068 1202
rect 11002 1190 11009 1201
rect 10661 1160 11009 1190
rect 10661 1149 10668 1160
rect 10602 1148 10668 1149
rect 11002 1149 11009 1160
rect 11061 1190 11068 1201
rect 11402 1201 11468 1202
rect 11402 1190 11409 1201
rect 11061 1160 11409 1190
rect 11061 1149 11068 1160
rect 11002 1148 11068 1149
rect 11402 1149 11409 1160
rect 11461 1190 11468 1201
rect 11802 1201 11868 1202
rect 11802 1190 11809 1201
rect 11461 1160 11809 1190
rect 11461 1149 11468 1160
rect 11402 1148 11468 1149
rect 11802 1149 11809 1160
rect 11861 1190 11868 1201
rect 12202 1201 12268 1202
rect 12202 1190 12209 1201
rect 11861 1160 12209 1190
rect 11861 1149 11868 1160
rect 11802 1148 11868 1149
rect 12202 1149 12209 1160
rect 12261 1190 12268 1201
rect 12602 1201 12668 1202
rect 12602 1190 12609 1201
rect 12261 1160 12609 1190
rect 12261 1149 12268 1160
rect 12202 1148 12268 1149
rect 12602 1149 12609 1160
rect 12661 1190 12668 1201
rect 13104 1201 13170 1202
rect 13104 1190 13111 1201
rect 12661 1160 13111 1190
rect 12661 1149 12668 1160
rect 12602 1148 12668 1149
rect 13104 1149 13111 1160
rect 13163 1149 13170 1201
rect 13104 1148 13170 1149
rect 2 1131 68 1132
rect 2 1120 9 1131
rect 0 1090 9 1120
rect 2 1079 9 1090
rect 61 1120 68 1131
rect 402 1131 468 1132
rect 402 1120 409 1131
rect 61 1090 409 1120
rect 61 1079 68 1090
rect 2 1078 68 1079
rect 402 1079 409 1090
rect 461 1120 468 1131
rect 802 1131 868 1132
rect 802 1120 809 1131
rect 461 1090 809 1120
rect 461 1079 468 1090
rect 402 1078 468 1079
rect 802 1079 809 1090
rect 861 1120 868 1131
rect 1202 1131 1268 1132
rect 1202 1120 1209 1131
rect 861 1090 1209 1120
rect 861 1079 868 1090
rect 802 1078 868 1079
rect 1202 1079 1209 1090
rect 1261 1120 1268 1131
rect 1602 1131 1668 1132
rect 1602 1120 1609 1131
rect 1261 1090 1609 1120
rect 1261 1079 1268 1090
rect 1202 1078 1268 1079
rect 1602 1079 1609 1090
rect 1661 1120 1668 1131
rect 2002 1131 2068 1132
rect 2002 1120 2009 1131
rect 1661 1090 2009 1120
rect 1661 1079 1668 1090
rect 1602 1078 1668 1079
rect 2002 1079 2009 1090
rect 2061 1120 2068 1131
rect 2402 1131 2468 1132
rect 2402 1120 2409 1131
rect 2061 1090 2409 1120
rect 2061 1079 2068 1090
rect 2002 1078 2068 1079
rect 2402 1079 2409 1090
rect 2461 1120 2468 1131
rect 2802 1131 2868 1132
rect 2802 1120 2809 1131
rect 2461 1090 2809 1120
rect 2461 1079 2468 1090
rect 2402 1078 2468 1079
rect 2802 1079 2809 1090
rect 2861 1120 2868 1131
rect 3202 1131 3268 1132
rect 3202 1120 3209 1131
rect 2861 1090 3209 1120
rect 2861 1079 2868 1090
rect 2802 1078 2868 1079
rect 3202 1079 3209 1090
rect 3261 1120 3268 1131
rect 3602 1131 3668 1132
rect 3602 1120 3609 1131
rect 3261 1090 3609 1120
rect 3261 1079 3268 1090
rect 3202 1078 3268 1079
rect 3602 1079 3609 1090
rect 3661 1120 3668 1131
rect 4002 1131 4068 1132
rect 4002 1120 4009 1131
rect 3661 1090 4009 1120
rect 3661 1079 3668 1090
rect 3602 1078 3668 1079
rect 4002 1079 4009 1090
rect 4061 1120 4068 1131
rect 4402 1131 4468 1132
rect 4402 1120 4409 1131
rect 4061 1090 4409 1120
rect 4061 1079 4068 1090
rect 4002 1078 4068 1079
rect 4402 1079 4409 1090
rect 4461 1120 4468 1131
rect 4802 1131 4868 1132
rect 4802 1120 4809 1131
rect 4461 1090 4809 1120
rect 4461 1079 4468 1090
rect 4402 1078 4468 1079
rect 4802 1079 4809 1090
rect 4861 1120 4868 1131
rect 5202 1131 5268 1132
rect 5202 1120 5209 1131
rect 4861 1090 5209 1120
rect 4861 1079 4868 1090
rect 4802 1078 4868 1079
rect 5202 1079 5209 1090
rect 5261 1120 5268 1131
rect 5602 1131 5668 1132
rect 5602 1120 5609 1131
rect 5261 1090 5609 1120
rect 5261 1079 5268 1090
rect 5202 1078 5268 1079
rect 5602 1079 5609 1090
rect 5661 1120 5668 1131
rect 6002 1131 6068 1132
rect 6002 1120 6009 1131
rect 5661 1090 6009 1120
rect 5661 1079 5668 1090
rect 5602 1078 5668 1079
rect 6002 1079 6009 1090
rect 6061 1120 6068 1131
rect 6402 1131 6468 1132
rect 6402 1120 6409 1131
rect 6061 1090 6409 1120
rect 6061 1079 6068 1090
rect 6002 1078 6068 1079
rect 6402 1079 6409 1090
rect 6461 1120 6468 1131
rect 6802 1131 6868 1132
rect 6802 1120 6809 1131
rect 6461 1090 6809 1120
rect 6461 1079 6468 1090
rect 6402 1078 6468 1079
rect 6802 1079 6809 1090
rect 6861 1120 6868 1131
rect 7202 1131 7268 1132
rect 7202 1120 7209 1131
rect 6861 1090 7209 1120
rect 6861 1079 6868 1090
rect 6802 1078 6868 1079
rect 7202 1079 7209 1090
rect 7261 1120 7268 1131
rect 7602 1131 7668 1132
rect 7602 1120 7609 1131
rect 7261 1090 7609 1120
rect 7261 1079 7268 1090
rect 7202 1078 7268 1079
rect 7602 1079 7609 1090
rect 7661 1120 7668 1131
rect 8002 1131 8068 1132
rect 8002 1120 8009 1131
rect 7661 1090 8009 1120
rect 7661 1079 7668 1090
rect 7602 1078 7668 1079
rect 8002 1079 8009 1090
rect 8061 1120 8068 1131
rect 8402 1131 8468 1132
rect 8402 1120 8409 1131
rect 8061 1090 8409 1120
rect 8061 1079 8068 1090
rect 8002 1078 8068 1079
rect 8402 1079 8409 1090
rect 8461 1120 8468 1131
rect 8802 1131 8868 1132
rect 8802 1120 8809 1131
rect 8461 1090 8809 1120
rect 8461 1079 8468 1090
rect 8402 1078 8468 1079
rect 8802 1079 8809 1090
rect 8861 1120 8868 1131
rect 9202 1131 9268 1132
rect 9202 1120 9209 1131
rect 8861 1090 9209 1120
rect 8861 1079 8868 1090
rect 8802 1078 8868 1079
rect 9202 1079 9209 1090
rect 9261 1120 9268 1131
rect 9602 1131 9668 1132
rect 9602 1120 9609 1131
rect 9261 1090 9609 1120
rect 9261 1079 9268 1090
rect 9202 1078 9268 1079
rect 9602 1079 9609 1090
rect 9661 1120 9668 1131
rect 10002 1131 10068 1132
rect 10002 1120 10009 1131
rect 9661 1090 10009 1120
rect 9661 1079 9668 1090
rect 9602 1078 9668 1079
rect 10002 1079 10009 1090
rect 10061 1120 10068 1131
rect 10402 1131 10468 1132
rect 10402 1120 10409 1131
rect 10061 1090 10409 1120
rect 10061 1079 10068 1090
rect 10002 1078 10068 1079
rect 10402 1079 10409 1090
rect 10461 1120 10468 1131
rect 10802 1131 10868 1132
rect 10802 1120 10809 1131
rect 10461 1090 10809 1120
rect 10461 1079 10468 1090
rect 10402 1078 10468 1079
rect 10802 1079 10809 1090
rect 10861 1120 10868 1131
rect 11202 1131 11268 1132
rect 11202 1120 11209 1131
rect 10861 1090 11209 1120
rect 10861 1079 10868 1090
rect 10802 1078 10868 1079
rect 11202 1079 11209 1090
rect 11261 1120 11268 1131
rect 11602 1131 11668 1132
rect 11602 1120 11609 1131
rect 11261 1090 11609 1120
rect 11261 1079 11268 1090
rect 11202 1078 11268 1079
rect 11602 1079 11609 1090
rect 11661 1120 11668 1131
rect 12002 1131 12068 1132
rect 12002 1120 12009 1131
rect 11661 1090 12009 1120
rect 11661 1079 11668 1090
rect 11602 1078 11668 1079
rect 12002 1079 12009 1090
rect 12061 1120 12068 1131
rect 12402 1131 12468 1132
rect 12402 1120 12409 1131
rect 12061 1090 12409 1120
rect 12061 1079 12068 1090
rect 12002 1078 12068 1079
rect 12402 1079 12409 1090
rect 12461 1120 12468 1131
rect 12802 1131 12868 1132
rect 12802 1120 12809 1131
rect 12461 1090 12809 1120
rect 12461 1079 12468 1090
rect 12402 1078 12468 1079
rect 12802 1079 12809 1090
rect 12861 1120 12868 1131
rect 12900 1131 12966 1132
rect 12900 1120 12907 1131
rect 12861 1090 12907 1120
rect 12861 1079 12868 1090
rect 12802 1078 12868 1079
rect 12900 1079 12907 1090
rect 12959 1079 12966 1131
rect 12900 1078 12966 1079
rect 202 1061 268 1062
rect 202 1050 209 1061
rect 0 1020 209 1050
rect 202 1009 209 1020
rect 261 1050 268 1061
rect 602 1061 668 1062
rect 602 1050 609 1061
rect 261 1020 609 1050
rect 261 1009 268 1020
rect 202 1008 268 1009
rect 602 1009 609 1020
rect 661 1050 668 1061
rect 1002 1061 1068 1062
rect 1002 1050 1009 1061
rect 661 1020 1009 1050
rect 661 1009 668 1020
rect 602 1008 668 1009
rect 1002 1009 1009 1020
rect 1061 1050 1068 1061
rect 1402 1061 1468 1062
rect 1402 1050 1409 1061
rect 1061 1020 1409 1050
rect 1061 1009 1068 1020
rect 1002 1008 1068 1009
rect 1402 1009 1409 1020
rect 1461 1050 1468 1061
rect 1802 1061 1868 1062
rect 1802 1050 1809 1061
rect 1461 1020 1809 1050
rect 1461 1009 1468 1020
rect 1402 1008 1468 1009
rect 1802 1009 1809 1020
rect 1861 1050 1868 1061
rect 2202 1061 2268 1062
rect 2202 1050 2209 1061
rect 1861 1020 2209 1050
rect 1861 1009 1868 1020
rect 1802 1008 1868 1009
rect 2202 1009 2209 1020
rect 2261 1050 2268 1061
rect 2602 1061 2668 1062
rect 2602 1050 2609 1061
rect 2261 1020 2609 1050
rect 2261 1009 2268 1020
rect 2202 1008 2268 1009
rect 2602 1009 2609 1020
rect 2661 1050 2668 1061
rect 3002 1061 3068 1062
rect 3002 1050 3009 1061
rect 2661 1020 3009 1050
rect 2661 1009 2668 1020
rect 2602 1008 2668 1009
rect 3002 1009 3009 1020
rect 3061 1050 3068 1061
rect 3402 1061 3468 1062
rect 3402 1050 3409 1061
rect 3061 1020 3409 1050
rect 3061 1009 3068 1020
rect 3002 1008 3068 1009
rect 3402 1009 3409 1020
rect 3461 1050 3468 1061
rect 3802 1061 3868 1062
rect 3802 1050 3809 1061
rect 3461 1020 3809 1050
rect 3461 1009 3468 1020
rect 3402 1008 3468 1009
rect 3802 1009 3809 1020
rect 3861 1050 3868 1061
rect 4202 1061 4268 1062
rect 4202 1050 4209 1061
rect 3861 1020 4209 1050
rect 3861 1009 3868 1020
rect 3802 1008 3868 1009
rect 4202 1009 4209 1020
rect 4261 1050 4268 1061
rect 4602 1061 4668 1062
rect 4602 1050 4609 1061
rect 4261 1020 4609 1050
rect 4261 1009 4268 1020
rect 4202 1008 4268 1009
rect 4602 1009 4609 1020
rect 4661 1050 4668 1061
rect 5002 1061 5068 1062
rect 5002 1050 5009 1061
rect 4661 1020 5009 1050
rect 4661 1009 4668 1020
rect 4602 1008 4668 1009
rect 5002 1009 5009 1020
rect 5061 1050 5068 1061
rect 5402 1061 5468 1062
rect 5402 1050 5409 1061
rect 5061 1020 5409 1050
rect 5061 1009 5068 1020
rect 5002 1008 5068 1009
rect 5402 1009 5409 1020
rect 5461 1050 5468 1061
rect 5802 1061 5868 1062
rect 5802 1050 5809 1061
rect 5461 1020 5809 1050
rect 5461 1009 5468 1020
rect 5402 1008 5468 1009
rect 5802 1009 5809 1020
rect 5861 1050 5868 1061
rect 6202 1061 6268 1062
rect 6202 1050 6209 1061
rect 5861 1020 6209 1050
rect 5861 1009 5868 1020
rect 5802 1008 5868 1009
rect 6202 1009 6209 1020
rect 6261 1050 6268 1061
rect 6602 1061 6668 1062
rect 6602 1050 6609 1061
rect 6261 1020 6609 1050
rect 6261 1009 6268 1020
rect 6202 1008 6268 1009
rect 6602 1009 6609 1020
rect 6661 1050 6668 1061
rect 7002 1061 7068 1062
rect 7002 1050 7009 1061
rect 6661 1020 7009 1050
rect 6661 1009 6668 1020
rect 6602 1008 6668 1009
rect 7002 1009 7009 1020
rect 7061 1050 7068 1061
rect 7402 1061 7468 1062
rect 7402 1050 7409 1061
rect 7061 1020 7409 1050
rect 7061 1009 7068 1020
rect 7002 1008 7068 1009
rect 7402 1009 7409 1020
rect 7461 1050 7468 1061
rect 7802 1061 7868 1062
rect 7802 1050 7809 1061
rect 7461 1020 7809 1050
rect 7461 1009 7468 1020
rect 7402 1008 7468 1009
rect 7802 1009 7809 1020
rect 7861 1050 7868 1061
rect 8202 1061 8268 1062
rect 8202 1050 8209 1061
rect 7861 1020 8209 1050
rect 7861 1009 7868 1020
rect 7802 1008 7868 1009
rect 8202 1009 8209 1020
rect 8261 1050 8268 1061
rect 8602 1061 8668 1062
rect 8602 1050 8609 1061
rect 8261 1020 8609 1050
rect 8261 1009 8268 1020
rect 8202 1008 8268 1009
rect 8602 1009 8609 1020
rect 8661 1050 8668 1061
rect 9002 1061 9068 1062
rect 9002 1050 9009 1061
rect 8661 1020 9009 1050
rect 8661 1009 8668 1020
rect 8602 1008 8668 1009
rect 9002 1009 9009 1020
rect 9061 1050 9068 1061
rect 9402 1061 9468 1062
rect 9402 1050 9409 1061
rect 9061 1020 9409 1050
rect 9061 1009 9068 1020
rect 9002 1008 9068 1009
rect 9402 1009 9409 1020
rect 9461 1050 9468 1061
rect 9802 1061 9868 1062
rect 9802 1050 9809 1061
rect 9461 1020 9809 1050
rect 9461 1009 9468 1020
rect 9402 1008 9468 1009
rect 9802 1009 9809 1020
rect 9861 1050 9868 1061
rect 10202 1061 10268 1062
rect 10202 1050 10209 1061
rect 9861 1020 10209 1050
rect 9861 1009 9868 1020
rect 9802 1008 9868 1009
rect 10202 1009 10209 1020
rect 10261 1050 10268 1061
rect 10602 1061 10668 1062
rect 10602 1050 10609 1061
rect 10261 1020 10609 1050
rect 10261 1009 10268 1020
rect 10202 1008 10268 1009
rect 10602 1009 10609 1020
rect 10661 1050 10668 1061
rect 11002 1061 11068 1062
rect 11002 1050 11009 1061
rect 10661 1020 11009 1050
rect 10661 1009 10668 1020
rect 10602 1008 10668 1009
rect 11002 1009 11009 1020
rect 11061 1050 11068 1061
rect 11402 1061 11468 1062
rect 11402 1050 11409 1061
rect 11061 1020 11409 1050
rect 11061 1009 11068 1020
rect 11002 1008 11068 1009
rect 11402 1009 11409 1020
rect 11461 1050 11468 1061
rect 11802 1061 11868 1062
rect 11802 1050 11809 1061
rect 11461 1020 11809 1050
rect 11461 1009 11468 1020
rect 11402 1008 11468 1009
rect 11802 1009 11809 1020
rect 11861 1050 11868 1061
rect 12202 1061 12268 1062
rect 12202 1050 12209 1061
rect 11861 1020 12209 1050
rect 11861 1009 11868 1020
rect 11802 1008 11868 1009
rect 12202 1009 12209 1020
rect 12261 1050 12268 1061
rect 12602 1061 12668 1062
rect 12602 1050 12609 1061
rect 12261 1020 12609 1050
rect 12261 1009 12268 1020
rect 12202 1008 12268 1009
rect 12602 1009 12609 1020
rect 12661 1050 12668 1061
rect 13104 1061 13170 1062
rect 13104 1050 13111 1061
rect 12661 1020 13111 1050
rect 12661 1009 12668 1020
rect 12602 1008 12668 1009
rect 13104 1009 13111 1020
rect 13163 1009 13170 1061
rect 13104 1008 13170 1009
rect 2 991 68 992
rect 2 980 9 991
rect 0 950 9 980
rect 2 939 9 950
rect 61 980 68 991
rect 402 991 468 992
rect 402 980 409 991
rect 61 950 409 980
rect 61 939 68 950
rect 2 938 68 939
rect 402 939 409 950
rect 461 980 468 991
rect 802 991 868 992
rect 802 980 809 991
rect 461 950 809 980
rect 461 939 468 950
rect 402 938 468 939
rect 802 939 809 950
rect 861 980 868 991
rect 1202 991 1268 992
rect 1202 980 1209 991
rect 861 950 1209 980
rect 861 939 868 950
rect 802 938 868 939
rect 1202 939 1209 950
rect 1261 980 1268 991
rect 1602 991 1668 992
rect 1602 980 1609 991
rect 1261 950 1609 980
rect 1261 939 1268 950
rect 1202 938 1268 939
rect 1602 939 1609 950
rect 1661 980 1668 991
rect 2002 991 2068 992
rect 2002 980 2009 991
rect 1661 950 2009 980
rect 1661 939 1668 950
rect 1602 938 1668 939
rect 2002 939 2009 950
rect 2061 980 2068 991
rect 2402 991 2468 992
rect 2402 980 2409 991
rect 2061 950 2409 980
rect 2061 939 2068 950
rect 2002 938 2068 939
rect 2402 939 2409 950
rect 2461 980 2468 991
rect 2802 991 2868 992
rect 2802 980 2809 991
rect 2461 950 2809 980
rect 2461 939 2468 950
rect 2402 938 2468 939
rect 2802 939 2809 950
rect 2861 980 2868 991
rect 3202 991 3268 992
rect 3202 980 3209 991
rect 2861 950 3209 980
rect 2861 939 2868 950
rect 2802 938 2868 939
rect 3202 939 3209 950
rect 3261 980 3268 991
rect 3602 991 3668 992
rect 3602 980 3609 991
rect 3261 950 3609 980
rect 3261 939 3268 950
rect 3202 938 3268 939
rect 3602 939 3609 950
rect 3661 980 3668 991
rect 4002 991 4068 992
rect 4002 980 4009 991
rect 3661 950 4009 980
rect 3661 939 3668 950
rect 3602 938 3668 939
rect 4002 939 4009 950
rect 4061 980 4068 991
rect 4402 991 4468 992
rect 4402 980 4409 991
rect 4061 950 4409 980
rect 4061 939 4068 950
rect 4002 938 4068 939
rect 4402 939 4409 950
rect 4461 980 4468 991
rect 4802 991 4868 992
rect 4802 980 4809 991
rect 4461 950 4809 980
rect 4461 939 4468 950
rect 4402 938 4468 939
rect 4802 939 4809 950
rect 4861 980 4868 991
rect 5202 991 5268 992
rect 5202 980 5209 991
rect 4861 950 5209 980
rect 4861 939 4868 950
rect 4802 938 4868 939
rect 5202 939 5209 950
rect 5261 980 5268 991
rect 5602 991 5668 992
rect 5602 980 5609 991
rect 5261 950 5609 980
rect 5261 939 5268 950
rect 5202 938 5268 939
rect 5602 939 5609 950
rect 5661 980 5668 991
rect 6002 991 6068 992
rect 6002 980 6009 991
rect 5661 950 6009 980
rect 5661 939 5668 950
rect 5602 938 5668 939
rect 6002 939 6009 950
rect 6061 980 6068 991
rect 6402 991 6468 992
rect 6402 980 6409 991
rect 6061 950 6409 980
rect 6061 939 6068 950
rect 6002 938 6068 939
rect 6402 939 6409 950
rect 6461 980 6468 991
rect 6802 991 6868 992
rect 6802 980 6809 991
rect 6461 950 6809 980
rect 6461 939 6468 950
rect 6402 938 6468 939
rect 6802 939 6809 950
rect 6861 980 6868 991
rect 7202 991 7268 992
rect 7202 980 7209 991
rect 6861 950 7209 980
rect 6861 939 6868 950
rect 6802 938 6868 939
rect 7202 939 7209 950
rect 7261 980 7268 991
rect 7602 991 7668 992
rect 7602 980 7609 991
rect 7261 950 7609 980
rect 7261 939 7268 950
rect 7202 938 7268 939
rect 7602 939 7609 950
rect 7661 980 7668 991
rect 8002 991 8068 992
rect 8002 980 8009 991
rect 7661 950 8009 980
rect 7661 939 7668 950
rect 7602 938 7668 939
rect 8002 939 8009 950
rect 8061 980 8068 991
rect 8402 991 8468 992
rect 8402 980 8409 991
rect 8061 950 8409 980
rect 8061 939 8068 950
rect 8002 938 8068 939
rect 8402 939 8409 950
rect 8461 980 8468 991
rect 8802 991 8868 992
rect 8802 980 8809 991
rect 8461 950 8809 980
rect 8461 939 8468 950
rect 8402 938 8468 939
rect 8802 939 8809 950
rect 8861 980 8868 991
rect 9202 991 9268 992
rect 9202 980 9209 991
rect 8861 950 9209 980
rect 8861 939 8868 950
rect 8802 938 8868 939
rect 9202 939 9209 950
rect 9261 980 9268 991
rect 9602 991 9668 992
rect 9602 980 9609 991
rect 9261 950 9609 980
rect 9261 939 9268 950
rect 9202 938 9268 939
rect 9602 939 9609 950
rect 9661 980 9668 991
rect 10002 991 10068 992
rect 10002 980 10009 991
rect 9661 950 10009 980
rect 9661 939 9668 950
rect 9602 938 9668 939
rect 10002 939 10009 950
rect 10061 980 10068 991
rect 10402 991 10468 992
rect 10402 980 10409 991
rect 10061 950 10409 980
rect 10061 939 10068 950
rect 10002 938 10068 939
rect 10402 939 10409 950
rect 10461 980 10468 991
rect 10802 991 10868 992
rect 10802 980 10809 991
rect 10461 950 10809 980
rect 10461 939 10468 950
rect 10402 938 10468 939
rect 10802 939 10809 950
rect 10861 980 10868 991
rect 11202 991 11268 992
rect 11202 980 11209 991
rect 10861 950 11209 980
rect 10861 939 10868 950
rect 10802 938 10868 939
rect 11202 939 11209 950
rect 11261 980 11268 991
rect 11602 991 11668 992
rect 11602 980 11609 991
rect 11261 950 11609 980
rect 11261 939 11268 950
rect 11202 938 11268 939
rect 11602 939 11609 950
rect 11661 980 11668 991
rect 12002 991 12068 992
rect 12002 980 12009 991
rect 11661 950 12009 980
rect 11661 939 11668 950
rect 11602 938 11668 939
rect 12002 939 12009 950
rect 12061 980 12068 991
rect 12402 991 12468 992
rect 12402 980 12409 991
rect 12061 950 12409 980
rect 12061 939 12068 950
rect 12002 938 12068 939
rect 12402 939 12409 950
rect 12461 980 12468 991
rect 12802 991 12868 992
rect 12802 980 12809 991
rect 12461 950 12809 980
rect 12461 939 12468 950
rect 12402 938 12468 939
rect 12802 939 12809 950
rect 12861 980 12868 991
rect 12900 991 12966 992
rect 12900 980 12907 991
rect 12861 950 12907 980
rect 12861 939 12868 950
rect 12802 938 12868 939
rect 12900 939 12907 950
rect 12959 939 12966 991
rect 12900 938 12966 939
rect 202 921 268 922
rect 202 910 209 921
rect 0 880 209 910
rect 202 869 209 880
rect 261 910 268 921
rect 602 921 668 922
rect 602 910 609 921
rect 261 880 609 910
rect 261 869 268 880
rect 202 868 268 869
rect 602 869 609 880
rect 661 910 668 921
rect 1002 921 1068 922
rect 1002 910 1009 921
rect 661 880 1009 910
rect 661 869 668 880
rect 602 868 668 869
rect 1002 869 1009 880
rect 1061 910 1068 921
rect 1402 921 1468 922
rect 1402 910 1409 921
rect 1061 880 1409 910
rect 1061 869 1068 880
rect 1002 868 1068 869
rect 1402 869 1409 880
rect 1461 910 1468 921
rect 1802 921 1868 922
rect 1802 910 1809 921
rect 1461 880 1809 910
rect 1461 869 1468 880
rect 1402 868 1468 869
rect 1802 869 1809 880
rect 1861 910 1868 921
rect 2202 921 2268 922
rect 2202 910 2209 921
rect 1861 880 2209 910
rect 1861 869 1868 880
rect 1802 868 1868 869
rect 2202 869 2209 880
rect 2261 910 2268 921
rect 2602 921 2668 922
rect 2602 910 2609 921
rect 2261 880 2609 910
rect 2261 869 2268 880
rect 2202 868 2268 869
rect 2602 869 2609 880
rect 2661 910 2668 921
rect 3002 921 3068 922
rect 3002 910 3009 921
rect 2661 880 3009 910
rect 2661 869 2668 880
rect 2602 868 2668 869
rect 3002 869 3009 880
rect 3061 910 3068 921
rect 3402 921 3468 922
rect 3402 910 3409 921
rect 3061 880 3409 910
rect 3061 869 3068 880
rect 3002 868 3068 869
rect 3402 869 3409 880
rect 3461 910 3468 921
rect 3802 921 3868 922
rect 3802 910 3809 921
rect 3461 880 3809 910
rect 3461 869 3468 880
rect 3402 868 3468 869
rect 3802 869 3809 880
rect 3861 910 3868 921
rect 4202 921 4268 922
rect 4202 910 4209 921
rect 3861 880 4209 910
rect 3861 869 3868 880
rect 3802 868 3868 869
rect 4202 869 4209 880
rect 4261 910 4268 921
rect 4602 921 4668 922
rect 4602 910 4609 921
rect 4261 880 4609 910
rect 4261 869 4268 880
rect 4202 868 4268 869
rect 4602 869 4609 880
rect 4661 910 4668 921
rect 5002 921 5068 922
rect 5002 910 5009 921
rect 4661 880 5009 910
rect 4661 869 4668 880
rect 4602 868 4668 869
rect 5002 869 5009 880
rect 5061 910 5068 921
rect 5402 921 5468 922
rect 5402 910 5409 921
rect 5061 880 5409 910
rect 5061 869 5068 880
rect 5002 868 5068 869
rect 5402 869 5409 880
rect 5461 910 5468 921
rect 5802 921 5868 922
rect 5802 910 5809 921
rect 5461 880 5809 910
rect 5461 869 5468 880
rect 5402 868 5468 869
rect 5802 869 5809 880
rect 5861 910 5868 921
rect 6202 921 6268 922
rect 6202 910 6209 921
rect 5861 880 6209 910
rect 5861 869 5868 880
rect 5802 868 5868 869
rect 6202 869 6209 880
rect 6261 910 6268 921
rect 6602 921 6668 922
rect 6602 910 6609 921
rect 6261 880 6609 910
rect 6261 869 6268 880
rect 6202 868 6268 869
rect 6602 869 6609 880
rect 6661 910 6668 921
rect 7002 921 7068 922
rect 7002 910 7009 921
rect 6661 880 7009 910
rect 6661 869 6668 880
rect 6602 868 6668 869
rect 7002 869 7009 880
rect 7061 910 7068 921
rect 7402 921 7468 922
rect 7402 910 7409 921
rect 7061 880 7409 910
rect 7061 869 7068 880
rect 7002 868 7068 869
rect 7402 869 7409 880
rect 7461 910 7468 921
rect 7802 921 7868 922
rect 7802 910 7809 921
rect 7461 880 7809 910
rect 7461 869 7468 880
rect 7402 868 7468 869
rect 7802 869 7809 880
rect 7861 910 7868 921
rect 8202 921 8268 922
rect 8202 910 8209 921
rect 7861 880 8209 910
rect 7861 869 7868 880
rect 7802 868 7868 869
rect 8202 869 8209 880
rect 8261 910 8268 921
rect 8602 921 8668 922
rect 8602 910 8609 921
rect 8261 880 8609 910
rect 8261 869 8268 880
rect 8202 868 8268 869
rect 8602 869 8609 880
rect 8661 910 8668 921
rect 9002 921 9068 922
rect 9002 910 9009 921
rect 8661 880 9009 910
rect 8661 869 8668 880
rect 8602 868 8668 869
rect 9002 869 9009 880
rect 9061 910 9068 921
rect 9402 921 9468 922
rect 9402 910 9409 921
rect 9061 880 9409 910
rect 9061 869 9068 880
rect 9002 868 9068 869
rect 9402 869 9409 880
rect 9461 910 9468 921
rect 9802 921 9868 922
rect 9802 910 9809 921
rect 9461 880 9809 910
rect 9461 869 9468 880
rect 9402 868 9468 869
rect 9802 869 9809 880
rect 9861 910 9868 921
rect 10202 921 10268 922
rect 10202 910 10209 921
rect 9861 880 10209 910
rect 9861 869 9868 880
rect 9802 868 9868 869
rect 10202 869 10209 880
rect 10261 910 10268 921
rect 10602 921 10668 922
rect 10602 910 10609 921
rect 10261 880 10609 910
rect 10261 869 10268 880
rect 10202 868 10268 869
rect 10602 869 10609 880
rect 10661 910 10668 921
rect 11002 921 11068 922
rect 11002 910 11009 921
rect 10661 880 11009 910
rect 10661 869 10668 880
rect 10602 868 10668 869
rect 11002 869 11009 880
rect 11061 910 11068 921
rect 11402 921 11468 922
rect 11402 910 11409 921
rect 11061 880 11409 910
rect 11061 869 11068 880
rect 11002 868 11068 869
rect 11402 869 11409 880
rect 11461 910 11468 921
rect 11802 921 11868 922
rect 11802 910 11809 921
rect 11461 880 11809 910
rect 11461 869 11468 880
rect 11402 868 11468 869
rect 11802 869 11809 880
rect 11861 910 11868 921
rect 12202 921 12268 922
rect 12202 910 12209 921
rect 11861 880 12209 910
rect 11861 869 11868 880
rect 11802 868 11868 869
rect 12202 869 12209 880
rect 12261 910 12268 921
rect 12602 921 12668 922
rect 12602 910 12609 921
rect 12261 880 12609 910
rect 12261 869 12268 880
rect 12202 868 12268 869
rect 12602 869 12609 880
rect 12661 910 12668 921
rect 13104 921 13170 922
rect 13104 910 13111 921
rect 12661 880 13111 910
rect 12661 869 12668 880
rect 12602 868 12668 869
rect 13104 869 13111 880
rect 13163 869 13170 921
rect 13104 868 13170 869
rect 2 851 68 852
rect 2 840 9 851
rect 0 810 9 840
rect 2 799 9 810
rect 61 840 68 851
rect 402 851 468 852
rect 402 840 409 851
rect 61 810 409 840
rect 61 799 68 810
rect 2 798 68 799
rect 402 799 409 810
rect 461 840 468 851
rect 802 851 868 852
rect 802 840 809 851
rect 461 810 809 840
rect 461 799 468 810
rect 402 798 468 799
rect 802 799 809 810
rect 861 840 868 851
rect 1202 851 1268 852
rect 1202 840 1209 851
rect 861 810 1209 840
rect 861 799 868 810
rect 802 798 868 799
rect 1202 799 1209 810
rect 1261 840 1268 851
rect 1602 851 1668 852
rect 1602 840 1609 851
rect 1261 810 1609 840
rect 1261 799 1268 810
rect 1202 798 1268 799
rect 1602 799 1609 810
rect 1661 840 1668 851
rect 2002 851 2068 852
rect 2002 840 2009 851
rect 1661 810 2009 840
rect 1661 799 1668 810
rect 1602 798 1668 799
rect 2002 799 2009 810
rect 2061 840 2068 851
rect 2402 851 2468 852
rect 2402 840 2409 851
rect 2061 810 2409 840
rect 2061 799 2068 810
rect 2002 798 2068 799
rect 2402 799 2409 810
rect 2461 840 2468 851
rect 2802 851 2868 852
rect 2802 840 2809 851
rect 2461 810 2809 840
rect 2461 799 2468 810
rect 2402 798 2468 799
rect 2802 799 2809 810
rect 2861 840 2868 851
rect 3202 851 3268 852
rect 3202 840 3209 851
rect 2861 810 3209 840
rect 2861 799 2868 810
rect 2802 798 2868 799
rect 3202 799 3209 810
rect 3261 840 3268 851
rect 3602 851 3668 852
rect 3602 840 3609 851
rect 3261 810 3609 840
rect 3261 799 3268 810
rect 3202 798 3268 799
rect 3602 799 3609 810
rect 3661 840 3668 851
rect 4002 851 4068 852
rect 4002 840 4009 851
rect 3661 810 4009 840
rect 3661 799 3668 810
rect 3602 798 3668 799
rect 4002 799 4009 810
rect 4061 840 4068 851
rect 4402 851 4468 852
rect 4402 840 4409 851
rect 4061 810 4409 840
rect 4061 799 4068 810
rect 4002 798 4068 799
rect 4402 799 4409 810
rect 4461 840 4468 851
rect 4802 851 4868 852
rect 4802 840 4809 851
rect 4461 810 4809 840
rect 4461 799 4468 810
rect 4402 798 4468 799
rect 4802 799 4809 810
rect 4861 840 4868 851
rect 5202 851 5268 852
rect 5202 840 5209 851
rect 4861 810 5209 840
rect 4861 799 4868 810
rect 4802 798 4868 799
rect 5202 799 5209 810
rect 5261 840 5268 851
rect 5602 851 5668 852
rect 5602 840 5609 851
rect 5261 810 5609 840
rect 5261 799 5268 810
rect 5202 798 5268 799
rect 5602 799 5609 810
rect 5661 840 5668 851
rect 6002 851 6068 852
rect 6002 840 6009 851
rect 5661 810 6009 840
rect 5661 799 5668 810
rect 5602 798 5668 799
rect 6002 799 6009 810
rect 6061 840 6068 851
rect 6402 851 6468 852
rect 6402 840 6409 851
rect 6061 810 6409 840
rect 6061 799 6068 810
rect 6002 798 6068 799
rect 6402 799 6409 810
rect 6461 840 6468 851
rect 6802 851 6868 852
rect 6802 840 6809 851
rect 6461 810 6809 840
rect 6461 799 6468 810
rect 6402 798 6468 799
rect 6802 799 6809 810
rect 6861 840 6868 851
rect 7202 851 7268 852
rect 7202 840 7209 851
rect 6861 810 7209 840
rect 6861 799 6868 810
rect 6802 798 6868 799
rect 7202 799 7209 810
rect 7261 840 7268 851
rect 7602 851 7668 852
rect 7602 840 7609 851
rect 7261 810 7609 840
rect 7261 799 7268 810
rect 7202 798 7268 799
rect 7602 799 7609 810
rect 7661 840 7668 851
rect 8002 851 8068 852
rect 8002 840 8009 851
rect 7661 810 8009 840
rect 7661 799 7668 810
rect 7602 798 7668 799
rect 8002 799 8009 810
rect 8061 840 8068 851
rect 8402 851 8468 852
rect 8402 840 8409 851
rect 8061 810 8409 840
rect 8061 799 8068 810
rect 8002 798 8068 799
rect 8402 799 8409 810
rect 8461 840 8468 851
rect 8802 851 8868 852
rect 8802 840 8809 851
rect 8461 810 8809 840
rect 8461 799 8468 810
rect 8402 798 8468 799
rect 8802 799 8809 810
rect 8861 840 8868 851
rect 9202 851 9268 852
rect 9202 840 9209 851
rect 8861 810 9209 840
rect 8861 799 8868 810
rect 8802 798 8868 799
rect 9202 799 9209 810
rect 9261 840 9268 851
rect 9602 851 9668 852
rect 9602 840 9609 851
rect 9261 810 9609 840
rect 9261 799 9268 810
rect 9202 798 9268 799
rect 9602 799 9609 810
rect 9661 840 9668 851
rect 10002 851 10068 852
rect 10002 840 10009 851
rect 9661 810 10009 840
rect 9661 799 9668 810
rect 9602 798 9668 799
rect 10002 799 10009 810
rect 10061 840 10068 851
rect 10402 851 10468 852
rect 10402 840 10409 851
rect 10061 810 10409 840
rect 10061 799 10068 810
rect 10002 798 10068 799
rect 10402 799 10409 810
rect 10461 840 10468 851
rect 10802 851 10868 852
rect 10802 840 10809 851
rect 10461 810 10809 840
rect 10461 799 10468 810
rect 10402 798 10468 799
rect 10802 799 10809 810
rect 10861 840 10868 851
rect 11202 851 11268 852
rect 11202 840 11209 851
rect 10861 810 11209 840
rect 10861 799 10868 810
rect 10802 798 10868 799
rect 11202 799 11209 810
rect 11261 840 11268 851
rect 11602 851 11668 852
rect 11602 840 11609 851
rect 11261 810 11609 840
rect 11261 799 11268 810
rect 11202 798 11268 799
rect 11602 799 11609 810
rect 11661 840 11668 851
rect 12002 851 12068 852
rect 12002 840 12009 851
rect 11661 810 12009 840
rect 11661 799 11668 810
rect 11602 798 11668 799
rect 12002 799 12009 810
rect 12061 840 12068 851
rect 12402 851 12468 852
rect 12402 840 12409 851
rect 12061 810 12409 840
rect 12061 799 12068 810
rect 12002 798 12068 799
rect 12402 799 12409 810
rect 12461 840 12468 851
rect 12802 851 12868 852
rect 12802 840 12809 851
rect 12461 810 12809 840
rect 12461 799 12468 810
rect 12402 798 12468 799
rect 12802 799 12809 810
rect 12861 840 12868 851
rect 12900 851 12966 852
rect 12900 840 12907 851
rect 12861 810 12907 840
rect 12861 799 12868 810
rect 12802 798 12868 799
rect 12900 799 12907 810
rect 12959 799 12966 851
rect 12900 798 12966 799
rect 202 781 268 782
rect 202 770 209 781
rect 0 740 209 770
rect 202 729 209 740
rect 261 770 268 781
rect 602 781 668 782
rect 602 770 609 781
rect 261 740 609 770
rect 261 729 268 740
rect 202 728 268 729
rect 602 729 609 740
rect 661 770 668 781
rect 1002 781 1068 782
rect 1002 770 1009 781
rect 661 740 1009 770
rect 661 729 668 740
rect 602 728 668 729
rect 1002 729 1009 740
rect 1061 770 1068 781
rect 1402 781 1468 782
rect 1402 770 1409 781
rect 1061 740 1409 770
rect 1061 729 1068 740
rect 1002 728 1068 729
rect 1402 729 1409 740
rect 1461 770 1468 781
rect 1802 781 1868 782
rect 1802 770 1809 781
rect 1461 740 1809 770
rect 1461 729 1468 740
rect 1402 728 1468 729
rect 1802 729 1809 740
rect 1861 770 1868 781
rect 2202 781 2268 782
rect 2202 770 2209 781
rect 1861 740 2209 770
rect 1861 729 1868 740
rect 1802 728 1868 729
rect 2202 729 2209 740
rect 2261 770 2268 781
rect 2602 781 2668 782
rect 2602 770 2609 781
rect 2261 740 2609 770
rect 2261 729 2268 740
rect 2202 728 2268 729
rect 2602 729 2609 740
rect 2661 770 2668 781
rect 3002 781 3068 782
rect 3002 770 3009 781
rect 2661 740 3009 770
rect 2661 729 2668 740
rect 2602 728 2668 729
rect 3002 729 3009 740
rect 3061 770 3068 781
rect 3402 781 3468 782
rect 3402 770 3409 781
rect 3061 740 3409 770
rect 3061 729 3068 740
rect 3002 728 3068 729
rect 3402 729 3409 740
rect 3461 770 3468 781
rect 3802 781 3868 782
rect 3802 770 3809 781
rect 3461 740 3809 770
rect 3461 729 3468 740
rect 3402 728 3468 729
rect 3802 729 3809 740
rect 3861 770 3868 781
rect 4202 781 4268 782
rect 4202 770 4209 781
rect 3861 740 4209 770
rect 3861 729 3868 740
rect 3802 728 3868 729
rect 4202 729 4209 740
rect 4261 770 4268 781
rect 4602 781 4668 782
rect 4602 770 4609 781
rect 4261 740 4609 770
rect 4261 729 4268 740
rect 4202 728 4268 729
rect 4602 729 4609 740
rect 4661 770 4668 781
rect 5002 781 5068 782
rect 5002 770 5009 781
rect 4661 740 5009 770
rect 4661 729 4668 740
rect 4602 728 4668 729
rect 5002 729 5009 740
rect 5061 770 5068 781
rect 5402 781 5468 782
rect 5402 770 5409 781
rect 5061 740 5409 770
rect 5061 729 5068 740
rect 5002 728 5068 729
rect 5402 729 5409 740
rect 5461 770 5468 781
rect 5802 781 5868 782
rect 5802 770 5809 781
rect 5461 740 5809 770
rect 5461 729 5468 740
rect 5402 728 5468 729
rect 5802 729 5809 740
rect 5861 770 5868 781
rect 6202 781 6268 782
rect 6202 770 6209 781
rect 5861 740 6209 770
rect 5861 729 5868 740
rect 5802 728 5868 729
rect 6202 729 6209 740
rect 6261 770 6268 781
rect 6602 781 6668 782
rect 6602 770 6609 781
rect 6261 740 6609 770
rect 6261 729 6268 740
rect 6202 728 6268 729
rect 6602 729 6609 740
rect 6661 770 6668 781
rect 7002 781 7068 782
rect 7002 770 7009 781
rect 6661 740 7009 770
rect 6661 729 6668 740
rect 6602 728 6668 729
rect 7002 729 7009 740
rect 7061 770 7068 781
rect 7402 781 7468 782
rect 7402 770 7409 781
rect 7061 740 7409 770
rect 7061 729 7068 740
rect 7002 728 7068 729
rect 7402 729 7409 740
rect 7461 770 7468 781
rect 7802 781 7868 782
rect 7802 770 7809 781
rect 7461 740 7809 770
rect 7461 729 7468 740
rect 7402 728 7468 729
rect 7802 729 7809 740
rect 7861 770 7868 781
rect 8202 781 8268 782
rect 8202 770 8209 781
rect 7861 740 8209 770
rect 7861 729 7868 740
rect 7802 728 7868 729
rect 8202 729 8209 740
rect 8261 770 8268 781
rect 8602 781 8668 782
rect 8602 770 8609 781
rect 8261 740 8609 770
rect 8261 729 8268 740
rect 8202 728 8268 729
rect 8602 729 8609 740
rect 8661 770 8668 781
rect 9002 781 9068 782
rect 9002 770 9009 781
rect 8661 740 9009 770
rect 8661 729 8668 740
rect 8602 728 8668 729
rect 9002 729 9009 740
rect 9061 770 9068 781
rect 9402 781 9468 782
rect 9402 770 9409 781
rect 9061 740 9409 770
rect 9061 729 9068 740
rect 9002 728 9068 729
rect 9402 729 9409 740
rect 9461 770 9468 781
rect 9802 781 9868 782
rect 9802 770 9809 781
rect 9461 740 9809 770
rect 9461 729 9468 740
rect 9402 728 9468 729
rect 9802 729 9809 740
rect 9861 770 9868 781
rect 10202 781 10268 782
rect 10202 770 10209 781
rect 9861 740 10209 770
rect 9861 729 9868 740
rect 9802 728 9868 729
rect 10202 729 10209 740
rect 10261 770 10268 781
rect 10602 781 10668 782
rect 10602 770 10609 781
rect 10261 740 10609 770
rect 10261 729 10268 740
rect 10202 728 10268 729
rect 10602 729 10609 740
rect 10661 770 10668 781
rect 11002 781 11068 782
rect 11002 770 11009 781
rect 10661 740 11009 770
rect 10661 729 10668 740
rect 10602 728 10668 729
rect 11002 729 11009 740
rect 11061 770 11068 781
rect 11402 781 11468 782
rect 11402 770 11409 781
rect 11061 740 11409 770
rect 11061 729 11068 740
rect 11002 728 11068 729
rect 11402 729 11409 740
rect 11461 770 11468 781
rect 11802 781 11868 782
rect 11802 770 11809 781
rect 11461 740 11809 770
rect 11461 729 11468 740
rect 11402 728 11468 729
rect 11802 729 11809 740
rect 11861 770 11868 781
rect 12202 781 12268 782
rect 12202 770 12209 781
rect 11861 740 12209 770
rect 11861 729 11868 740
rect 11802 728 11868 729
rect 12202 729 12209 740
rect 12261 770 12268 781
rect 12602 781 12668 782
rect 12602 770 12609 781
rect 12261 740 12609 770
rect 12261 729 12268 740
rect 12202 728 12268 729
rect 12602 729 12609 740
rect 12661 770 12668 781
rect 13104 781 13170 782
rect 13104 770 13111 781
rect 12661 740 13111 770
rect 12661 729 12668 740
rect 12602 728 12668 729
rect 13104 729 13111 740
rect 13163 729 13170 781
rect 13104 728 13170 729
rect 2 711 68 712
rect 2 700 9 711
rect 0 670 9 700
rect 2 659 9 670
rect 61 700 68 711
rect 402 711 468 712
rect 402 700 409 711
rect 61 670 409 700
rect 61 659 68 670
rect 2 658 68 659
rect 402 659 409 670
rect 461 700 468 711
rect 802 711 868 712
rect 802 700 809 711
rect 461 670 809 700
rect 461 659 468 670
rect 402 658 468 659
rect 802 659 809 670
rect 861 700 868 711
rect 1202 711 1268 712
rect 1202 700 1209 711
rect 861 670 1209 700
rect 861 659 868 670
rect 802 658 868 659
rect 1202 659 1209 670
rect 1261 700 1268 711
rect 1602 711 1668 712
rect 1602 700 1609 711
rect 1261 670 1609 700
rect 1261 659 1268 670
rect 1202 658 1268 659
rect 1602 659 1609 670
rect 1661 700 1668 711
rect 2002 711 2068 712
rect 2002 700 2009 711
rect 1661 670 2009 700
rect 1661 659 1668 670
rect 1602 658 1668 659
rect 2002 659 2009 670
rect 2061 700 2068 711
rect 2402 711 2468 712
rect 2402 700 2409 711
rect 2061 670 2409 700
rect 2061 659 2068 670
rect 2002 658 2068 659
rect 2402 659 2409 670
rect 2461 700 2468 711
rect 2802 711 2868 712
rect 2802 700 2809 711
rect 2461 670 2809 700
rect 2461 659 2468 670
rect 2402 658 2468 659
rect 2802 659 2809 670
rect 2861 700 2868 711
rect 3202 711 3268 712
rect 3202 700 3209 711
rect 2861 670 3209 700
rect 2861 659 2868 670
rect 2802 658 2868 659
rect 3202 659 3209 670
rect 3261 700 3268 711
rect 3602 711 3668 712
rect 3602 700 3609 711
rect 3261 670 3609 700
rect 3261 659 3268 670
rect 3202 658 3268 659
rect 3602 659 3609 670
rect 3661 700 3668 711
rect 4002 711 4068 712
rect 4002 700 4009 711
rect 3661 670 4009 700
rect 3661 659 3668 670
rect 3602 658 3668 659
rect 4002 659 4009 670
rect 4061 700 4068 711
rect 4402 711 4468 712
rect 4402 700 4409 711
rect 4061 670 4409 700
rect 4061 659 4068 670
rect 4002 658 4068 659
rect 4402 659 4409 670
rect 4461 700 4468 711
rect 4802 711 4868 712
rect 4802 700 4809 711
rect 4461 670 4809 700
rect 4461 659 4468 670
rect 4402 658 4468 659
rect 4802 659 4809 670
rect 4861 700 4868 711
rect 5202 711 5268 712
rect 5202 700 5209 711
rect 4861 670 5209 700
rect 4861 659 4868 670
rect 4802 658 4868 659
rect 5202 659 5209 670
rect 5261 700 5268 711
rect 5602 711 5668 712
rect 5602 700 5609 711
rect 5261 670 5609 700
rect 5261 659 5268 670
rect 5202 658 5268 659
rect 5602 659 5609 670
rect 5661 700 5668 711
rect 6002 711 6068 712
rect 6002 700 6009 711
rect 5661 670 6009 700
rect 5661 659 5668 670
rect 5602 658 5668 659
rect 6002 659 6009 670
rect 6061 700 6068 711
rect 6402 711 6468 712
rect 6402 700 6409 711
rect 6061 670 6409 700
rect 6061 659 6068 670
rect 6002 658 6068 659
rect 6402 659 6409 670
rect 6461 700 6468 711
rect 6802 711 6868 712
rect 6802 700 6809 711
rect 6461 670 6809 700
rect 6461 659 6468 670
rect 6402 658 6468 659
rect 6802 659 6809 670
rect 6861 700 6868 711
rect 7202 711 7268 712
rect 7202 700 7209 711
rect 6861 670 7209 700
rect 6861 659 6868 670
rect 6802 658 6868 659
rect 7202 659 7209 670
rect 7261 700 7268 711
rect 7602 711 7668 712
rect 7602 700 7609 711
rect 7261 670 7609 700
rect 7261 659 7268 670
rect 7202 658 7268 659
rect 7602 659 7609 670
rect 7661 700 7668 711
rect 8002 711 8068 712
rect 8002 700 8009 711
rect 7661 670 8009 700
rect 7661 659 7668 670
rect 7602 658 7668 659
rect 8002 659 8009 670
rect 8061 700 8068 711
rect 8402 711 8468 712
rect 8402 700 8409 711
rect 8061 670 8409 700
rect 8061 659 8068 670
rect 8002 658 8068 659
rect 8402 659 8409 670
rect 8461 700 8468 711
rect 8802 711 8868 712
rect 8802 700 8809 711
rect 8461 670 8809 700
rect 8461 659 8468 670
rect 8402 658 8468 659
rect 8802 659 8809 670
rect 8861 700 8868 711
rect 9202 711 9268 712
rect 9202 700 9209 711
rect 8861 670 9209 700
rect 8861 659 8868 670
rect 8802 658 8868 659
rect 9202 659 9209 670
rect 9261 700 9268 711
rect 9602 711 9668 712
rect 9602 700 9609 711
rect 9261 670 9609 700
rect 9261 659 9268 670
rect 9202 658 9268 659
rect 9602 659 9609 670
rect 9661 700 9668 711
rect 10002 711 10068 712
rect 10002 700 10009 711
rect 9661 670 10009 700
rect 9661 659 9668 670
rect 9602 658 9668 659
rect 10002 659 10009 670
rect 10061 700 10068 711
rect 10402 711 10468 712
rect 10402 700 10409 711
rect 10061 670 10409 700
rect 10061 659 10068 670
rect 10002 658 10068 659
rect 10402 659 10409 670
rect 10461 700 10468 711
rect 10802 711 10868 712
rect 10802 700 10809 711
rect 10461 670 10809 700
rect 10461 659 10468 670
rect 10402 658 10468 659
rect 10802 659 10809 670
rect 10861 700 10868 711
rect 11202 711 11268 712
rect 11202 700 11209 711
rect 10861 670 11209 700
rect 10861 659 10868 670
rect 10802 658 10868 659
rect 11202 659 11209 670
rect 11261 700 11268 711
rect 11602 711 11668 712
rect 11602 700 11609 711
rect 11261 670 11609 700
rect 11261 659 11268 670
rect 11202 658 11268 659
rect 11602 659 11609 670
rect 11661 700 11668 711
rect 12002 711 12068 712
rect 12002 700 12009 711
rect 11661 670 12009 700
rect 11661 659 11668 670
rect 11602 658 11668 659
rect 12002 659 12009 670
rect 12061 700 12068 711
rect 12402 711 12468 712
rect 12402 700 12409 711
rect 12061 670 12409 700
rect 12061 659 12068 670
rect 12002 658 12068 659
rect 12402 659 12409 670
rect 12461 700 12468 711
rect 12802 711 12868 712
rect 12802 700 12809 711
rect 12461 670 12809 700
rect 12461 659 12468 670
rect 12402 658 12468 659
rect 12802 659 12809 670
rect 12861 700 12868 711
rect 12900 711 12966 712
rect 12900 700 12907 711
rect 12861 670 12907 700
rect 12861 659 12868 670
rect 12802 658 12868 659
rect 12900 659 12907 670
rect 12959 659 12966 711
rect 12900 658 12966 659
rect 202 641 268 642
rect 202 630 209 641
rect 0 600 209 630
rect 202 589 209 600
rect 261 630 268 641
rect 602 641 668 642
rect 602 630 609 641
rect 261 600 609 630
rect 261 589 268 600
rect 202 588 268 589
rect 602 589 609 600
rect 661 630 668 641
rect 1002 641 1068 642
rect 1002 630 1009 641
rect 661 600 1009 630
rect 661 589 668 600
rect 602 588 668 589
rect 1002 589 1009 600
rect 1061 630 1068 641
rect 1402 641 1468 642
rect 1402 630 1409 641
rect 1061 600 1409 630
rect 1061 589 1068 600
rect 1002 588 1068 589
rect 1402 589 1409 600
rect 1461 630 1468 641
rect 1802 641 1868 642
rect 1802 630 1809 641
rect 1461 600 1809 630
rect 1461 589 1468 600
rect 1402 588 1468 589
rect 1802 589 1809 600
rect 1861 630 1868 641
rect 2202 641 2268 642
rect 2202 630 2209 641
rect 1861 600 2209 630
rect 1861 589 1868 600
rect 1802 588 1868 589
rect 2202 589 2209 600
rect 2261 630 2268 641
rect 2602 641 2668 642
rect 2602 630 2609 641
rect 2261 600 2609 630
rect 2261 589 2268 600
rect 2202 588 2268 589
rect 2602 589 2609 600
rect 2661 630 2668 641
rect 3002 641 3068 642
rect 3002 630 3009 641
rect 2661 600 3009 630
rect 2661 589 2668 600
rect 2602 588 2668 589
rect 3002 589 3009 600
rect 3061 630 3068 641
rect 3402 641 3468 642
rect 3402 630 3409 641
rect 3061 600 3409 630
rect 3061 589 3068 600
rect 3002 588 3068 589
rect 3402 589 3409 600
rect 3461 630 3468 641
rect 3802 641 3868 642
rect 3802 630 3809 641
rect 3461 600 3809 630
rect 3461 589 3468 600
rect 3402 588 3468 589
rect 3802 589 3809 600
rect 3861 630 3868 641
rect 4202 641 4268 642
rect 4202 630 4209 641
rect 3861 600 4209 630
rect 3861 589 3868 600
rect 3802 588 3868 589
rect 4202 589 4209 600
rect 4261 630 4268 641
rect 4602 641 4668 642
rect 4602 630 4609 641
rect 4261 600 4609 630
rect 4261 589 4268 600
rect 4202 588 4268 589
rect 4602 589 4609 600
rect 4661 630 4668 641
rect 5002 641 5068 642
rect 5002 630 5009 641
rect 4661 600 5009 630
rect 4661 589 4668 600
rect 4602 588 4668 589
rect 5002 589 5009 600
rect 5061 630 5068 641
rect 5402 641 5468 642
rect 5402 630 5409 641
rect 5061 600 5409 630
rect 5061 589 5068 600
rect 5002 588 5068 589
rect 5402 589 5409 600
rect 5461 630 5468 641
rect 5802 641 5868 642
rect 5802 630 5809 641
rect 5461 600 5809 630
rect 5461 589 5468 600
rect 5402 588 5468 589
rect 5802 589 5809 600
rect 5861 630 5868 641
rect 6202 641 6268 642
rect 6202 630 6209 641
rect 5861 600 6209 630
rect 5861 589 5868 600
rect 5802 588 5868 589
rect 6202 589 6209 600
rect 6261 630 6268 641
rect 6602 641 6668 642
rect 6602 630 6609 641
rect 6261 600 6609 630
rect 6261 589 6268 600
rect 6202 588 6268 589
rect 6602 589 6609 600
rect 6661 630 6668 641
rect 7002 641 7068 642
rect 7002 630 7009 641
rect 6661 600 7009 630
rect 6661 589 6668 600
rect 6602 588 6668 589
rect 7002 589 7009 600
rect 7061 630 7068 641
rect 7402 641 7468 642
rect 7402 630 7409 641
rect 7061 600 7409 630
rect 7061 589 7068 600
rect 7002 588 7068 589
rect 7402 589 7409 600
rect 7461 630 7468 641
rect 7802 641 7868 642
rect 7802 630 7809 641
rect 7461 600 7809 630
rect 7461 589 7468 600
rect 7402 588 7468 589
rect 7802 589 7809 600
rect 7861 630 7868 641
rect 8202 641 8268 642
rect 8202 630 8209 641
rect 7861 600 8209 630
rect 7861 589 7868 600
rect 7802 588 7868 589
rect 8202 589 8209 600
rect 8261 630 8268 641
rect 8602 641 8668 642
rect 8602 630 8609 641
rect 8261 600 8609 630
rect 8261 589 8268 600
rect 8202 588 8268 589
rect 8602 589 8609 600
rect 8661 630 8668 641
rect 9002 641 9068 642
rect 9002 630 9009 641
rect 8661 600 9009 630
rect 8661 589 8668 600
rect 8602 588 8668 589
rect 9002 589 9009 600
rect 9061 630 9068 641
rect 9402 641 9468 642
rect 9402 630 9409 641
rect 9061 600 9409 630
rect 9061 589 9068 600
rect 9002 588 9068 589
rect 9402 589 9409 600
rect 9461 630 9468 641
rect 9802 641 9868 642
rect 9802 630 9809 641
rect 9461 600 9809 630
rect 9461 589 9468 600
rect 9402 588 9468 589
rect 9802 589 9809 600
rect 9861 630 9868 641
rect 10202 641 10268 642
rect 10202 630 10209 641
rect 9861 600 10209 630
rect 9861 589 9868 600
rect 9802 588 9868 589
rect 10202 589 10209 600
rect 10261 630 10268 641
rect 10602 641 10668 642
rect 10602 630 10609 641
rect 10261 600 10609 630
rect 10261 589 10268 600
rect 10202 588 10268 589
rect 10602 589 10609 600
rect 10661 630 10668 641
rect 11002 641 11068 642
rect 11002 630 11009 641
rect 10661 600 11009 630
rect 10661 589 10668 600
rect 10602 588 10668 589
rect 11002 589 11009 600
rect 11061 630 11068 641
rect 11402 641 11468 642
rect 11402 630 11409 641
rect 11061 600 11409 630
rect 11061 589 11068 600
rect 11002 588 11068 589
rect 11402 589 11409 600
rect 11461 630 11468 641
rect 11802 641 11868 642
rect 11802 630 11809 641
rect 11461 600 11809 630
rect 11461 589 11468 600
rect 11402 588 11468 589
rect 11802 589 11809 600
rect 11861 630 11868 641
rect 12202 641 12268 642
rect 12202 630 12209 641
rect 11861 600 12209 630
rect 11861 589 11868 600
rect 11802 588 11868 589
rect 12202 589 12209 600
rect 12261 630 12268 641
rect 12602 641 12668 642
rect 12602 630 12609 641
rect 12261 600 12609 630
rect 12261 589 12268 600
rect 12202 588 12268 589
rect 12602 589 12609 600
rect 12661 630 12668 641
rect 13104 641 13170 642
rect 13104 630 13111 641
rect 12661 600 13111 630
rect 12661 589 12668 600
rect 12602 588 12668 589
rect 13104 589 13111 600
rect 13163 589 13170 641
rect 13104 588 13170 589
rect 2 571 68 572
rect 2 560 9 571
rect 0 530 9 560
rect 2 519 9 530
rect 61 560 68 571
rect 402 571 468 572
rect 402 560 409 571
rect 61 530 409 560
rect 61 519 68 530
rect 2 518 68 519
rect 402 519 409 530
rect 461 560 468 571
rect 802 571 868 572
rect 802 560 809 571
rect 461 530 809 560
rect 461 519 468 530
rect 402 518 468 519
rect 802 519 809 530
rect 861 560 868 571
rect 1202 571 1268 572
rect 1202 560 1209 571
rect 861 530 1209 560
rect 861 519 868 530
rect 802 518 868 519
rect 1202 519 1209 530
rect 1261 560 1268 571
rect 1602 571 1668 572
rect 1602 560 1609 571
rect 1261 530 1609 560
rect 1261 519 1268 530
rect 1202 518 1268 519
rect 1602 519 1609 530
rect 1661 560 1668 571
rect 2002 571 2068 572
rect 2002 560 2009 571
rect 1661 530 2009 560
rect 1661 519 1668 530
rect 1602 518 1668 519
rect 2002 519 2009 530
rect 2061 560 2068 571
rect 2402 571 2468 572
rect 2402 560 2409 571
rect 2061 530 2409 560
rect 2061 519 2068 530
rect 2002 518 2068 519
rect 2402 519 2409 530
rect 2461 560 2468 571
rect 2802 571 2868 572
rect 2802 560 2809 571
rect 2461 530 2809 560
rect 2461 519 2468 530
rect 2402 518 2468 519
rect 2802 519 2809 530
rect 2861 560 2868 571
rect 3202 571 3268 572
rect 3202 560 3209 571
rect 2861 530 3209 560
rect 2861 519 2868 530
rect 2802 518 2868 519
rect 3202 519 3209 530
rect 3261 560 3268 571
rect 3602 571 3668 572
rect 3602 560 3609 571
rect 3261 530 3609 560
rect 3261 519 3268 530
rect 3202 518 3268 519
rect 3602 519 3609 530
rect 3661 560 3668 571
rect 4002 571 4068 572
rect 4002 560 4009 571
rect 3661 530 4009 560
rect 3661 519 3668 530
rect 3602 518 3668 519
rect 4002 519 4009 530
rect 4061 560 4068 571
rect 4402 571 4468 572
rect 4402 560 4409 571
rect 4061 530 4409 560
rect 4061 519 4068 530
rect 4002 518 4068 519
rect 4402 519 4409 530
rect 4461 560 4468 571
rect 4802 571 4868 572
rect 4802 560 4809 571
rect 4461 530 4809 560
rect 4461 519 4468 530
rect 4402 518 4468 519
rect 4802 519 4809 530
rect 4861 560 4868 571
rect 5202 571 5268 572
rect 5202 560 5209 571
rect 4861 530 5209 560
rect 4861 519 4868 530
rect 4802 518 4868 519
rect 5202 519 5209 530
rect 5261 560 5268 571
rect 5602 571 5668 572
rect 5602 560 5609 571
rect 5261 530 5609 560
rect 5261 519 5268 530
rect 5202 518 5268 519
rect 5602 519 5609 530
rect 5661 560 5668 571
rect 6002 571 6068 572
rect 6002 560 6009 571
rect 5661 530 6009 560
rect 5661 519 5668 530
rect 5602 518 5668 519
rect 6002 519 6009 530
rect 6061 560 6068 571
rect 6402 571 6468 572
rect 6402 560 6409 571
rect 6061 530 6409 560
rect 6061 519 6068 530
rect 6002 518 6068 519
rect 6402 519 6409 530
rect 6461 560 6468 571
rect 6802 571 6868 572
rect 6802 560 6809 571
rect 6461 530 6809 560
rect 6461 519 6468 530
rect 6402 518 6468 519
rect 6802 519 6809 530
rect 6861 560 6868 571
rect 7202 571 7268 572
rect 7202 560 7209 571
rect 6861 530 7209 560
rect 6861 519 6868 530
rect 6802 518 6868 519
rect 7202 519 7209 530
rect 7261 560 7268 571
rect 7602 571 7668 572
rect 7602 560 7609 571
rect 7261 530 7609 560
rect 7261 519 7268 530
rect 7202 518 7268 519
rect 7602 519 7609 530
rect 7661 560 7668 571
rect 8002 571 8068 572
rect 8002 560 8009 571
rect 7661 530 8009 560
rect 7661 519 7668 530
rect 7602 518 7668 519
rect 8002 519 8009 530
rect 8061 560 8068 571
rect 8402 571 8468 572
rect 8402 560 8409 571
rect 8061 530 8409 560
rect 8061 519 8068 530
rect 8002 518 8068 519
rect 8402 519 8409 530
rect 8461 560 8468 571
rect 8802 571 8868 572
rect 8802 560 8809 571
rect 8461 530 8809 560
rect 8461 519 8468 530
rect 8402 518 8468 519
rect 8802 519 8809 530
rect 8861 560 8868 571
rect 9202 571 9268 572
rect 9202 560 9209 571
rect 8861 530 9209 560
rect 8861 519 8868 530
rect 8802 518 8868 519
rect 9202 519 9209 530
rect 9261 560 9268 571
rect 9602 571 9668 572
rect 9602 560 9609 571
rect 9261 530 9609 560
rect 9261 519 9268 530
rect 9202 518 9268 519
rect 9602 519 9609 530
rect 9661 560 9668 571
rect 10002 571 10068 572
rect 10002 560 10009 571
rect 9661 530 10009 560
rect 9661 519 9668 530
rect 9602 518 9668 519
rect 10002 519 10009 530
rect 10061 560 10068 571
rect 10402 571 10468 572
rect 10402 560 10409 571
rect 10061 530 10409 560
rect 10061 519 10068 530
rect 10002 518 10068 519
rect 10402 519 10409 530
rect 10461 560 10468 571
rect 10802 571 10868 572
rect 10802 560 10809 571
rect 10461 530 10809 560
rect 10461 519 10468 530
rect 10402 518 10468 519
rect 10802 519 10809 530
rect 10861 560 10868 571
rect 11202 571 11268 572
rect 11202 560 11209 571
rect 10861 530 11209 560
rect 10861 519 10868 530
rect 10802 518 10868 519
rect 11202 519 11209 530
rect 11261 560 11268 571
rect 11602 571 11668 572
rect 11602 560 11609 571
rect 11261 530 11609 560
rect 11261 519 11268 530
rect 11202 518 11268 519
rect 11602 519 11609 530
rect 11661 560 11668 571
rect 12002 571 12068 572
rect 12002 560 12009 571
rect 11661 530 12009 560
rect 11661 519 11668 530
rect 11602 518 11668 519
rect 12002 519 12009 530
rect 12061 560 12068 571
rect 12402 571 12468 572
rect 12402 560 12409 571
rect 12061 530 12409 560
rect 12061 519 12068 530
rect 12002 518 12068 519
rect 12402 519 12409 530
rect 12461 560 12468 571
rect 12802 571 12868 572
rect 12802 560 12809 571
rect 12461 530 12809 560
rect 12461 519 12468 530
rect 12402 518 12468 519
rect 12802 519 12809 530
rect 12861 560 12868 571
rect 12900 571 12966 572
rect 12900 560 12907 571
rect 12861 530 12907 560
rect 12861 519 12868 530
rect 12802 518 12868 519
rect 12900 519 12907 530
rect 12959 519 12966 571
rect 12900 518 12966 519
rect 202 501 268 502
rect 202 490 209 501
rect 0 460 209 490
rect 202 449 209 460
rect 261 490 268 501
rect 602 501 668 502
rect 602 490 609 501
rect 261 460 609 490
rect 261 449 268 460
rect 202 448 268 449
rect 602 449 609 460
rect 661 490 668 501
rect 1002 501 1068 502
rect 1002 490 1009 501
rect 661 460 1009 490
rect 661 449 668 460
rect 602 448 668 449
rect 1002 449 1009 460
rect 1061 490 1068 501
rect 1402 501 1468 502
rect 1402 490 1409 501
rect 1061 460 1409 490
rect 1061 449 1068 460
rect 1002 448 1068 449
rect 1402 449 1409 460
rect 1461 490 1468 501
rect 1802 501 1868 502
rect 1802 490 1809 501
rect 1461 460 1809 490
rect 1461 449 1468 460
rect 1402 448 1468 449
rect 1802 449 1809 460
rect 1861 490 1868 501
rect 2202 501 2268 502
rect 2202 490 2209 501
rect 1861 460 2209 490
rect 1861 449 1868 460
rect 1802 448 1868 449
rect 2202 449 2209 460
rect 2261 490 2268 501
rect 2602 501 2668 502
rect 2602 490 2609 501
rect 2261 460 2609 490
rect 2261 449 2268 460
rect 2202 448 2268 449
rect 2602 449 2609 460
rect 2661 490 2668 501
rect 3002 501 3068 502
rect 3002 490 3009 501
rect 2661 460 3009 490
rect 2661 449 2668 460
rect 2602 448 2668 449
rect 3002 449 3009 460
rect 3061 490 3068 501
rect 3402 501 3468 502
rect 3402 490 3409 501
rect 3061 460 3409 490
rect 3061 449 3068 460
rect 3002 448 3068 449
rect 3402 449 3409 460
rect 3461 490 3468 501
rect 3802 501 3868 502
rect 3802 490 3809 501
rect 3461 460 3809 490
rect 3461 449 3468 460
rect 3402 448 3468 449
rect 3802 449 3809 460
rect 3861 490 3868 501
rect 4202 501 4268 502
rect 4202 490 4209 501
rect 3861 460 4209 490
rect 3861 449 3868 460
rect 3802 448 3868 449
rect 4202 449 4209 460
rect 4261 490 4268 501
rect 4602 501 4668 502
rect 4602 490 4609 501
rect 4261 460 4609 490
rect 4261 449 4268 460
rect 4202 448 4268 449
rect 4602 449 4609 460
rect 4661 490 4668 501
rect 5002 501 5068 502
rect 5002 490 5009 501
rect 4661 460 5009 490
rect 4661 449 4668 460
rect 4602 448 4668 449
rect 5002 449 5009 460
rect 5061 490 5068 501
rect 5402 501 5468 502
rect 5402 490 5409 501
rect 5061 460 5409 490
rect 5061 449 5068 460
rect 5002 448 5068 449
rect 5402 449 5409 460
rect 5461 490 5468 501
rect 5802 501 5868 502
rect 5802 490 5809 501
rect 5461 460 5809 490
rect 5461 449 5468 460
rect 5402 448 5468 449
rect 5802 449 5809 460
rect 5861 490 5868 501
rect 6202 501 6268 502
rect 6202 490 6209 501
rect 5861 460 6209 490
rect 5861 449 5868 460
rect 5802 448 5868 449
rect 6202 449 6209 460
rect 6261 490 6268 501
rect 6602 501 6668 502
rect 6602 490 6609 501
rect 6261 460 6609 490
rect 6261 449 6268 460
rect 6202 448 6268 449
rect 6602 449 6609 460
rect 6661 490 6668 501
rect 7002 501 7068 502
rect 7002 490 7009 501
rect 6661 460 7009 490
rect 6661 449 6668 460
rect 6602 448 6668 449
rect 7002 449 7009 460
rect 7061 490 7068 501
rect 7402 501 7468 502
rect 7402 490 7409 501
rect 7061 460 7409 490
rect 7061 449 7068 460
rect 7002 448 7068 449
rect 7402 449 7409 460
rect 7461 490 7468 501
rect 7802 501 7868 502
rect 7802 490 7809 501
rect 7461 460 7809 490
rect 7461 449 7468 460
rect 7402 448 7468 449
rect 7802 449 7809 460
rect 7861 490 7868 501
rect 8202 501 8268 502
rect 8202 490 8209 501
rect 7861 460 8209 490
rect 7861 449 7868 460
rect 7802 448 7868 449
rect 8202 449 8209 460
rect 8261 490 8268 501
rect 8602 501 8668 502
rect 8602 490 8609 501
rect 8261 460 8609 490
rect 8261 449 8268 460
rect 8202 448 8268 449
rect 8602 449 8609 460
rect 8661 490 8668 501
rect 9002 501 9068 502
rect 9002 490 9009 501
rect 8661 460 9009 490
rect 8661 449 8668 460
rect 8602 448 8668 449
rect 9002 449 9009 460
rect 9061 490 9068 501
rect 9402 501 9468 502
rect 9402 490 9409 501
rect 9061 460 9409 490
rect 9061 449 9068 460
rect 9002 448 9068 449
rect 9402 449 9409 460
rect 9461 490 9468 501
rect 9802 501 9868 502
rect 9802 490 9809 501
rect 9461 460 9809 490
rect 9461 449 9468 460
rect 9402 448 9468 449
rect 9802 449 9809 460
rect 9861 490 9868 501
rect 10202 501 10268 502
rect 10202 490 10209 501
rect 9861 460 10209 490
rect 9861 449 9868 460
rect 9802 448 9868 449
rect 10202 449 10209 460
rect 10261 490 10268 501
rect 10602 501 10668 502
rect 10602 490 10609 501
rect 10261 460 10609 490
rect 10261 449 10268 460
rect 10202 448 10268 449
rect 10602 449 10609 460
rect 10661 490 10668 501
rect 11002 501 11068 502
rect 11002 490 11009 501
rect 10661 460 11009 490
rect 10661 449 10668 460
rect 10602 448 10668 449
rect 11002 449 11009 460
rect 11061 490 11068 501
rect 11402 501 11468 502
rect 11402 490 11409 501
rect 11061 460 11409 490
rect 11061 449 11068 460
rect 11002 448 11068 449
rect 11402 449 11409 460
rect 11461 490 11468 501
rect 11802 501 11868 502
rect 11802 490 11809 501
rect 11461 460 11809 490
rect 11461 449 11468 460
rect 11402 448 11468 449
rect 11802 449 11809 460
rect 11861 490 11868 501
rect 12202 501 12268 502
rect 12202 490 12209 501
rect 11861 460 12209 490
rect 11861 449 11868 460
rect 11802 448 11868 449
rect 12202 449 12209 460
rect 12261 490 12268 501
rect 12602 501 12668 502
rect 12602 490 12609 501
rect 12261 460 12609 490
rect 12261 449 12268 460
rect 12202 448 12268 449
rect 12602 449 12609 460
rect 12661 490 12668 501
rect 13104 501 13170 502
rect 13104 490 13111 501
rect 12661 460 13111 490
rect 12661 449 12668 460
rect 12602 448 12668 449
rect 13104 449 13111 460
rect 13163 449 13170 501
rect 13104 448 13170 449
rect 2 431 68 432
rect 2 420 9 431
rect 0 390 9 420
rect 2 379 9 390
rect 61 420 68 431
rect 402 431 468 432
rect 402 420 409 431
rect 61 390 409 420
rect 61 379 68 390
rect 2 378 68 379
rect 402 379 409 390
rect 461 420 468 431
rect 802 431 868 432
rect 802 420 809 431
rect 461 390 809 420
rect 461 379 468 390
rect 402 378 468 379
rect 802 379 809 390
rect 861 420 868 431
rect 1202 431 1268 432
rect 1202 420 1209 431
rect 861 390 1209 420
rect 861 379 868 390
rect 802 378 868 379
rect 1202 379 1209 390
rect 1261 420 1268 431
rect 1602 431 1668 432
rect 1602 420 1609 431
rect 1261 390 1609 420
rect 1261 379 1268 390
rect 1202 378 1268 379
rect 1602 379 1609 390
rect 1661 420 1668 431
rect 2002 431 2068 432
rect 2002 420 2009 431
rect 1661 390 2009 420
rect 1661 379 1668 390
rect 1602 378 1668 379
rect 2002 379 2009 390
rect 2061 420 2068 431
rect 2402 431 2468 432
rect 2402 420 2409 431
rect 2061 390 2409 420
rect 2061 379 2068 390
rect 2002 378 2068 379
rect 2402 379 2409 390
rect 2461 420 2468 431
rect 2802 431 2868 432
rect 2802 420 2809 431
rect 2461 390 2809 420
rect 2461 379 2468 390
rect 2402 378 2468 379
rect 2802 379 2809 390
rect 2861 420 2868 431
rect 3202 431 3268 432
rect 3202 420 3209 431
rect 2861 390 3209 420
rect 2861 379 2868 390
rect 2802 378 2868 379
rect 3202 379 3209 390
rect 3261 420 3268 431
rect 3602 431 3668 432
rect 3602 420 3609 431
rect 3261 390 3609 420
rect 3261 379 3268 390
rect 3202 378 3268 379
rect 3602 379 3609 390
rect 3661 420 3668 431
rect 4002 431 4068 432
rect 4002 420 4009 431
rect 3661 390 4009 420
rect 3661 379 3668 390
rect 3602 378 3668 379
rect 4002 379 4009 390
rect 4061 420 4068 431
rect 4402 431 4468 432
rect 4402 420 4409 431
rect 4061 390 4409 420
rect 4061 379 4068 390
rect 4002 378 4068 379
rect 4402 379 4409 390
rect 4461 420 4468 431
rect 4802 431 4868 432
rect 4802 420 4809 431
rect 4461 390 4809 420
rect 4461 379 4468 390
rect 4402 378 4468 379
rect 4802 379 4809 390
rect 4861 420 4868 431
rect 5202 431 5268 432
rect 5202 420 5209 431
rect 4861 390 5209 420
rect 4861 379 4868 390
rect 4802 378 4868 379
rect 5202 379 5209 390
rect 5261 420 5268 431
rect 5602 431 5668 432
rect 5602 420 5609 431
rect 5261 390 5609 420
rect 5261 379 5268 390
rect 5202 378 5268 379
rect 5602 379 5609 390
rect 5661 420 5668 431
rect 6002 431 6068 432
rect 6002 420 6009 431
rect 5661 390 6009 420
rect 5661 379 5668 390
rect 5602 378 5668 379
rect 6002 379 6009 390
rect 6061 420 6068 431
rect 6402 431 6468 432
rect 6402 420 6409 431
rect 6061 390 6409 420
rect 6061 379 6068 390
rect 6002 378 6068 379
rect 6402 379 6409 390
rect 6461 420 6468 431
rect 6802 431 6868 432
rect 6802 420 6809 431
rect 6461 390 6809 420
rect 6461 379 6468 390
rect 6402 378 6468 379
rect 6802 379 6809 390
rect 6861 420 6868 431
rect 7202 431 7268 432
rect 7202 420 7209 431
rect 6861 390 7209 420
rect 6861 379 6868 390
rect 6802 378 6868 379
rect 7202 379 7209 390
rect 7261 420 7268 431
rect 7602 431 7668 432
rect 7602 420 7609 431
rect 7261 390 7609 420
rect 7261 379 7268 390
rect 7202 378 7268 379
rect 7602 379 7609 390
rect 7661 420 7668 431
rect 8002 431 8068 432
rect 8002 420 8009 431
rect 7661 390 8009 420
rect 7661 379 7668 390
rect 7602 378 7668 379
rect 8002 379 8009 390
rect 8061 420 8068 431
rect 8402 431 8468 432
rect 8402 420 8409 431
rect 8061 390 8409 420
rect 8061 379 8068 390
rect 8002 378 8068 379
rect 8402 379 8409 390
rect 8461 420 8468 431
rect 8802 431 8868 432
rect 8802 420 8809 431
rect 8461 390 8809 420
rect 8461 379 8468 390
rect 8402 378 8468 379
rect 8802 379 8809 390
rect 8861 420 8868 431
rect 9202 431 9268 432
rect 9202 420 9209 431
rect 8861 390 9209 420
rect 8861 379 8868 390
rect 8802 378 8868 379
rect 9202 379 9209 390
rect 9261 420 9268 431
rect 9602 431 9668 432
rect 9602 420 9609 431
rect 9261 390 9609 420
rect 9261 379 9268 390
rect 9202 378 9268 379
rect 9602 379 9609 390
rect 9661 420 9668 431
rect 10002 431 10068 432
rect 10002 420 10009 431
rect 9661 390 10009 420
rect 9661 379 9668 390
rect 9602 378 9668 379
rect 10002 379 10009 390
rect 10061 420 10068 431
rect 10402 431 10468 432
rect 10402 420 10409 431
rect 10061 390 10409 420
rect 10061 379 10068 390
rect 10002 378 10068 379
rect 10402 379 10409 390
rect 10461 420 10468 431
rect 10802 431 10868 432
rect 10802 420 10809 431
rect 10461 390 10809 420
rect 10461 379 10468 390
rect 10402 378 10468 379
rect 10802 379 10809 390
rect 10861 420 10868 431
rect 11202 431 11268 432
rect 11202 420 11209 431
rect 10861 390 11209 420
rect 10861 379 10868 390
rect 10802 378 10868 379
rect 11202 379 11209 390
rect 11261 420 11268 431
rect 11602 431 11668 432
rect 11602 420 11609 431
rect 11261 390 11609 420
rect 11261 379 11268 390
rect 11202 378 11268 379
rect 11602 379 11609 390
rect 11661 420 11668 431
rect 12002 431 12068 432
rect 12002 420 12009 431
rect 11661 390 12009 420
rect 11661 379 11668 390
rect 11602 378 11668 379
rect 12002 379 12009 390
rect 12061 420 12068 431
rect 12402 431 12468 432
rect 12402 420 12409 431
rect 12061 390 12409 420
rect 12061 379 12068 390
rect 12002 378 12068 379
rect 12402 379 12409 390
rect 12461 420 12468 431
rect 12802 431 12868 432
rect 12802 420 12809 431
rect 12461 390 12809 420
rect 12461 379 12468 390
rect 12402 378 12468 379
rect 12802 379 12809 390
rect 12861 420 12868 431
rect 12900 431 12966 432
rect 12900 420 12907 431
rect 12861 390 12907 420
rect 12861 379 12868 390
rect 12802 378 12868 379
rect 12900 379 12907 390
rect 12959 379 12966 431
rect 12900 378 12966 379
rect 202 361 268 362
rect 202 350 209 361
rect 0 320 209 350
rect 202 309 209 320
rect 261 350 268 361
rect 602 361 668 362
rect 602 350 609 361
rect 261 320 609 350
rect 261 309 268 320
rect 202 308 268 309
rect 602 309 609 320
rect 661 350 668 361
rect 1002 361 1068 362
rect 1002 350 1009 361
rect 661 320 1009 350
rect 661 309 668 320
rect 602 308 668 309
rect 1002 309 1009 320
rect 1061 350 1068 361
rect 1402 361 1468 362
rect 1402 350 1409 361
rect 1061 320 1409 350
rect 1061 309 1068 320
rect 1002 308 1068 309
rect 1402 309 1409 320
rect 1461 350 1468 361
rect 1802 361 1868 362
rect 1802 350 1809 361
rect 1461 320 1809 350
rect 1461 309 1468 320
rect 1402 308 1468 309
rect 1802 309 1809 320
rect 1861 350 1868 361
rect 2202 361 2268 362
rect 2202 350 2209 361
rect 1861 320 2209 350
rect 1861 309 1868 320
rect 1802 308 1868 309
rect 2202 309 2209 320
rect 2261 350 2268 361
rect 2602 361 2668 362
rect 2602 350 2609 361
rect 2261 320 2609 350
rect 2261 309 2268 320
rect 2202 308 2268 309
rect 2602 309 2609 320
rect 2661 350 2668 361
rect 3002 361 3068 362
rect 3002 350 3009 361
rect 2661 320 3009 350
rect 2661 309 2668 320
rect 2602 308 2668 309
rect 3002 309 3009 320
rect 3061 350 3068 361
rect 3402 361 3468 362
rect 3402 350 3409 361
rect 3061 320 3409 350
rect 3061 309 3068 320
rect 3002 308 3068 309
rect 3402 309 3409 320
rect 3461 350 3468 361
rect 3802 361 3868 362
rect 3802 350 3809 361
rect 3461 320 3809 350
rect 3461 309 3468 320
rect 3402 308 3468 309
rect 3802 309 3809 320
rect 3861 350 3868 361
rect 4202 361 4268 362
rect 4202 350 4209 361
rect 3861 320 4209 350
rect 3861 309 3868 320
rect 3802 308 3868 309
rect 4202 309 4209 320
rect 4261 350 4268 361
rect 4602 361 4668 362
rect 4602 350 4609 361
rect 4261 320 4609 350
rect 4261 309 4268 320
rect 4202 308 4268 309
rect 4602 309 4609 320
rect 4661 350 4668 361
rect 5002 361 5068 362
rect 5002 350 5009 361
rect 4661 320 5009 350
rect 4661 309 4668 320
rect 4602 308 4668 309
rect 5002 309 5009 320
rect 5061 350 5068 361
rect 5402 361 5468 362
rect 5402 350 5409 361
rect 5061 320 5409 350
rect 5061 309 5068 320
rect 5002 308 5068 309
rect 5402 309 5409 320
rect 5461 350 5468 361
rect 5802 361 5868 362
rect 5802 350 5809 361
rect 5461 320 5809 350
rect 5461 309 5468 320
rect 5402 308 5468 309
rect 5802 309 5809 320
rect 5861 350 5868 361
rect 6202 361 6268 362
rect 6202 350 6209 361
rect 5861 320 6209 350
rect 5861 309 5868 320
rect 5802 308 5868 309
rect 6202 309 6209 320
rect 6261 350 6268 361
rect 6602 361 6668 362
rect 6602 350 6609 361
rect 6261 320 6609 350
rect 6261 309 6268 320
rect 6202 308 6268 309
rect 6602 309 6609 320
rect 6661 350 6668 361
rect 7002 361 7068 362
rect 7002 350 7009 361
rect 6661 320 7009 350
rect 6661 309 6668 320
rect 6602 308 6668 309
rect 7002 309 7009 320
rect 7061 350 7068 361
rect 7402 361 7468 362
rect 7402 350 7409 361
rect 7061 320 7409 350
rect 7061 309 7068 320
rect 7002 308 7068 309
rect 7402 309 7409 320
rect 7461 350 7468 361
rect 7802 361 7868 362
rect 7802 350 7809 361
rect 7461 320 7809 350
rect 7461 309 7468 320
rect 7402 308 7468 309
rect 7802 309 7809 320
rect 7861 350 7868 361
rect 8202 361 8268 362
rect 8202 350 8209 361
rect 7861 320 8209 350
rect 7861 309 7868 320
rect 7802 308 7868 309
rect 8202 309 8209 320
rect 8261 350 8268 361
rect 8602 361 8668 362
rect 8602 350 8609 361
rect 8261 320 8609 350
rect 8261 309 8268 320
rect 8202 308 8268 309
rect 8602 309 8609 320
rect 8661 350 8668 361
rect 9002 361 9068 362
rect 9002 350 9009 361
rect 8661 320 9009 350
rect 8661 309 8668 320
rect 8602 308 8668 309
rect 9002 309 9009 320
rect 9061 350 9068 361
rect 9402 361 9468 362
rect 9402 350 9409 361
rect 9061 320 9409 350
rect 9061 309 9068 320
rect 9002 308 9068 309
rect 9402 309 9409 320
rect 9461 350 9468 361
rect 9802 361 9868 362
rect 9802 350 9809 361
rect 9461 320 9809 350
rect 9461 309 9468 320
rect 9402 308 9468 309
rect 9802 309 9809 320
rect 9861 350 9868 361
rect 10202 361 10268 362
rect 10202 350 10209 361
rect 9861 320 10209 350
rect 9861 309 9868 320
rect 9802 308 9868 309
rect 10202 309 10209 320
rect 10261 350 10268 361
rect 10602 361 10668 362
rect 10602 350 10609 361
rect 10261 320 10609 350
rect 10261 309 10268 320
rect 10202 308 10268 309
rect 10602 309 10609 320
rect 10661 350 10668 361
rect 11002 361 11068 362
rect 11002 350 11009 361
rect 10661 320 11009 350
rect 10661 309 10668 320
rect 10602 308 10668 309
rect 11002 309 11009 320
rect 11061 350 11068 361
rect 11402 361 11468 362
rect 11402 350 11409 361
rect 11061 320 11409 350
rect 11061 309 11068 320
rect 11002 308 11068 309
rect 11402 309 11409 320
rect 11461 350 11468 361
rect 11802 361 11868 362
rect 11802 350 11809 361
rect 11461 320 11809 350
rect 11461 309 11468 320
rect 11402 308 11468 309
rect 11802 309 11809 320
rect 11861 350 11868 361
rect 12202 361 12268 362
rect 12202 350 12209 361
rect 11861 320 12209 350
rect 11861 309 11868 320
rect 11802 308 11868 309
rect 12202 309 12209 320
rect 12261 350 12268 361
rect 12602 361 12668 362
rect 12602 350 12609 361
rect 12261 320 12609 350
rect 12261 309 12268 320
rect 12202 308 12268 309
rect 12602 309 12609 320
rect 12661 350 12668 361
rect 13104 361 13170 362
rect 13104 350 13111 361
rect 12661 320 13111 350
rect 12661 309 12668 320
rect 12602 308 12668 309
rect 13104 309 13111 320
rect 13163 309 13170 361
rect 13104 308 13170 309
rect 2 291 68 292
rect 2 280 9 291
rect 0 250 9 280
rect 2 239 9 250
rect 61 280 68 291
rect 402 291 468 292
rect 402 280 409 291
rect 61 250 409 280
rect 61 239 68 250
rect 2 238 68 239
rect 402 239 409 250
rect 461 280 468 291
rect 802 291 868 292
rect 802 280 809 291
rect 461 250 809 280
rect 461 239 468 250
rect 402 238 468 239
rect 802 239 809 250
rect 861 280 868 291
rect 1202 291 1268 292
rect 1202 280 1209 291
rect 861 250 1209 280
rect 861 239 868 250
rect 802 238 868 239
rect 1202 239 1209 250
rect 1261 280 1268 291
rect 1602 291 1668 292
rect 1602 280 1609 291
rect 1261 250 1609 280
rect 1261 239 1268 250
rect 1202 238 1268 239
rect 1602 239 1609 250
rect 1661 280 1668 291
rect 2002 291 2068 292
rect 2002 280 2009 291
rect 1661 250 2009 280
rect 1661 239 1668 250
rect 1602 238 1668 239
rect 2002 239 2009 250
rect 2061 280 2068 291
rect 2402 291 2468 292
rect 2402 280 2409 291
rect 2061 250 2409 280
rect 2061 239 2068 250
rect 2002 238 2068 239
rect 2402 239 2409 250
rect 2461 280 2468 291
rect 2802 291 2868 292
rect 2802 280 2809 291
rect 2461 250 2809 280
rect 2461 239 2468 250
rect 2402 238 2468 239
rect 2802 239 2809 250
rect 2861 280 2868 291
rect 3202 291 3268 292
rect 3202 280 3209 291
rect 2861 250 3209 280
rect 2861 239 2868 250
rect 2802 238 2868 239
rect 3202 239 3209 250
rect 3261 280 3268 291
rect 3602 291 3668 292
rect 3602 280 3609 291
rect 3261 250 3609 280
rect 3261 239 3268 250
rect 3202 238 3268 239
rect 3602 239 3609 250
rect 3661 280 3668 291
rect 4002 291 4068 292
rect 4002 280 4009 291
rect 3661 250 4009 280
rect 3661 239 3668 250
rect 3602 238 3668 239
rect 4002 239 4009 250
rect 4061 280 4068 291
rect 4402 291 4468 292
rect 4402 280 4409 291
rect 4061 250 4409 280
rect 4061 239 4068 250
rect 4002 238 4068 239
rect 4402 239 4409 250
rect 4461 280 4468 291
rect 4802 291 4868 292
rect 4802 280 4809 291
rect 4461 250 4809 280
rect 4461 239 4468 250
rect 4402 238 4468 239
rect 4802 239 4809 250
rect 4861 280 4868 291
rect 5202 291 5268 292
rect 5202 280 5209 291
rect 4861 250 5209 280
rect 4861 239 4868 250
rect 4802 238 4868 239
rect 5202 239 5209 250
rect 5261 280 5268 291
rect 5602 291 5668 292
rect 5602 280 5609 291
rect 5261 250 5609 280
rect 5261 239 5268 250
rect 5202 238 5268 239
rect 5602 239 5609 250
rect 5661 280 5668 291
rect 6002 291 6068 292
rect 6002 280 6009 291
rect 5661 250 6009 280
rect 5661 239 5668 250
rect 5602 238 5668 239
rect 6002 239 6009 250
rect 6061 280 6068 291
rect 6402 291 6468 292
rect 6402 280 6409 291
rect 6061 250 6409 280
rect 6061 239 6068 250
rect 6002 238 6068 239
rect 6402 239 6409 250
rect 6461 280 6468 291
rect 6802 291 6868 292
rect 6802 280 6809 291
rect 6461 250 6809 280
rect 6461 239 6468 250
rect 6402 238 6468 239
rect 6802 239 6809 250
rect 6861 280 6868 291
rect 7202 291 7268 292
rect 7202 280 7209 291
rect 6861 250 7209 280
rect 6861 239 6868 250
rect 6802 238 6868 239
rect 7202 239 7209 250
rect 7261 280 7268 291
rect 7602 291 7668 292
rect 7602 280 7609 291
rect 7261 250 7609 280
rect 7261 239 7268 250
rect 7202 238 7268 239
rect 7602 239 7609 250
rect 7661 280 7668 291
rect 8002 291 8068 292
rect 8002 280 8009 291
rect 7661 250 8009 280
rect 7661 239 7668 250
rect 7602 238 7668 239
rect 8002 239 8009 250
rect 8061 280 8068 291
rect 8402 291 8468 292
rect 8402 280 8409 291
rect 8061 250 8409 280
rect 8061 239 8068 250
rect 8002 238 8068 239
rect 8402 239 8409 250
rect 8461 280 8468 291
rect 8802 291 8868 292
rect 8802 280 8809 291
rect 8461 250 8809 280
rect 8461 239 8468 250
rect 8402 238 8468 239
rect 8802 239 8809 250
rect 8861 280 8868 291
rect 9202 291 9268 292
rect 9202 280 9209 291
rect 8861 250 9209 280
rect 8861 239 8868 250
rect 8802 238 8868 239
rect 9202 239 9209 250
rect 9261 280 9268 291
rect 9602 291 9668 292
rect 9602 280 9609 291
rect 9261 250 9609 280
rect 9261 239 9268 250
rect 9202 238 9268 239
rect 9602 239 9609 250
rect 9661 280 9668 291
rect 10002 291 10068 292
rect 10002 280 10009 291
rect 9661 250 10009 280
rect 9661 239 9668 250
rect 9602 238 9668 239
rect 10002 239 10009 250
rect 10061 280 10068 291
rect 10402 291 10468 292
rect 10402 280 10409 291
rect 10061 250 10409 280
rect 10061 239 10068 250
rect 10002 238 10068 239
rect 10402 239 10409 250
rect 10461 280 10468 291
rect 10802 291 10868 292
rect 10802 280 10809 291
rect 10461 250 10809 280
rect 10461 239 10468 250
rect 10402 238 10468 239
rect 10802 239 10809 250
rect 10861 280 10868 291
rect 11202 291 11268 292
rect 11202 280 11209 291
rect 10861 250 11209 280
rect 10861 239 10868 250
rect 10802 238 10868 239
rect 11202 239 11209 250
rect 11261 280 11268 291
rect 11602 291 11668 292
rect 11602 280 11609 291
rect 11261 250 11609 280
rect 11261 239 11268 250
rect 11202 238 11268 239
rect 11602 239 11609 250
rect 11661 280 11668 291
rect 12002 291 12068 292
rect 12002 280 12009 291
rect 11661 250 12009 280
rect 11661 239 11668 250
rect 11602 238 11668 239
rect 12002 239 12009 250
rect 12061 280 12068 291
rect 12402 291 12468 292
rect 12402 280 12409 291
rect 12061 250 12409 280
rect 12061 239 12068 250
rect 12002 238 12068 239
rect 12402 239 12409 250
rect 12461 280 12468 291
rect 12802 291 12868 292
rect 12802 280 12809 291
rect 12461 250 12809 280
rect 12461 239 12468 250
rect 12402 238 12468 239
rect 12802 239 12809 250
rect 12861 280 12868 291
rect 12900 291 12966 292
rect 12900 280 12907 291
rect 12861 250 12907 280
rect 12861 239 12868 250
rect 12802 238 12868 239
rect 12900 239 12907 250
rect 12959 239 12966 291
rect 12900 238 12966 239
rect 202 221 268 222
rect 202 210 209 221
rect 0 180 209 210
rect 202 169 209 180
rect 261 210 268 221
rect 602 221 668 222
rect 602 210 609 221
rect 261 180 609 210
rect 261 169 268 180
rect 202 168 268 169
rect 602 169 609 180
rect 661 210 668 221
rect 1002 221 1068 222
rect 1002 210 1009 221
rect 661 180 1009 210
rect 661 169 668 180
rect 602 168 668 169
rect 1002 169 1009 180
rect 1061 210 1068 221
rect 1402 221 1468 222
rect 1402 210 1409 221
rect 1061 180 1409 210
rect 1061 169 1068 180
rect 1002 168 1068 169
rect 1402 169 1409 180
rect 1461 210 1468 221
rect 1802 221 1868 222
rect 1802 210 1809 221
rect 1461 180 1809 210
rect 1461 169 1468 180
rect 1402 168 1468 169
rect 1802 169 1809 180
rect 1861 210 1868 221
rect 2202 221 2268 222
rect 2202 210 2209 221
rect 1861 180 2209 210
rect 1861 169 1868 180
rect 1802 168 1868 169
rect 2202 169 2209 180
rect 2261 210 2268 221
rect 2602 221 2668 222
rect 2602 210 2609 221
rect 2261 180 2609 210
rect 2261 169 2268 180
rect 2202 168 2268 169
rect 2602 169 2609 180
rect 2661 210 2668 221
rect 3002 221 3068 222
rect 3002 210 3009 221
rect 2661 180 3009 210
rect 2661 169 2668 180
rect 2602 168 2668 169
rect 3002 169 3009 180
rect 3061 210 3068 221
rect 3402 221 3468 222
rect 3402 210 3409 221
rect 3061 180 3409 210
rect 3061 169 3068 180
rect 3002 168 3068 169
rect 3402 169 3409 180
rect 3461 210 3468 221
rect 3802 221 3868 222
rect 3802 210 3809 221
rect 3461 180 3809 210
rect 3461 169 3468 180
rect 3402 168 3468 169
rect 3802 169 3809 180
rect 3861 210 3868 221
rect 4202 221 4268 222
rect 4202 210 4209 221
rect 3861 180 4209 210
rect 3861 169 3868 180
rect 3802 168 3868 169
rect 4202 169 4209 180
rect 4261 210 4268 221
rect 4602 221 4668 222
rect 4602 210 4609 221
rect 4261 180 4609 210
rect 4261 169 4268 180
rect 4202 168 4268 169
rect 4602 169 4609 180
rect 4661 210 4668 221
rect 5002 221 5068 222
rect 5002 210 5009 221
rect 4661 180 5009 210
rect 4661 169 4668 180
rect 4602 168 4668 169
rect 5002 169 5009 180
rect 5061 210 5068 221
rect 5402 221 5468 222
rect 5402 210 5409 221
rect 5061 180 5409 210
rect 5061 169 5068 180
rect 5002 168 5068 169
rect 5402 169 5409 180
rect 5461 210 5468 221
rect 5802 221 5868 222
rect 5802 210 5809 221
rect 5461 180 5809 210
rect 5461 169 5468 180
rect 5402 168 5468 169
rect 5802 169 5809 180
rect 5861 210 5868 221
rect 6202 221 6268 222
rect 6202 210 6209 221
rect 5861 180 6209 210
rect 5861 169 5868 180
rect 5802 168 5868 169
rect 6202 169 6209 180
rect 6261 210 6268 221
rect 6602 221 6668 222
rect 6602 210 6609 221
rect 6261 180 6609 210
rect 6261 169 6268 180
rect 6202 168 6268 169
rect 6602 169 6609 180
rect 6661 210 6668 221
rect 7002 221 7068 222
rect 7002 210 7009 221
rect 6661 180 7009 210
rect 6661 169 6668 180
rect 6602 168 6668 169
rect 7002 169 7009 180
rect 7061 210 7068 221
rect 7402 221 7468 222
rect 7402 210 7409 221
rect 7061 180 7409 210
rect 7061 169 7068 180
rect 7002 168 7068 169
rect 7402 169 7409 180
rect 7461 210 7468 221
rect 7802 221 7868 222
rect 7802 210 7809 221
rect 7461 180 7809 210
rect 7461 169 7468 180
rect 7402 168 7468 169
rect 7802 169 7809 180
rect 7861 210 7868 221
rect 8202 221 8268 222
rect 8202 210 8209 221
rect 7861 180 8209 210
rect 7861 169 7868 180
rect 7802 168 7868 169
rect 8202 169 8209 180
rect 8261 210 8268 221
rect 8602 221 8668 222
rect 8602 210 8609 221
rect 8261 180 8609 210
rect 8261 169 8268 180
rect 8202 168 8268 169
rect 8602 169 8609 180
rect 8661 210 8668 221
rect 9002 221 9068 222
rect 9002 210 9009 221
rect 8661 180 9009 210
rect 8661 169 8668 180
rect 8602 168 8668 169
rect 9002 169 9009 180
rect 9061 210 9068 221
rect 9402 221 9468 222
rect 9402 210 9409 221
rect 9061 180 9409 210
rect 9061 169 9068 180
rect 9002 168 9068 169
rect 9402 169 9409 180
rect 9461 210 9468 221
rect 9802 221 9868 222
rect 9802 210 9809 221
rect 9461 180 9809 210
rect 9461 169 9468 180
rect 9402 168 9468 169
rect 9802 169 9809 180
rect 9861 210 9868 221
rect 10202 221 10268 222
rect 10202 210 10209 221
rect 9861 180 10209 210
rect 9861 169 9868 180
rect 9802 168 9868 169
rect 10202 169 10209 180
rect 10261 210 10268 221
rect 10602 221 10668 222
rect 10602 210 10609 221
rect 10261 180 10609 210
rect 10261 169 10268 180
rect 10202 168 10268 169
rect 10602 169 10609 180
rect 10661 210 10668 221
rect 11002 221 11068 222
rect 11002 210 11009 221
rect 10661 180 11009 210
rect 10661 169 10668 180
rect 10602 168 10668 169
rect 11002 169 11009 180
rect 11061 210 11068 221
rect 11402 221 11468 222
rect 11402 210 11409 221
rect 11061 180 11409 210
rect 11061 169 11068 180
rect 11002 168 11068 169
rect 11402 169 11409 180
rect 11461 210 11468 221
rect 11802 221 11868 222
rect 11802 210 11809 221
rect 11461 180 11809 210
rect 11461 169 11468 180
rect 11402 168 11468 169
rect 11802 169 11809 180
rect 11861 210 11868 221
rect 12202 221 12268 222
rect 12202 210 12209 221
rect 11861 180 12209 210
rect 11861 169 11868 180
rect 11802 168 11868 169
rect 12202 169 12209 180
rect 12261 210 12268 221
rect 12602 221 12668 222
rect 12602 210 12609 221
rect 12261 180 12609 210
rect 12261 169 12268 180
rect 12202 168 12268 169
rect 12602 169 12609 180
rect 12661 210 12668 221
rect 13104 221 13170 222
rect 13104 210 13111 221
rect 12661 180 13111 210
rect 12661 169 12668 180
rect 12602 168 12668 169
rect 13104 169 13111 180
rect 13163 169 13170 221
rect 13104 168 13170 169
rect 2 151 68 152
rect 2 140 9 151
rect 0 110 9 140
rect 2 99 9 110
rect 61 140 68 151
rect 402 151 468 152
rect 402 140 409 151
rect 61 110 409 140
rect 61 99 68 110
rect 2 98 68 99
rect 402 99 409 110
rect 461 140 468 151
rect 802 151 868 152
rect 802 140 809 151
rect 461 110 809 140
rect 461 99 468 110
rect 402 98 468 99
rect 802 99 809 110
rect 861 140 868 151
rect 1202 151 1268 152
rect 1202 140 1209 151
rect 861 110 1209 140
rect 861 99 868 110
rect 802 98 868 99
rect 1202 99 1209 110
rect 1261 140 1268 151
rect 1602 151 1668 152
rect 1602 140 1609 151
rect 1261 110 1609 140
rect 1261 99 1268 110
rect 1202 98 1268 99
rect 1602 99 1609 110
rect 1661 140 1668 151
rect 2002 151 2068 152
rect 2002 140 2009 151
rect 1661 110 2009 140
rect 1661 99 1668 110
rect 1602 98 1668 99
rect 2002 99 2009 110
rect 2061 140 2068 151
rect 2402 151 2468 152
rect 2402 140 2409 151
rect 2061 110 2409 140
rect 2061 99 2068 110
rect 2002 98 2068 99
rect 2402 99 2409 110
rect 2461 140 2468 151
rect 2802 151 2868 152
rect 2802 140 2809 151
rect 2461 110 2809 140
rect 2461 99 2468 110
rect 2402 98 2468 99
rect 2802 99 2809 110
rect 2861 140 2868 151
rect 3202 151 3268 152
rect 3202 140 3209 151
rect 2861 110 3209 140
rect 2861 99 2868 110
rect 2802 98 2868 99
rect 3202 99 3209 110
rect 3261 140 3268 151
rect 3602 151 3668 152
rect 3602 140 3609 151
rect 3261 110 3609 140
rect 3261 99 3268 110
rect 3202 98 3268 99
rect 3602 99 3609 110
rect 3661 140 3668 151
rect 4002 151 4068 152
rect 4002 140 4009 151
rect 3661 110 4009 140
rect 3661 99 3668 110
rect 3602 98 3668 99
rect 4002 99 4009 110
rect 4061 140 4068 151
rect 4402 151 4468 152
rect 4402 140 4409 151
rect 4061 110 4409 140
rect 4061 99 4068 110
rect 4002 98 4068 99
rect 4402 99 4409 110
rect 4461 140 4468 151
rect 4802 151 4868 152
rect 4802 140 4809 151
rect 4461 110 4809 140
rect 4461 99 4468 110
rect 4402 98 4468 99
rect 4802 99 4809 110
rect 4861 140 4868 151
rect 5202 151 5268 152
rect 5202 140 5209 151
rect 4861 110 5209 140
rect 4861 99 4868 110
rect 4802 98 4868 99
rect 5202 99 5209 110
rect 5261 140 5268 151
rect 5602 151 5668 152
rect 5602 140 5609 151
rect 5261 110 5609 140
rect 5261 99 5268 110
rect 5202 98 5268 99
rect 5602 99 5609 110
rect 5661 140 5668 151
rect 6002 151 6068 152
rect 6002 140 6009 151
rect 5661 110 6009 140
rect 5661 99 5668 110
rect 5602 98 5668 99
rect 6002 99 6009 110
rect 6061 140 6068 151
rect 6402 151 6468 152
rect 6402 140 6409 151
rect 6061 110 6409 140
rect 6061 99 6068 110
rect 6002 98 6068 99
rect 6402 99 6409 110
rect 6461 140 6468 151
rect 6802 151 6868 152
rect 6802 140 6809 151
rect 6461 110 6809 140
rect 6461 99 6468 110
rect 6402 98 6468 99
rect 6802 99 6809 110
rect 6861 140 6868 151
rect 7202 151 7268 152
rect 7202 140 7209 151
rect 6861 110 7209 140
rect 6861 99 6868 110
rect 6802 98 6868 99
rect 7202 99 7209 110
rect 7261 140 7268 151
rect 7602 151 7668 152
rect 7602 140 7609 151
rect 7261 110 7609 140
rect 7261 99 7268 110
rect 7202 98 7268 99
rect 7602 99 7609 110
rect 7661 140 7668 151
rect 8002 151 8068 152
rect 8002 140 8009 151
rect 7661 110 8009 140
rect 7661 99 7668 110
rect 7602 98 7668 99
rect 8002 99 8009 110
rect 8061 140 8068 151
rect 8402 151 8468 152
rect 8402 140 8409 151
rect 8061 110 8409 140
rect 8061 99 8068 110
rect 8002 98 8068 99
rect 8402 99 8409 110
rect 8461 140 8468 151
rect 8802 151 8868 152
rect 8802 140 8809 151
rect 8461 110 8809 140
rect 8461 99 8468 110
rect 8402 98 8468 99
rect 8802 99 8809 110
rect 8861 140 8868 151
rect 9202 151 9268 152
rect 9202 140 9209 151
rect 8861 110 9209 140
rect 8861 99 8868 110
rect 8802 98 8868 99
rect 9202 99 9209 110
rect 9261 140 9268 151
rect 9602 151 9668 152
rect 9602 140 9609 151
rect 9261 110 9609 140
rect 9261 99 9268 110
rect 9202 98 9268 99
rect 9602 99 9609 110
rect 9661 140 9668 151
rect 10002 151 10068 152
rect 10002 140 10009 151
rect 9661 110 10009 140
rect 9661 99 9668 110
rect 9602 98 9668 99
rect 10002 99 10009 110
rect 10061 140 10068 151
rect 10402 151 10468 152
rect 10402 140 10409 151
rect 10061 110 10409 140
rect 10061 99 10068 110
rect 10002 98 10068 99
rect 10402 99 10409 110
rect 10461 140 10468 151
rect 10802 151 10868 152
rect 10802 140 10809 151
rect 10461 110 10809 140
rect 10461 99 10468 110
rect 10402 98 10468 99
rect 10802 99 10809 110
rect 10861 140 10868 151
rect 11202 151 11268 152
rect 11202 140 11209 151
rect 10861 110 11209 140
rect 10861 99 10868 110
rect 10802 98 10868 99
rect 11202 99 11209 110
rect 11261 140 11268 151
rect 11602 151 11668 152
rect 11602 140 11609 151
rect 11261 110 11609 140
rect 11261 99 11268 110
rect 11202 98 11268 99
rect 11602 99 11609 110
rect 11661 140 11668 151
rect 12002 151 12068 152
rect 12002 140 12009 151
rect 11661 110 12009 140
rect 11661 99 11668 110
rect 11602 98 11668 99
rect 12002 99 12009 110
rect 12061 140 12068 151
rect 12402 151 12468 152
rect 12402 140 12409 151
rect 12061 110 12409 140
rect 12061 99 12068 110
rect 12002 98 12068 99
rect 12402 99 12409 110
rect 12461 140 12468 151
rect 12802 151 12868 152
rect 12802 140 12809 151
rect 12461 110 12809 140
rect 12461 99 12468 110
rect 12402 98 12468 99
rect 12802 99 12809 110
rect 12861 140 12868 151
rect 12900 151 12966 152
rect 12900 140 12907 151
rect 12861 110 12907 140
rect 12861 99 12868 110
rect 12802 98 12868 99
rect 12900 99 12907 110
rect 12959 99 12966 151
rect 12900 98 12966 99
rect 196 81 274 82
rect -4 65 74 66
rect -4 9 7 65
rect 63 9 74 65
rect 196 25 207 81
rect 263 25 274 81
rect 596 81 674 82
rect 196 24 274 25
rect 396 65 474 66
rect -4 8 74 9
rect -93 -15 -37 0
rect -93 -67 -91 -15
rect -39 -67 -37 -15
rect -93 -79 -37 -67
rect -93 -110 -91 -79
rect -138 -131 -91 -110
rect -39 -110 -37 -79
rect 7 -16 63 8
rect 7 -74 9 -72
rect 61 -74 63 -72
rect 7 -81 63 -74
rect 107 -15 163 0
rect 107 -67 109 -15
rect 161 -67 163 -15
rect 107 -79 163 -67
rect 107 -110 109 -79
rect -39 -131 109 -110
rect 161 -110 163 -79
rect 207 -16 263 24
rect 396 9 407 65
rect 463 9 474 65
rect 596 25 607 81
rect 663 25 674 81
rect 996 81 1074 82
rect 596 24 674 25
rect 796 65 874 66
rect 396 8 474 9
rect 207 -74 209 -72
rect 261 -74 263 -72
rect 207 -81 263 -74
rect 307 -15 363 0
rect 307 -67 309 -15
rect 361 -67 363 -15
rect 307 -79 363 -67
rect 307 -110 309 -79
rect 161 -131 309 -110
rect 361 -110 363 -79
rect 407 -16 463 8
rect 407 -74 409 -72
rect 461 -74 463 -72
rect 407 -81 463 -74
rect 507 -15 563 0
rect 507 -67 509 -15
rect 561 -67 563 -15
rect 507 -79 563 -67
rect 507 -110 509 -79
rect 361 -131 509 -110
rect 561 -110 563 -79
rect 607 -16 663 24
rect 796 9 807 65
rect 863 9 874 65
rect 996 25 1007 81
rect 1063 25 1074 81
rect 1396 81 1474 82
rect 996 24 1074 25
rect 1196 65 1274 66
rect 796 8 874 9
rect 607 -74 609 -72
rect 661 -74 663 -72
rect 607 -81 663 -74
rect 707 -15 763 0
rect 707 -67 709 -15
rect 761 -67 763 -15
rect 707 -79 763 -67
rect 707 -110 709 -79
rect 561 -131 709 -110
rect 761 -110 763 -79
rect 807 -16 863 8
rect 807 -74 809 -72
rect 861 -74 863 -72
rect 807 -81 863 -74
rect 907 -15 963 0
rect 907 -67 909 -15
rect 961 -67 963 -15
rect 907 -79 963 -67
rect 907 -110 909 -79
rect 761 -131 909 -110
rect 961 -110 963 -79
rect 1007 -16 1063 24
rect 1196 9 1207 65
rect 1263 9 1274 65
rect 1396 25 1407 81
rect 1463 25 1474 81
rect 1796 81 1874 82
rect 1396 24 1474 25
rect 1596 65 1674 66
rect 1196 8 1274 9
rect 1007 -74 1009 -72
rect 1061 -74 1063 -72
rect 1007 -81 1063 -74
rect 1107 -15 1163 0
rect 1107 -67 1109 -15
rect 1161 -67 1163 -15
rect 1107 -79 1163 -67
rect 1107 -110 1109 -79
rect 961 -131 1109 -110
rect 1161 -110 1163 -79
rect 1207 -16 1263 8
rect 1207 -74 1209 -72
rect 1261 -74 1263 -72
rect 1207 -81 1263 -74
rect 1307 -15 1363 0
rect 1307 -67 1309 -15
rect 1361 -67 1363 -15
rect 1307 -79 1363 -67
rect 1307 -110 1309 -79
rect 1161 -131 1309 -110
rect 1361 -110 1363 -79
rect 1407 -16 1463 24
rect 1596 9 1607 65
rect 1663 9 1674 65
rect 1796 25 1807 81
rect 1863 25 1874 81
rect 2196 81 2274 82
rect 1796 24 1874 25
rect 1996 65 2074 66
rect 1596 8 1674 9
rect 1407 -74 1409 -72
rect 1461 -74 1463 -72
rect 1407 -81 1463 -74
rect 1507 -15 1563 0
rect 1507 -67 1509 -15
rect 1561 -67 1563 -15
rect 1507 -79 1563 -67
rect 1507 -110 1509 -79
rect 1361 -131 1509 -110
rect 1561 -110 1563 -79
rect 1607 -16 1663 8
rect 1607 -74 1609 -72
rect 1661 -74 1663 -72
rect 1607 -81 1663 -74
rect 1707 -15 1763 0
rect 1707 -67 1709 -15
rect 1761 -67 1763 -15
rect 1707 -79 1763 -67
rect 1707 -110 1709 -79
rect 1561 -131 1709 -110
rect 1761 -110 1763 -79
rect 1807 -16 1863 24
rect 1996 9 2007 65
rect 2063 9 2074 65
rect 2196 25 2207 81
rect 2263 25 2274 81
rect 2596 81 2674 82
rect 2196 24 2274 25
rect 2396 65 2474 66
rect 1996 8 2074 9
rect 1807 -74 1809 -72
rect 1861 -74 1863 -72
rect 1807 -81 1863 -74
rect 1907 -15 1963 0
rect 1907 -67 1909 -15
rect 1961 -67 1963 -15
rect 1907 -79 1963 -67
rect 1907 -110 1909 -79
rect 1761 -131 1909 -110
rect 1961 -110 1963 -79
rect 2007 -16 2063 8
rect 2007 -74 2009 -72
rect 2061 -74 2063 -72
rect 2007 -81 2063 -74
rect 2107 -15 2163 0
rect 2107 -67 2109 -15
rect 2161 -67 2163 -15
rect 2107 -79 2163 -67
rect 2107 -110 2109 -79
rect 1961 -131 2109 -110
rect 2161 -110 2163 -79
rect 2207 -16 2263 24
rect 2396 9 2407 65
rect 2463 9 2474 65
rect 2596 25 2607 81
rect 2663 25 2674 81
rect 2996 81 3074 82
rect 2596 24 2674 25
rect 2796 65 2874 66
rect 2396 8 2474 9
rect 2207 -74 2209 -72
rect 2261 -74 2263 -72
rect 2207 -81 2263 -74
rect 2307 -15 2363 0
rect 2307 -67 2309 -15
rect 2361 -67 2363 -15
rect 2307 -79 2363 -67
rect 2307 -110 2309 -79
rect 2161 -131 2309 -110
rect 2361 -110 2363 -79
rect 2407 -16 2463 8
rect 2407 -74 2409 -72
rect 2461 -74 2463 -72
rect 2407 -81 2463 -74
rect 2507 -15 2563 0
rect 2507 -67 2509 -15
rect 2561 -67 2563 -15
rect 2507 -79 2563 -67
rect 2507 -110 2509 -79
rect 2361 -131 2509 -110
rect 2561 -110 2563 -79
rect 2607 -16 2663 24
rect 2796 9 2807 65
rect 2863 9 2874 65
rect 2996 25 3007 81
rect 3063 25 3074 81
rect 3396 81 3474 82
rect 2996 24 3074 25
rect 3196 65 3274 66
rect 2796 8 2874 9
rect 2607 -74 2609 -72
rect 2661 -74 2663 -72
rect 2607 -81 2663 -74
rect 2707 -15 2763 0
rect 2707 -67 2709 -15
rect 2761 -67 2763 -15
rect 2707 -79 2763 -67
rect 2707 -110 2709 -79
rect 2561 -131 2709 -110
rect 2761 -110 2763 -79
rect 2807 -16 2863 8
rect 2807 -74 2809 -72
rect 2861 -74 2863 -72
rect 2807 -81 2863 -74
rect 2907 -15 2963 0
rect 2907 -67 2909 -15
rect 2961 -67 2963 -15
rect 2907 -79 2963 -67
rect 2907 -110 2909 -79
rect 2761 -131 2909 -110
rect 2961 -110 2963 -79
rect 3007 -16 3063 24
rect 3196 9 3207 65
rect 3263 9 3274 65
rect 3396 25 3407 81
rect 3463 25 3474 81
rect 3796 81 3874 82
rect 3396 24 3474 25
rect 3596 65 3674 66
rect 3196 8 3274 9
rect 3007 -74 3009 -72
rect 3061 -74 3063 -72
rect 3007 -81 3063 -74
rect 3107 -15 3163 0
rect 3107 -67 3109 -15
rect 3161 -67 3163 -15
rect 3107 -79 3163 -67
rect 3107 -110 3109 -79
rect 2961 -131 3109 -110
rect 3161 -110 3163 -79
rect 3207 -16 3263 8
rect 3207 -74 3209 -72
rect 3261 -74 3263 -72
rect 3207 -81 3263 -74
rect 3307 -15 3363 0
rect 3307 -67 3309 -15
rect 3361 -67 3363 -15
rect 3307 -79 3363 -67
rect 3307 -110 3309 -79
rect 3161 -131 3309 -110
rect 3361 -110 3363 -79
rect 3407 -16 3463 24
rect 3596 9 3607 65
rect 3663 9 3674 65
rect 3796 25 3807 81
rect 3863 25 3874 81
rect 4196 81 4274 82
rect 3796 24 3874 25
rect 3996 65 4074 66
rect 3596 8 3674 9
rect 3407 -74 3409 -72
rect 3461 -74 3463 -72
rect 3407 -81 3463 -74
rect 3507 -15 3563 0
rect 3507 -67 3509 -15
rect 3561 -67 3563 -15
rect 3507 -79 3563 -67
rect 3507 -110 3509 -79
rect 3361 -131 3509 -110
rect 3561 -110 3563 -79
rect 3607 -16 3663 8
rect 3607 -74 3609 -72
rect 3661 -74 3663 -72
rect 3607 -81 3663 -74
rect 3707 -15 3763 0
rect 3707 -67 3709 -15
rect 3761 -67 3763 -15
rect 3707 -79 3763 -67
rect 3707 -110 3709 -79
rect 3561 -131 3709 -110
rect 3761 -110 3763 -79
rect 3807 -16 3863 24
rect 3996 9 4007 65
rect 4063 9 4074 65
rect 4196 25 4207 81
rect 4263 25 4274 81
rect 4596 81 4674 82
rect 4196 24 4274 25
rect 4396 65 4474 66
rect 3996 8 4074 9
rect 3807 -74 3809 -72
rect 3861 -74 3863 -72
rect 3807 -81 3863 -74
rect 3907 -15 3963 0
rect 3907 -67 3909 -15
rect 3961 -67 3963 -15
rect 3907 -79 3963 -67
rect 3907 -110 3909 -79
rect 3761 -131 3909 -110
rect 3961 -110 3963 -79
rect 4007 -16 4063 8
rect 4007 -74 4009 -72
rect 4061 -74 4063 -72
rect 4007 -81 4063 -74
rect 4107 -15 4163 0
rect 4107 -67 4109 -15
rect 4161 -67 4163 -15
rect 4107 -79 4163 -67
rect 4107 -110 4109 -79
rect 3961 -131 4109 -110
rect 4161 -110 4163 -79
rect 4207 -16 4263 24
rect 4396 9 4407 65
rect 4463 9 4474 65
rect 4596 25 4607 81
rect 4663 25 4674 81
rect 4996 81 5074 82
rect 4596 24 4674 25
rect 4796 65 4874 66
rect 4396 8 4474 9
rect 4207 -74 4209 -72
rect 4261 -74 4263 -72
rect 4207 -81 4263 -74
rect 4307 -15 4363 0
rect 4307 -67 4309 -15
rect 4361 -67 4363 -15
rect 4307 -79 4363 -67
rect 4307 -110 4309 -79
rect 4161 -131 4309 -110
rect 4361 -110 4363 -79
rect 4407 -16 4463 8
rect 4407 -74 4409 -72
rect 4461 -74 4463 -72
rect 4407 -81 4463 -74
rect 4507 -15 4563 0
rect 4507 -67 4509 -15
rect 4561 -67 4563 -15
rect 4507 -79 4563 -67
rect 4507 -110 4509 -79
rect 4361 -131 4509 -110
rect 4561 -110 4563 -79
rect 4607 -16 4663 24
rect 4796 9 4807 65
rect 4863 9 4874 65
rect 4996 25 5007 81
rect 5063 25 5074 81
rect 5396 81 5474 82
rect 4996 24 5074 25
rect 5196 65 5274 66
rect 4796 8 4874 9
rect 4607 -74 4609 -72
rect 4661 -74 4663 -72
rect 4607 -81 4663 -74
rect 4707 -15 4763 0
rect 4707 -67 4709 -15
rect 4761 -67 4763 -15
rect 4707 -79 4763 -67
rect 4707 -110 4709 -79
rect 4561 -131 4709 -110
rect 4761 -110 4763 -79
rect 4807 -16 4863 8
rect 4807 -74 4809 -72
rect 4861 -74 4863 -72
rect 4807 -81 4863 -74
rect 4907 -15 4963 0
rect 4907 -67 4909 -15
rect 4961 -67 4963 -15
rect 4907 -79 4963 -67
rect 4907 -110 4909 -79
rect 4761 -131 4909 -110
rect 4961 -110 4963 -79
rect 5007 -16 5063 24
rect 5196 9 5207 65
rect 5263 9 5274 65
rect 5396 25 5407 81
rect 5463 25 5474 81
rect 5796 81 5874 82
rect 5396 24 5474 25
rect 5596 65 5674 66
rect 5196 8 5274 9
rect 5007 -74 5009 -72
rect 5061 -74 5063 -72
rect 5007 -81 5063 -74
rect 5107 -15 5163 0
rect 5107 -67 5109 -15
rect 5161 -67 5163 -15
rect 5107 -79 5163 -67
rect 5107 -110 5109 -79
rect 4961 -131 5109 -110
rect 5161 -110 5163 -79
rect 5207 -16 5263 8
rect 5207 -74 5209 -72
rect 5261 -74 5263 -72
rect 5207 -81 5263 -74
rect 5307 -15 5363 0
rect 5307 -67 5309 -15
rect 5361 -67 5363 -15
rect 5307 -79 5363 -67
rect 5307 -110 5309 -79
rect 5161 -131 5309 -110
rect 5361 -110 5363 -79
rect 5407 -16 5463 24
rect 5596 9 5607 65
rect 5663 9 5674 65
rect 5796 25 5807 81
rect 5863 25 5874 81
rect 6196 81 6274 82
rect 5796 24 5874 25
rect 5996 65 6074 66
rect 5596 8 5674 9
rect 5407 -74 5409 -72
rect 5461 -74 5463 -72
rect 5407 -81 5463 -74
rect 5507 -15 5563 0
rect 5507 -67 5509 -15
rect 5561 -67 5563 -15
rect 5507 -79 5563 -67
rect 5507 -110 5509 -79
rect 5361 -131 5509 -110
rect 5561 -110 5563 -79
rect 5607 -16 5663 8
rect 5607 -74 5609 -72
rect 5661 -74 5663 -72
rect 5607 -81 5663 -74
rect 5707 -15 5763 0
rect 5707 -67 5709 -15
rect 5761 -67 5763 -15
rect 5707 -79 5763 -67
rect 5707 -110 5709 -79
rect 5561 -131 5709 -110
rect 5761 -110 5763 -79
rect 5807 -16 5863 24
rect 5996 9 6007 65
rect 6063 9 6074 65
rect 6196 25 6207 81
rect 6263 25 6274 81
rect 6596 81 6674 82
rect 6196 24 6274 25
rect 6396 65 6474 66
rect 5996 8 6074 9
rect 5807 -74 5809 -72
rect 5861 -74 5863 -72
rect 5807 -81 5863 -74
rect 5907 -15 5963 0
rect 5907 -67 5909 -15
rect 5961 -67 5963 -15
rect 5907 -79 5963 -67
rect 5907 -110 5909 -79
rect 5761 -131 5909 -110
rect 5961 -110 5963 -79
rect 6007 -16 6063 8
rect 6007 -74 6009 -72
rect 6061 -74 6063 -72
rect 6007 -81 6063 -74
rect 6107 -15 6163 0
rect 6107 -67 6109 -15
rect 6161 -67 6163 -15
rect 6107 -79 6163 -67
rect 6107 -110 6109 -79
rect 5961 -131 6109 -110
rect 6161 -110 6163 -79
rect 6207 -16 6263 24
rect 6396 9 6407 65
rect 6463 9 6474 65
rect 6596 25 6607 81
rect 6663 25 6674 81
rect 6996 81 7074 82
rect 6596 24 6674 25
rect 6796 65 6874 66
rect 6396 8 6474 9
rect 6207 -74 6209 -72
rect 6261 -74 6263 -72
rect 6207 -81 6263 -74
rect 6307 -15 6363 0
rect 6307 -67 6309 -15
rect 6361 -67 6363 -15
rect 6307 -79 6363 -67
rect 6307 -110 6309 -79
rect 6161 -131 6309 -110
rect 6361 -110 6363 -79
rect 6407 -16 6463 8
rect 6407 -74 6409 -72
rect 6461 -74 6463 -72
rect 6407 -81 6463 -74
rect 6507 -15 6563 0
rect 6507 -67 6509 -15
rect 6561 -67 6563 -15
rect 6507 -79 6563 -67
rect 6507 -110 6509 -79
rect 6361 -131 6509 -110
rect 6561 -110 6563 -79
rect 6607 -16 6663 24
rect 6796 9 6807 65
rect 6863 9 6874 65
rect 6996 25 7007 81
rect 7063 25 7074 81
rect 7396 81 7474 82
rect 6996 24 7074 25
rect 7196 65 7274 66
rect 6796 8 6874 9
rect 6607 -74 6609 -72
rect 6661 -74 6663 -72
rect 6607 -81 6663 -74
rect 6707 -15 6763 0
rect 6707 -67 6709 -15
rect 6761 -67 6763 -15
rect 6707 -79 6763 -67
rect 6707 -110 6709 -79
rect 6561 -131 6709 -110
rect 6761 -110 6763 -79
rect 6807 -16 6863 8
rect 6807 -74 6809 -72
rect 6861 -74 6863 -72
rect 6807 -81 6863 -74
rect 6907 -15 6963 0
rect 6907 -67 6909 -15
rect 6961 -67 6963 -15
rect 6907 -79 6963 -67
rect 6907 -110 6909 -79
rect 6761 -131 6909 -110
rect 6961 -110 6963 -79
rect 7007 -16 7063 24
rect 7196 9 7207 65
rect 7263 9 7274 65
rect 7396 25 7407 81
rect 7463 25 7474 81
rect 7796 81 7874 82
rect 7396 24 7474 25
rect 7596 65 7674 66
rect 7196 8 7274 9
rect 7007 -74 7009 -72
rect 7061 -74 7063 -72
rect 7007 -81 7063 -74
rect 7107 -15 7163 0
rect 7107 -67 7109 -15
rect 7161 -67 7163 -15
rect 7107 -79 7163 -67
rect 7107 -110 7109 -79
rect 6961 -131 7109 -110
rect 7161 -110 7163 -79
rect 7207 -16 7263 8
rect 7207 -74 7209 -72
rect 7261 -74 7263 -72
rect 7207 -81 7263 -74
rect 7307 -15 7363 0
rect 7307 -67 7309 -15
rect 7361 -67 7363 -15
rect 7307 -79 7363 -67
rect 7307 -110 7309 -79
rect 7161 -131 7309 -110
rect 7361 -110 7363 -79
rect 7407 -16 7463 24
rect 7596 9 7607 65
rect 7663 9 7674 65
rect 7796 25 7807 81
rect 7863 25 7874 81
rect 8196 81 8274 82
rect 7796 24 7874 25
rect 7996 65 8074 66
rect 7596 8 7674 9
rect 7407 -74 7409 -72
rect 7461 -74 7463 -72
rect 7407 -81 7463 -74
rect 7507 -15 7563 0
rect 7507 -67 7509 -15
rect 7561 -67 7563 -15
rect 7507 -79 7563 -67
rect 7507 -110 7509 -79
rect 7361 -131 7509 -110
rect 7561 -110 7563 -79
rect 7607 -16 7663 8
rect 7607 -74 7609 -72
rect 7661 -74 7663 -72
rect 7607 -81 7663 -74
rect 7707 -15 7763 0
rect 7707 -67 7709 -15
rect 7761 -67 7763 -15
rect 7707 -79 7763 -67
rect 7707 -110 7709 -79
rect 7561 -131 7709 -110
rect 7761 -110 7763 -79
rect 7807 -16 7863 24
rect 7996 9 8007 65
rect 8063 9 8074 65
rect 8196 25 8207 81
rect 8263 25 8274 81
rect 8596 81 8674 82
rect 8196 24 8274 25
rect 8396 65 8474 66
rect 7996 8 8074 9
rect 7807 -74 7809 -72
rect 7861 -74 7863 -72
rect 7807 -81 7863 -74
rect 7907 -15 7963 0
rect 7907 -67 7909 -15
rect 7961 -67 7963 -15
rect 7907 -79 7963 -67
rect 7907 -110 7909 -79
rect 7761 -131 7909 -110
rect 7961 -110 7963 -79
rect 8007 -16 8063 8
rect 8007 -74 8009 -72
rect 8061 -74 8063 -72
rect 8007 -81 8063 -74
rect 8107 -15 8163 0
rect 8107 -67 8109 -15
rect 8161 -67 8163 -15
rect 8107 -79 8163 -67
rect 8107 -110 8109 -79
rect 7961 -131 8109 -110
rect 8161 -110 8163 -79
rect 8207 -16 8263 24
rect 8396 9 8407 65
rect 8463 9 8474 65
rect 8596 25 8607 81
rect 8663 25 8674 81
rect 8996 81 9074 82
rect 8596 24 8674 25
rect 8796 65 8874 66
rect 8396 8 8474 9
rect 8207 -74 8209 -72
rect 8261 -74 8263 -72
rect 8207 -81 8263 -74
rect 8307 -15 8363 0
rect 8307 -67 8309 -15
rect 8361 -67 8363 -15
rect 8307 -79 8363 -67
rect 8307 -110 8309 -79
rect 8161 -131 8309 -110
rect 8361 -110 8363 -79
rect 8407 -16 8463 8
rect 8407 -74 8409 -72
rect 8461 -74 8463 -72
rect 8407 -81 8463 -74
rect 8507 -15 8563 0
rect 8507 -67 8509 -15
rect 8561 -67 8563 -15
rect 8507 -79 8563 -67
rect 8507 -110 8509 -79
rect 8361 -131 8509 -110
rect 8561 -110 8563 -79
rect 8607 -16 8663 24
rect 8796 9 8807 65
rect 8863 9 8874 65
rect 8996 25 9007 81
rect 9063 25 9074 81
rect 9396 81 9474 82
rect 8996 24 9074 25
rect 9196 65 9274 66
rect 8796 8 8874 9
rect 8607 -74 8609 -72
rect 8661 -74 8663 -72
rect 8607 -81 8663 -74
rect 8707 -15 8763 0
rect 8707 -67 8709 -15
rect 8761 -67 8763 -15
rect 8707 -79 8763 -67
rect 8707 -110 8709 -79
rect 8561 -131 8709 -110
rect 8761 -110 8763 -79
rect 8807 -16 8863 8
rect 8807 -74 8809 -72
rect 8861 -74 8863 -72
rect 8807 -81 8863 -74
rect 8907 -15 8963 0
rect 8907 -67 8909 -15
rect 8961 -67 8963 -15
rect 8907 -79 8963 -67
rect 8907 -110 8909 -79
rect 8761 -131 8909 -110
rect 8961 -110 8963 -79
rect 9007 -16 9063 24
rect 9196 9 9207 65
rect 9263 9 9274 65
rect 9396 25 9407 81
rect 9463 25 9474 81
rect 9796 81 9874 82
rect 9396 24 9474 25
rect 9596 65 9674 66
rect 9196 8 9274 9
rect 9007 -74 9009 -72
rect 9061 -74 9063 -72
rect 9007 -81 9063 -74
rect 9107 -15 9163 0
rect 9107 -67 9109 -15
rect 9161 -67 9163 -15
rect 9107 -79 9163 -67
rect 9107 -110 9109 -79
rect 8961 -131 9109 -110
rect 9161 -110 9163 -79
rect 9207 -16 9263 8
rect 9207 -74 9209 -72
rect 9261 -74 9263 -72
rect 9207 -81 9263 -74
rect 9307 -15 9363 0
rect 9307 -67 9309 -15
rect 9361 -67 9363 -15
rect 9307 -79 9363 -67
rect 9307 -110 9309 -79
rect 9161 -131 9309 -110
rect 9361 -110 9363 -79
rect 9407 -16 9463 24
rect 9596 9 9607 65
rect 9663 9 9674 65
rect 9796 25 9807 81
rect 9863 25 9874 81
rect 10196 81 10274 82
rect 9796 24 9874 25
rect 9996 65 10074 66
rect 9596 8 9674 9
rect 9407 -74 9409 -72
rect 9461 -74 9463 -72
rect 9407 -81 9463 -74
rect 9507 -15 9563 0
rect 9507 -67 9509 -15
rect 9561 -67 9563 -15
rect 9507 -79 9563 -67
rect 9507 -110 9509 -79
rect 9361 -131 9509 -110
rect 9561 -110 9563 -79
rect 9607 -16 9663 8
rect 9607 -74 9609 -72
rect 9661 -74 9663 -72
rect 9607 -81 9663 -74
rect 9707 -15 9763 0
rect 9707 -67 9709 -15
rect 9761 -67 9763 -15
rect 9707 -79 9763 -67
rect 9707 -110 9709 -79
rect 9561 -131 9709 -110
rect 9761 -110 9763 -79
rect 9807 -16 9863 24
rect 9996 9 10007 65
rect 10063 9 10074 65
rect 10196 25 10207 81
rect 10263 25 10274 81
rect 10596 81 10674 82
rect 10196 24 10274 25
rect 10396 65 10474 66
rect 9996 8 10074 9
rect 9807 -74 9809 -72
rect 9861 -74 9863 -72
rect 9807 -81 9863 -74
rect 9907 -15 9963 0
rect 9907 -67 9909 -15
rect 9961 -67 9963 -15
rect 9907 -79 9963 -67
rect 9907 -110 9909 -79
rect 9761 -131 9909 -110
rect 9961 -110 9963 -79
rect 10007 -16 10063 8
rect 10007 -74 10009 -72
rect 10061 -74 10063 -72
rect 10007 -81 10063 -74
rect 10107 -15 10163 0
rect 10107 -67 10109 -15
rect 10161 -67 10163 -15
rect 10107 -79 10163 -67
rect 10107 -110 10109 -79
rect 9961 -131 10109 -110
rect 10161 -110 10163 -79
rect 10207 -16 10263 24
rect 10396 9 10407 65
rect 10463 9 10474 65
rect 10596 25 10607 81
rect 10663 25 10674 81
rect 10996 81 11074 82
rect 10596 24 10674 25
rect 10796 65 10874 66
rect 10396 8 10474 9
rect 10207 -74 10209 -72
rect 10261 -74 10263 -72
rect 10207 -81 10263 -74
rect 10307 -15 10363 0
rect 10307 -67 10309 -15
rect 10361 -67 10363 -15
rect 10307 -79 10363 -67
rect 10307 -110 10309 -79
rect 10161 -131 10309 -110
rect 10361 -110 10363 -79
rect 10407 -16 10463 8
rect 10407 -74 10409 -72
rect 10461 -74 10463 -72
rect 10407 -81 10463 -74
rect 10507 -15 10563 0
rect 10507 -67 10509 -15
rect 10561 -67 10563 -15
rect 10507 -79 10563 -67
rect 10507 -110 10509 -79
rect 10361 -131 10509 -110
rect 10561 -110 10563 -79
rect 10607 -16 10663 24
rect 10796 9 10807 65
rect 10863 9 10874 65
rect 10996 25 11007 81
rect 11063 25 11074 81
rect 11396 81 11474 82
rect 10996 24 11074 25
rect 11196 65 11274 66
rect 10796 8 10874 9
rect 10607 -74 10609 -72
rect 10661 -74 10663 -72
rect 10607 -81 10663 -74
rect 10707 -15 10763 0
rect 10707 -67 10709 -15
rect 10761 -67 10763 -15
rect 10707 -79 10763 -67
rect 10707 -110 10709 -79
rect 10561 -131 10709 -110
rect 10761 -110 10763 -79
rect 10807 -16 10863 8
rect 10807 -74 10809 -72
rect 10861 -74 10863 -72
rect 10807 -81 10863 -74
rect 10907 -15 10963 0
rect 10907 -67 10909 -15
rect 10961 -67 10963 -15
rect 10907 -79 10963 -67
rect 10907 -110 10909 -79
rect 10761 -131 10909 -110
rect 10961 -110 10963 -79
rect 11007 -16 11063 24
rect 11196 9 11207 65
rect 11263 9 11274 65
rect 11396 25 11407 81
rect 11463 25 11474 81
rect 11796 81 11874 82
rect 11396 24 11474 25
rect 11596 65 11674 66
rect 11196 8 11274 9
rect 11007 -74 11009 -72
rect 11061 -74 11063 -72
rect 11007 -81 11063 -74
rect 11107 -15 11163 0
rect 11107 -67 11109 -15
rect 11161 -67 11163 -15
rect 11107 -79 11163 -67
rect 11107 -110 11109 -79
rect 10961 -131 11109 -110
rect 11161 -110 11163 -79
rect 11207 -16 11263 8
rect 11207 -74 11209 -72
rect 11261 -74 11263 -72
rect 11207 -81 11263 -74
rect 11307 -15 11363 0
rect 11307 -67 11309 -15
rect 11361 -67 11363 -15
rect 11307 -79 11363 -67
rect 11307 -110 11309 -79
rect 11161 -131 11309 -110
rect 11361 -110 11363 -79
rect 11407 -16 11463 24
rect 11596 9 11607 65
rect 11663 9 11674 65
rect 11796 25 11807 81
rect 11863 25 11874 81
rect 12196 81 12274 82
rect 11796 24 11874 25
rect 11996 65 12074 66
rect 11596 8 11674 9
rect 11407 -74 11409 -72
rect 11461 -74 11463 -72
rect 11407 -81 11463 -74
rect 11507 -15 11563 0
rect 11507 -67 11509 -15
rect 11561 -67 11563 -15
rect 11507 -79 11563 -67
rect 11507 -110 11509 -79
rect 11361 -131 11509 -110
rect 11561 -110 11563 -79
rect 11607 -16 11663 8
rect 11607 -74 11609 -72
rect 11661 -74 11663 -72
rect 11607 -81 11663 -74
rect 11707 -15 11763 0
rect 11707 -67 11709 -15
rect 11761 -67 11763 -15
rect 11707 -79 11763 -67
rect 11707 -110 11709 -79
rect 11561 -131 11709 -110
rect 11761 -110 11763 -79
rect 11807 -16 11863 24
rect 11996 9 12007 65
rect 12063 9 12074 65
rect 12196 25 12207 81
rect 12263 25 12274 81
rect 12596 81 12674 82
rect 12196 24 12274 25
rect 12396 65 12474 66
rect 11996 8 12074 9
rect 11807 -74 11809 -72
rect 11861 -74 11863 -72
rect 11807 -81 11863 -74
rect 11907 -15 11963 0
rect 11907 -67 11909 -15
rect 11961 -67 11963 -15
rect 11907 -79 11963 -67
rect 11907 -110 11909 -79
rect 11761 -131 11909 -110
rect 11961 -110 11963 -79
rect 12007 -16 12063 8
rect 12007 -74 12009 -72
rect 12061 -74 12063 -72
rect 12007 -81 12063 -74
rect 12107 -15 12163 0
rect 12107 -67 12109 -15
rect 12161 -67 12163 -15
rect 12107 -79 12163 -67
rect 12107 -110 12109 -79
rect 11961 -131 12109 -110
rect 12161 -110 12163 -79
rect 12207 -16 12263 24
rect 12396 9 12407 65
rect 12463 9 12474 65
rect 12596 25 12607 81
rect 12663 25 12674 81
rect 12596 24 12674 25
rect 12396 8 12474 9
rect 12207 -74 12209 -72
rect 12261 -74 12263 -72
rect 12207 -81 12263 -74
rect 12307 -15 12363 0
rect 12307 -67 12309 -15
rect 12361 -67 12363 -15
rect 12307 -79 12363 -67
rect 12307 -110 12309 -79
rect 12161 -131 12309 -110
rect 12361 -110 12363 -79
rect 12407 -16 12463 8
rect 12407 -74 12409 -72
rect 12461 -74 12463 -72
rect 12407 -81 12463 -74
rect 12507 -15 12563 0
rect 12507 -67 12509 -15
rect 12561 -67 12563 -15
rect 12507 -79 12563 -67
rect 12507 -110 12509 -79
rect 12361 -131 12509 -110
rect 12561 -110 12563 -79
rect 12607 -16 12663 24
rect 12607 -74 12609 -72
rect 12661 -74 12663 -72
rect 12607 -81 12663 -74
rect 12707 -15 12763 0
rect 12707 -67 12709 -15
rect 12761 -67 12763 -15
rect 12707 -79 12763 -67
rect 12707 -110 12709 -79
rect 12561 -131 12709 -110
rect 12761 -110 12763 -79
rect 12761 -131 12808 -110
rect -138 -143 12808 -131
rect -138 -145 -91 -143
rect -39 -145 109 -143
rect 161 -145 309 -143
rect 361 -145 509 -143
rect 561 -145 709 -143
rect 761 -145 909 -143
rect 961 -145 1109 -143
rect 1161 -145 1309 -143
rect 1361 -145 1509 -143
rect 1561 -145 1709 -143
rect 1761 -145 1909 -143
rect 1961 -145 2109 -143
rect 2161 -145 2309 -143
rect 2361 -145 2509 -143
rect 2561 -145 2709 -143
rect 2761 -145 2909 -143
rect 2961 -145 3109 -143
rect 3161 -145 3309 -143
rect 3361 -145 3509 -143
rect 3561 -145 3709 -143
rect 3761 -145 3909 -143
rect 3961 -145 4109 -143
rect 4161 -145 4309 -143
rect 4361 -145 4509 -143
rect 4561 -145 4709 -143
rect 4761 -145 4909 -143
rect 4961 -145 5109 -143
rect 5161 -145 5309 -143
rect 5361 -145 5509 -143
rect 5561 -145 5709 -143
rect 5761 -145 5909 -143
rect 5961 -145 6109 -143
rect 6161 -145 6309 -143
rect 6361 -145 6509 -143
rect 6561 -145 6709 -143
rect 6761 -145 6909 -143
rect 6961 -145 7109 -143
rect 7161 -145 7309 -143
rect 7361 -145 7509 -143
rect 7561 -145 7709 -143
rect 7761 -145 7909 -143
rect 7961 -145 8109 -143
rect 8161 -145 8309 -143
rect 8361 -145 8509 -143
rect 8561 -145 8709 -143
rect 8761 -145 8909 -143
rect 8961 -145 9109 -143
rect 9161 -145 9309 -143
rect 9361 -145 9509 -143
rect 9561 -145 9709 -143
rect 9761 -145 9909 -143
rect 9961 -145 10109 -143
rect 10161 -145 10309 -143
rect 10361 -145 10509 -143
rect 10561 -145 10709 -143
rect 10761 -145 10909 -143
rect 10961 -145 11109 -143
rect 11161 -145 11309 -143
rect 11361 -145 11509 -143
rect 11561 -145 11709 -143
rect 11761 -145 11909 -143
rect 11961 -145 12109 -143
rect 12161 -145 12309 -143
rect 12361 -145 12509 -143
rect 12561 -145 12709 -143
rect 12761 -145 12808 -143
rect -138 -201 -133 -145
rect -77 -201 -53 -195
rect 3 -201 67 -145
rect 123 -201 147 -195
rect 203 -201 267 -145
rect 323 -201 347 -195
rect 403 -201 467 -145
rect 523 -201 547 -195
rect 603 -201 667 -145
rect 723 -201 747 -195
rect 803 -201 867 -145
rect 923 -201 947 -195
rect 1003 -201 1067 -145
rect 1123 -201 1147 -195
rect 1203 -201 1267 -145
rect 1323 -201 1347 -195
rect 1403 -201 1467 -145
rect 1523 -201 1547 -195
rect 1603 -201 1667 -145
rect 1723 -201 1747 -195
rect 1803 -201 1867 -145
rect 1923 -201 1947 -195
rect 2003 -201 2067 -145
rect 2123 -201 2147 -195
rect 2203 -201 2267 -145
rect 2323 -201 2347 -195
rect 2403 -201 2467 -145
rect 2523 -201 2547 -195
rect 2603 -201 2667 -145
rect 2723 -201 2747 -195
rect 2803 -201 2867 -145
rect 2923 -201 2947 -195
rect 3003 -201 3067 -145
rect 3123 -201 3147 -195
rect 3203 -201 3267 -145
rect 3323 -201 3347 -195
rect 3403 -201 3467 -145
rect 3523 -201 3547 -195
rect 3603 -201 3667 -145
rect 3723 -201 3747 -195
rect 3803 -201 3867 -145
rect 3923 -201 3947 -195
rect 4003 -201 4067 -145
rect 4123 -201 4147 -195
rect 4203 -201 4267 -145
rect 4323 -201 4347 -195
rect 4403 -201 4467 -145
rect 4523 -201 4547 -195
rect 4603 -201 4667 -145
rect 4723 -201 4747 -195
rect 4803 -201 4867 -145
rect 4923 -201 4947 -195
rect 5003 -201 5067 -145
rect 5123 -201 5147 -195
rect 5203 -201 5267 -145
rect 5323 -201 5347 -195
rect 5403 -201 5467 -145
rect 5523 -201 5547 -195
rect 5603 -201 5667 -145
rect 5723 -201 5747 -195
rect 5803 -201 5867 -145
rect 5923 -201 5947 -195
rect 6003 -201 6067 -145
rect 6123 -201 6147 -195
rect 6203 -201 6267 -145
rect 6323 -201 6347 -195
rect 6403 -201 6467 -145
rect 6523 -201 6547 -195
rect 6603 -201 6667 -145
rect 6723 -201 6747 -195
rect 6803 -201 6867 -145
rect 6923 -201 6947 -195
rect 7003 -201 7067 -145
rect 7123 -201 7147 -195
rect 7203 -201 7267 -145
rect 7323 -201 7347 -195
rect 7403 -201 7467 -145
rect 7523 -201 7547 -195
rect 7603 -201 7667 -145
rect 7723 -201 7747 -195
rect 7803 -201 7867 -145
rect 7923 -201 7947 -195
rect 8003 -201 8067 -145
rect 8123 -201 8147 -195
rect 8203 -201 8267 -145
rect 8323 -201 8347 -195
rect 8403 -201 8467 -145
rect 8523 -201 8547 -195
rect 8603 -201 8667 -145
rect 8723 -201 8747 -195
rect 8803 -201 8867 -145
rect 8923 -201 8947 -195
rect 9003 -201 9067 -145
rect 9123 -201 9147 -195
rect 9203 -201 9267 -145
rect 9323 -201 9347 -195
rect 9403 -201 9467 -145
rect 9523 -201 9547 -195
rect 9603 -201 9667 -145
rect 9723 -201 9747 -195
rect 9803 -201 9867 -145
rect 9923 -201 9947 -195
rect 10003 -201 10067 -145
rect 10123 -201 10147 -195
rect 10203 -201 10267 -145
rect 10323 -201 10347 -195
rect 10403 -201 10467 -145
rect 10523 -201 10547 -195
rect 10603 -201 10667 -145
rect 10723 -201 10747 -195
rect 10803 -201 10867 -145
rect 10923 -201 10947 -195
rect 11003 -201 11067 -145
rect 11123 -201 11147 -195
rect 11203 -201 11267 -145
rect 11323 -201 11347 -195
rect 11403 -201 11467 -145
rect 11523 -201 11547 -195
rect 11603 -201 11667 -145
rect 11723 -201 11747 -195
rect 11803 -201 11867 -145
rect 11923 -201 11947 -195
rect 12003 -201 12067 -145
rect 12123 -201 12147 -195
rect 12203 -201 12267 -145
rect 12323 -201 12347 -195
rect 12403 -201 12467 -145
rect 12523 -201 12547 -195
rect 12603 -201 12667 -145
rect 12723 -201 12747 -195
rect 12803 -201 12808 -145
rect -138 -210 12808 -201
rect 14526 -197 14697 -188
rect -81 -291 -75 -239
rect -23 -291 61 -239
rect 119 -291 125 -239
rect 177 -291 261 -239
rect 319 -291 325 -239
rect 377 -291 461 -239
rect 519 -291 525 -239
rect 577 -291 661 -239
rect 719 -291 725 -239
rect 777 -291 861 -239
rect 919 -291 925 -239
rect 977 -291 1061 -239
rect 1119 -291 1125 -239
rect 1177 -291 1261 -239
rect 1319 -291 1325 -239
rect 1377 -291 1461 -239
rect 1519 -291 1525 -239
rect 1577 -291 1661 -239
rect 1719 -291 1725 -239
rect 1777 -291 1861 -239
rect 1919 -291 1925 -239
rect 1977 -291 2061 -239
rect 2119 -291 2125 -239
rect 2177 -291 2261 -239
rect 2319 -291 2325 -239
rect 2377 -291 2461 -239
rect 2519 -291 2525 -239
rect 2577 -291 2661 -239
rect 2719 -291 2725 -239
rect 2777 -291 2861 -239
rect 2919 -291 2925 -239
rect 2977 -291 3061 -239
rect 3119 -291 3125 -239
rect 3177 -291 3261 -239
rect 3319 -291 3325 -239
rect 3377 -291 3461 -239
rect 3519 -291 3525 -239
rect 3577 -291 3661 -239
rect 3719 -291 3725 -239
rect 3777 -291 3861 -239
rect 3919 -291 3925 -239
rect 3977 -291 4061 -239
rect 4119 -291 4125 -239
rect 4177 -291 4261 -239
rect 4319 -291 4325 -239
rect 4377 -291 4461 -239
rect 4519 -291 4525 -239
rect 4577 -291 4661 -239
rect 4719 -291 4725 -239
rect 4777 -291 4861 -239
rect 4919 -291 4925 -239
rect 4977 -291 5061 -239
rect 5119 -291 5125 -239
rect 5177 -291 5261 -239
rect 5319 -291 5325 -239
rect 5377 -291 5461 -239
rect 5519 -291 5525 -239
rect 5577 -291 5661 -239
rect 5719 -291 5725 -239
rect 5777 -291 5861 -239
rect 5919 -291 5925 -239
rect 5977 -291 6061 -239
rect 6119 -291 6125 -239
rect 6177 -291 6261 -239
rect 6319 -291 6325 -239
rect 6377 -291 6461 -239
rect 6519 -291 6525 -239
rect 6577 -291 6661 -239
rect 6719 -291 6725 -239
rect 6777 -291 6861 -239
rect 6919 -291 6925 -239
rect 6977 -291 7061 -239
rect 7119 -291 7125 -239
rect 7177 -291 7261 -239
rect 7319 -291 7325 -239
rect 7377 -291 7461 -239
rect 7519 -291 7525 -239
rect 7577 -291 7661 -239
rect 7719 -291 7725 -239
rect 7777 -291 7861 -239
rect 7919 -291 7925 -239
rect 7977 -291 8061 -239
rect 8119 -291 8125 -239
rect 8177 -291 8261 -239
rect 8319 -291 8325 -239
rect 8377 -291 8461 -239
rect 8519 -291 8525 -239
rect 8577 -291 8661 -239
rect 8719 -291 8725 -239
rect 8777 -291 8861 -239
rect 8919 -291 8925 -239
rect 8977 -291 9061 -239
rect 9119 -291 9125 -239
rect 9177 -291 9261 -239
rect 9319 -291 9325 -239
rect 9377 -291 9461 -239
rect 9519 -291 9525 -239
rect 9577 -291 9661 -239
rect 9719 -291 9725 -239
rect 9777 -291 9861 -239
rect 9919 -291 9925 -239
rect 9977 -291 10061 -239
rect 10119 -291 10125 -239
rect 10177 -291 10261 -239
rect 10319 -291 10325 -239
rect 10377 -291 10461 -239
rect 10519 -291 10525 -239
rect 10577 -291 10661 -239
rect 10719 -291 10725 -239
rect 10777 -291 10861 -239
rect 10919 -291 10925 -239
rect 10977 -291 11061 -239
rect 11119 -291 11125 -239
rect 11177 -291 11261 -239
rect 11319 -291 11325 -239
rect 11377 -291 11461 -239
rect 11519 -291 11525 -239
rect 11577 -291 11661 -239
rect 11719 -291 11725 -239
rect 11777 -291 11861 -239
rect 11919 -291 11925 -239
rect 11977 -291 12061 -239
rect 12119 -291 12125 -239
rect 12177 -291 12261 -239
rect 12319 -291 12325 -239
rect 12377 -291 12461 -239
rect 12519 -291 12525 -239
rect 12577 -291 12661 -239
rect 14526 -253 14543 -197
rect 14599 -199 14623 -197
rect 14605 -251 14617 -199
rect 14599 -253 14623 -251
rect 14679 -253 14697 -197
rect 14526 -262 14697 -253
rect 14805 -197 15136 -188
rect 14805 -199 14822 -197
rect 14878 -199 14902 -197
rect 14958 -199 14982 -197
rect 15038 -199 15062 -197
rect 15118 -199 15136 -197
rect 14805 -251 14816 -199
rect 14878 -251 14880 -199
rect 15060 -251 15062 -199
rect 15124 -251 15136 -199
rect 14805 -253 14822 -251
rect 14878 -253 14902 -251
rect 14958 -253 14982 -251
rect 15038 -253 15062 -251
rect 15118 -253 15136 -251
rect 14805 -262 15136 -253
rect 15206 -197 15537 -188
rect 15206 -199 15223 -197
rect 15279 -199 15303 -197
rect 15359 -199 15383 -197
rect 15439 -199 15463 -197
rect 15519 -199 15537 -197
rect 15206 -251 15217 -199
rect 15279 -251 15281 -199
rect 15461 -251 15463 -199
rect 15525 -251 15537 -199
rect 15206 -253 15223 -251
rect 15279 -253 15303 -251
rect 15359 -253 15383 -251
rect 15439 -253 15463 -251
rect 15519 -253 15537 -251
rect 15206 -262 15537 -253
rect 15645 -197 15816 -188
rect 15645 -253 15662 -197
rect 15718 -199 15742 -197
rect 15724 -251 15736 -199
rect 15718 -253 15742 -251
rect 15798 -253 15816 -197
rect 15645 -262 15816 -253
rect -93 -326 -37 -320
rect -93 -348 -91 -326
rect -39 -348 -37 -326
rect -93 -428 -91 -404
rect -39 -428 -37 -404
rect -93 -506 -91 -484
rect -39 -506 -37 -484
rect -93 -512 -37 -506
rect 9 -828 61 -291
rect 107 -326 163 -320
rect 107 -348 109 -326
rect 161 -348 163 -326
rect 107 -428 109 -404
rect 161 -428 163 -404
rect 107 -506 109 -484
rect 161 -506 163 -484
rect 107 -512 163 -506
rect 209 -828 261 -291
rect 307 -326 363 -320
rect 307 -348 309 -326
rect 361 -348 363 -326
rect 307 -428 309 -404
rect 361 -428 363 -404
rect 307 -506 309 -484
rect 361 -506 363 -484
rect 307 -512 363 -506
rect 409 -828 461 -291
rect 507 -326 563 -320
rect 507 -348 509 -326
rect 561 -348 563 -326
rect 507 -428 509 -404
rect 561 -428 563 -404
rect 507 -506 509 -484
rect 561 -506 563 -484
rect 507 -512 563 -506
rect 609 -828 661 -291
rect 707 -326 763 -320
rect 707 -348 709 -326
rect 761 -348 763 -326
rect 707 -428 709 -404
rect 761 -428 763 -404
rect 707 -506 709 -484
rect 761 -506 763 -484
rect 707 -512 763 -506
rect 809 -828 861 -291
rect 907 -326 963 -320
rect 907 -348 909 -326
rect 961 -348 963 -326
rect 907 -428 909 -404
rect 961 -428 963 -404
rect 907 -506 909 -484
rect 961 -506 963 -484
rect 907 -512 963 -506
rect 1009 -828 1061 -291
rect 1107 -326 1163 -320
rect 1107 -348 1109 -326
rect 1161 -348 1163 -326
rect 1107 -428 1109 -404
rect 1161 -428 1163 -404
rect 1107 -506 1109 -484
rect 1161 -506 1163 -484
rect 1107 -512 1163 -506
rect 1209 -828 1261 -291
rect 1307 -326 1363 -320
rect 1307 -348 1309 -326
rect 1361 -348 1363 -326
rect 1307 -428 1309 -404
rect 1361 -428 1363 -404
rect 1307 -506 1309 -484
rect 1361 -506 1363 -484
rect 1307 -512 1363 -506
rect 1409 -828 1461 -291
rect 1507 -326 1563 -320
rect 1507 -348 1509 -326
rect 1561 -348 1563 -326
rect 1507 -428 1509 -404
rect 1561 -428 1563 -404
rect 1507 -506 1509 -484
rect 1561 -506 1563 -484
rect 1507 -512 1563 -506
rect 1609 -828 1661 -291
rect 1707 -326 1763 -320
rect 1707 -348 1709 -326
rect 1761 -348 1763 -326
rect 1707 -428 1709 -404
rect 1761 -428 1763 -404
rect 1707 -506 1709 -484
rect 1761 -506 1763 -484
rect 1707 -512 1763 -506
rect 1809 -828 1861 -291
rect 1907 -326 1963 -320
rect 1907 -348 1909 -326
rect 1961 -348 1963 -326
rect 1907 -428 1909 -404
rect 1961 -428 1963 -404
rect 1907 -506 1909 -484
rect 1961 -506 1963 -484
rect 1907 -512 1963 -506
rect 2009 -828 2061 -291
rect 2107 -326 2163 -320
rect 2107 -348 2109 -326
rect 2161 -348 2163 -326
rect 2107 -428 2109 -404
rect 2161 -428 2163 -404
rect 2107 -506 2109 -484
rect 2161 -506 2163 -484
rect 2107 -512 2163 -506
rect 2209 -828 2261 -291
rect 2307 -326 2363 -320
rect 2307 -348 2309 -326
rect 2361 -348 2363 -326
rect 2307 -428 2309 -404
rect 2361 -428 2363 -404
rect 2307 -506 2309 -484
rect 2361 -506 2363 -484
rect 2307 -512 2363 -506
rect 2409 -828 2461 -291
rect 2507 -326 2563 -320
rect 2507 -348 2509 -326
rect 2561 -348 2563 -326
rect 2507 -428 2509 -404
rect 2561 -428 2563 -404
rect 2507 -506 2509 -484
rect 2561 -506 2563 -484
rect 2507 -512 2563 -506
rect 2609 -828 2661 -291
rect 2707 -326 2763 -320
rect 2707 -348 2709 -326
rect 2761 -348 2763 -326
rect 2707 -428 2709 -404
rect 2761 -428 2763 -404
rect 2707 -506 2709 -484
rect 2761 -506 2763 -484
rect 2707 -512 2763 -506
rect 2809 -828 2861 -291
rect 2907 -326 2963 -320
rect 2907 -348 2909 -326
rect 2961 -348 2963 -326
rect 2907 -428 2909 -404
rect 2961 -428 2963 -404
rect 2907 -506 2909 -484
rect 2961 -506 2963 -484
rect 2907 -512 2963 -506
rect 3009 -828 3061 -291
rect 3107 -326 3163 -320
rect 3107 -348 3109 -326
rect 3161 -348 3163 -326
rect 3107 -428 3109 -404
rect 3161 -428 3163 -404
rect 3107 -506 3109 -484
rect 3161 -506 3163 -484
rect 3107 -512 3163 -506
rect 3209 -828 3261 -291
rect 3307 -326 3363 -320
rect 3307 -348 3309 -326
rect 3361 -348 3363 -326
rect 3307 -428 3309 -404
rect 3361 -428 3363 -404
rect 3307 -506 3309 -484
rect 3361 -506 3363 -484
rect 3307 -512 3363 -506
rect 3409 -828 3461 -291
rect 3507 -326 3563 -320
rect 3507 -348 3509 -326
rect 3561 -348 3563 -326
rect 3507 -428 3509 -404
rect 3561 -428 3563 -404
rect 3507 -506 3509 -484
rect 3561 -506 3563 -484
rect 3507 -512 3563 -506
rect 3609 -828 3661 -291
rect 3707 -326 3763 -320
rect 3707 -348 3709 -326
rect 3761 -348 3763 -326
rect 3707 -428 3709 -404
rect 3761 -428 3763 -404
rect 3707 -506 3709 -484
rect 3761 -506 3763 -484
rect 3707 -512 3763 -506
rect 3809 -828 3861 -291
rect 3907 -326 3963 -320
rect 3907 -348 3909 -326
rect 3961 -348 3963 -326
rect 3907 -428 3909 -404
rect 3961 -428 3963 -404
rect 3907 -506 3909 -484
rect 3961 -506 3963 -484
rect 3907 -512 3963 -506
rect 4009 -828 4061 -291
rect 4107 -326 4163 -320
rect 4107 -348 4109 -326
rect 4161 -348 4163 -326
rect 4107 -428 4109 -404
rect 4161 -428 4163 -404
rect 4107 -506 4109 -484
rect 4161 -506 4163 -484
rect 4107 -512 4163 -506
rect 4209 -828 4261 -291
rect 4307 -326 4363 -320
rect 4307 -348 4309 -326
rect 4361 -348 4363 -326
rect 4307 -428 4309 -404
rect 4361 -428 4363 -404
rect 4307 -506 4309 -484
rect 4361 -506 4363 -484
rect 4307 -512 4363 -506
rect 4409 -828 4461 -291
rect 4507 -326 4563 -320
rect 4507 -348 4509 -326
rect 4561 -348 4563 -326
rect 4507 -428 4509 -404
rect 4561 -428 4563 -404
rect 4507 -506 4509 -484
rect 4561 -506 4563 -484
rect 4507 -512 4563 -506
rect 4609 -828 4661 -291
rect 4707 -326 4763 -320
rect 4707 -348 4709 -326
rect 4761 -348 4763 -326
rect 4707 -428 4709 -404
rect 4761 -428 4763 -404
rect 4707 -506 4709 -484
rect 4761 -506 4763 -484
rect 4707 -512 4763 -506
rect 4809 -828 4861 -291
rect 4907 -326 4963 -320
rect 4907 -348 4909 -326
rect 4961 -348 4963 -326
rect 4907 -428 4909 -404
rect 4961 -428 4963 -404
rect 4907 -506 4909 -484
rect 4961 -506 4963 -484
rect 4907 -512 4963 -506
rect 5009 -828 5061 -291
rect 5107 -326 5163 -320
rect 5107 -348 5109 -326
rect 5161 -348 5163 -326
rect 5107 -428 5109 -404
rect 5161 -428 5163 -404
rect 5107 -506 5109 -484
rect 5161 -506 5163 -484
rect 5107 -512 5163 -506
rect 5209 -828 5261 -291
rect 5307 -326 5363 -320
rect 5307 -348 5309 -326
rect 5361 -348 5363 -326
rect 5307 -428 5309 -404
rect 5361 -428 5363 -404
rect 5307 -506 5309 -484
rect 5361 -506 5363 -484
rect 5307 -512 5363 -506
rect 5409 -828 5461 -291
rect 5507 -326 5563 -320
rect 5507 -348 5509 -326
rect 5561 -348 5563 -326
rect 5507 -428 5509 -404
rect 5561 -428 5563 -404
rect 5507 -506 5509 -484
rect 5561 -506 5563 -484
rect 5507 -512 5563 -506
rect 5609 -828 5661 -291
rect 5707 -326 5763 -320
rect 5707 -348 5709 -326
rect 5761 -348 5763 -326
rect 5707 -428 5709 -404
rect 5761 -428 5763 -404
rect 5707 -506 5709 -484
rect 5761 -506 5763 -484
rect 5707 -512 5763 -506
rect 5809 -828 5861 -291
rect 5907 -326 5963 -320
rect 5907 -348 5909 -326
rect 5961 -348 5963 -326
rect 5907 -428 5909 -404
rect 5961 -428 5963 -404
rect 5907 -506 5909 -484
rect 5961 -506 5963 -484
rect 5907 -512 5963 -506
rect 6009 -828 6061 -291
rect 6107 -326 6163 -320
rect 6107 -348 6109 -326
rect 6161 -348 6163 -326
rect 6107 -428 6109 -404
rect 6161 -428 6163 -404
rect 6107 -506 6109 -484
rect 6161 -506 6163 -484
rect 6107 -512 6163 -506
rect 6209 -828 6261 -291
rect 6307 -326 6363 -320
rect 6307 -348 6309 -326
rect 6361 -348 6363 -326
rect 6307 -428 6309 -404
rect 6361 -428 6363 -404
rect 6307 -506 6309 -484
rect 6361 -506 6363 -484
rect 6307 -512 6363 -506
rect 6409 -828 6461 -291
rect 6507 -326 6563 -320
rect 6507 -348 6509 -326
rect 6561 -348 6563 -326
rect 6507 -428 6509 -404
rect 6561 -428 6563 -404
rect 6507 -506 6509 -484
rect 6561 -506 6563 -484
rect 6507 -512 6563 -506
rect 6609 -828 6661 -291
rect 6707 -326 6763 -320
rect 6707 -348 6709 -326
rect 6761 -348 6763 -326
rect 6707 -428 6709 -404
rect 6761 -428 6763 -404
rect 6707 -506 6709 -484
rect 6761 -506 6763 -484
rect 6707 -512 6763 -506
rect 6809 -828 6861 -291
rect 6907 -326 6963 -320
rect 6907 -348 6909 -326
rect 6961 -348 6963 -326
rect 6907 -428 6909 -404
rect 6961 -428 6963 -404
rect 6907 -506 6909 -484
rect 6961 -506 6963 -484
rect 6907 -512 6963 -506
rect 7009 -828 7061 -291
rect 7107 -326 7163 -320
rect 7107 -348 7109 -326
rect 7161 -348 7163 -326
rect 7107 -428 7109 -404
rect 7161 -428 7163 -404
rect 7107 -506 7109 -484
rect 7161 -506 7163 -484
rect 7107 -512 7163 -506
rect 7209 -828 7261 -291
rect 7307 -326 7363 -320
rect 7307 -348 7309 -326
rect 7361 -348 7363 -326
rect 7307 -428 7309 -404
rect 7361 -428 7363 -404
rect 7307 -506 7309 -484
rect 7361 -506 7363 -484
rect 7307 -512 7363 -506
rect 7409 -828 7461 -291
rect 7507 -326 7563 -320
rect 7507 -348 7509 -326
rect 7561 -348 7563 -326
rect 7507 -428 7509 -404
rect 7561 -428 7563 -404
rect 7507 -506 7509 -484
rect 7561 -506 7563 -484
rect 7507 -512 7563 -506
rect 7609 -828 7661 -291
rect 7707 -326 7763 -320
rect 7707 -348 7709 -326
rect 7761 -348 7763 -326
rect 7707 -428 7709 -404
rect 7761 -428 7763 -404
rect 7707 -506 7709 -484
rect 7761 -506 7763 -484
rect 7707 -512 7763 -506
rect 7809 -828 7861 -291
rect 7907 -326 7963 -320
rect 7907 -348 7909 -326
rect 7961 -348 7963 -326
rect 7907 -428 7909 -404
rect 7961 -428 7963 -404
rect 7907 -506 7909 -484
rect 7961 -506 7963 -484
rect 7907 -512 7963 -506
rect 8009 -828 8061 -291
rect 8107 -326 8163 -320
rect 8107 -348 8109 -326
rect 8161 -348 8163 -326
rect 8107 -428 8109 -404
rect 8161 -428 8163 -404
rect 8107 -506 8109 -484
rect 8161 -506 8163 -484
rect 8107 -512 8163 -506
rect 8209 -828 8261 -291
rect 8307 -326 8363 -320
rect 8307 -348 8309 -326
rect 8361 -348 8363 -326
rect 8307 -428 8309 -404
rect 8361 -428 8363 -404
rect 8307 -506 8309 -484
rect 8361 -506 8363 -484
rect 8307 -512 8363 -506
rect 8409 -828 8461 -291
rect 8507 -326 8563 -320
rect 8507 -348 8509 -326
rect 8561 -348 8563 -326
rect 8507 -428 8509 -404
rect 8561 -428 8563 -404
rect 8507 -506 8509 -484
rect 8561 -506 8563 -484
rect 8507 -512 8563 -506
rect 8609 -828 8661 -291
rect 8707 -326 8763 -320
rect 8707 -348 8709 -326
rect 8761 -348 8763 -326
rect 8707 -428 8709 -404
rect 8761 -428 8763 -404
rect 8707 -506 8709 -484
rect 8761 -506 8763 -484
rect 8707 -512 8763 -506
rect 8809 -828 8861 -291
rect 8907 -326 8963 -320
rect 8907 -348 8909 -326
rect 8961 -348 8963 -326
rect 8907 -428 8909 -404
rect 8961 -428 8963 -404
rect 8907 -506 8909 -484
rect 8961 -506 8963 -484
rect 8907 -512 8963 -506
rect 9009 -828 9061 -291
rect 9107 -326 9163 -320
rect 9107 -348 9109 -326
rect 9161 -348 9163 -326
rect 9107 -428 9109 -404
rect 9161 -428 9163 -404
rect 9107 -506 9109 -484
rect 9161 -506 9163 -484
rect 9107 -512 9163 -506
rect 9209 -828 9261 -291
rect 9307 -326 9363 -320
rect 9307 -348 9309 -326
rect 9361 -348 9363 -326
rect 9307 -428 9309 -404
rect 9361 -428 9363 -404
rect 9307 -506 9309 -484
rect 9361 -506 9363 -484
rect 9307 -512 9363 -506
rect 9409 -828 9461 -291
rect 9507 -326 9563 -320
rect 9507 -348 9509 -326
rect 9561 -348 9563 -326
rect 9507 -428 9509 -404
rect 9561 -428 9563 -404
rect 9507 -506 9509 -484
rect 9561 -506 9563 -484
rect 9507 -512 9563 -506
rect 9609 -828 9661 -291
rect 9707 -326 9763 -320
rect 9707 -348 9709 -326
rect 9761 -348 9763 -326
rect 9707 -428 9709 -404
rect 9761 -428 9763 -404
rect 9707 -506 9709 -484
rect 9761 -506 9763 -484
rect 9707 -512 9763 -506
rect 9809 -828 9861 -291
rect 9907 -326 9963 -320
rect 9907 -348 9909 -326
rect 9961 -348 9963 -326
rect 9907 -428 9909 -404
rect 9961 -428 9963 -404
rect 9907 -506 9909 -484
rect 9961 -506 9963 -484
rect 9907 -512 9963 -506
rect 10009 -828 10061 -291
rect 10107 -326 10163 -320
rect 10107 -348 10109 -326
rect 10161 -348 10163 -326
rect 10107 -428 10109 -404
rect 10161 -428 10163 -404
rect 10107 -506 10109 -484
rect 10161 -506 10163 -484
rect 10107 -512 10163 -506
rect 10209 -828 10261 -291
rect 10307 -326 10363 -320
rect 10307 -348 10309 -326
rect 10361 -348 10363 -326
rect 10307 -428 10309 -404
rect 10361 -428 10363 -404
rect 10307 -506 10309 -484
rect 10361 -506 10363 -484
rect 10307 -512 10363 -506
rect 10409 -828 10461 -291
rect 10507 -326 10563 -320
rect 10507 -348 10509 -326
rect 10561 -348 10563 -326
rect 10507 -428 10509 -404
rect 10561 -428 10563 -404
rect 10507 -506 10509 -484
rect 10561 -506 10563 -484
rect 10507 -512 10563 -506
rect 10609 -828 10661 -291
rect 10707 -326 10763 -320
rect 10707 -348 10709 -326
rect 10761 -348 10763 -326
rect 10707 -428 10709 -404
rect 10761 -428 10763 -404
rect 10707 -506 10709 -484
rect 10761 -506 10763 -484
rect 10707 -512 10763 -506
rect 10809 -828 10861 -291
rect 10907 -326 10963 -320
rect 10907 -348 10909 -326
rect 10961 -348 10963 -326
rect 10907 -428 10909 -404
rect 10961 -428 10963 -404
rect 10907 -506 10909 -484
rect 10961 -506 10963 -484
rect 10907 -512 10963 -506
rect 11009 -828 11061 -291
rect 11107 -326 11163 -320
rect 11107 -348 11109 -326
rect 11161 -348 11163 -326
rect 11107 -428 11109 -404
rect 11161 -428 11163 -404
rect 11107 -506 11109 -484
rect 11161 -506 11163 -484
rect 11107 -512 11163 -506
rect 11209 -828 11261 -291
rect 11307 -326 11363 -320
rect 11307 -348 11309 -326
rect 11361 -348 11363 -326
rect 11307 -428 11309 -404
rect 11361 -428 11363 -404
rect 11307 -506 11309 -484
rect 11361 -506 11363 -484
rect 11307 -512 11363 -506
rect 11409 -828 11461 -291
rect 11507 -326 11563 -320
rect 11507 -348 11509 -326
rect 11561 -348 11563 -326
rect 11507 -428 11509 -404
rect 11561 -428 11563 -404
rect 11507 -506 11509 -484
rect 11561 -506 11563 -484
rect 11507 -512 11563 -506
rect 11609 -828 11661 -291
rect 11707 -326 11763 -320
rect 11707 -348 11709 -326
rect 11761 -348 11763 -326
rect 11707 -428 11709 -404
rect 11761 -428 11763 -404
rect 11707 -506 11709 -484
rect 11761 -506 11763 -484
rect 11707 -512 11763 -506
rect 11809 -828 11861 -291
rect 11907 -326 11963 -320
rect 11907 -348 11909 -326
rect 11961 -348 11963 -326
rect 11907 -428 11909 -404
rect 11961 -428 11963 -404
rect 11907 -506 11909 -484
rect 11961 -506 11963 -484
rect 11907 -512 11963 -506
rect 12009 -828 12061 -291
rect 12107 -326 12163 -320
rect 12107 -348 12109 -326
rect 12161 -348 12163 -326
rect 12107 -428 12109 -404
rect 12161 -428 12163 -404
rect 12107 -506 12109 -484
rect 12161 -506 12163 -484
rect 12107 -512 12163 -506
rect 12209 -828 12261 -291
rect 12307 -326 12363 -320
rect 12307 -348 12309 -326
rect 12361 -348 12363 -326
rect 12307 -428 12309 -404
rect 12361 -428 12363 -404
rect 12307 -506 12309 -484
rect 12361 -506 12363 -484
rect 12307 -512 12363 -506
rect 12409 -828 12461 -291
rect 12507 -326 12563 -320
rect 12507 -348 12509 -326
rect 12561 -348 12563 -326
rect 12507 -428 12509 -404
rect 12561 -428 12563 -404
rect 12507 -506 12509 -484
rect 12561 -506 12563 -484
rect 12507 -512 12563 -506
rect 12609 -828 12661 -291
rect 12707 -326 12763 -320
rect 12707 -348 12709 -326
rect 12761 -348 12763 -326
rect 12707 -428 12709 -404
rect 12761 -428 12763 -404
rect 14440 -351 15212 -299
rect 15264 -351 15270 -299
rect 15565 -351 15840 -299
rect 14440 -399 14492 -351
rect 14440 -457 14492 -451
rect 14526 -397 14697 -388
rect 14526 -453 14543 -397
rect 14599 -399 14623 -397
rect 14605 -451 14617 -399
rect 14599 -453 14623 -451
rect 14679 -453 14697 -397
rect 14526 -462 14697 -453
rect 14725 -399 14777 -351
rect 14725 -457 14777 -451
rect 14805 -397 15136 -388
rect 14805 -399 14822 -397
rect 14878 -399 14902 -397
rect 14958 -399 14982 -397
rect 15038 -399 15062 -397
rect 15118 -399 15136 -397
rect 14805 -451 14816 -399
rect 14878 -451 14880 -399
rect 15060 -451 15062 -399
rect 15124 -451 15136 -399
rect 14805 -453 14822 -451
rect 14878 -453 14902 -451
rect 14958 -453 14982 -451
rect 15038 -453 15062 -451
rect 15118 -453 15136 -451
rect 14805 -462 15136 -453
rect 15206 -397 15537 -388
rect 15206 -399 15223 -397
rect 15279 -399 15303 -397
rect 15359 -399 15383 -397
rect 15439 -399 15463 -397
rect 15519 -399 15537 -397
rect 15206 -451 15217 -399
rect 15279 -451 15281 -399
rect 15461 -451 15463 -399
rect 15525 -451 15537 -399
rect 15206 -453 15223 -451
rect 15279 -453 15303 -451
rect 15359 -453 15383 -451
rect 15439 -453 15463 -451
rect 15519 -453 15537 -451
rect 15206 -462 15537 -453
rect 15565 -399 15617 -351
rect 15565 -457 15617 -451
rect 15645 -397 15816 -388
rect 15645 -453 15662 -397
rect 15718 -399 15742 -397
rect 15724 -451 15736 -399
rect 15718 -453 15742 -451
rect 15798 -453 15816 -397
rect 15645 -462 15816 -453
rect 12707 -506 12709 -484
rect 12761 -506 12763 -484
rect 12707 -512 12763 -506
rect 14440 -551 15212 -499
rect 15264 -551 15270 -499
rect 15565 -551 15840 -499
rect 14440 -599 14492 -551
rect 14440 -657 14492 -651
rect 14526 -597 14697 -588
rect 14526 -653 14543 -597
rect 14599 -599 14623 -597
rect 14605 -651 14617 -599
rect 14599 -653 14623 -651
rect 14679 -653 14697 -597
rect 14526 -662 14697 -653
rect 14725 -599 14777 -551
rect 14725 -657 14777 -651
rect 14805 -597 15136 -588
rect 14805 -599 14822 -597
rect 14878 -599 14902 -597
rect 14958 -599 14982 -597
rect 15038 -599 15062 -597
rect 15118 -599 15136 -597
rect 14805 -651 14816 -599
rect 14878 -651 14880 -599
rect 15060 -651 15062 -599
rect 15124 -651 15136 -599
rect 14805 -653 14822 -651
rect 14878 -653 14902 -651
rect 14958 -653 14982 -651
rect 15038 -653 15062 -651
rect 15118 -653 15136 -651
rect 14805 -662 15136 -653
rect 15206 -597 15537 -588
rect 15206 -599 15223 -597
rect 15279 -599 15303 -597
rect 15359 -599 15383 -597
rect 15439 -599 15463 -597
rect 15519 -599 15537 -597
rect 15206 -651 15217 -599
rect 15279 -651 15281 -599
rect 15461 -651 15463 -599
rect 15525 -651 15537 -599
rect 15206 -653 15223 -651
rect 15279 -653 15303 -651
rect 15359 -653 15383 -651
rect 15439 -653 15463 -651
rect 15519 -653 15537 -651
rect 15206 -662 15537 -653
rect 15565 -599 15617 -551
rect 15565 -657 15617 -651
rect 15645 -597 15816 -588
rect 15645 -653 15662 -597
rect 15718 -599 15742 -597
rect 15724 -651 15736 -599
rect 15718 -653 15742 -651
rect 15798 -653 15816 -597
rect 15645 -662 15816 -653
rect 14440 -751 15212 -699
rect 15264 -751 15270 -699
rect 15565 -751 15840 -699
rect 14440 -799 14492 -751
rect -18 -880 -9 -828
rect 43 -880 55 -828
rect 107 -880 116 -828
rect 154 -880 163 -828
rect 215 -880 227 -828
rect 279 -880 288 -828
rect 382 -880 391 -828
rect 443 -880 455 -828
rect 507 -880 516 -828
rect 554 -880 563 -828
rect 615 -880 627 -828
rect 679 -880 688 -828
rect 782 -880 791 -828
rect 843 -880 855 -828
rect 907 -880 916 -828
rect 954 -880 963 -828
rect 1015 -880 1027 -828
rect 1079 -880 1088 -828
rect 1182 -880 1191 -828
rect 1243 -880 1255 -828
rect 1307 -880 1316 -828
rect 1354 -880 1363 -828
rect 1415 -880 1427 -828
rect 1479 -880 1488 -828
rect 1582 -880 1591 -828
rect 1643 -880 1655 -828
rect 1707 -880 1716 -828
rect 1754 -880 1763 -828
rect 1815 -880 1827 -828
rect 1879 -880 1888 -828
rect 1982 -880 1991 -828
rect 2043 -880 2055 -828
rect 2107 -880 2116 -828
rect 2154 -880 2163 -828
rect 2215 -880 2227 -828
rect 2279 -880 2288 -828
rect 2382 -880 2391 -828
rect 2443 -880 2455 -828
rect 2507 -880 2516 -828
rect 2554 -880 2563 -828
rect 2615 -880 2627 -828
rect 2679 -880 2688 -828
rect 2782 -880 2791 -828
rect 2843 -880 2855 -828
rect 2907 -880 2916 -828
rect 2954 -880 2963 -828
rect 3015 -880 3027 -828
rect 3079 -880 3088 -828
rect 3182 -880 3191 -828
rect 3243 -880 3255 -828
rect 3307 -880 3316 -828
rect 3354 -880 3363 -828
rect 3415 -880 3427 -828
rect 3479 -880 3488 -828
rect 3582 -880 3591 -828
rect 3643 -880 3655 -828
rect 3707 -880 3716 -828
rect 3754 -880 3763 -828
rect 3815 -880 3827 -828
rect 3879 -880 3888 -828
rect 3982 -880 3991 -828
rect 4043 -880 4055 -828
rect 4107 -880 4116 -828
rect 4154 -880 4163 -828
rect 4215 -880 4227 -828
rect 4279 -880 4288 -828
rect 4382 -880 4391 -828
rect 4443 -880 4455 -828
rect 4507 -880 4516 -828
rect 4554 -880 4563 -828
rect 4615 -880 4627 -828
rect 4679 -880 4688 -828
rect 4782 -880 4791 -828
rect 4843 -880 4855 -828
rect 4907 -880 4916 -828
rect 4954 -880 4963 -828
rect 5015 -880 5027 -828
rect 5079 -880 5088 -828
rect 5182 -880 5191 -828
rect 5243 -880 5255 -828
rect 5307 -880 5316 -828
rect 5354 -880 5363 -828
rect 5415 -880 5427 -828
rect 5479 -880 5488 -828
rect 5582 -880 5591 -828
rect 5643 -880 5655 -828
rect 5707 -880 5716 -828
rect 5754 -880 5763 -828
rect 5815 -880 5827 -828
rect 5879 -880 5888 -828
rect 5982 -880 5991 -828
rect 6043 -880 6055 -828
rect 6107 -880 6116 -828
rect 6154 -880 6163 -828
rect 6215 -880 6227 -828
rect 6279 -880 6288 -828
rect 6382 -880 6391 -828
rect 6443 -880 6455 -828
rect 6507 -880 6516 -828
rect 6554 -880 6563 -828
rect 6615 -880 6627 -828
rect 6679 -880 6688 -828
rect 6782 -880 6791 -828
rect 6843 -880 6855 -828
rect 6907 -880 6916 -828
rect 6954 -880 6963 -828
rect 7015 -880 7027 -828
rect 7079 -880 7088 -828
rect 7182 -880 7191 -828
rect 7243 -880 7255 -828
rect 7307 -880 7316 -828
rect 7354 -880 7363 -828
rect 7415 -880 7427 -828
rect 7479 -880 7488 -828
rect 7582 -880 7591 -828
rect 7643 -880 7655 -828
rect 7707 -880 7716 -828
rect 7754 -880 7763 -828
rect 7815 -880 7827 -828
rect 7879 -880 7888 -828
rect 7982 -880 7991 -828
rect 8043 -880 8055 -828
rect 8107 -880 8116 -828
rect 8154 -880 8163 -828
rect 8215 -880 8227 -828
rect 8279 -880 8288 -828
rect 8382 -880 8391 -828
rect 8443 -880 8455 -828
rect 8507 -880 8516 -828
rect 8554 -880 8563 -828
rect 8615 -880 8627 -828
rect 8679 -880 8688 -828
rect 8782 -880 8791 -828
rect 8843 -880 8855 -828
rect 8907 -880 8916 -828
rect 8954 -880 8963 -828
rect 9015 -880 9027 -828
rect 9079 -880 9088 -828
rect 9182 -880 9191 -828
rect 9243 -880 9255 -828
rect 9307 -880 9316 -828
rect 9354 -880 9363 -828
rect 9415 -880 9427 -828
rect 9479 -880 9488 -828
rect 9582 -880 9591 -828
rect 9643 -880 9655 -828
rect 9707 -880 9716 -828
rect 9754 -880 9763 -828
rect 9815 -880 9827 -828
rect 9879 -880 9888 -828
rect 9982 -880 9991 -828
rect 10043 -880 10055 -828
rect 10107 -880 10116 -828
rect 10154 -880 10163 -828
rect 10215 -880 10227 -828
rect 10279 -880 10288 -828
rect 10382 -880 10391 -828
rect 10443 -880 10455 -828
rect 10507 -880 10516 -828
rect 10554 -880 10563 -828
rect 10615 -880 10627 -828
rect 10679 -880 10688 -828
rect 10782 -880 10791 -828
rect 10843 -880 10855 -828
rect 10907 -880 10916 -828
rect 10954 -880 10963 -828
rect 11015 -880 11027 -828
rect 11079 -880 11088 -828
rect 11182 -880 11191 -828
rect 11243 -880 11255 -828
rect 11307 -880 11316 -828
rect 11354 -880 11363 -828
rect 11415 -880 11427 -828
rect 11479 -880 11488 -828
rect 11582 -880 11591 -828
rect 11643 -880 11655 -828
rect 11707 -880 11716 -828
rect 11754 -880 11763 -828
rect 11815 -880 11827 -828
rect 11879 -880 11888 -828
rect 11982 -880 11991 -828
rect 12043 -880 12055 -828
rect 12107 -880 12116 -828
rect 12154 -880 12163 -828
rect 12215 -880 12227 -828
rect 12279 -880 12288 -828
rect 12382 -880 12391 -828
rect 12443 -880 12455 -828
rect 12507 -880 12516 -828
rect 12554 -880 12563 -828
rect 12615 -880 12627 -828
rect 12679 -880 12688 -828
rect 14440 -857 14492 -851
rect 14526 -797 14697 -788
rect 14526 -853 14543 -797
rect 14599 -799 14623 -797
rect 14605 -851 14617 -799
rect 14599 -853 14623 -851
rect 14679 -853 14697 -797
rect 14526 -862 14697 -853
rect 14725 -799 14777 -751
rect 14725 -857 14777 -851
rect 14805 -797 15136 -788
rect 14805 -799 14822 -797
rect 14878 -799 14902 -797
rect 14958 -799 14982 -797
rect 15038 -799 15062 -797
rect 15118 -799 15136 -797
rect 14805 -851 14816 -799
rect 14878 -851 14880 -799
rect 15060 -851 15062 -799
rect 15124 -851 15136 -799
rect 14805 -853 14822 -851
rect 14878 -853 14902 -851
rect 14958 -853 14982 -851
rect 15038 -853 15062 -851
rect 15118 -853 15136 -851
rect 14805 -862 15136 -853
rect 15206 -797 15537 -788
rect 15206 -799 15223 -797
rect 15279 -799 15303 -797
rect 15359 -799 15383 -797
rect 15439 -799 15463 -797
rect 15519 -799 15537 -797
rect 15206 -851 15217 -799
rect 15279 -851 15281 -799
rect 15461 -851 15463 -799
rect 15525 -851 15537 -799
rect 15206 -853 15223 -851
rect 15279 -853 15303 -851
rect 15359 -853 15383 -851
rect 15439 -853 15463 -851
rect 15519 -853 15537 -851
rect 15206 -862 15537 -853
rect 15565 -799 15617 -751
rect 15565 -857 15617 -851
rect 15645 -797 15816 -788
rect 15645 -853 15662 -797
rect 15718 -799 15742 -797
rect 15724 -851 15736 -799
rect 15718 -853 15742 -851
rect 15798 -853 15816 -797
rect 15645 -862 15816 -853
rect 14440 -951 15212 -899
rect 15264 -951 15270 -899
rect 15565 -951 15840 -899
rect 14440 -999 14492 -951
rect 14440 -1057 14492 -1051
rect 14526 -997 14697 -988
rect 14526 -1053 14543 -997
rect 14599 -999 14623 -997
rect 14605 -1051 14617 -999
rect 14599 -1053 14623 -1051
rect 14679 -1053 14697 -997
rect 14526 -1062 14697 -1053
rect 14725 -999 14777 -951
rect 14725 -1057 14777 -1051
rect 14805 -997 15136 -988
rect 14805 -999 14822 -997
rect 14878 -999 14902 -997
rect 14958 -999 14982 -997
rect 15038 -999 15062 -997
rect 15118 -999 15136 -997
rect 14805 -1051 14816 -999
rect 14878 -1051 14880 -999
rect 15060 -1051 15062 -999
rect 15124 -1051 15136 -999
rect 14805 -1053 14822 -1051
rect 14878 -1053 14902 -1051
rect 14958 -1053 14982 -1051
rect 15038 -1053 15062 -1051
rect 15118 -1053 15136 -1051
rect 14805 -1062 15136 -1053
rect 15206 -997 15537 -988
rect 15206 -999 15223 -997
rect 15279 -999 15303 -997
rect 15359 -999 15383 -997
rect 15439 -999 15463 -997
rect 15519 -999 15537 -997
rect 15206 -1051 15217 -999
rect 15279 -1051 15281 -999
rect 15461 -1051 15463 -999
rect 15525 -1051 15537 -999
rect 15206 -1053 15223 -1051
rect 15279 -1053 15303 -1051
rect 15359 -1053 15383 -1051
rect 15439 -1053 15463 -1051
rect 15519 -1053 15537 -1051
rect 15206 -1062 15537 -1053
rect 15565 -999 15617 -951
rect 15565 -1057 15617 -1051
rect 15645 -997 15816 -988
rect 15645 -1053 15662 -997
rect 15718 -999 15742 -997
rect 15724 -1051 15736 -999
rect 15718 -1053 15742 -1051
rect 15798 -1053 15816 -997
rect 15645 -1062 15816 -1053
rect 14440 -1151 15212 -1099
rect 15264 -1151 15270 -1099
rect 15565 -1151 15840 -1099
rect 14440 -1199 14492 -1151
rect 14440 -1257 14492 -1251
rect 14526 -1197 14697 -1188
rect 14526 -1253 14543 -1197
rect 14599 -1199 14623 -1197
rect 14605 -1251 14617 -1199
rect 14599 -1253 14623 -1251
rect 14679 -1253 14697 -1197
rect 14526 -1262 14697 -1253
rect 14725 -1199 14777 -1151
rect 14725 -1257 14777 -1251
rect 14805 -1197 15136 -1188
rect 14805 -1199 14822 -1197
rect 14878 -1199 14902 -1197
rect 14958 -1199 14982 -1197
rect 15038 -1199 15062 -1197
rect 15118 -1199 15136 -1197
rect 14805 -1251 14816 -1199
rect 14878 -1251 14880 -1199
rect 15060 -1251 15062 -1199
rect 15124 -1251 15136 -1199
rect 14805 -1253 14822 -1251
rect 14878 -1253 14902 -1251
rect 14958 -1253 14982 -1251
rect 15038 -1253 15062 -1251
rect 15118 -1253 15136 -1251
rect 14805 -1262 15136 -1253
rect 15206 -1197 15537 -1188
rect 15206 -1199 15223 -1197
rect 15279 -1199 15303 -1197
rect 15359 -1199 15383 -1197
rect 15439 -1199 15463 -1197
rect 15519 -1199 15537 -1197
rect 15206 -1251 15217 -1199
rect 15279 -1251 15281 -1199
rect 15461 -1251 15463 -1199
rect 15525 -1251 15537 -1199
rect 15206 -1253 15223 -1251
rect 15279 -1253 15303 -1251
rect 15359 -1253 15383 -1251
rect 15439 -1253 15463 -1251
rect 15519 -1253 15537 -1251
rect 15206 -1262 15537 -1253
rect 15565 -1199 15617 -1151
rect 15565 -1257 15617 -1251
rect 15645 -1197 15816 -1188
rect 15645 -1253 15662 -1197
rect 15718 -1199 15742 -1197
rect 15724 -1251 15736 -1199
rect 15718 -1253 15742 -1251
rect 15798 -1253 15816 -1197
rect 15645 -1262 15816 -1253
rect 14440 -1351 15212 -1299
rect 15264 -1351 15270 -1299
rect 15565 -1351 15840 -1299
rect 14440 -1399 14492 -1351
rect 14440 -1457 14492 -1451
rect 14526 -1397 14697 -1388
rect 14526 -1453 14543 -1397
rect 14599 -1399 14623 -1397
rect 14605 -1451 14617 -1399
rect 14599 -1453 14623 -1451
rect 14679 -1453 14697 -1397
rect 14526 -1462 14697 -1453
rect 14725 -1399 14777 -1351
rect 14725 -1457 14777 -1451
rect 14805 -1397 15136 -1388
rect 14805 -1399 14822 -1397
rect 14878 -1399 14902 -1397
rect 14958 -1399 14982 -1397
rect 15038 -1399 15062 -1397
rect 15118 -1399 15136 -1397
rect 14805 -1451 14816 -1399
rect 14878 -1451 14880 -1399
rect 15060 -1451 15062 -1399
rect 15124 -1451 15136 -1399
rect 14805 -1453 14822 -1451
rect 14878 -1453 14902 -1451
rect 14958 -1453 14982 -1451
rect 15038 -1453 15062 -1451
rect 15118 -1453 15136 -1451
rect 14805 -1462 15136 -1453
rect 15206 -1397 15537 -1388
rect 15206 -1399 15223 -1397
rect 15279 -1399 15303 -1397
rect 15359 -1399 15383 -1397
rect 15439 -1399 15463 -1397
rect 15519 -1399 15537 -1397
rect 15206 -1451 15217 -1399
rect 15279 -1451 15281 -1399
rect 15461 -1451 15463 -1399
rect 15525 -1451 15537 -1399
rect 15206 -1453 15223 -1451
rect 15279 -1453 15303 -1451
rect 15359 -1453 15383 -1451
rect 15439 -1453 15463 -1451
rect 15519 -1453 15537 -1451
rect 15206 -1462 15537 -1453
rect 15565 -1399 15617 -1351
rect 15565 -1457 15617 -1451
rect 15645 -1397 15816 -1388
rect 15645 -1453 15662 -1397
rect 15718 -1399 15742 -1397
rect 15724 -1451 15736 -1399
rect 15718 -1453 15742 -1451
rect 15798 -1453 15816 -1397
rect 15645 -1462 15816 -1453
rect 14440 -1551 15212 -1499
rect 15264 -1551 15270 -1499
rect 15565 -1551 15840 -1499
rect 14440 -1599 14492 -1551
rect 14440 -1657 14492 -1651
rect 14526 -1597 14697 -1588
rect 14526 -1653 14543 -1597
rect 14599 -1599 14623 -1597
rect 14605 -1651 14617 -1599
rect 14599 -1653 14623 -1651
rect 14679 -1653 14697 -1597
rect 14526 -1662 14697 -1653
rect 14725 -1599 14777 -1551
rect 14725 -1657 14777 -1651
rect 14805 -1597 15136 -1588
rect 14805 -1599 14822 -1597
rect 14878 -1599 14902 -1597
rect 14958 -1599 14982 -1597
rect 15038 -1599 15062 -1597
rect 15118 -1599 15136 -1597
rect 14805 -1651 14816 -1599
rect 14878 -1651 14880 -1599
rect 15060 -1651 15062 -1599
rect 15124 -1651 15136 -1599
rect 14805 -1653 14822 -1651
rect 14878 -1653 14902 -1651
rect 14958 -1653 14982 -1651
rect 15038 -1653 15062 -1651
rect 15118 -1653 15136 -1651
rect 14805 -1662 15136 -1653
rect 15206 -1597 15537 -1588
rect 15206 -1599 15223 -1597
rect 15279 -1599 15303 -1597
rect 15359 -1599 15383 -1597
rect 15439 -1599 15463 -1597
rect 15519 -1599 15537 -1597
rect 15206 -1651 15217 -1599
rect 15279 -1651 15281 -1599
rect 15461 -1651 15463 -1599
rect 15525 -1651 15537 -1599
rect 15206 -1653 15223 -1651
rect 15279 -1653 15303 -1651
rect 15359 -1653 15383 -1651
rect 15439 -1653 15463 -1651
rect 15519 -1653 15537 -1651
rect 15206 -1662 15537 -1653
rect 15565 -1599 15617 -1551
rect 15565 -1657 15617 -1651
rect 15645 -1597 15816 -1588
rect 15645 -1653 15662 -1597
rect 15718 -1599 15742 -1597
rect 15724 -1651 15736 -1599
rect 15718 -1653 15742 -1651
rect 15798 -1653 15816 -1597
rect 15645 -1662 15816 -1653
rect 14440 -1751 15212 -1699
rect 15264 -1751 15270 -1699
rect 15565 -1751 15840 -1699
rect 14440 -1799 14492 -1751
rect 14440 -1857 14492 -1851
rect 14526 -1797 14697 -1788
rect 14526 -1853 14543 -1797
rect 14599 -1799 14623 -1797
rect 14605 -1851 14617 -1799
rect 14599 -1853 14623 -1851
rect 14679 -1853 14697 -1797
rect 14526 -1862 14697 -1853
rect 14725 -1799 14777 -1751
rect 14725 -1857 14777 -1851
rect 14805 -1797 15136 -1788
rect 14805 -1799 14822 -1797
rect 14878 -1799 14902 -1797
rect 14958 -1799 14982 -1797
rect 15038 -1799 15062 -1797
rect 15118 -1799 15136 -1797
rect 14805 -1851 14816 -1799
rect 14878 -1851 14880 -1799
rect 15060 -1851 15062 -1799
rect 15124 -1851 15136 -1799
rect 14805 -1853 14822 -1851
rect 14878 -1853 14902 -1851
rect 14958 -1853 14982 -1851
rect 15038 -1853 15062 -1851
rect 15118 -1853 15136 -1851
rect 14805 -1862 15136 -1853
rect 15206 -1797 15537 -1788
rect 15206 -1799 15223 -1797
rect 15279 -1799 15303 -1797
rect 15359 -1799 15383 -1797
rect 15439 -1799 15463 -1797
rect 15519 -1799 15537 -1797
rect 15206 -1851 15217 -1799
rect 15279 -1851 15281 -1799
rect 15461 -1851 15463 -1799
rect 15525 -1851 15537 -1799
rect 15206 -1853 15223 -1851
rect 15279 -1853 15303 -1851
rect 15359 -1853 15383 -1851
rect 15439 -1853 15463 -1851
rect 15519 -1853 15537 -1851
rect 15206 -1862 15537 -1853
rect 15565 -1799 15617 -1751
rect 15565 -1857 15617 -1851
rect 15645 -1797 15816 -1788
rect 15645 -1853 15662 -1797
rect 15718 -1799 15742 -1797
rect 15724 -1851 15736 -1799
rect 15718 -1853 15742 -1851
rect 15798 -1853 15816 -1797
rect 15645 -1862 15816 -1853
rect 14440 -1951 15212 -1899
rect 15264 -1951 15270 -1899
rect 15565 -1951 15840 -1899
rect 14440 -1999 14492 -1951
rect 14440 -2057 14492 -2051
rect 14526 -1997 14697 -1988
rect 14526 -2053 14543 -1997
rect 14599 -1999 14623 -1997
rect 14605 -2051 14617 -1999
rect 14599 -2053 14623 -2051
rect 14679 -2053 14697 -1997
rect 14526 -2062 14697 -2053
rect 14725 -1999 14777 -1951
rect 14725 -2057 14777 -2051
rect 14805 -1997 15136 -1988
rect 14805 -1999 14822 -1997
rect 14878 -1999 14902 -1997
rect 14958 -1999 14982 -1997
rect 15038 -1999 15062 -1997
rect 15118 -1999 15136 -1997
rect 14805 -2051 14816 -1999
rect 14878 -2051 14880 -1999
rect 15060 -2051 15062 -1999
rect 15124 -2051 15136 -1999
rect 14805 -2053 14822 -2051
rect 14878 -2053 14902 -2051
rect 14958 -2053 14982 -2051
rect 15038 -2053 15062 -2051
rect 15118 -2053 15136 -2051
rect 14805 -2062 15136 -2053
rect 15206 -1997 15537 -1988
rect 15206 -1999 15223 -1997
rect 15279 -1999 15303 -1997
rect 15359 -1999 15383 -1997
rect 15439 -1999 15463 -1997
rect 15519 -1999 15537 -1997
rect 15206 -2051 15217 -1999
rect 15279 -2051 15281 -1999
rect 15461 -2051 15463 -1999
rect 15525 -2051 15537 -1999
rect 15206 -2053 15223 -2051
rect 15279 -2053 15303 -2051
rect 15359 -2053 15383 -2051
rect 15439 -2053 15463 -2051
rect 15519 -2053 15537 -2051
rect 15206 -2062 15537 -2053
rect 15565 -1999 15617 -1951
rect 15565 -2057 15617 -2051
rect 15645 -1997 15816 -1988
rect 15645 -2053 15662 -1997
rect 15718 -1999 15742 -1997
rect 15724 -2051 15736 -1999
rect 15718 -2053 15742 -2051
rect 15798 -2053 15816 -1997
rect 15645 -2062 15816 -2053
<< via2 >>
rect 7 4903 63 4905
rect 7 4851 9 4903
rect 9 4851 61 4903
rect 61 4851 63 4903
rect 7 4849 63 4851
rect 207 4919 263 4921
rect 207 4867 209 4919
rect 209 4867 261 4919
rect 261 4867 263 4919
rect 207 4865 263 4867
rect 407 4903 463 4905
rect 407 4851 409 4903
rect 409 4851 461 4903
rect 461 4851 463 4903
rect 407 4849 463 4851
rect 607 4919 663 4921
rect 607 4867 609 4919
rect 609 4867 661 4919
rect 661 4867 663 4919
rect 607 4865 663 4867
rect 807 4903 863 4905
rect 807 4851 809 4903
rect 809 4851 861 4903
rect 861 4851 863 4903
rect 807 4849 863 4851
rect 1007 4919 1063 4921
rect 1007 4867 1009 4919
rect 1009 4867 1061 4919
rect 1061 4867 1063 4919
rect 1007 4865 1063 4867
rect 1207 4903 1263 4905
rect 1207 4851 1209 4903
rect 1209 4851 1261 4903
rect 1261 4851 1263 4903
rect 1207 4849 1263 4851
rect 1407 4919 1463 4921
rect 1407 4867 1409 4919
rect 1409 4867 1461 4919
rect 1461 4867 1463 4919
rect 1407 4865 1463 4867
rect 1607 4903 1663 4905
rect 1607 4851 1609 4903
rect 1609 4851 1661 4903
rect 1661 4851 1663 4903
rect 1607 4849 1663 4851
rect 1807 4919 1863 4921
rect 1807 4867 1809 4919
rect 1809 4867 1861 4919
rect 1861 4867 1863 4919
rect 1807 4865 1863 4867
rect 2007 4903 2063 4905
rect 2007 4851 2009 4903
rect 2009 4851 2061 4903
rect 2061 4851 2063 4903
rect 2007 4849 2063 4851
rect 2207 4919 2263 4921
rect 2207 4867 2209 4919
rect 2209 4867 2261 4919
rect 2261 4867 2263 4919
rect 2207 4865 2263 4867
rect 2407 4903 2463 4905
rect 2407 4851 2409 4903
rect 2409 4851 2461 4903
rect 2461 4851 2463 4903
rect 2407 4849 2463 4851
rect 2607 4919 2663 4921
rect 2607 4867 2609 4919
rect 2609 4867 2661 4919
rect 2661 4867 2663 4919
rect 2607 4865 2663 4867
rect 2807 4903 2863 4905
rect 2807 4851 2809 4903
rect 2809 4851 2861 4903
rect 2861 4851 2863 4903
rect 2807 4849 2863 4851
rect 3007 4919 3063 4921
rect 3007 4867 3009 4919
rect 3009 4867 3061 4919
rect 3061 4867 3063 4919
rect 3007 4865 3063 4867
rect 3207 4903 3263 4905
rect 3207 4851 3209 4903
rect 3209 4851 3261 4903
rect 3261 4851 3263 4903
rect 3207 4849 3263 4851
rect 3407 4919 3463 4921
rect 3407 4867 3409 4919
rect 3409 4867 3461 4919
rect 3461 4867 3463 4919
rect 3407 4865 3463 4867
rect 3607 4903 3663 4905
rect 3607 4851 3609 4903
rect 3609 4851 3661 4903
rect 3661 4851 3663 4903
rect 3607 4849 3663 4851
rect 3807 4919 3863 4921
rect 3807 4867 3809 4919
rect 3809 4867 3861 4919
rect 3861 4867 3863 4919
rect 3807 4865 3863 4867
rect 4007 4903 4063 4905
rect 4007 4851 4009 4903
rect 4009 4851 4061 4903
rect 4061 4851 4063 4903
rect 4007 4849 4063 4851
rect 4207 4919 4263 4921
rect 4207 4867 4209 4919
rect 4209 4867 4261 4919
rect 4261 4867 4263 4919
rect 4207 4865 4263 4867
rect 4407 4903 4463 4905
rect 4407 4851 4409 4903
rect 4409 4851 4461 4903
rect 4461 4851 4463 4903
rect 4407 4849 4463 4851
rect 4607 4919 4663 4921
rect 4607 4867 4609 4919
rect 4609 4867 4661 4919
rect 4661 4867 4663 4919
rect 4607 4865 4663 4867
rect 4807 4903 4863 4905
rect 4807 4851 4809 4903
rect 4809 4851 4861 4903
rect 4861 4851 4863 4903
rect 4807 4849 4863 4851
rect 5007 4919 5063 4921
rect 5007 4867 5009 4919
rect 5009 4867 5061 4919
rect 5061 4867 5063 4919
rect 5007 4865 5063 4867
rect 5207 4903 5263 4905
rect 5207 4851 5209 4903
rect 5209 4851 5261 4903
rect 5261 4851 5263 4903
rect 5207 4849 5263 4851
rect 5407 4919 5463 4921
rect 5407 4867 5409 4919
rect 5409 4867 5461 4919
rect 5461 4867 5463 4919
rect 5407 4865 5463 4867
rect 5607 4903 5663 4905
rect 5607 4851 5609 4903
rect 5609 4851 5661 4903
rect 5661 4851 5663 4903
rect 5607 4849 5663 4851
rect 5807 4919 5863 4921
rect 5807 4867 5809 4919
rect 5809 4867 5861 4919
rect 5861 4867 5863 4919
rect 5807 4865 5863 4867
rect 6007 4903 6063 4905
rect 6007 4851 6009 4903
rect 6009 4851 6061 4903
rect 6061 4851 6063 4903
rect 6007 4849 6063 4851
rect 6207 4919 6263 4921
rect 6207 4867 6209 4919
rect 6209 4867 6261 4919
rect 6261 4867 6263 4919
rect 6207 4865 6263 4867
rect 6407 4903 6463 4905
rect 6407 4851 6409 4903
rect 6409 4851 6461 4903
rect 6461 4851 6463 4903
rect 6407 4849 6463 4851
rect 6607 4919 6663 4921
rect 6607 4867 6609 4919
rect 6609 4867 6661 4919
rect 6661 4867 6663 4919
rect 6607 4865 6663 4867
rect 6807 4903 6863 4905
rect 6807 4851 6809 4903
rect 6809 4851 6861 4903
rect 6861 4851 6863 4903
rect 6807 4849 6863 4851
rect 7007 4919 7063 4921
rect 7007 4867 7009 4919
rect 7009 4867 7061 4919
rect 7061 4867 7063 4919
rect 7007 4865 7063 4867
rect 7207 4903 7263 4905
rect 7207 4851 7209 4903
rect 7209 4851 7261 4903
rect 7261 4851 7263 4903
rect 7207 4849 7263 4851
rect 7407 4919 7463 4921
rect 7407 4867 7409 4919
rect 7409 4867 7461 4919
rect 7461 4867 7463 4919
rect 7407 4865 7463 4867
rect 7607 4903 7663 4905
rect 7607 4851 7609 4903
rect 7609 4851 7661 4903
rect 7661 4851 7663 4903
rect 7607 4849 7663 4851
rect 7807 4919 7863 4921
rect 7807 4867 7809 4919
rect 7809 4867 7861 4919
rect 7861 4867 7863 4919
rect 7807 4865 7863 4867
rect 8007 4903 8063 4905
rect 8007 4851 8009 4903
rect 8009 4851 8061 4903
rect 8061 4851 8063 4903
rect 8007 4849 8063 4851
rect 8207 4919 8263 4921
rect 8207 4867 8209 4919
rect 8209 4867 8261 4919
rect 8261 4867 8263 4919
rect 8207 4865 8263 4867
rect 8407 4903 8463 4905
rect 8407 4851 8409 4903
rect 8409 4851 8461 4903
rect 8461 4851 8463 4903
rect 8407 4849 8463 4851
rect 8607 4919 8663 4921
rect 8607 4867 8609 4919
rect 8609 4867 8661 4919
rect 8661 4867 8663 4919
rect 8607 4865 8663 4867
rect 8807 4903 8863 4905
rect 8807 4851 8809 4903
rect 8809 4851 8861 4903
rect 8861 4851 8863 4903
rect 8807 4849 8863 4851
rect 9007 4919 9063 4921
rect 9007 4867 9009 4919
rect 9009 4867 9061 4919
rect 9061 4867 9063 4919
rect 9007 4865 9063 4867
rect 9207 4903 9263 4905
rect 9207 4851 9209 4903
rect 9209 4851 9261 4903
rect 9261 4851 9263 4903
rect 9207 4849 9263 4851
rect 9407 4919 9463 4921
rect 9407 4867 9409 4919
rect 9409 4867 9461 4919
rect 9461 4867 9463 4919
rect 9407 4865 9463 4867
rect 9607 4903 9663 4905
rect 9607 4851 9609 4903
rect 9609 4851 9661 4903
rect 9661 4851 9663 4903
rect 9607 4849 9663 4851
rect 9807 4919 9863 4921
rect 9807 4867 9809 4919
rect 9809 4867 9861 4919
rect 9861 4867 9863 4919
rect 9807 4865 9863 4867
rect 10007 4903 10063 4905
rect 10007 4851 10009 4903
rect 10009 4851 10061 4903
rect 10061 4851 10063 4903
rect 10007 4849 10063 4851
rect 10207 4919 10263 4921
rect 10207 4867 10209 4919
rect 10209 4867 10261 4919
rect 10261 4867 10263 4919
rect 10207 4865 10263 4867
rect 10407 4903 10463 4905
rect 10407 4851 10409 4903
rect 10409 4851 10461 4903
rect 10461 4851 10463 4903
rect 10407 4849 10463 4851
rect 10607 4919 10663 4921
rect 10607 4867 10609 4919
rect 10609 4867 10661 4919
rect 10661 4867 10663 4919
rect 10607 4865 10663 4867
rect 10807 4903 10863 4905
rect 10807 4851 10809 4903
rect 10809 4851 10861 4903
rect 10861 4851 10863 4903
rect 10807 4849 10863 4851
rect 11007 4919 11063 4921
rect 11007 4867 11009 4919
rect 11009 4867 11061 4919
rect 11061 4867 11063 4919
rect 11007 4865 11063 4867
rect 11207 4903 11263 4905
rect 11207 4851 11209 4903
rect 11209 4851 11261 4903
rect 11261 4851 11263 4903
rect 11207 4849 11263 4851
rect 11407 4919 11463 4921
rect 11407 4867 11409 4919
rect 11409 4867 11461 4919
rect 11461 4867 11463 4919
rect 11407 4865 11463 4867
rect 11607 4903 11663 4905
rect 11607 4851 11609 4903
rect 11609 4851 11661 4903
rect 11661 4851 11663 4903
rect 11607 4849 11663 4851
rect 11807 4919 11863 4921
rect 11807 4867 11809 4919
rect 11809 4867 11861 4919
rect 11861 4867 11863 4919
rect 11807 4865 11863 4867
rect 12007 4903 12063 4905
rect 12007 4851 12009 4903
rect 12009 4851 12061 4903
rect 12061 4851 12063 4903
rect 12007 4849 12063 4851
rect 12207 4919 12263 4921
rect 12207 4867 12209 4919
rect 12209 4867 12261 4919
rect 12261 4867 12263 4919
rect 12207 4865 12263 4867
rect 12407 4903 12463 4905
rect 12407 4851 12409 4903
rect 12409 4851 12461 4903
rect 12461 4851 12463 4903
rect 12407 4849 12463 4851
rect 12607 4919 12663 4921
rect 12607 4867 12609 4919
rect 12609 4867 12661 4919
rect 12661 4867 12663 4919
rect 12607 4865 12663 4867
rect 7 3693 63 3695
rect 7 3641 9 3693
rect 9 3641 61 3693
rect 61 3641 63 3693
rect 7 3639 63 3641
rect 207 3709 263 3711
rect 207 3657 209 3709
rect 209 3657 261 3709
rect 261 3657 263 3709
rect 207 3655 263 3657
rect 407 3693 463 3695
rect 407 3641 409 3693
rect 409 3641 461 3693
rect 461 3641 463 3693
rect 407 3639 463 3641
rect 607 3709 663 3711
rect 607 3657 609 3709
rect 609 3657 661 3709
rect 661 3657 663 3709
rect 607 3655 663 3657
rect 807 3693 863 3695
rect 807 3641 809 3693
rect 809 3641 861 3693
rect 861 3641 863 3693
rect 807 3639 863 3641
rect 1007 3709 1063 3711
rect 1007 3657 1009 3709
rect 1009 3657 1061 3709
rect 1061 3657 1063 3709
rect 1007 3655 1063 3657
rect 1207 3693 1263 3695
rect 1207 3641 1209 3693
rect 1209 3641 1261 3693
rect 1261 3641 1263 3693
rect 1207 3639 1263 3641
rect 1407 3709 1463 3711
rect 1407 3657 1409 3709
rect 1409 3657 1461 3709
rect 1461 3657 1463 3709
rect 1407 3655 1463 3657
rect 1607 3693 1663 3695
rect 1607 3641 1609 3693
rect 1609 3641 1661 3693
rect 1661 3641 1663 3693
rect 1607 3639 1663 3641
rect 1807 3709 1863 3711
rect 1807 3657 1809 3709
rect 1809 3657 1861 3709
rect 1861 3657 1863 3709
rect 1807 3655 1863 3657
rect 2007 3693 2063 3695
rect 2007 3641 2009 3693
rect 2009 3641 2061 3693
rect 2061 3641 2063 3693
rect 2007 3639 2063 3641
rect 2207 3709 2263 3711
rect 2207 3657 2209 3709
rect 2209 3657 2261 3709
rect 2261 3657 2263 3709
rect 2207 3655 2263 3657
rect 2407 3693 2463 3695
rect 2407 3641 2409 3693
rect 2409 3641 2461 3693
rect 2461 3641 2463 3693
rect 2407 3639 2463 3641
rect 2607 3709 2663 3711
rect 2607 3657 2609 3709
rect 2609 3657 2661 3709
rect 2661 3657 2663 3709
rect 2607 3655 2663 3657
rect 2807 3693 2863 3695
rect 2807 3641 2809 3693
rect 2809 3641 2861 3693
rect 2861 3641 2863 3693
rect 2807 3639 2863 3641
rect 3007 3709 3063 3711
rect 3007 3657 3009 3709
rect 3009 3657 3061 3709
rect 3061 3657 3063 3709
rect 3007 3655 3063 3657
rect 3207 3693 3263 3695
rect 3207 3641 3209 3693
rect 3209 3641 3261 3693
rect 3261 3641 3263 3693
rect 3207 3639 3263 3641
rect 3407 3709 3463 3711
rect 3407 3657 3409 3709
rect 3409 3657 3461 3709
rect 3461 3657 3463 3709
rect 3407 3655 3463 3657
rect 3607 3693 3663 3695
rect 3607 3641 3609 3693
rect 3609 3641 3661 3693
rect 3661 3641 3663 3693
rect 3607 3639 3663 3641
rect 3807 3709 3863 3711
rect 3807 3657 3809 3709
rect 3809 3657 3861 3709
rect 3861 3657 3863 3709
rect 3807 3655 3863 3657
rect 4007 3693 4063 3695
rect 4007 3641 4009 3693
rect 4009 3641 4061 3693
rect 4061 3641 4063 3693
rect 4007 3639 4063 3641
rect 4207 3709 4263 3711
rect 4207 3657 4209 3709
rect 4209 3657 4261 3709
rect 4261 3657 4263 3709
rect 4207 3655 4263 3657
rect 4407 3693 4463 3695
rect 4407 3641 4409 3693
rect 4409 3641 4461 3693
rect 4461 3641 4463 3693
rect 4407 3639 4463 3641
rect 4607 3709 4663 3711
rect 4607 3657 4609 3709
rect 4609 3657 4661 3709
rect 4661 3657 4663 3709
rect 4607 3655 4663 3657
rect 4807 3693 4863 3695
rect 4807 3641 4809 3693
rect 4809 3641 4861 3693
rect 4861 3641 4863 3693
rect 4807 3639 4863 3641
rect 5007 3709 5063 3711
rect 5007 3657 5009 3709
rect 5009 3657 5061 3709
rect 5061 3657 5063 3709
rect 5007 3655 5063 3657
rect 5207 3693 5263 3695
rect 5207 3641 5209 3693
rect 5209 3641 5261 3693
rect 5261 3641 5263 3693
rect 5207 3639 5263 3641
rect 5407 3709 5463 3711
rect 5407 3657 5409 3709
rect 5409 3657 5461 3709
rect 5461 3657 5463 3709
rect 5407 3655 5463 3657
rect 5607 3693 5663 3695
rect 5607 3641 5609 3693
rect 5609 3641 5661 3693
rect 5661 3641 5663 3693
rect 5607 3639 5663 3641
rect 5807 3709 5863 3711
rect 5807 3657 5809 3709
rect 5809 3657 5861 3709
rect 5861 3657 5863 3709
rect 5807 3655 5863 3657
rect 6007 3693 6063 3695
rect 6007 3641 6009 3693
rect 6009 3641 6061 3693
rect 6061 3641 6063 3693
rect 6007 3639 6063 3641
rect 6207 3709 6263 3711
rect 6207 3657 6209 3709
rect 6209 3657 6261 3709
rect 6261 3657 6263 3709
rect 6207 3655 6263 3657
rect 6407 3693 6463 3695
rect 6407 3641 6409 3693
rect 6409 3641 6461 3693
rect 6461 3641 6463 3693
rect 6407 3639 6463 3641
rect 6607 3709 6663 3711
rect 6607 3657 6609 3709
rect 6609 3657 6661 3709
rect 6661 3657 6663 3709
rect 6607 3655 6663 3657
rect 6807 3693 6863 3695
rect 6807 3641 6809 3693
rect 6809 3641 6861 3693
rect 6861 3641 6863 3693
rect 6807 3639 6863 3641
rect 7007 3709 7063 3711
rect 7007 3657 7009 3709
rect 7009 3657 7061 3709
rect 7061 3657 7063 3709
rect 7007 3655 7063 3657
rect 7207 3693 7263 3695
rect 7207 3641 7209 3693
rect 7209 3641 7261 3693
rect 7261 3641 7263 3693
rect 7207 3639 7263 3641
rect 7407 3709 7463 3711
rect 7407 3657 7409 3709
rect 7409 3657 7461 3709
rect 7461 3657 7463 3709
rect 7407 3655 7463 3657
rect 7607 3693 7663 3695
rect 7607 3641 7609 3693
rect 7609 3641 7661 3693
rect 7661 3641 7663 3693
rect 7607 3639 7663 3641
rect 7807 3709 7863 3711
rect 7807 3657 7809 3709
rect 7809 3657 7861 3709
rect 7861 3657 7863 3709
rect 7807 3655 7863 3657
rect 8007 3693 8063 3695
rect 8007 3641 8009 3693
rect 8009 3641 8061 3693
rect 8061 3641 8063 3693
rect 8007 3639 8063 3641
rect 8207 3709 8263 3711
rect 8207 3657 8209 3709
rect 8209 3657 8261 3709
rect 8261 3657 8263 3709
rect 8207 3655 8263 3657
rect 8407 3693 8463 3695
rect 8407 3641 8409 3693
rect 8409 3641 8461 3693
rect 8461 3641 8463 3693
rect 8407 3639 8463 3641
rect 8607 3709 8663 3711
rect 8607 3657 8609 3709
rect 8609 3657 8661 3709
rect 8661 3657 8663 3709
rect 8607 3655 8663 3657
rect 8807 3693 8863 3695
rect 8807 3641 8809 3693
rect 8809 3641 8861 3693
rect 8861 3641 8863 3693
rect 8807 3639 8863 3641
rect 9007 3709 9063 3711
rect 9007 3657 9009 3709
rect 9009 3657 9061 3709
rect 9061 3657 9063 3709
rect 9007 3655 9063 3657
rect 9207 3693 9263 3695
rect 9207 3641 9209 3693
rect 9209 3641 9261 3693
rect 9261 3641 9263 3693
rect 9207 3639 9263 3641
rect 9407 3709 9463 3711
rect 9407 3657 9409 3709
rect 9409 3657 9461 3709
rect 9461 3657 9463 3709
rect 9407 3655 9463 3657
rect 9607 3693 9663 3695
rect 9607 3641 9609 3693
rect 9609 3641 9661 3693
rect 9661 3641 9663 3693
rect 9607 3639 9663 3641
rect 9807 3709 9863 3711
rect 9807 3657 9809 3709
rect 9809 3657 9861 3709
rect 9861 3657 9863 3709
rect 9807 3655 9863 3657
rect 10007 3693 10063 3695
rect 10007 3641 10009 3693
rect 10009 3641 10061 3693
rect 10061 3641 10063 3693
rect 10007 3639 10063 3641
rect 10207 3709 10263 3711
rect 10207 3657 10209 3709
rect 10209 3657 10261 3709
rect 10261 3657 10263 3709
rect 10207 3655 10263 3657
rect 10407 3693 10463 3695
rect 10407 3641 10409 3693
rect 10409 3641 10461 3693
rect 10461 3641 10463 3693
rect 10407 3639 10463 3641
rect 10607 3709 10663 3711
rect 10607 3657 10609 3709
rect 10609 3657 10661 3709
rect 10661 3657 10663 3709
rect 10607 3655 10663 3657
rect 10807 3693 10863 3695
rect 10807 3641 10809 3693
rect 10809 3641 10861 3693
rect 10861 3641 10863 3693
rect 10807 3639 10863 3641
rect 11007 3709 11063 3711
rect 11007 3657 11009 3709
rect 11009 3657 11061 3709
rect 11061 3657 11063 3709
rect 11007 3655 11063 3657
rect 11207 3693 11263 3695
rect 11207 3641 11209 3693
rect 11209 3641 11261 3693
rect 11261 3641 11263 3693
rect 11207 3639 11263 3641
rect 11407 3709 11463 3711
rect 11407 3657 11409 3709
rect 11409 3657 11461 3709
rect 11461 3657 11463 3709
rect 11407 3655 11463 3657
rect 11607 3693 11663 3695
rect 11607 3641 11609 3693
rect 11609 3641 11661 3693
rect 11661 3641 11663 3693
rect 11607 3639 11663 3641
rect 11807 3709 11863 3711
rect 11807 3657 11809 3709
rect 11809 3657 11861 3709
rect 11861 3657 11863 3709
rect 11807 3655 11863 3657
rect 12007 3693 12063 3695
rect 12007 3641 12009 3693
rect 12009 3641 12061 3693
rect 12061 3641 12063 3693
rect 12007 3639 12063 3641
rect 12207 3709 12263 3711
rect 12207 3657 12209 3709
rect 12209 3657 12261 3709
rect 12261 3657 12263 3709
rect 12207 3655 12263 3657
rect 12407 3693 12463 3695
rect 12407 3641 12409 3693
rect 12409 3641 12461 3693
rect 12461 3641 12463 3693
rect 12407 3639 12463 3641
rect 12607 3709 12663 3711
rect 12607 3657 12609 3709
rect 12609 3657 12661 3709
rect 12661 3657 12663 3709
rect 12607 3655 12663 3657
rect 7 2483 63 2485
rect 7 2431 9 2483
rect 9 2431 61 2483
rect 61 2431 63 2483
rect 7 2429 63 2431
rect 207 2499 263 2501
rect 207 2447 209 2499
rect 209 2447 261 2499
rect 261 2447 263 2499
rect 207 2445 263 2447
rect 407 2483 463 2485
rect 407 2431 409 2483
rect 409 2431 461 2483
rect 461 2431 463 2483
rect 407 2429 463 2431
rect 607 2499 663 2501
rect 607 2447 609 2499
rect 609 2447 661 2499
rect 661 2447 663 2499
rect 607 2445 663 2447
rect 807 2483 863 2485
rect 807 2431 809 2483
rect 809 2431 861 2483
rect 861 2431 863 2483
rect 807 2429 863 2431
rect 1007 2499 1063 2501
rect 1007 2447 1009 2499
rect 1009 2447 1061 2499
rect 1061 2447 1063 2499
rect 1007 2445 1063 2447
rect 1207 2483 1263 2485
rect 1207 2431 1209 2483
rect 1209 2431 1261 2483
rect 1261 2431 1263 2483
rect 1207 2429 1263 2431
rect 1407 2499 1463 2501
rect 1407 2447 1409 2499
rect 1409 2447 1461 2499
rect 1461 2447 1463 2499
rect 1407 2445 1463 2447
rect 1607 2483 1663 2485
rect 1607 2431 1609 2483
rect 1609 2431 1661 2483
rect 1661 2431 1663 2483
rect 1607 2429 1663 2431
rect 1807 2499 1863 2501
rect 1807 2447 1809 2499
rect 1809 2447 1861 2499
rect 1861 2447 1863 2499
rect 1807 2445 1863 2447
rect 2007 2483 2063 2485
rect 2007 2431 2009 2483
rect 2009 2431 2061 2483
rect 2061 2431 2063 2483
rect 2007 2429 2063 2431
rect 2207 2499 2263 2501
rect 2207 2447 2209 2499
rect 2209 2447 2261 2499
rect 2261 2447 2263 2499
rect 2207 2445 2263 2447
rect 2407 2483 2463 2485
rect 2407 2431 2409 2483
rect 2409 2431 2461 2483
rect 2461 2431 2463 2483
rect 2407 2429 2463 2431
rect 2607 2499 2663 2501
rect 2607 2447 2609 2499
rect 2609 2447 2661 2499
rect 2661 2447 2663 2499
rect 2607 2445 2663 2447
rect 2807 2483 2863 2485
rect 2807 2431 2809 2483
rect 2809 2431 2861 2483
rect 2861 2431 2863 2483
rect 2807 2429 2863 2431
rect 3007 2499 3063 2501
rect 3007 2447 3009 2499
rect 3009 2447 3061 2499
rect 3061 2447 3063 2499
rect 3007 2445 3063 2447
rect 3207 2483 3263 2485
rect 3207 2431 3209 2483
rect 3209 2431 3261 2483
rect 3261 2431 3263 2483
rect 3207 2429 3263 2431
rect 3407 2499 3463 2501
rect 3407 2447 3409 2499
rect 3409 2447 3461 2499
rect 3461 2447 3463 2499
rect 3407 2445 3463 2447
rect 3607 2483 3663 2485
rect 3607 2431 3609 2483
rect 3609 2431 3661 2483
rect 3661 2431 3663 2483
rect 3607 2429 3663 2431
rect 3807 2499 3863 2501
rect 3807 2447 3809 2499
rect 3809 2447 3861 2499
rect 3861 2447 3863 2499
rect 3807 2445 3863 2447
rect 4007 2483 4063 2485
rect 4007 2431 4009 2483
rect 4009 2431 4061 2483
rect 4061 2431 4063 2483
rect 4007 2429 4063 2431
rect 4207 2499 4263 2501
rect 4207 2447 4209 2499
rect 4209 2447 4261 2499
rect 4261 2447 4263 2499
rect 4207 2445 4263 2447
rect 4407 2483 4463 2485
rect 4407 2431 4409 2483
rect 4409 2431 4461 2483
rect 4461 2431 4463 2483
rect 4407 2429 4463 2431
rect 4607 2499 4663 2501
rect 4607 2447 4609 2499
rect 4609 2447 4661 2499
rect 4661 2447 4663 2499
rect 4607 2445 4663 2447
rect 4807 2483 4863 2485
rect 4807 2431 4809 2483
rect 4809 2431 4861 2483
rect 4861 2431 4863 2483
rect 4807 2429 4863 2431
rect 5007 2499 5063 2501
rect 5007 2447 5009 2499
rect 5009 2447 5061 2499
rect 5061 2447 5063 2499
rect 5007 2445 5063 2447
rect 5207 2483 5263 2485
rect 5207 2431 5209 2483
rect 5209 2431 5261 2483
rect 5261 2431 5263 2483
rect 5207 2429 5263 2431
rect 5407 2499 5463 2501
rect 5407 2447 5409 2499
rect 5409 2447 5461 2499
rect 5461 2447 5463 2499
rect 5407 2445 5463 2447
rect 5607 2483 5663 2485
rect 5607 2431 5609 2483
rect 5609 2431 5661 2483
rect 5661 2431 5663 2483
rect 5607 2429 5663 2431
rect 5807 2499 5863 2501
rect 5807 2447 5809 2499
rect 5809 2447 5861 2499
rect 5861 2447 5863 2499
rect 5807 2445 5863 2447
rect 6007 2483 6063 2485
rect 6007 2431 6009 2483
rect 6009 2431 6061 2483
rect 6061 2431 6063 2483
rect 6007 2429 6063 2431
rect 6207 2499 6263 2501
rect 6207 2447 6209 2499
rect 6209 2447 6261 2499
rect 6261 2447 6263 2499
rect 6207 2445 6263 2447
rect 6407 2483 6463 2485
rect 6407 2431 6409 2483
rect 6409 2431 6461 2483
rect 6461 2431 6463 2483
rect 6407 2429 6463 2431
rect 6607 2499 6663 2501
rect 6607 2447 6609 2499
rect 6609 2447 6661 2499
rect 6661 2447 6663 2499
rect 6607 2445 6663 2447
rect 6807 2483 6863 2485
rect 6807 2431 6809 2483
rect 6809 2431 6861 2483
rect 6861 2431 6863 2483
rect 6807 2429 6863 2431
rect 7007 2499 7063 2501
rect 7007 2447 7009 2499
rect 7009 2447 7061 2499
rect 7061 2447 7063 2499
rect 7007 2445 7063 2447
rect 7207 2483 7263 2485
rect 7207 2431 7209 2483
rect 7209 2431 7261 2483
rect 7261 2431 7263 2483
rect 7207 2429 7263 2431
rect 7407 2499 7463 2501
rect 7407 2447 7409 2499
rect 7409 2447 7461 2499
rect 7461 2447 7463 2499
rect 7407 2445 7463 2447
rect 7607 2483 7663 2485
rect 7607 2431 7609 2483
rect 7609 2431 7661 2483
rect 7661 2431 7663 2483
rect 7607 2429 7663 2431
rect 7807 2499 7863 2501
rect 7807 2447 7809 2499
rect 7809 2447 7861 2499
rect 7861 2447 7863 2499
rect 7807 2445 7863 2447
rect 8007 2483 8063 2485
rect 8007 2431 8009 2483
rect 8009 2431 8061 2483
rect 8061 2431 8063 2483
rect 8007 2429 8063 2431
rect 8207 2499 8263 2501
rect 8207 2447 8209 2499
rect 8209 2447 8261 2499
rect 8261 2447 8263 2499
rect 8207 2445 8263 2447
rect 8407 2483 8463 2485
rect 8407 2431 8409 2483
rect 8409 2431 8461 2483
rect 8461 2431 8463 2483
rect 8407 2429 8463 2431
rect 8607 2499 8663 2501
rect 8607 2447 8609 2499
rect 8609 2447 8661 2499
rect 8661 2447 8663 2499
rect 8607 2445 8663 2447
rect 8807 2483 8863 2485
rect 8807 2431 8809 2483
rect 8809 2431 8861 2483
rect 8861 2431 8863 2483
rect 8807 2429 8863 2431
rect 9007 2499 9063 2501
rect 9007 2447 9009 2499
rect 9009 2447 9061 2499
rect 9061 2447 9063 2499
rect 9007 2445 9063 2447
rect 9207 2483 9263 2485
rect 9207 2431 9209 2483
rect 9209 2431 9261 2483
rect 9261 2431 9263 2483
rect 9207 2429 9263 2431
rect 9407 2499 9463 2501
rect 9407 2447 9409 2499
rect 9409 2447 9461 2499
rect 9461 2447 9463 2499
rect 9407 2445 9463 2447
rect 9607 2483 9663 2485
rect 9607 2431 9609 2483
rect 9609 2431 9661 2483
rect 9661 2431 9663 2483
rect 9607 2429 9663 2431
rect 9807 2499 9863 2501
rect 9807 2447 9809 2499
rect 9809 2447 9861 2499
rect 9861 2447 9863 2499
rect 9807 2445 9863 2447
rect 10007 2483 10063 2485
rect 10007 2431 10009 2483
rect 10009 2431 10061 2483
rect 10061 2431 10063 2483
rect 10007 2429 10063 2431
rect 10207 2499 10263 2501
rect 10207 2447 10209 2499
rect 10209 2447 10261 2499
rect 10261 2447 10263 2499
rect 10207 2445 10263 2447
rect 10407 2483 10463 2485
rect 10407 2431 10409 2483
rect 10409 2431 10461 2483
rect 10461 2431 10463 2483
rect 10407 2429 10463 2431
rect 10607 2499 10663 2501
rect 10607 2447 10609 2499
rect 10609 2447 10661 2499
rect 10661 2447 10663 2499
rect 10607 2445 10663 2447
rect 10807 2483 10863 2485
rect 10807 2431 10809 2483
rect 10809 2431 10861 2483
rect 10861 2431 10863 2483
rect 10807 2429 10863 2431
rect 11007 2499 11063 2501
rect 11007 2447 11009 2499
rect 11009 2447 11061 2499
rect 11061 2447 11063 2499
rect 11007 2445 11063 2447
rect 11207 2483 11263 2485
rect 11207 2431 11209 2483
rect 11209 2431 11261 2483
rect 11261 2431 11263 2483
rect 11207 2429 11263 2431
rect 11407 2499 11463 2501
rect 11407 2447 11409 2499
rect 11409 2447 11461 2499
rect 11461 2447 11463 2499
rect 11407 2445 11463 2447
rect 11607 2483 11663 2485
rect 11607 2431 11609 2483
rect 11609 2431 11661 2483
rect 11661 2431 11663 2483
rect 11607 2429 11663 2431
rect 11807 2499 11863 2501
rect 11807 2447 11809 2499
rect 11809 2447 11861 2499
rect 11861 2447 11863 2499
rect 11807 2445 11863 2447
rect 12007 2483 12063 2485
rect 12007 2431 12009 2483
rect 12009 2431 12061 2483
rect 12061 2431 12063 2483
rect 12007 2429 12063 2431
rect 12207 2499 12263 2501
rect 12207 2447 12209 2499
rect 12209 2447 12261 2499
rect 12261 2447 12263 2499
rect 12207 2445 12263 2447
rect 12407 2483 12463 2485
rect 12407 2431 12409 2483
rect 12409 2431 12461 2483
rect 12461 2431 12463 2483
rect 12407 2429 12463 2431
rect 12607 2499 12663 2501
rect 12607 2447 12609 2499
rect 12609 2447 12661 2499
rect 12661 2447 12663 2499
rect 12607 2445 12663 2447
rect 7 1273 63 1275
rect 7 1221 9 1273
rect 9 1221 61 1273
rect 61 1221 63 1273
rect 7 1219 63 1221
rect 207 1289 263 1291
rect 207 1237 209 1289
rect 209 1237 261 1289
rect 261 1237 263 1289
rect 207 1235 263 1237
rect 407 1273 463 1275
rect 407 1221 409 1273
rect 409 1221 461 1273
rect 461 1221 463 1273
rect 407 1219 463 1221
rect 607 1289 663 1291
rect 607 1237 609 1289
rect 609 1237 661 1289
rect 661 1237 663 1289
rect 607 1235 663 1237
rect 807 1273 863 1275
rect 807 1221 809 1273
rect 809 1221 861 1273
rect 861 1221 863 1273
rect 807 1219 863 1221
rect 1007 1289 1063 1291
rect 1007 1237 1009 1289
rect 1009 1237 1061 1289
rect 1061 1237 1063 1289
rect 1007 1235 1063 1237
rect 1207 1273 1263 1275
rect 1207 1221 1209 1273
rect 1209 1221 1261 1273
rect 1261 1221 1263 1273
rect 1207 1219 1263 1221
rect 1407 1289 1463 1291
rect 1407 1237 1409 1289
rect 1409 1237 1461 1289
rect 1461 1237 1463 1289
rect 1407 1235 1463 1237
rect 1607 1273 1663 1275
rect 1607 1221 1609 1273
rect 1609 1221 1661 1273
rect 1661 1221 1663 1273
rect 1607 1219 1663 1221
rect 1807 1289 1863 1291
rect 1807 1237 1809 1289
rect 1809 1237 1861 1289
rect 1861 1237 1863 1289
rect 1807 1235 1863 1237
rect 2007 1273 2063 1275
rect 2007 1221 2009 1273
rect 2009 1221 2061 1273
rect 2061 1221 2063 1273
rect 2007 1219 2063 1221
rect 2207 1289 2263 1291
rect 2207 1237 2209 1289
rect 2209 1237 2261 1289
rect 2261 1237 2263 1289
rect 2207 1235 2263 1237
rect 2407 1273 2463 1275
rect 2407 1221 2409 1273
rect 2409 1221 2461 1273
rect 2461 1221 2463 1273
rect 2407 1219 2463 1221
rect 2607 1289 2663 1291
rect 2607 1237 2609 1289
rect 2609 1237 2661 1289
rect 2661 1237 2663 1289
rect 2607 1235 2663 1237
rect 2807 1273 2863 1275
rect 2807 1221 2809 1273
rect 2809 1221 2861 1273
rect 2861 1221 2863 1273
rect 2807 1219 2863 1221
rect 3007 1289 3063 1291
rect 3007 1237 3009 1289
rect 3009 1237 3061 1289
rect 3061 1237 3063 1289
rect 3007 1235 3063 1237
rect 3207 1273 3263 1275
rect 3207 1221 3209 1273
rect 3209 1221 3261 1273
rect 3261 1221 3263 1273
rect 3207 1219 3263 1221
rect 3407 1289 3463 1291
rect 3407 1237 3409 1289
rect 3409 1237 3461 1289
rect 3461 1237 3463 1289
rect 3407 1235 3463 1237
rect 3607 1273 3663 1275
rect 3607 1221 3609 1273
rect 3609 1221 3661 1273
rect 3661 1221 3663 1273
rect 3607 1219 3663 1221
rect 3807 1289 3863 1291
rect 3807 1237 3809 1289
rect 3809 1237 3861 1289
rect 3861 1237 3863 1289
rect 3807 1235 3863 1237
rect 4007 1273 4063 1275
rect 4007 1221 4009 1273
rect 4009 1221 4061 1273
rect 4061 1221 4063 1273
rect 4007 1219 4063 1221
rect 4207 1289 4263 1291
rect 4207 1237 4209 1289
rect 4209 1237 4261 1289
rect 4261 1237 4263 1289
rect 4207 1235 4263 1237
rect 4407 1273 4463 1275
rect 4407 1221 4409 1273
rect 4409 1221 4461 1273
rect 4461 1221 4463 1273
rect 4407 1219 4463 1221
rect 4607 1289 4663 1291
rect 4607 1237 4609 1289
rect 4609 1237 4661 1289
rect 4661 1237 4663 1289
rect 4607 1235 4663 1237
rect 4807 1273 4863 1275
rect 4807 1221 4809 1273
rect 4809 1221 4861 1273
rect 4861 1221 4863 1273
rect 4807 1219 4863 1221
rect 5007 1289 5063 1291
rect 5007 1237 5009 1289
rect 5009 1237 5061 1289
rect 5061 1237 5063 1289
rect 5007 1235 5063 1237
rect 5207 1273 5263 1275
rect 5207 1221 5209 1273
rect 5209 1221 5261 1273
rect 5261 1221 5263 1273
rect 5207 1219 5263 1221
rect 5407 1289 5463 1291
rect 5407 1237 5409 1289
rect 5409 1237 5461 1289
rect 5461 1237 5463 1289
rect 5407 1235 5463 1237
rect 5607 1273 5663 1275
rect 5607 1221 5609 1273
rect 5609 1221 5661 1273
rect 5661 1221 5663 1273
rect 5607 1219 5663 1221
rect 5807 1289 5863 1291
rect 5807 1237 5809 1289
rect 5809 1237 5861 1289
rect 5861 1237 5863 1289
rect 5807 1235 5863 1237
rect 6007 1273 6063 1275
rect 6007 1221 6009 1273
rect 6009 1221 6061 1273
rect 6061 1221 6063 1273
rect 6007 1219 6063 1221
rect 6207 1289 6263 1291
rect 6207 1237 6209 1289
rect 6209 1237 6261 1289
rect 6261 1237 6263 1289
rect 6207 1235 6263 1237
rect 6407 1273 6463 1275
rect 6407 1221 6409 1273
rect 6409 1221 6461 1273
rect 6461 1221 6463 1273
rect 6407 1219 6463 1221
rect 6607 1289 6663 1291
rect 6607 1237 6609 1289
rect 6609 1237 6661 1289
rect 6661 1237 6663 1289
rect 6607 1235 6663 1237
rect 6807 1273 6863 1275
rect 6807 1221 6809 1273
rect 6809 1221 6861 1273
rect 6861 1221 6863 1273
rect 6807 1219 6863 1221
rect 7007 1289 7063 1291
rect 7007 1237 7009 1289
rect 7009 1237 7061 1289
rect 7061 1237 7063 1289
rect 7007 1235 7063 1237
rect 7207 1273 7263 1275
rect 7207 1221 7209 1273
rect 7209 1221 7261 1273
rect 7261 1221 7263 1273
rect 7207 1219 7263 1221
rect 7407 1289 7463 1291
rect 7407 1237 7409 1289
rect 7409 1237 7461 1289
rect 7461 1237 7463 1289
rect 7407 1235 7463 1237
rect 7607 1273 7663 1275
rect 7607 1221 7609 1273
rect 7609 1221 7661 1273
rect 7661 1221 7663 1273
rect 7607 1219 7663 1221
rect 7807 1289 7863 1291
rect 7807 1237 7809 1289
rect 7809 1237 7861 1289
rect 7861 1237 7863 1289
rect 7807 1235 7863 1237
rect 8007 1273 8063 1275
rect 8007 1221 8009 1273
rect 8009 1221 8061 1273
rect 8061 1221 8063 1273
rect 8007 1219 8063 1221
rect 8207 1289 8263 1291
rect 8207 1237 8209 1289
rect 8209 1237 8261 1289
rect 8261 1237 8263 1289
rect 8207 1235 8263 1237
rect 8407 1273 8463 1275
rect 8407 1221 8409 1273
rect 8409 1221 8461 1273
rect 8461 1221 8463 1273
rect 8407 1219 8463 1221
rect 8607 1289 8663 1291
rect 8607 1237 8609 1289
rect 8609 1237 8661 1289
rect 8661 1237 8663 1289
rect 8607 1235 8663 1237
rect 8807 1273 8863 1275
rect 8807 1221 8809 1273
rect 8809 1221 8861 1273
rect 8861 1221 8863 1273
rect 8807 1219 8863 1221
rect 9007 1289 9063 1291
rect 9007 1237 9009 1289
rect 9009 1237 9061 1289
rect 9061 1237 9063 1289
rect 9007 1235 9063 1237
rect 9207 1273 9263 1275
rect 9207 1221 9209 1273
rect 9209 1221 9261 1273
rect 9261 1221 9263 1273
rect 9207 1219 9263 1221
rect 9407 1289 9463 1291
rect 9407 1237 9409 1289
rect 9409 1237 9461 1289
rect 9461 1237 9463 1289
rect 9407 1235 9463 1237
rect 9607 1273 9663 1275
rect 9607 1221 9609 1273
rect 9609 1221 9661 1273
rect 9661 1221 9663 1273
rect 9607 1219 9663 1221
rect 9807 1289 9863 1291
rect 9807 1237 9809 1289
rect 9809 1237 9861 1289
rect 9861 1237 9863 1289
rect 9807 1235 9863 1237
rect 10007 1273 10063 1275
rect 10007 1221 10009 1273
rect 10009 1221 10061 1273
rect 10061 1221 10063 1273
rect 10007 1219 10063 1221
rect 10207 1289 10263 1291
rect 10207 1237 10209 1289
rect 10209 1237 10261 1289
rect 10261 1237 10263 1289
rect 10207 1235 10263 1237
rect 10407 1273 10463 1275
rect 10407 1221 10409 1273
rect 10409 1221 10461 1273
rect 10461 1221 10463 1273
rect 10407 1219 10463 1221
rect 10607 1289 10663 1291
rect 10607 1237 10609 1289
rect 10609 1237 10661 1289
rect 10661 1237 10663 1289
rect 10607 1235 10663 1237
rect 10807 1273 10863 1275
rect 10807 1221 10809 1273
rect 10809 1221 10861 1273
rect 10861 1221 10863 1273
rect 10807 1219 10863 1221
rect 11007 1289 11063 1291
rect 11007 1237 11009 1289
rect 11009 1237 11061 1289
rect 11061 1237 11063 1289
rect 11007 1235 11063 1237
rect 11207 1273 11263 1275
rect 11207 1221 11209 1273
rect 11209 1221 11261 1273
rect 11261 1221 11263 1273
rect 11207 1219 11263 1221
rect 11407 1289 11463 1291
rect 11407 1237 11409 1289
rect 11409 1237 11461 1289
rect 11461 1237 11463 1289
rect 11407 1235 11463 1237
rect 11607 1273 11663 1275
rect 11607 1221 11609 1273
rect 11609 1221 11661 1273
rect 11661 1221 11663 1273
rect 11607 1219 11663 1221
rect 11807 1289 11863 1291
rect 11807 1237 11809 1289
rect 11809 1237 11861 1289
rect 11861 1237 11863 1289
rect 11807 1235 11863 1237
rect 12007 1273 12063 1275
rect 12007 1221 12009 1273
rect 12009 1221 12061 1273
rect 12061 1221 12063 1273
rect 12007 1219 12063 1221
rect 12207 1289 12263 1291
rect 12207 1237 12209 1289
rect 12209 1237 12261 1289
rect 12261 1237 12263 1289
rect 12207 1235 12263 1237
rect 12407 1273 12463 1275
rect 12407 1221 12409 1273
rect 12409 1221 12461 1273
rect 12461 1221 12463 1273
rect 12407 1219 12463 1221
rect 12607 1289 12663 1291
rect 12607 1237 12609 1289
rect 12609 1237 12661 1289
rect 12661 1237 12663 1289
rect 12607 1235 12663 1237
rect 7 63 63 65
rect 7 11 9 63
rect 9 11 61 63
rect 61 11 63 63
rect 7 9 63 11
rect 207 79 263 81
rect 207 27 209 79
rect 209 27 261 79
rect 261 27 263 79
rect 207 25 263 27
rect 7 -22 63 -16
rect 7 -72 9 -22
rect 9 -72 61 -22
rect 61 -72 63 -22
rect 407 63 463 65
rect 407 11 409 63
rect 409 11 461 63
rect 461 11 463 63
rect 407 9 463 11
rect 607 79 663 81
rect 607 27 609 79
rect 609 27 661 79
rect 661 27 663 79
rect 607 25 663 27
rect 207 -22 263 -16
rect 207 -72 209 -22
rect 209 -72 261 -22
rect 261 -72 263 -22
rect 407 -22 463 -16
rect 407 -72 409 -22
rect 409 -72 461 -22
rect 461 -72 463 -22
rect 807 63 863 65
rect 807 11 809 63
rect 809 11 861 63
rect 861 11 863 63
rect 807 9 863 11
rect 1007 79 1063 81
rect 1007 27 1009 79
rect 1009 27 1061 79
rect 1061 27 1063 79
rect 1007 25 1063 27
rect 607 -22 663 -16
rect 607 -72 609 -22
rect 609 -72 661 -22
rect 661 -72 663 -22
rect 807 -22 863 -16
rect 807 -72 809 -22
rect 809 -72 861 -22
rect 861 -72 863 -22
rect 1207 63 1263 65
rect 1207 11 1209 63
rect 1209 11 1261 63
rect 1261 11 1263 63
rect 1207 9 1263 11
rect 1407 79 1463 81
rect 1407 27 1409 79
rect 1409 27 1461 79
rect 1461 27 1463 79
rect 1407 25 1463 27
rect 1007 -22 1063 -16
rect 1007 -72 1009 -22
rect 1009 -72 1061 -22
rect 1061 -72 1063 -22
rect 1207 -22 1263 -16
rect 1207 -72 1209 -22
rect 1209 -72 1261 -22
rect 1261 -72 1263 -22
rect 1607 63 1663 65
rect 1607 11 1609 63
rect 1609 11 1661 63
rect 1661 11 1663 63
rect 1607 9 1663 11
rect 1807 79 1863 81
rect 1807 27 1809 79
rect 1809 27 1861 79
rect 1861 27 1863 79
rect 1807 25 1863 27
rect 1407 -22 1463 -16
rect 1407 -72 1409 -22
rect 1409 -72 1461 -22
rect 1461 -72 1463 -22
rect 1607 -22 1663 -16
rect 1607 -72 1609 -22
rect 1609 -72 1661 -22
rect 1661 -72 1663 -22
rect 2007 63 2063 65
rect 2007 11 2009 63
rect 2009 11 2061 63
rect 2061 11 2063 63
rect 2007 9 2063 11
rect 2207 79 2263 81
rect 2207 27 2209 79
rect 2209 27 2261 79
rect 2261 27 2263 79
rect 2207 25 2263 27
rect 1807 -22 1863 -16
rect 1807 -72 1809 -22
rect 1809 -72 1861 -22
rect 1861 -72 1863 -22
rect 2007 -22 2063 -16
rect 2007 -72 2009 -22
rect 2009 -72 2061 -22
rect 2061 -72 2063 -22
rect 2407 63 2463 65
rect 2407 11 2409 63
rect 2409 11 2461 63
rect 2461 11 2463 63
rect 2407 9 2463 11
rect 2607 79 2663 81
rect 2607 27 2609 79
rect 2609 27 2661 79
rect 2661 27 2663 79
rect 2607 25 2663 27
rect 2207 -22 2263 -16
rect 2207 -72 2209 -22
rect 2209 -72 2261 -22
rect 2261 -72 2263 -22
rect 2407 -22 2463 -16
rect 2407 -72 2409 -22
rect 2409 -72 2461 -22
rect 2461 -72 2463 -22
rect 2807 63 2863 65
rect 2807 11 2809 63
rect 2809 11 2861 63
rect 2861 11 2863 63
rect 2807 9 2863 11
rect 3007 79 3063 81
rect 3007 27 3009 79
rect 3009 27 3061 79
rect 3061 27 3063 79
rect 3007 25 3063 27
rect 2607 -22 2663 -16
rect 2607 -72 2609 -22
rect 2609 -72 2661 -22
rect 2661 -72 2663 -22
rect 2807 -22 2863 -16
rect 2807 -72 2809 -22
rect 2809 -72 2861 -22
rect 2861 -72 2863 -22
rect 3207 63 3263 65
rect 3207 11 3209 63
rect 3209 11 3261 63
rect 3261 11 3263 63
rect 3207 9 3263 11
rect 3407 79 3463 81
rect 3407 27 3409 79
rect 3409 27 3461 79
rect 3461 27 3463 79
rect 3407 25 3463 27
rect 3007 -22 3063 -16
rect 3007 -72 3009 -22
rect 3009 -72 3061 -22
rect 3061 -72 3063 -22
rect 3207 -22 3263 -16
rect 3207 -72 3209 -22
rect 3209 -72 3261 -22
rect 3261 -72 3263 -22
rect 3607 63 3663 65
rect 3607 11 3609 63
rect 3609 11 3661 63
rect 3661 11 3663 63
rect 3607 9 3663 11
rect 3807 79 3863 81
rect 3807 27 3809 79
rect 3809 27 3861 79
rect 3861 27 3863 79
rect 3807 25 3863 27
rect 3407 -22 3463 -16
rect 3407 -72 3409 -22
rect 3409 -72 3461 -22
rect 3461 -72 3463 -22
rect 3607 -22 3663 -16
rect 3607 -72 3609 -22
rect 3609 -72 3661 -22
rect 3661 -72 3663 -22
rect 4007 63 4063 65
rect 4007 11 4009 63
rect 4009 11 4061 63
rect 4061 11 4063 63
rect 4007 9 4063 11
rect 4207 79 4263 81
rect 4207 27 4209 79
rect 4209 27 4261 79
rect 4261 27 4263 79
rect 4207 25 4263 27
rect 3807 -22 3863 -16
rect 3807 -72 3809 -22
rect 3809 -72 3861 -22
rect 3861 -72 3863 -22
rect 4007 -22 4063 -16
rect 4007 -72 4009 -22
rect 4009 -72 4061 -22
rect 4061 -72 4063 -22
rect 4407 63 4463 65
rect 4407 11 4409 63
rect 4409 11 4461 63
rect 4461 11 4463 63
rect 4407 9 4463 11
rect 4607 79 4663 81
rect 4607 27 4609 79
rect 4609 27 4661 79
rect 4661 27 4663 79
rect 4607 25 4663 27
rect 4207 -22 4263 -16
rect 4207 -72 4209 -22
rect 4209 -72 4261 -22
rect 4261 -72 4263 -22
rect 4407 -22 4463 -16
rect 4407 -72 4409 -22
rect 4409 -72 4461 -22
rect 4461 -72 4463 -22
rect 4807 63 4863 65
rect 4807 11 4809 63
rect 4809 11 4861 63
rect 4861 11 4863 63
rect 4807 9 4863 11
rect 5007 79 5063 81
rect 5007 27 5009 79
rect 5009 27 5061 79
rect 5061 27 5063 79
rect 5007 25 5063 27
rect 4607 -22 4663 -16
rect 4607 -72 4609 -22
rect 4609 -72 4661 -22
rect 4661 -72 4663 -22
rect 4807 -22 4863 -16
rect 4807 -72 4809 -22
rect 4809 -72 4861 -22
rect 4861 -72 4863 -22
rect 5207 63 5263 65
rect 5207 11 5209 63
rect 5209 11 5261 63
rect 5261 11 5263 63
rect 5207 9 5263 11
rect 5407 79 5463 81
rect 5407 27 5409 79
rect 5409 27 5461 79
rect 5461 27 5463 79
rect 5407 25 5463 27
rect 5007 -22 5063 -16
rect 5007 -72 5009 -22
rect 5009 -72 5061 -22
rect 5061 -72 5063 -22
rect 5207 -22 5263 -16
rect 5207 -72 5209 -22
rect 5209 -72 5261 -22
rect 5261 -72 5263 -22
rect 5607 63 5663 65
rect 5607 11 5609 63
rect 5609 11 5661 63
rect 5661 11 5663 63
rect 5607 9 5663 11
rect 5807 79 5863 81
rect 5807 27 5809 79
rect 5809 27 5861 79
rect 5861 27 5863 79
rect 5807 25 5863 27
rect 5407 -22 5463 -16
rect 5407 -72 5409 -22
rect 5409 -72 5461 -22
rect 5461 -72 5463 -22
rect 5607 -22 5663 -16
rect 5607 -72 5609 -22
rect 5609 -72 5661 -22
rect 5661 -72 5663 -22
rect 6007 63 6063 65
rect 6007 11 6009 63
rect 6009 11 6061 63
rect 6061 11 6063 63
rect 6007 9 6063 11
rect 6207 79 6263 81
rect 6207 27 6209 79
rect 6209 27 6261 79
rect 6261 27 6263 79
rect 6207 25 6263 27
rect 5807 -22 5863 -16
rect 5807 -72 5809 -22
rect 5809 -72 5861 -22
rect 5861 -72 5863 -22
rect 6007 -22 6063 -16
rect 6007 -72 6009 -22
rect 6009 -72 6061 -22
rect 6061 -72 6063 -22
rect 6407 63 6463 65
rect 6407 11 6409 63
rect 6409 11 6461 63
rect 6461 11 6463 63
rect 6407 9 6463 11
rect 6607 79 6663 81
rect 6607 27 6609 79
rect 6609 27 6661 79
rect 6661 27 6663 79
rect 6607 25 6663 27
rect 6207 -22 6263 -16
rect 6207 -72 6209 -22
rect 6209 -72 6261 -22
rect 6261 -72 6263 -22
rect 6407 -22 6463 -16
rect 6407 -72 6409 -22
rect 6409 -72 6461 -22
rect 6461 -72 6463 -22
rect 6807 63 6863 65
rect 6807 11 6809 63
rect 6809 11 6861 63
rect 6861 11 6863 63
rect 6807 9 6863 11
rect 7007 79 7063 81
rect 7007 27 7009 79
rect 7009 27 7061 79
rect 7061 27 7063 79
rect 7007 25 7063 27
rect 6607 -22 6663 -16
rect 6607 -72 6609 -22
rect 6609 -72 6661 -22
rect 6661 -72 6663 -22
rect 6807 -22 6863 -16
rect 6807 -72 6809 -22
rect 6809 -72 6861 -22
rect 6861 -72 6863 -22
rect 7207 63 7263 65
rect 7207 11 7209 63
rect 7209 11 7261 63
rect 7261 11 7263 63
rect 7207 9 7263 11
rect 7407 79 7463 81
rect 7407 27 7409 79
rect 7409 27 7461 79
rect 7461 27 7463 79
rect 7407 25 7463 27
rect 7007 -22 7063 -16
rect 7007 -72 7009 -22
rect 7009 -72 7061 -22
rect 7061 -72 7063 -22
rect 7207 -22 7263 -16
rect 7207 -72 7209 -22
rect 7209 -72 7261 -22
rect 7261 -72 7263 -22
rect 7607 63 7663 65
rect 7607 11 7609 63
rect 7609 11 7661 63
rect 7661 11 7663 63
rect 7607 9 7663 11
rect 7807 79 7863 81
rect 7807 27 7809 79
rect 7809 27 7861 79
rect 7861 27 7863 79
rect 7807 25 7863 27
rect 7407 -22 7463 -16
rect 7407 -72 7409 -22
rect 7409 -72 7461 -22
rect 7461 -72 7463 -22
rect 7607 -22 7663 -16
rect 7607 -72 7609 -22
rect 7609 -72 7661 -22
rect 7661 -72 7663 -22
rect 8007 63 8063 65
rect 8007 11 8009 63
rect 8009 11 8061 63
rect 8061 11 8063 63
rect 8007 9 8063 11
rect 8207 79 8263 81
rect 8207 27 8209 79
rect 8209 27 8261 79
rect 8261 27 8263 79
rect 8207 25 8263 27
rect 7807 -22 7863 -16
rect 7807 -72 7809 -22
rect 7809 -72 7861 -22
rect 7861 -72 7863 -22
rect 8007 -22 8063 -16
rect 8007 -72 8009 -22
rect 8009 -72 8061 -22
rect 8061 -72 8063 -22
rect 8407 63 8463 65
rect 8407 11 8409 63
rect 8409 11 8461 63
rect 8461 11 8463 63
rect 8407 9 8463 11
rect 8607 79 8663 81
rect 8607 27 8609 79
rect 8609 27 8661 79
rect 8661 27 8663 79
rect 8607 25 8663 27
rect 8207 -22 8263 -16
rect 8207 -72 8209 -22
rect 8209 -72 8261 -22
rect 8261 -72 8263 -22
rect 8407 -22 8463 -16
rect 8407 -72 8409 -22
rect 8409 -72 8461 -22
rect 8461 -72 8463 -22
rect 8807 63 8863 65
rect 8807 11 8809 63
rect 8809 11 8861 63
rect 8861 11 8863 63
rect 8807 9 8863 11
rect 9007 79 9063 81
rect 9007 27 9009 79
rect 9009 27 9061 79
rect 9061 27 9063 79
rect 9007 25 9063 27
rect 8607 -22 8663 -16
rect 8607 -72 8609 -22
rect 8609 -72 8661 -22
rect 8661 -72 8663 -22
rect 8807 -22 8863 -16
rect 8807 -72 8809 -22
rect 8809 -72 8861 -22
rect 8861 -72 8863 -22
rect 9207 63 9263 65
rect 9207 11 9209 63
rect 9209 11 9261 63
rect 9261 11 9263 63
rect 9207 9 9263 11
rect 9407 79 9463 81
rect 9407 27 9409 79
rect 9409 27 9461 79
rect 9461 27 9463 79
rect 9407 25 9463 27
rect 9007 -22 9063 -16
rect 9007 -72 9009 -22
rect 9009 -72 9061 -22
rect 9061 -72 9063 -22
rect 9207 -22 9263 -16
rect 9207 -72 9209 -22
rect 9209 -72 9261 -22
rect 9261 -72 9263 -22
rect 9607 63 9663 65
rect 9607 11 9609 63
rect 9609 11 9661 63
rect 9661 11 9663 63
rect 9607 9 9663 11
rect 9807 79 9863 81
rect 9807 27 9809 79
rect 9809 27 9861 79
rect 9861 27 9863 79
rect 9807 25 9863 27
rect 9407 -22 9463 -16
rect 9407 -72 9409 -22
rect 9409 -72 9461 -22
rect 9461 -72 9463 -22
rect 9607 -22 9663 -16
rect 9607 -72 9609 -22
rect 9609 -72 9661 -22
rect 9661 -72 9663 -22
rect 10007 63 10063 65
rect 10007 11 10009 63
rect 10009 11 10061 63
rect 10061 11 10063 63
rect 10007 9 10063 11
rect 10207 79 10263 81
rect 10207 27 10209 79
rect 10209 27 10261 79
rect 10261 27 10263 79
rect 10207 25 10263 27
rect 9807 -22 9863 -16
rect 9807 -72 9809 -22
rect 9809 -72 9861 -22
rect 9861 -72 9863 -22
rect 10007 -22 10063 -16
rect 10007 -72 10009 -22
rect 10009 -72 10061 -22
rect 10061 -72 10063 -22
rect 10407 63 10463 65
rect 10407 11 10409 63
rect 10409 11 10461 63
rect 10461 11 10463 63
rect 10407 9 10463 11
rect 10607 79 10663 81
rect 10607 27 10609 79
rect 10609 27 10661 79
rect 10661 27 10663 79
rect 10607 25 10663 27
rect 10207 -22 10263 -16
rect 10207 -72 10209 -22
rect 10209 -72 10261 -22
rect 10261 -72 10263 -22
rect 10407 -22 10463 -16
rect 10407 -72 10409 -22
rect 10409 -72 10461 -22
rect 10461 -72 10463 -22
rect 10807 63 10863 65
rect 10807 11 10809 63
rect 10809 11 10861 63
rect 10861 11 10863 63
rect 10807 9 10863 11
rect 11007 79 11063 81
rect 11007 27 11009 79
rect 11009 27 11061 79
rect 11061 27 11063 79
rect 11007 25 11063 27
rect 10607 -22 10663 -16
rect 10607 -72 10609 -22
rect 10609 -72 10661 -22
rect 10661 -72 10663 -22
rect 10807 -22 10863 -16
rect 10807 -72 10809 -22
rect 10809 -72 10861 -22
rect 10861 -72 10863 -22
rect 11207 63 11263 65
rect 11207 11 11209 63
rect 11209 11 11261 63
rect 11261 11 11263 63
rect 11207 9 11263 11
rect 11407 79 11463 81
rect 11407 27 11409 79
rect 11409 27 11461 79
rect 11461 27 11463 79
rect 11407 25 11463 27
rect 11007 -22 11063 -16
rect 11007 -72 11009 -22
rect 11009 -72 11061 -22
rect 11061 -72 11063 -22
rect 11207 -22 11263 -16
rect 11207 -72 11209 -22
rect 11209 -72 11261 -22
rect 11261 -72 11263 -22
rect 11607 63 11663 65
rect 11607 11 11609 63
rect 11609 11 11661 63
rect 11661 11 11663 63
rect 11607 9 11663 11
rect 11807 79 11863 81
rect 11807 27 11809 79
rect 11809 27 11861 79
rect 11861 27 11863 79
rect 11807 25 11863 27
rect 11407 -22 11463 -16
rect 11407 -72 11409 -22
rect 11409 -72 11461 -22
rect 11461 -72 11463 -22
rect 11607 -22 11663 -16
rect 11607 -72 11609 -22
rect 11609 -72 11661 -22
rect 11661 -72 11663 -22
rect 12007 63 12063 65
rect 12007 11 12009 63
rect 12009 11 12061 63
rect 12061 11 12063 63
rect 12007 9 12063 11
rect 12207 79 12263 81
rect 12207 27 12209 79
rect 12209 27 12261 79
rect 12261 27 12263 79
rect 12207 25 12263 27
rect 11807 -22 11863 -16
rect 11807 -72 11809 -22
rect 11809 -72 11861 -22
rect 11861 -72 11863 -22
rect 12007 -22 12063 -16
rect 12007 -72 12009 -22
rect 12009 -72 12061 -22
rect 12061 -72 12063 -22
rect 12407 63 12463 65
rect 12407 11 12409 63
rect 12409 11 12461 63
rect 12461 11 12463 63
rect 12407 9 12463 11
rect 12607 79 12663 81
rect 12607 27 12609 79
rect 12609 27 12661 79
rect 12661 27 12663 79
rect 12607 25 12663 27
rect 12207 -22 12263 -16
rect 12207 -72 12209 -22
rect 12209 -72 12261 -22
rect 12261 -72 12263 -22
rect 12407 -22 12463 -16
rect 12407 -72 12409 -22
rect 12409 -72 12461 -22
rect 12461 -72 12463 -22
rect 12607 -22 12663 -16
rect 12607 -72 12609 -22
rect 12609 -72 12661 -22
rect 12661 -72 12663 -22
rect -133 -195 -91 -145
rect -91 -195 -77 -145
rect -53 -195 -39 -145
rect -39 -195 3 -145
rect -133 -201 -77 -195
rect -53 -201 3 -195
rect 67 -195 109 -145
rect 109 -195 123 -145
rect 147 -195 161 -145
rect 161 -195 203 -145
rect 67 -201 123 -195
rect 147 -201 203 -195
rect 267 -195 309 -145
rect 309 -195 323 -145
rect 347 -195 361 -145
rect 361 -195 403 -145
rect 267 -201 323 -195
rect 347 -201 403 -195
rect 467 -195 509 -145
rect 509 -195 523 -145
rect 547 -195 561 -145
rect 561 -195 603 -145
rect 467 -201 523 -195
rect 547 -201 603 -195
rect 667 -195 709 -145
rect 709 -195 723 -145
rect 747 -195 761 -145
rect 761 -195 803 -145
rect 667 -201 723 -195
rect 747 -201 803 -195
rect 867 -195 909 -145
rect 909 -195 923 -145
rect 947 -195 961 -145
rect 961 -195 1003 -145
rect 867 -201 923 -195
rect 947 -201 1003 -195
rect 1067 -195 1109 -145
rect 1109 -195 1123 -145
rect 1147 -195 1161 -145
rect 1161 -195 1203 -145
rect 1067 -201 1123 -195
rect 1147 -201 1203 -195
rect 1267 -195 1309 -145
rect 1309 -195 1323 -145
rect 1347 -195 1361 -145
rect 1361 -195 1403 -145
rect 1267 -201 1323 -195
rect 1347 -201 1403 -195
rect 1467 -195 1509 -145
rect 1509 -195 1523 -145
rect 1547 -195 1561 -145
rect 1561 -195 1603 -145
rect 1467 -201 1523 -195
rect 1547 -201 1603 -195
rect 1667 -195 1709 -145
rect 1709 -195 1723 -145
rect 1747 -195 1761 -145
rect 1761 -195 1803 -145
rect 1667 -201 1723 -195
rect 1747 -201 1803 -195
rect 1867 -195 1909 -145
rect 1909 -195 1923 -145
rect 1947 -195 1961 -145
rect 1961 -195 2003 -145
rect 1867 -201 1923 -195
rect 1947 -201 2003 -195
rect 2067 -195 2109 -145
rect 2109 -195 2123 -145
rect 2147 -195 2161 -145
rect 2161 -195 2203 -145
rect 2067 -201 2123 -195
rect 2147 -201 2203 -195
rect 2267 -195 2309 -145
rect 2309 -195 2323 -145
rect 2347 -195 2361 -145
rect 2361 -195 2403 -145
rect 2267 -201 2323 -195
rect 2347 -201 2403 -195
rect 2467 -195 2509 -145
rect 2509 -195 2523 -145
rect 2547 -195 2561 -145
rect 2561 -195 2603 -145
rect 2467 -201 2523 -195
rect 2547 -201 2603 -195
rect 2667 -195 2709 -145
rect 2709 -195 2723 -145
rect 2747 -195 2761 -145
rect 2761 -195 2803 -145
rect 2667 -201 2723 -195
rect 2747 -201 2803 -195
rect 2867 -195 2909 -145
rect 2909 -195 2923 -145
rect 2947 -195 2961 -145
rect 2961 -195 3003 -145
rect 2867 -201 2923 -195
rect 2947 -201 3003 -195
rect 3067 -195 3109 -145
rect 3109 -195 3123 -145
rect 3147 -195 3161 -145
rect 3161 -195 3203 -145
rect 3067 -201 3123 -195
rect 3147 -201 3203 -195
rect 3267 -195 3309 -145
rect 3309 -195 3323 -145
rect 3347 -195 3361 -145
rect 3361 -195 3403 -145
rect 3267 -201 3323 -195
rect 3347 -201 3403 -195
rect 3467 -195 3509 -145
rect 3509 -195 3523 -145
rect 3547 -195 3561 -145
rect 3561 -195 3603 -145
rect 3467 -201 3523 -195
rect 3547 -201 3603 -195
rect 3667 -195 3709 -145
rect 3709 -195 3723 -145
rect 3747 -195 3761 -145
rect 3761 -195 3803 -145
rect 3667 -201 3723 -195
rect 3747 -201 3803 -195
rect 3867 -195 3909 -145
rect 3909 -195 3923 -145
rect 3947 -195 3961 -145
rect 3961 -195 4003 -145
rect 3867 -201 3923 -195
rect 3947 -201 4003 -195
rect 4067 -195 4109 -145
rect 4109 -195 4123 -145
rect 4147 -195 4161 -145
rect 4161 -195 4203 -145
rect 4067 -201 4123 -195
rect 4147 -201 4203 -195
rect 4267 -195 4309 -145
rect 4309 -195 4323 -145
rect 4347 -195 4361 -145
rect 4361 -195 4403 -145
rect 4267 -201 4323 -195
rect 4347 -201 4403 -195
rect 4467 -195 4509 -145
rect 4509 -195 4523 -145
rect 4547 -195 4561 -145
rect 4561 -195 4603 -145
rect 4467 -201 4523 -195
rect 4547 -201 4603 -195
rect 4667 -195 4709 -145
rect 4709 -195 4723 -145
rect 4747 -195 4761 -145
rect 4761 -195 4803 -145
rect 4667 -201 4723 -195
rect 4747 -201 4803 -195
rect 4867 -195 4909 -145
rect 4909 -195 4923 -145
rect 4947 -195 4961 -145
rect 4961 -195 5003 -145
rect 4867 -201 4923 -195
rect 4947 -201 5003 -195
rect 5067 -195 5109 -145
rect 5109 -195 5123 -145
rect 5147 -195 5161 -145
rect 5161 -195 5203 -145
rect 5067 -201 5123 -195
rect 5147 -201 5203 -195
rect 5267 -195 5309 -145
rect 5309 -195 5323 -145
rect 5347 -195 5361 -145
rect 5361 -195 5403 -145
rect 5267 -201 5323 -195
rect 5347 -201 5403 -195
rect 5467 -195 5509 -145
rect 5509 -195 5523 -145
rect 5547 -195 5561 -145
rect 5561 -195 5603 -145
rect 5467 -201 5523 -195
rect 5547 -201 5603 -195
rect 5667 -195 5709 -145
rect 5709 -195 5723 -145
rect 5747 -195 5761 -145
rect 5761 -195 5803 -145
rect 5667 -201 5723 -195
rect 5747 -201 5803 -195
rect 5867 -195 5909 -145
rect 5909 -195 5923 -145
rect 5947 -195 5961 -145
rect 5961 -195 6003 -145
rect 5867 -201 5923 -195
rect 5947 -201 6003 -195
rect 6067 -195 6109 -145
rect 6109 -195 6123 -145
rect 6147 -195 6161 -145
rect 6161 -195 6203 -145
rect 6067 -201 6123 -195
rect 6147 -201 6203 -195
rect 6267 -195 6309 -145
rect 6309 -195 6323 -145
rect 6347 -195 6361 -145
rect 6361 -195 6403 -145
rect 6267 -201 6323 -195
rect 6347 -201 6403 -195
rect 6467 -195 6509 -145
rect 6509 -195 6523 -145
rect 6547 -195 6561 -145
rect 6561 -195 6603 -145
rect 6467 -201 6523 -195
rect 6547 -201 6603 -195
rect 6667 -195 6709 -145
rect 6709 -195 6723 -145
rect 6747 -195 6761 -145
rect 6761 -195 6803 -145
rect 6667 -201 6723 -195
rect 6747 -201 6803 -195
rect 6867 -195 6909 -145
rect 6909 -195 6923 -145
rect 6947 -195 6961 -145
rect 6961 -195 7003 -145
rect 6867 -201 6923 -195
rect 6947 -201 7003 -195
rect 7067 -195 7109 -145
rect 7109 -195 7123 -145
rect 7147 -195 7161 -145
rect 7161 -195 7203 -145
rect 7067 -201 7123 -195
rect 7147 -201 7203 -195
rect 7267 -195 7309 -145
rect 7309 -195 7323 -145
rect 7347 -195 7361 -145
rect 7361 -195 7403 -145
rect 7267 -201 7323 -195
rect 7347 -201 7403 -195
rect 7467 -195 7509 -145
rect 7509 -195 7523 -145
rect 7547 -195 7561 -145
rect 7561 -195 7603 -145
rect 7467 -201 7523 -195
rect 7547 -201 7603 -195
rect 7667 -195 7709 -145
rect 7709 -195 7723 -145
rect 7747 -195 7761 -145
rect 7761 -195 7803 -145
rect 7667 -201 7723 -195
rect 7747 -201 7803 -195
rect 7867 -195 7909 -145
rect 7909 -195 7923 -145
rect 7947 -195 7961 -145
rect 7961 -195 8003 -145
rect 7867 -201 7923 -195
rect 7947 -201 8003 -195
rect 8067 -195 8109 -145
rect 8109 -195 8123 -145
rect 8147 -195 8161 -145
rect 8161 -195 8203 -145
rect 8067 -201 8123 -195
rect 8147 -201 8203 -195
rect 8267 -195 8309 -145
rect 8309 -195 8323 -145
rect 8347 -195 8361 -145
rect 8361 -195 8403 -145
rect 8267 -201 8323 -195
rect 8347 -201 8403 -195
rect 8467 -195 8509 -145
rect 8509 -195 8523 -145
rect 8547 -195 8561 -145
rect 8561 -195 8603 -145
rect 8467 -201 8523 -195
rect 8547 -201 8603 -195
rect 8667 -195 8709 -145
rect 8709 -195 8723 -145
rect 8747 -195 8761 -145
rect 8761 -195 8803 -145
rect 8667 -201 8723 -195
rect 8747 -201 8803 -195
rect 8867 -195 8909 -145
rect 8909 -195 8923 -145
rect 8947 -195 8961 -145
rect 8961 -195 9003 -145
rect 8867 -201 8923 -195
rect 8947 -201 9003 -195
rect 9067 -195 9109 -145
rect 9109 -195 9123 -145
rect 9147 -195 9161 -145
rect 9161 -195 9203 -145
rect 9067 -201 9123 -195
rect 9147 -201 9203 -195
rect 9267 -195 9309 -145
rect 9309 -195 9323 -145
rect 9347 -195 9361 -145
rect 9361 -195 9403 -145
rect 9267 -201 9323 -195
rect 9347 -201 9403 -195
rect 9467 -195 9509 -145
rect 9509 -195 9523 -145
rect 9547 -195 9561 -145
rect 9561 -195 9603 -145
rect 9467 -201 9523 -195
rect 9547 -201 9603 -195
rect 9667 -195 9709 -145
rect 9709 -195 9723 -145
rect 9747 -195 9761 -145
rect 9761 -195 9803 -145
rect 9667 -201 9723 -195
rect 9747 -201 9803 -195
rect 9867 -195 9909 -145
rect 9909 -195 9923 -145
rect 9947 -195 9961 -145
rect 9961 -195 10003 -145
rect 9867 -201 9923 -195
rect 9947 -201 10003 -195
rect 10067 -195 10109 -145
rect 10109 -195 10123 -145
rect 10147 -195 10161 -145
rect 10161 -195 10203 -145
rect 10067 -201 10123 -195
rect 10147 -201 10203 -195
rect 10267 -195 10309 -145
rect 10309 -195 10323 -145
rect 10347 -195 10361 -145
rect 10361 -195 10403 -145
rect 10267 -201 10323 -195
rect 10347 -201 10403 -195
rect 10467 -195 10509 -145
rect 10509 -195 10523 -145
rect 10547 -195 10561 -145
rect 10561 -195 10603 -145
rect 10467 -201 10523 -195
rect 10547 -201 10603 -195
rect 10667 -195 10709 -145
rect 10709 -195 10723 -145
rect 10747 -195 10761 -145
rect 10761 -195 10803 -145
rect 10667 -201 10723 -195
rect 10747 -201 10803 -195
rect 10867 -195 10909 -145
rect 10909 -195 10923 -145
rect 10947 -195 10961 -145
rect 10961 -195 11003 -145
rect 10867 -201 10923 -195
rect 10947 -201 11003 -195
rect 11067 -195 11109 -145
rect 11109 -195 11123 -145
rect 11147 -195 11161 -145
rect 11161 -195 11203 -145
rect 11067 -201 11123 -195
rect 11147 -201 11203 -195
rect 11267 -195 11309 -145
rect 11309 -195 11323 -145
rect 11347 -195 11361 -145
rect 11361 -195 11403 -145
rect 11267 -201 11323 -195
rect 11347 -201 11403 -195
rect 11467 -195 11509 -145
rect 11509 -195 11523 -145
rect 11547 -195 11561 -145
rect 11561 -195 11603 -145
rect 11467 -201 11523 -195
rect 11547 -201 11603 -195
rect 11667 -195 11709 -145
rect 11709 -195 11723 -145
rect 11747 -195 11761 -145
rect 11761 -195 11803 -145
rect 11667 -201 11723 -195
rect 11747 -201 11803 -195
rect 11867 -195 11909 -145
rect 11909 -195 11923 -145
rect 11947 -195 11961 -145
rect 11961 -195 12003 -145
rect 11867 -201 11923 -195
rect 11947 -201 12003 -195
rect 12067 -195 12109 -145
rect 12109 -195 12123 -145
rect 12147 -195 12161 -145
rect 12161 -195 12203 -145
rect 12067 -201 12123 -195
rect 12147 -201 12203 -195
rect 12267 -195 12309 -145
rect 12309 -195 12323 -145
rect 12347 -195 12361 -145
rect 12361 -195 12403 -145
rect 12267 -201 12323 -195
rect 12347 -201 12403 -195
rect 12467 -195 12509 -145
rect 12509 -195 12523 -145
rect 12547 -195 12561 -145
rect 12561 -195 12603 -145
rect 12467 -201 12523 -195
rect 12547 -201 12603 -195
rect 12667 -195 12709 -145
rect 12709 -195 12723 -145
rect 12747 -195 12761 -145
rect 12761 -195 12803 -145
rect 12667 -201 12723 -195
rect 12747 -201 12803 -195
rect 14543 -199 14599 -197
rect 14623 -199 14679 -197
rect 14543 -251 14553 -199
rect 14553 -251 14599 -199
rect 14623 -251 14669 -199
rect 14669 -251 14679 -199
rect 14543 -253 14599 -251
rect 14623 -253 14679 -251
rect 14822 -199 14878 -197
rect 14902 -199 14958 -197
rect 14982 -199 15038 -197
rect 15062 -199 15118 -197
rect 14822 -251 14868 -199
rect 14868 -251 14878 -199
rect 14902 -251 14932 -199
rect 14932 -251 14944 -199
rect 14944 -251 14958 -199
rect 14982 -251 14996 -199
rect 14996 -251 15008 -199
rect 15008 -251 15038 -199
rect 15062 -251 15072 -199
rect 15072 -251 15118 -199
rect 14822 -253 14878 -251
rect 14902 -253 14958 -251
rect 14982 -253 15038 -251
rect 15062 -253 15118 -251
rect 15223 -199 15279 -197
rect 15303 -199 15359 -197
rect 15383 -199 15439 -197
rect 15463 -199 15519 -197
rect 15223 -251 15269 -199
rect 15269 -251 15279 -199
rect 15303 -251 15333 -199
rect 15333 -251 15345 -199
rect 15345 -251 15359 -199
rect 15383 -251 15397 -199
rect 15397 -251 15409 -199
rect 15409 -251 15439 -199
rect 15463 -251 15473 -199
rect 15473 -251 15519 -199
rect 15223 -253 15279 -251
rect 15303 -253 15359 -251
rect 15383 -253 15439 -251
rect 15463 -253 15519 -251
rect 15662 -199 15718 -197
rect 15742 -199 15798 -197
rect 15662 -251 15672 -199
rect 15672 -251 15718 -199
rect 15742 -251 15788 -199
rect 15788 -251 15798 -199
rect 15662 -253 15718 -251
rect 15742 -253 15798 -251
rect -93 -378 -91 -348
rect -91 -378 -39 -348
rect -39 -378 -37 -348
rect -93 -390 -37 -378
rect -93 -404 -91 -390
rect -91 -404 -39 -390
rect -39 -404 -37 -390
rect -93 -442 -91 -428
rect -91 -442 -39 -428
rect -39 -442 -37 -428
rect -93 -454 -37 -442
rect -93 -484 -91 -454
rect -91 -484 -39 -454
rect -39 -484 -37 -454
rect 107 -378 109 -348
rect 109 -378 161 -348
rect 161 -378 163 -348
rect 107 -390 163 -378
rect 107 -404 109 -390
rect 109 -404 161 -390
rect 161 -404 163 -390
rect 107 -442 109 -428
rect 109 -442 161 -428
rect 161 -442 163 -428
rect 107 -454 163 -442
rect 107 -484 109 -454
rect 109 -484 161 -454
rect 161 -484 163 -454
rect 307 -378 309 -348
rect 309 -378 361 -348
rect 361 -378 363 -348
rect 307 -390 363 -378
rect 307 -404 309 -390
rect 309 -404 361 -390
rect 361 -404 363 -390
rect 307 -442 309 -428
rect 309 -442 361 -428
rect 361 -442 363 -428
rect 307 -454 363 -442
rect 307 -484 309 -454
rect 309 -484 361 -454
rect 361 -484 363 -454
rect 507 -378 509 -348
rect 509 -378 561 -348
rect 561 -378 563 -348
rect 507 -390 563 -378
rect 507 -404 509 -390
rect 509 -404 561 -390
rect 561 -404 563 -390
rect 507 -442 509 -428
rect 509 -442 561 -428
rect 561 -442 563 -428
rect 507 -454 563 -442
rect 507 -484 509 -454
rect 509 -484 561 -454
rect 561 -484 563 -454
rect 707 -378 709 -348
rect 709 -378 761 -348
rect 761 -378 763 -348
rect 707 -390 763 -378
rect 707 -404 709 -390
rect 709 -404 761 -390
rect 761 -404 763 -390
rect 707 -442 709 -428
rect 709 -442 761 -428
rect 761 -442 763 -428
rect 707 -454 763 -442
rect 707 -484 709 -454
rect 709 -484 761 -454
rect 761 -484 763 -454
rect 907 -378 909 -348
rect 909 -378 961 -348
rect 961 -378 963 -348
rect 907 -390 963 -378
rect 907 -404 909 -390
rect 909 -404 961 -390
rect 961 -404 963 -390
rect 907 -442 909 -428
rect 909 -442 961 -428
rect 961 -442 963 -428
rect 907 -454 963 -442
rect 907 -484 909 -454
rect 909 -484 961 -454
rect 961 -484 963 -454
rect 1107 -378 1109 -348
rect 1109 -378 1161 -348
rect 1161 -378 1163 -348
rect 1107 -390 1163 -378
rect 1107 -404 1109 -390
rect 1109 -404 1161 -390
rect 1161 -404 1163 -390
rect 1107 -442 1109 -428
rect 1109 -442 1161 -428
rect 1161 -442 1163 -428
rect 1107 -454 1163 -442
rect 1107 -484 1109 -454
rect 1109 -484 1161 -454
rect 1161 -484 1163 -454
rect 1307 -378 1309 -348
rect 1309 -378 1361 -348
rect 1361 -378 1363 -348
rect 1307 -390 1363 -378
rect 1307 -404 1309 -390
rect 1309 -404 1361 -390
rect 1361 -404 1363 -390
rect 1307 -442 1309 -428
rect 1309 -442 1361 -428
rect 1361 -442 1363 -428
rect 1307 -454 1363 -442
rect 1307 -484 1309 -454
rect 1309 -484 1361 -454
rect 1361 -484 1363 -454
rect 1507 -378 1509 -348
rect 1509 -378 1561 -348
rect 1561 -378 1563 -348
rect 1507 -390 1563 -378
rect 1507 -404 1509 -390
rect 1509 -404 1561 -390
rect 1561 -404 1563 -390
rect 1507 -442 1509 -428
rect 1509 -442 1561 -428
rect 1561 -442 1563 -428
rect 1507 -454 1563 -442
rect 1507 -484 1509 -454
rect 1509 -484 1561 -454
rect 1561 -484 1563 -454
rect 1707 -378 1709 -348
rect 1709 -378 1761 -348
rect 1761 -378 1763 -348
rect 1707 -390 1763 -378
rect 1707 -404 1709 -390
rect 1709 -404 1761 -390
rect 1761 -404 1763 -390
rect 1707 -442 1709 -428
rect 1709 -442 1761 -428
rect 1761 -442 1763 -428
rect 1707 -454 1763 -442
rect 1707 -484 1709 -454
rect 1709 -484 1761 -454
rect 1761 -484 1763 -454
rect 1907 -378 1909 -348
rect 1909 -378 1961 -348
rect 1961 -378 1963 -348
rect 1907 -390 1963 -378
rect 1907 -404 1909 -390
rect 1909 -404 1961 -390
rect 1961 -404 1963 -390
rect 1907 -442 1909 -428
rect 1909 -442 1961 -428
rect 1961 -442 1963 -428
rect 1907 -454 1963 -442
rect 1907 -484 1909 -454
rect 1909 -484 1961 -454
rect 1961 -484 1963 -454
rect 2107 -378 2109 -348
rect 2109 -378 2161 -348
rect 2161 -378 2163 -348
rect 2107 -390 2163 -378
rect 2107 -404 2109 -390
rect 2109 -404 2161 -390
rect 2161 -404 2163 -390
rect 2107 -442 2109 -428
rect 2109 -442 2161 -428
rect 2161 -442 2163 -428
rect 2107 -454 2163 -442
rect 2107 -484 2109 -454
rect 2109 -484 2161 -454
rect 2161 -484 2163 -454
rect 2307 -378 2309 -348
rect 2309 -378 2361 -348
rect 2361 -378 2363 -348
rect 2307 -390 2363 -378
rect 2307 -404 2309 -390
rect 2309 -404 2361 -390
rect 2361 -404 2363 -390
rect 2307 -442 2309 -428
rect 2309 -442 2361 -428
rect 2361 -442 2363 -428
rect 2307 -454 2363 -442
rect 2307 -484 2309 -454
rect 2309 -484 2361 -454
rect 2361 -484 2363 -454
rect 2507 -378 2509 -348
rect 2509 -378 2561 -348
rect 2561 -378 2563 -348
rect 2507 -390 2563 -378
rect 2507 -404 2509 -390
rect 2509 -404 2561 -390
rect 2561 -404 2563 -390
rect 2507 -442 2509 -428
rect 2509 -442 2561 -428
rect 2561 -442 2563 -428
rect 2507 -454 2563 -442
rect 2507 -484 2509 -454
rect 2509 -484 2561 -454
rect 2561 -484 2563 -454
rect 2707 -378 2709 -348
rect 2709 -378 2761 -348
rect 2761 -378 2763 -348
rect 2707 -390 2763 -378
rect 2707 -404 2709 -390
rect 2709 -404 2761 -390
rect 2761 -404 2763 -390
rect 2707 -442 2709 -428
rect 2709 -442 2761 -428
rect 2761 -442 2763 -428
rect 2707 -454 2763 -442
rect 2707 -484 2709 -454
rect 2709 -484 2761 -454
rect 2761 -484 2763 -454
rect 2907 -378 2909 -348
rect 2909 -378 2961 -348
rect 2961 -378 2963 -348
rect 2907 -390 2963 -378
rect 2907 -404 2909 -390
rect 2909 -404 2961 -390
rect 2961 -404 2963 -390
rect 2907 -442 2909 -428
rect 2909 -442 2961 -428
rect 2961 -442 2963 -428
rect 2907 -454 2963 -442
rect 2907 -484 2909 -454
rect 2909 -484 2961 -454
rect 2961 -484 2963 -454
rect 3107 -378 3109 -348
rect 3109 -378 3161 -348
rect 3161 -378 3163 -348
rect 3107 -390 3163 -378
rect 3107 -404 3109 -390
rect 3109 -404 3161 -390
rect 3161 -404 3163 -390
rect 3107 -442 3109 -428
rect 3109 -442 3161 -428
rect 3161 -442 3163 -428
rect 3107 -454 3163 -442
rect 3107 -484 3109 -454
rect 3109 -484 3161 -454
rect 3161 -484 3163 -454
rect 3307 -378 3309 -348
rect 3309 -378 3361 -348
rect 3361 -378 3363 -348
rect 3307 -390 3363 -378
rect 3307 -404 3309 -390
rect 3309 -404 3361 -390
rect 3361 -404 3363 -390
rect 3307 -442 3309 -428
rect 3309 -442 3361 -428
rect 3361 -442 3363 -428
rect 3307 -454 3363 -442
rect 3307 -484 3309 -454
rect 3309 -484 3361 -454
rect 3361 -484 3363 -454
rect 3507 -378 3509 -348
rect 3509 -378 3561 -348
rect 3561 -378 3563 -348
rect 3507 -390 3563 -378
rect 3507 -404 3509 -390
rect 3509 -404 3561 -390
rect 3561 -404 3563 -390
rect 3507 -442 3509 -428
rect 3509 -442 3561 -428
rect 3561 -442 3563 -428
rect 3507 -454 3563 -442
rect 3507 -484 3509 -454
rect 3509 -484 3561 -454
rect 3561 -484 3563 -454
rect 3707 -378 3709 -348
rect 3709 -378 3761 -348
rect 3761 -378 3763 -348
rect 3707 -390 3763 -378
rect 3707 -404 3709 -390
rect 3709 -404 3761 -390
rect 3761 -404 3763 -390
rect 3707 -442 3709 -428
rect 3709 -442 3761 -428
rect 3761 -442 3763 -428
rect 3707 -454 3763 -442
rect 3707 -484 3709 -454
rect 3709 -484 3761 -454
rect 3761 -484 3763 -454
rect 3907 -378 3909 -348
rect 3909 -378 3961 -348
rect 3961 -378 3963 -348
rect 3907 -390 3963 -378
rect 3907 -404 3909 -390
rect 3909 -404 3961 -390
rect 3961 -404 3963 -390
rect 3907 -442 3909 -428
rect 3909 -442 3961 -428
rect 3961 -442 3963 -428
rect 3907 -454 3963 -442
rect 3907 -484 3909 -454
rect 3909 -484 3961 -454
rect 3961 -484 3963 -454
rect 4107 -378 4109 -348
rect 4109 -378 4161 -348
rect 4161 -378 4163 -348
rect 4107 -390 4163 -378
rect 4107 -404 4109 -390
rect 4109 -404 4161 -390
rect 4161 -404 4163 -390
rect 4107 -442 4109 -428
rect 4109 -442 4161 -428
rect 4161 -442 4163 -428
rect 4107 -454 4163 -442
rect 4107 -484 4109 -454
rect 4109 -484 4161 -454
rect 4161 -484 4163 -454
rect 4307 -378 4309 -348
rect 4309 -378 4361 -348
rect 4361 -378 4363 -348
rect 4307 -390 4363 -378
rect 4307 -404 4309 -390
rect 4309 -404 4361 -390
rect 4361 -404 4363 -390
rect 4307 -442 4309 -428
rect 4309 -442 4361 -428
rect 4361 -442 4363 -428
rect 4307 -454 4363 -442
rect 4307 -484 4309 -454
rect 4309 -484 4361 -454
rect 4361 -484 4363 -454
rect 4507 -378 4509 -348
rect 4509 -378 4561 -348
rect 4561 -378 4563 -348
rect 4507 -390 4563 -378
rect 4507 -404 4509 -390
rect 4509 -404 4561 -390
rect 4561 -404 4563 -390
rect 4507 -442 4509 -428
rect 4509 -442 4561 -428
rect 4561 -442 4563 -428
rect 4507 -454 4563 -442
rect 4507 -484 4509 -454
rect 4509 -484 4561 -454
rect 4561 -484 4563 -454
rect 4707 -378 4709 -348
rect 4709 -378 4761 -348
rect 4761 -378 4763 -348
rect 4707 -390 4763 -378
rect 4707 -404 4709 -390
rect 4709 -404 4761 -390
rect 4761 -404 4763 -390
rect 4707 -442 4709 -428
rect 4709 -442 4761 -428
rect 4761 -442 4763 -428
rect 4707 -454 4763 -442
rect 4707 -484 4709 -454
rect 4709 -484 4761 -454
rect 4761 -484 4763 -454
rect 4907 -378 4909 -348
rect 4909 -378 4961 -348
rect 4961 -378 4963 -348
rect 4907 -390 4963 -378
rect 4907 -404 4909 -390
rect 4909 -404 4961 -390
rect 4961 -404 4963 -390
rect 4907 -442 4909 -428
rect 4909 -442 4961 -428
rect 4961 -442 4963 -428
rect 4907 -454 4963 -442
rect 4907 -484 4909 -454
rect 4909 -484 4961 -454
rect 4961 -484 4963 -454
rect 5107 -378 5109 -348
rect 5109 -378 5161 -348
rect 5161 -378 5163 -348
rect 5107 -390 5163 -378
rect 5107 -404 5109 -390
rect 5109 -404 5161 -390
rect 5161 -404 5163 -390
rect 5107 -442 5109 -428
rect 5109 -442 5161 -428
rect 5161 -442 5163 -428
rect 5107 -454 5163 -442
rect 5107 -484 5109 -454
rect 5109 -484 5161 -454
rect 5161 -484 5163 -454
rect 5307 -378 5309 -348
rect 5309 -378 5361 -348
rect 5361 -378 5363 -348
rect 5307 -390 5363 -378
rect 5307 -404 5309 -390
rect 5309 -404 5361 -390
rect 5361 -404 5363 -390
rect 5307 -442 5309 -428
rect 5309 -442 5361 -428
rect 5361 -442 5363 -428
rect 5307 -454 5363 -442
rect 5307 -484 5309 -454
rect 5309 -484 5361 -454
rect 5361 -484 5363 -454
rect 5507 -378 5509 -348
rect 5509 -378 5561 -348
rect 5561 -378 5563 -348
rect 5507 -390 5563 -378
rect 5507 -404 5509 -390
rect 5509 -404 5561 -390
rect 5561 -404 5563 -390
rect 5507 -442 5509 -428
rect 5509 -442 5561 -428
rect 5561 -442 5563 -428
rect 5507 -454 5563 -442
rect 5507 -484 5509 -454
rect 5509 -484 5561 -454
rect 5561 -484 5563 -454
rect 5707 -378 5709 -348
rect 5709 -378 5761 -348
rect 5761 -378 5763 -348
rect 5707 -390 5763 -378
rect 5707 -404 5709 -390
rect 5709 -404 5761 -390
rect 5761 -404 5763 -390
rect 5707 -442 5709 -428
rect 5709 -442 5761 -428
rect 5761 -442 5763 -428
rect 5707 -454 5763 -442
rect 5707 -484 5709 -454
rect 5709 -484 5761 -454
rect 5761 -484 5763 -454
rect 5907 -378 5909 -348
rect 5909 -378 5961 -348
rect 5961 -378 5963 -348
rect 5907 -390 5963 -378
rect 5907 -404 5909 -390
rect 5909 -404 5961 -390
rect 5961 -404 5963 -390
rect 5907 -442 5909 -428
rect 5909 -442 5961 -428
rect 5961 -442 5963 -428
rect 5907 -454 5963 -442
rect 5907 -484 5909 -454
rect 5909 -484 5961 -454
rect 5961 -484 5963 -454
rect 6107 -378 6109 -348
rect 6109 -378 6161 -348
rect 6161 -378 6163 -348
rect 6107 -390 6163 -378
rect 6107 -404 6109 -390
rect 6109 -404 6161 -390
rect 6161 -404 6163 -390
rect 6107 -442 6109 -428
rect 6109 -442 6161 -428
rect 6161 -442 6163 -428
rect 6107 -454 6163 -442
rect 6107 -484 6109 -454
rect 6109 -484 6161 -454
rect 6161 -484 6163 -454
rect 6307 -378 6309 -348
rect 6309 -378 6361 -348
rect 6361 -378 6363 -348
rect 6307 -390 6363 -378
rect 6307 -404 6309 -390
rect 6309 -404 6361 -390
rect 6361 -404 6363 -390
rect 6307 -442 6309 -428
rect 6309 -442 6361 -428
rect 6361 -442 6363 -428
rect 6307 -454 6363 -442
rect 6307 -484 6309 -454
rect 6309 -484 6361 -454
rect 6361 -484 6363 -454
rect 6507 -378 6509 -348
rect 6509 -378 6561 -348
rect 6561 -378 6563 -348
rect 6507 -390 6563 -378
rect 6507 -404 6509 -390
rect 6509 -404 6561 -390
rect 6561 -404 6563 -390
rect 6507 -442 6509 -428
rect 6509 -442 6561 -428
rect 6561 -442 6563 -428
rect 6507 -454 6563 -442
rect 6507 -484 6509 -454
rect 6509 -484 6561 -454
rect 6561 -484 6563 -454
rect 6707 -378 6709 -348
rect 6709 -378 6761 -348
rect 6761 -378 6763 -348
rect 6707 -390 6763 -378
rect 6707 -404 6709 -390
rect 6709 -404 6761 -390
rect 6761 -404 6763 -390
rect 6707 -442 6709 -428
rect 6709 -442 6761 -428
rect 6761 -442 6763 -428
rect 6707 -454 6763 -442
rect 6707 -484 6709 -454
rect 6709 -484 6761 -454
rect 6761 -484 6763 -454
rect 6907 -378 6909 -348
rect 6909 -378 6961 -348
rect 6961 -378 6963 -348
rect 6907 -390 6963 -378
rect 6907 -404 6909 -390
rect 6909 -404 6961 -390
rect 6961 -404 6963 -390
rect 6907 -442 6909 -428
rect 6909 -442 6961 -428
rect 6961 -442 6963 -428
rect 6907 -454 6963 -442
rect 6907 -484 6909 -454
rect 6909 -484 6961 -454
rect 6961 -484 6963 -454
rect 7107 -378 7109 -348
rect 7109 -378 7161 -348
rect 7161 -378 7163 -348
rect 7107 -390 7163 -378
rect 7107 -404 7109 -390
rect 7109 -404 7161 -390
rect 7161 -404 7163 -390
rect 7107 -442 7109 -428
rect 7109 -442 7161 -428
rect 7161 -442 7163 -428
rect 7107 -454 7163 -442
rect 7107 -484 7109 -454
rect 7109 -484 7161 -454
rect 7161 -484 7163 -454
rect 7307 -378 7309 -348
rect 7309 -378 7361 -348
rect 7361 -378 7363 -348
rect 7307 -390 7363 -378
rect 7307 -404 7309 -390
rect 7309 -404 7361 -390
rect 7361 -404 7363 -390
rect 7307 -442 7309 -428
rect 7309 -442 7361 -428
rect 7361 -442 7363 -428
rect 7307 -454 7363 -442
rect 7307 -484 7309 -454
rect 7309 -484 7361 -454
rect 7361 -484 7363 -454
rect 7507 -378 7509 -348
rect 7509 -378 7561 -348
rect 7561 -378 7563 -348
rect 7507 -390 7563 -378
rect 7507 -404 7509 -390
rect 7509 -404 7561 -390
rect 7561 -404 7563 -390
rect 7507 -442 7509 -428
rect 7509 -442 7561 -428
rect 7561 -442 7563 -428
rect 7507 -454 7563 -442
rect 7507 -484 7509 -454
rect 7509 -484 7561 -454
rect 7561 -484 7563 -454
rect 7707 -378 7709 -348
rect 7709 -378 7761 -348
rect 7761 -378 7763 -348
rect 7707 -390 7763 -378
rect 7707 -404 7709 -390
rect 7709 -404 7761 -390
rect 7761 -404 7763 -390
rect 7707 -442 7709 -428
rect 7709 -442 7761 -428
rect 7761 -442 7763 -428
rect 7707 -454 7763 -442
rect 7707 -484 7709 -454
rect 7709 -484 7761 -454
rect 7761 -484 7763 -454
rect 7907 -378 7909 -348
rect 7909 -378 7961 -348
rect 7961 -378 7963 -348
rect 7907 -390 7963 -378
rect 7907 -404 7909 -390
rect 7909 -404 7961 -390
rect 7961 -404 7963 -390
rect 7907 -442 7909 -428
rect 7909 -442 7961 -428
rect 7961 -442 7963 -428
rect 7907 -454 7963 -442
rect 7907 -484 7909 -454
rect 7909 -484 7961 -454
rect 7961 -484 7963 -454
rect 8107 -378 8109 -348
rect 8109 -378 8161 -348
rect 8161 -378 8163 -348
rect 8107 -390 8163 -378
rect 8107 -404 8109 -390
rect 8109 -404 8161 -390
rect 8161 -404 8163 -390
rect 8107 -442 8109 -428
rect 8109 -442 8161 -428
rect 8161 -442 8163 -428
rect 8107 -454 8163 -442
rect 8107 -484 8109 -454
rect 8109 -484 8161 -454
rect 8161 -484 8163 -454
rect 8307 -378 8309 -348
rect 8309 -378 8361 -348
rect 8361 -378 8363 -348
rect 8307 -390 8363 -378
rect 8307 -404 8309 -390
rect 8309 -404 8361 -390
rect 8361 -404 8363 -390
rect 8307 -442 8309 -428
rect 8309 -442 8361 -428
rect 8361 -442 8363 -428
rect 8307 -454 8363 -442
rect 8307 -484 8309 -454
rect 8309 -484 8361 -454
rect 8361 -484 8363 -454
rect 8507 -378 8509 -348
rect 8509 -378 8561 -348
rect 8561 -378 8563 -348
rect 8507 -390 8563 -378
rect 8507 -404 8509 -390
rect 8509 -404 8561 -390
rect 8561 -404 8563 -390
rect 8507 -442 8509 -428
rect 8509 -442 8561 -428
rect 8561 -442 8563 -428
rect 8507 -454 8563 -442
rect 8507 -484 8509 -454
rect 8509 -484 8561 -454
rect 8561 -484 8563 -454
rect 8707 -378 8709 -348
rect 8709 -378 8761 -348
rect 8761 -378 8763 -348
rect 8707 -390 8763 -378
rect 8707 -404 8709 -390
rect 8709 -404 8761 -390
rect 8761 -404 8763 -390
rect 8707 -442 8709 -428
rect 8709 -442 8761 -428
rect 8761 -442 8763 -428
rect 8707 -454 8763 -442
rect 8707 -484 8709 -454
rect 8709 -484 8761 -454
rect 8761 -484 8763 -454
rect 8907 -378 8909 -348
rect 8909 -378 8961 -348
rect 8961 -378 8963 -348
rect 8907 -390 8963 -378
rect 8907 -404 8909 -390
rect 8909 -404 8961 -390
rect 8961 -404 8963 -390
rect 8907 -442 8909 -428
rect 8909 -442 8961 -428
rect 8961 -442 8963 -428
rect 8907 -454 8963 -442
rect 8907 -484 8909 -454
rect 8909 -484 8961 -454
rect 8961 -484 8963 -454
rect 9107 -378 9109 -348
rect 9109 -378 9161 -348
rect 9161 -378 9163 -348
rect 9107 -390 9163 -378
rect 9107 -404 9109 -390
rect 9109 -404 9161 -390
rect 9161 -404 9163 -390
rect 9107 -442 9109 -428
rect 9109 -442 9161 -428
rect 9161 -442 9163 -428
rect 9107 -454 9163 -442
rect 9107 -484 9109 -454
rect 9109 -484 9161 -454
rect 9161 -484 9163 -454
rect 9307 -378 9309 -348
rect 9309 -378 9361 -348
rect 9361 -378 9363 -348
rect 9307 -390 9363 -378
rect 9307 -404 9309 -390
rect 9309 -404 9361 -390
rect 9361 -404 9363 -390
rect 9307 -442 9309 -428
rect 9309 -442 9361 -428
rect 9361 -442 9363 -428
rect 9307 -454 9363 -442
rect 9307 -484 9309 -454
rect 9309 -484 9361 -454
rect 9361 -484 9363 -454
rect 9507 -378 9509 -348
rect 9509 -378 9561 -348
rect 9561 -378 9563 -348
rect 9507 -390 9563 -378
rect 9507 -404 9509 -390
rect 9509 -404 9561 -390
rect 9561 -404 9563 -390
rect 9507 -442 9509 -428
rect 9509 -442 9561 -428
rect 9561 -442 9563 -428
rect 9507 -454 9563 -442
rect 9507 -484 9509 -454
rect 9509 -484 9561 -454
rect 9561 -484 9563 -454
rect 9707 -378 9709 -348
rect 9709 -378 9761 -348
rect 9761 -378 9763 -348
rect 9707 -390 9763 -378
rect 9707 -404 9709 -390
rect 9709 -404 9761 -390
rect 9761 -404 9763 -390
rect 9707 -442 9709 -428
rect 9709 -442 9761 -428
rect 9761 -442 9763 -428
rect 9707 -454 9763 -442
rect 9707 -484 9709 -454
rect 9709 -484 9761 -454
rect 9761 -484 9763 -454
rect 9907 -378 9909 -348
rect 9909 -378 9961 -348
rect 9961 -378 9963 -348
rect 9907 -390 9963 -378
rect 9907 -404 9909 -390
rect 9909 -404 9961 -390
rect 9961 -404 9963 -390
rect 9907 -442 9909 -428
rect 9909 -442 9961 -428
rect 9961 -442 9963 -428
rect 9907 -454 9963 -442
rect 9907 -484 9909 -454
rect 9909 -484 9961 -454
rect 9961 -484 9963 -454
rect 10107 -378 10109 -348
rect 10109 -378 10161 -348
rect 10161 -378 10163 -348
rect 10107 -390 10163 -378
rect 10107 -404 10109 -390
rect 10109 -404 10161 -390
rect 10161 -404 10163 -390
rect 10107 -442 10109 -428
rect 10109 -442 10161 -428
rect 10161 -442 10163 -428
rect 10107 -454 10163 -442
rect 10107 -484 10109 -454
rect 10109 -484 10161 -454
rect 10161 -484 10163 -454
rect 10307 -378 10309 -348
rect 10309 -378 10361 -348
rect 10361 -378 10363 -348
rect 10307 -390 10363 -378
rect 10307 -404 10309 -390
rect 10309 -404 10361 -390
rect 10361 -404 10363 -390
rect 10307 -442 10309 -428
rect 10309 -442 10361 -428
rect 10361 -442 10363 -428
rect 10307 -454 10363 -442
rect 10307 -484 10309 -454
rect 10309 -484 10361 -454
rect 10361 -484 10363 -454
rect 10507 -378 10509 -348
rect 10509 -378 10561 -348
rect 10561 -378 10563 -348
rect 10507 -390 10563 -378
rect 10507 -404 10509 -390
rect 10509 -404 10561 -390
rect 10561 -404 10563 -390
rect 10507 -442 10509 -428
rect 10509 -442 10561 -428
rect 10561 -442 10563 -428
rect 10507 -454 10563 -442
rect 10507 -484 10509 -454
rect 10509 -484 10561 -454
rect 10561 -484 10563 -454
rect 10707 -378 10709 -348
rect 10709 -378 10761 -348
rect 10761 -378 10763 -348
rect 10707 -390 10763 -378
rect 10707 -404 10709 -390
rect 10709 -404 10761 -390
rect 10761 -404 10763 -390
rect 10707 -442 10709 -428
rect 10709 -442 10761 -428
rect 10761 -442 10763 -428
rect 10707 -454 10763 -442
rect 10707 -484 10709 -454
rect 10709 -484 10761 -454
rect 10761 -484 10763 -454
rect 10907 -378 10909 -348
rect 10909 -378 10961 -348
rect 10961 -378 10963 -348
rect 10907 -390 10963 -378
rect 10907 -404 10909 -390
rect 10909 -404 10961 -390
rect 10961 -404 10963 -390
rect 10907 -442 10909 -428
rect 10909 -442 10961 -428
rect 10961 -442 10963 -428
rect 10907 -454 10963 -442
rect 10907 -484 10909 -454
rect 10909 -484 10961 -454
rect 10961 -484 10963 -454
rect 11107 -378 11109 -348
rect 11109 -378 11161 -348
rect 11161 -378 11163 -348
rect 11107 -390 11163 -378
rect 11107 -404 11109 -390
rect 11109 -404 11161 -390
rect 11161 -404 11163 -390
rect 11107 -442 11109 -428
rect 11109 -442 11161 -428
rect 11161 -442 11163 -428
rect 11107 -454 11163 -442
rect 11107 -484 11109 -454
rect 11109 -484 11161 -454
rect 11161 -484 11163 -454
rect 11307 -378 11309 -348
rect 11309 -378 11361 -348
rect 11361 -378 11363 -348
rect 11307 -390 11363 -378
rect 11307 -404 11309 -390
rect 11309 -404 11361 -390
rect 11361 -404 11363 -390
rect 11307 -442 11309 -428
rect 11309 -442 11361 -428
rect 11361 -442 11363 -428
rect 11307 -454 11363 -442
rect 11307 -484 11309 -454
rect 11309 -484 11361 -454
rect 11361 -484 11363 -454
rect 11507 -378 11509 -348
rect 11509 -378 11561 -348
rect 11561 -378 11563 -348
rect 11507 -390 11563 -378
rect 11507 -404 11509 -390
rect 11509 -404 11561 -390
rect 11561 -404 11563 -390
rect 11507 -442 11509 -428
rect 11509 -442 11561 -428
rect 11561 -442 11563 -428
rect 11507 -454 11563 -442
rect 11507 -484 11509 -454
rect 11509 -484 11561 -454
rect 11561 -484 11563 -454
rect 11707 -378 11709 -348
rect 11709 -378 11761 -348
rect 11761 -378 11763 -348
rect 11707 -390 11763 -378
rect 11707 -404 11709 -390
rect 11709 -404 11761 -390
rect 11761 -404 11763 -390
rect 11707 -442 11709 -428
rect 11709 -442 11761 -428
rect 11761 -442 11763 -428
rect 11707 -454 11763 -442
rect 11707 -484 11709 -454
rect 11709 -484 11761 -454
rect 11761 -484 11763 -454
rect 11907 -378 11909 -348
rect 11909 -378 11961 -348
rect 11961 -378 11963 -348
rect 11907 -390 11963 -378
rect 11907 -404 11909 -390
rect 11909 -404 11961 -390
rect 11961 -404 11963 -390
rect 11907 -442 11909 -428
rect 11909 -442 11961 -428
rect 11961 -442 11963 -428
rect 11907 -454 11963 -442
rect 11907 -484 11909 -454
rect 11909 -484 11961 -454
rect 11961 -484 11963 -454
rect 12107 -378 12109 -348
rect 12109 -378 12161 -348
rect 12161 -378 12163 -348
rect 12107 -390 12163 -378
rect 12107 -404 12109 -390
rect 12109 -404 12161 -390
rect 12161 -404 12163 -390
rect 12107 -442 12109 -428
rect 12109 -442 12161 -428
rect 12161 -442 12163 -428
rect 12107 -454 12163 -442
rect 12107 -484 12109 -454
rect 12109 -484 12161 -454
rect 12161 -484 12163 -454
rect 12307 -378 12309 -348
rect 12309 -378 12361 -348
rect 12361 -378 12363 -348
rect 12307 -390 12363 -378
rect 12307 -404 12309 -390
rect 12309 -404 12361 -390
rect 12361 -404 12363 -390
rect 12307 -442 12309 -428
rect 12309 -442 12361 -428
rect 12361 -442 12363 -428
rect 12307 -454 12363 -442
rect 12307 -484 12309 -454
rect 12309 -484 12361 -454
rect 12361 -484 12363 -454
rect 12507 -378 12509 -348
rect 12509 -378 12561 -348
rect 12561 -378 12563 -348
rect 12507 -390 12563 -378
rect 12507 -404 12509 -390
rect 12509 -404 12561 -390
rect 12561 -404 12563 -390
rect 12507 -442 12509 -428
rect 12509 -442 12561 -428
rect 12561 -442 12563 -428
rect 12507 -454 12563 -442
rect 12507 -484 12509 -454
rect 12509 -484 12561 -454
rect 12561 -484 12563 -454
rect 12707 -378 12709 -348
rect 12709 -378 12761 -348
rect 12761 -378 12763 -348
rect 12707 -390 12763 -378
rect 12707 -404 12709 -390
rect 12709 -404 12761 -390
rect 12761 -404 12763 -390
rect 12707 -442 12709 -428
rect 12709 -442 12761 -428
rect 12761 -442 12763 -428
rect 12707 -454 12763 -442
rect 12707 -484 12709 -454
rect 12709 -484 12761 -454
rect 12761 -484 12763 -454
rect 14543 -399 14599 -397
rect 14623 -399 14679 -397
rect 14543 -451 14553 -399
rect 14553 -451 14599 -399
rect 14623 -451 14669 -399
rect 14669 -451 14679 -399
rect 14543 -453 14599 -451
rect 14623 -453 14679 -451
rect 14822 -399 14878 -397
rect 14902 -399 14958 -397
rect 14982 -399 15038 -397
rect 15062 -399 15118 -397
rect 14822 -451 14868 -399
rect 14868 -451 14878 -399
rect 14902 -451 14932 -399
rect 14932 -451 14944 -399
rect 14944 -451 14958 -399
rect 14982 -451 14996 -399
rect 14996 -451 15008 -399
rect 15008 -451 15038 -399
rect 15062 -451 15072 -399
rect 15072 -451 15118 -399
rect 14822 -453 14878 -451
rect 14902 -453 14958 -451
rect 14982 -453 15038 -451
rect 15062 -453 15118 -451
rect 15223 -399 15279 -397
rect 15303 -399 15359 -397
rect 15383 -399 15439 -397
rect 15463 -399 15519 -397
rect 15223 -451 15269 -399
rect 15269 -451 15279 -399
rect 15303 -451 15333 -399
rect 15333 -451 15345 -399
rect 15345 -451 15359 -399
rect 15383 -451 15397 -399
rect 15397 -451 15409 -399
rect 15409 -451 15439 -399
rect 15463 -451 15473 -399
rect 15473 -451 15519 -399
rect 15223 -453 15279 -451
rect 15303 -453 15359 -451
rect 15383 -453 15439 -451
rect 15463 -453 15519 -451
rect 15662 -399 15718 -397
rect 15742 -399 15798 -397
rect 15662 -451 15672 -399
rect 15672 -451 15718 -399
rect 15742 -451 15788 -399
rect 15788 -451 15798 -399
rect 15662 -453 15718 -451
rect 15742 -453 15798 -451
rect 14543 -599 14599 -597
rect 14623 -599 14679 -597
rect 14543 -651 14553 -599
rect 14553 -651 14599 -599
rect 14623 -651 14669 -599
rect 14669 -651 14679 -599
rect 14543 -653 14599 -651
rect 14623 -653 14679 -651
rect 14822 -599 14878 -597
rect 14902 -599 14958 -597
rect 14982 -599 15038 -597
rect 15062 -599 15118 -597
rect 14822 -651 14868 -599
rect 14868 -651 14878 -599
rect 14902 -651 14932 -599
rect 14932 -651 14944 -599
rect 14944 -651 14958 -599
rect 14982 -651 14996 -599
rect 14996 -651 15008 -599
rect 15008 -651 15038 -599
rect 15062 -651 15072 -599
rect 15072 -651 15118 -599
rect 14822 -653 14878 -651
rect 14902 -653 14958 -651
rect 14982 -653 15038 -651
rect 15062 -653 15118 -651
rect 15223 -599 15279 -597
rect 15303 -599 15359 -597
rect 15383 -599 15439 -597
rect 15463 -599 15519 -597
rect 15223 -651 15269 -599
rect 15269 -651 15279 -599
rect 15303 -651 15333 -599
rect 15333 -651 15345 -599
rect 15345 -651 15359 -599
rect 15383 -651 15397 -599
rect 15397 -651 15409 -599
rect 15409 -651 15439 -599
rect 15463 -651 15473 -599
rect 15473 -651 15519 -599
rect 15223 -653 15279 -651
rect 15303 -653 15359 -651
rect 15383 -653 15439 -651
rect 15463 -653 15519 -651
rect 15662 -599 15718 -597
rect 15742 -599 15798 -597
rect 15662 -651 15672 -599
rect 15672 -651 15718 -599
rect 15742 -651 15788 -599
rect 15788 -651 15798 -599
rect 15662 -653 15718 -651
rect 15742 -653 15798 -651
rect 14543 -799 14599 -797
rect 14623 -799 14679 -797
rect 14543 -851 14553 -799
rect 14553 -851 14599 -799
rect 14623 -851 14669 -799
rect 14669 -851 14679 -799
rect 14543 -853 14599 -851
rect 14623 -853 14679 -851
rect 14822 -799 14878 -797
rect 14902 -799 14958 -797
rect 14982 -799 15038 -797
rect 15062 -799 15118 -797
rect 14822 -851 14868 -799
rect 14868 -851 14878 -799
rect 14902 -851 14932 -799
rect 14932 -851 14944 -799
rect 14944 -851 14958 -799
rect 14982 -851 14996 -799
rect 14996 -851 15008 -799
rect 15008 -851 15038 -799
rect 15062 -851 15072 -799
rect 15072 -851 15118 -799
rect 14822 -853 14878 -851
rect 14902 -853 14958 -851
rect 14982 -853 15038 -851
rect 15062 -853 15118 -851
rect 15223 -799 15279 -797
rect 15303 -799 15359 -797
rect 15383 -799 15439 -797
rect 15463 -799 15519 -797
rect 15223 -851 15269 -799
rect 15269 -851 15279 -799
rect 15303 -851 15333 -799
rect 15333 -851 15345 -799
rect 15345 -851 15359 -799
rect 15383 -851 15397 -799
rect 15397 -851 15409 -799
rect 15409 -851 15439 -799
rect 15463 -851 15473 -799
rect 15473 -851 15519 -799
rect 15223 -853 15279 -851
rect 15303 -853 15359 -851
rect 15383 -853 15439 -851
rect 15463 -853 15519 -851
rect 15662 -799 15718 -797
rect 15742 -799 15798 -797
rect 15662 -851 15672 -799
rect 15672 -851 15718 -799
rect 15742 -851 15788 -799
rect 15788 -851 15798 -799
rect 15662 -853 15718 -851
rect 15742 -853 15798 -851
rect 14543 -999 14599 -997
rect 14623 -999 14679 -997
rect 14543 -1051 14553 -999
rect 14553 -1051 14599 -999
rect 14623 -1051 14669 -999
rect 14669 -1051 14679 -999
rect 14543 -1053 14599 -1051
rect 14623 -1053 14679 -1051
rect 14822 -999 14878 -997
rect 14902 -999 14958 -997
rect 14982 -999 15038 -997
rect 15062 -999 15118 -997
rect 14822 -1051 14868 -999
rect 14868 -1051 14878 -999
rect 14902 -1051 14932 -999
rect 14932 -1051 14944 -999
rect 14944 -1051 14958 -999
rect 14982 -1051 14996 -999
rect 14996 -1051 15008 -999
rect 15008 -1051 15038 -999
rect 15062 -1051 15072 -999
rect 15072 -1051 15118 -999
rect 14822 -1053 14878 -1051
rect 14902 -1053 14958 -1051
rect 14982 -1053 15038 -1051
rect 15062 -1053 15118 -1051
rect 15223 -999 15279 -997
rect 15303 -999 15359 -997
rect 15383 -999 15439 -997
rect 15463 -999 15519 -997
rect 15223 -1051 15269 -999
rect 15269 -1051 15279 -999
rect 15303 -1051 15333 -999
rect 15333 -1051 15345 -999
rect 15345 -1051 15359 -999
rect 15383 -1051 15397 -999
rect 15397 -1051 15409 -999
rect 15409 -1051 15439 -999
rect 15463 -1051 15473 -999
rect 15473 -1051 15519 -999
rect 15223 -1053 15279 -1051
rect 15303 -1053 15359 -1051
rect 15383 -1053 15439 -1051
rect 15463 -1053 15519 -1051
rect 15662 -999 15718 -997
rect 15742 -999 15798 -997
rect 15662 -1051 15672 -999
rect 15672 -1051 15718 -999
rect 15742 -1051 15788 -999
rect 15788 -1051 15798 -999
rect 15662 -1053 15718 -1051
rect 15742 -1053 15798 -1051
rect 14543 -1199 14599 -1197
rect 14623 -1199 14679 -1197
rect 14543 -1251 14553 -1199
rect 14553 -1251 14599 -1199
rect 14623 -1251 14669 -1199
rect 14669 -1251 14679 -1199
rect 14543 -1253 14599 -1251
rect 14623 -1253 14679 -1251
rect 14822 -1199 14878 -1197
rect 14902 -1199 14958 -1197
rect 14982 -1199 15038 -1197
rect 15062 -1199 15118 -1197
rect 14822 -1251 14868 -1199
rect 14868 -1251 14878 -1199
rect 14902 -1251 14932 -1199
rect 14932 -1251 14944 -1199
rect 14944 -1251 14958 -1199
rect 14982 -1251 14996 -1199
rect 14996 -1251 15008 -1199
rect 15008 -1251 15038 -1199
rect 15062 -1251 15072 -1199
rect 15072 -1251 15118 -1199
rect 14822 -1253 14878 -1251
rect 14902 -1253 14958 -1251
rect 14982 -1253 15038 -1251
rect 15062 -1253 15118 -1251
rect 15223 -1199 15279 -1197
rect 15303 -1199 15359 -1197
rect 15383 -1199 15439 -1197
rect 15463 -1199 15519 -1197
rect 15223 -1251 15269 -1199
rect 15269 -1251 15279 -1199
rect 15303 -1251 15333 -1199
rect 15333 -1251 15345 -1199
rect 15345 -1251 15359 -1199
rect 15383 -1251 15397 -1199
rect 15397 -1251 15409 -1199
rect 15409 -1251 15439 -1199
rect 15463 -1251 15473 -1199
rect 15473 -1251 15519 -1199
rect 15223 -1253 15279 -1251
rect 15303 -1253 15359 -1251
rect 15383 -1253 15439 -1251
rect 15463 -1253 15519 -1251
rect 15662 -1199 15718 -1197
rect 15742 -1199 15798 -1197
rect 15662 -1251 15672 -1199
rect 15672 -1251 15718 -1199
rect 15742 -1251 15788 -1199
rect 15788 -1251 15798 -1199
rect 15662 -1253 15718 -1251
rect 15742 -1253 15798 -1251
rect 14543 -1399 14599 -1397
rect 14623 -1399 14679 -1397
rect 14543 -1451 14553 -1399
rect 14553 -1451 14599 -1399
rect 14623 -1451 14669 -1399
rect 14669 -1451 14679 -1399
rect 14543 -1453 14599 -1451
rect 14623 -1453 14679 -1451
rect 14822 -1399 14878 -1397
rect 14902 -1399 14958 -1397
rect 14982 -1399 15038 -1397
rect 15062 -1399 15118 -1397
rect 14822 -1451 14868 -1399
rect 14868 -1451 14878 -1399
rect 14902 -1451 14932 -1399
rect 14932 -1451 14944 -1399
rect 14944 -1451 14958 -1399
rect 14982 -1451 14996 -1399
rect 14996 -1451 15008 -1399
rect 15008 -1451 15038 -1399
rect 15062 -1451 15072 -1399
rect 15072 -1451 15118 -1399
rect 14822 -1453 14878 -1451
rect 14902 -1453 14958 -1451
rect 14982 -1453 15038 -1451
rect 15062 -1453 15118 -1451
rect 15223 -1399 15279 -1397
rect 15303 -1399 15359 -1397
rect 15383 -1399 15439 -1397
rect 15463 -1399 15519 -1397
rect 15223 -1451 15269 -1399
rect 15269 -1451 15279 -1399
rect 15303 -1451 15333 -1399
rect 15333 -1451 15345 -1399
rect 15345 -1451 15359 -1399
rect 15383 -1451 15397 -1399
rect 15397 -1451 15409 -1399
rect 15409 -1451 15439 -1399
rect 15463 -1451 15473 -1399
rect 15473 -1451 15519 -1399
rect 15223 -1453 15279 -1451
rect 15303 -1453 15359 -1451
rect 15383 -1453 15439 -1451
rect 15463 -1453 15519 -1451
rect 15662 -1399 15718 -1397
rect 15742 -1399 15798 -1397
rect 15662 -1451 15672 -1399
rect 15672 -1451 15718 -1399
rect 15742 -1451 15788 -1399
rect 15788 -1451 15798 -1399
rect 15662 -1453 15718 -1451
rect 15742 -1453 15798 -1451
rect 14543 -1599 14599 -1597
rect 14623 -1599 14679 -1597
rect 14543 -1651 14553 -1599
rect 14553 -1651 14599 -1599
rect 14623 -1651 14669 -1599
rect 14669 -1651 14679 -1599
rect 14543 -1653 14599 -1651
rect 14623 -1653 14679 -1651
rect 14822 -1599 14878 -1597
rect 14902 -1599 14958 -1597
rect 14982 -1599 15038 -1597
rect 15062 -1599 15118 -1597
rect 14822 -1651 14868 -1599
rect 14868 -1651 14878 -1599
rect 14902 -1651 14932 -1599
rect 14932 -1651 14944 -1599
rect 14944 -1651 14958 -1599
rect 14982 -1651 14996 -1599
rect 14996 -1651 15008 -1599
rect 15008 -1651 15038 -1599
rect 15062 -1651 15072 -1599
rect 15072 -1651 15118 -1599
rect 14822 -1653 14878 -1651
rect 14902 -1653 14958 -1651
rect 14982 -1653 15038 -1651
rect 15062 -1653 15118 -1651
rect 15223 -1599 15279 -1597
rect 15303 -1599 15359 -1597
rect 15383 -1599 15439 -1597
rect 15463 -1599 15519 -1597
rect 15223 -1651 15269 -1599
rect 15269 -1651 15279 -1599
rect 15303 -1651 15333 -1599
rect 15333 -1651 15345 -1599
rect 15345 -1651 15359 -1599
rect 15383 -1651 15397 -1599
rect 15397 -1651 15409 -1599
rect 15409 -1651 15439 -1599
rect 15463 -1651 15473 -1599
rect 15473 -1651 15519 -1599
rect 15223 -1653 15279 -1651
rect 15303 -1653 15359 -1651
rect 15383 -1653 15439 -1651
rect 15463 -1653 15519 -1651
rect 15662 -1599 15718 -1597
rect 15742 -1599 15798 -1597
rect 15662 -1651 15672 -1599
rect 15672 -1651 15718 -1599
rect 15742 -1651 15788 -1599
rect 15788 -1651 15798 -1599
rect 15662 -1653 15718 -1651
rect 15742 -1653 15798 -1651
rect 14543 -1799 14599 -1797
rect 14623 -1799 14679 -1797
rect 14543 -1851 14553 -1799
rect 14553 -1851 14599 -1799
rect 14623 -1851 14669 -1799
rect 14669 -1851 14679 -1799
rect 14543 -1853 14599 -1851
rect 14623 -1853 14679 -1851
rect 14822 -1799 14878 -1797
rect 14902 -1799 14958 -1797
rect 14982 -1799 15038 -1797
rect 15062 -1799 15118 -1797
rect 14822 -1851 14868 -1799
rect 14868 -1851 14878 -1799
rect 14902 -1851 14932 -1799
rect 14932 -1851 14944 -1799
rect 14944 -1851 14958 -1799
rect 14982 -1851 14996 -1799
rect 14996 -1851 15008 -1799
rect 15008 -1851 15038 -1799
rect 15062 -1851 15072 -1799
rect 15072 -1851 15118 -1799
rect 14822 -1853 14878 -1851
rect 14902 -1853 14958 -1851
rect 14982 -1853 15038 -1851
rect 15062 -1853 15118 -1851
rect 15223 -1799 15279 -1797
rect 15303 -1799 15359 -1797
rect 15383 -1799 15439 -1797
rect 15463 -1799 15519 -1797
rect 15223 -1851 15269 -1799
rect 15269 -1851 15279 -1799
rect 15303 -1851 15333 -1799
rect 15333 -1851 15345 -1799
rect 15345 -1851 15359 -1799
rect 15383 -1851 15397 -1799
rect 15397 -1851 15409 -1799
rect 15409 -1851 15439 -1799
rect 15463 -1851 15473 -1799
rect 15473 -1851 15519 -1799
rect 15223 -1853 15279 -1851
rect 15303 -1853 15359 -1851
rect 15383 -1853 15439 -1851
rect 15463 -1853 15519 -1851
rect 15662 -1799 15718 -1797
rect 15742 -1799 15798 -1797
rect 15662 -1851 15672 -1799
rect 15672 -1851 15718 -1799
rect 15742 -1851 15788 -1799
rect 15788 -1851 15798 -1799
rect 15662 -1853 15718 -1851
rect 15742 -1853 15798 -1851
rect 14543 -1999 14599 -1997
rect 14623 -1999 14679 -1997
rect 14543 -2051 14553 -1999
rect 14553 -2051 14599 -1999
rect 14623 -2051 14669 -1999
rect 14669 -2051 14679 -1999
rect 14543 -2053 14599 -2051
rect 14623 -2053 14679 -2051
rect 14822 -1999 14878 -1997
rect 14902 -1999 14958 -1997
rect 14982 -1999 15038 -1997
rect 15062 -1999 15118 -1997
rect 14822 -2051 14868 -1999
rect 14868 -2051 14878 -1999
rect 14902 -2051 14932 -1999
rect 14932 -2051 14944 -1999
rect 14944 -2051 14958 -1999
rect 14982 -2051 14996 -1999
rect 14996 -2051 15008 -1999
rect 15008 -2051 15038 -1999
rect 15062 -2051 15072 -1999
rect 15072 -2051 15118 -1999
rect 14822 -2053 14878 -2051
rect 14902 -2053 14958 -2051
rect 14982 -2053 15038 -2051
rect 15062 -2053 15118 -2051
rect 15223 -1999 15279 -1997
rect 15303 -1999 15359 -1997
rect 15383 -1999 15439 -1997
rect 15463 -1999 15519 -1997
rect 15223 -2051 15269 -1999
rect 15269 -2051 15279 -1999
rect 15303 -2051 15333 -1999
rect 15333 -2051 15345 -1999
rect 15345 -2051 15359 -1999
rect 15383 -2051 15397 -1999
rect 15397 -2051 15409 -1999
rect 15409 -2051 15439 -1999
rect 15463 -2051 15473 -1999
rect 15473 -2051 15519 -1999
rect 15223 -2053 15279 -2051
rect 15303 -2053 15359 -2051
rect 15383 -2053 15439 -2051
rect 15463 -2053 15519 -2051
rect 15662 -1999 15718 -1997
rect 15742 -1999 15798 -1997
rect 15662 -2051 15672 -1999
rect 15672 -2051 15718 -1999
rect 15742 -2051 15788 -1999
rect 15788 -2051 15798 -1999
rect 15662 -2053 15718 -2051
rect 15742 -2053 15798 -2051
<< metal3 >>
rect 0 4905 70 5070
rect 0 4849 7 4905
rect 63 4849 70 4905
rect 0 3695 70 4849
rect 0 3639 7 3695
rect 63 3639 70 3695
rect 0 2485 70 3639
rect 0 2429 7 2485
rect 63 2429 70 2485
rect 0 1275 70 2429
rect 0 1219 7 1275
rect 63 1219 70 1275
rect 0 65 70 1219
rect 0 9 7 65
rect 63 9 70 65
rect 0 -16 70 9
rect 0 -72 7 -16
rect 63 -72 70 -16
rect 0 -77 70 -72
rect 200 4921 270 5070
rect 200 4865 207 4921
rect 263 4865 270 4921
rect 200 3711 270 4865
rect 200 3655 207 3711
rect 263 3655 270 3711
rect 200 2501 270 3655
rect 200 2445 207 2501
rect 263 2445 270 2501
rect 200 1291 270 2445
rect 200 1235 207 1291
rect 263 1235 270 1291
rect 200 81 270 1235
rect 200 25 207 81
rect 263 25 270 81
rect 200 -16 270 25
rect 200 -72 207 -16
rect 263 -72 270 -16
rect 200 -77 270 -72
rect 400 4905 470 5070
rect 400 4849 407 4905
rect 463 4849 470 4905
rect 400 3695 470 4849
rect 400 3639 407 3695
rect 463 3639 470 3695
rect 400 2485 470 3639
rect 400 2429 407 2485
rect 463 2429 470 2485
rect 400 1275 470 2429
rect 400 1219 407 1275
rect 463 1219 470 1275
rect 400 65 470 1219
rect 400 9 407 65
rect 463 9 470 65
rect 400 -16 470 9
rect 400 -72 407 -16
rect 463 -72 470 -16
rect 400 -77 470 -72
rect 600 4921 670 5070
rect 600 4865 607 4921
rect 663 4865 670 4921
rect 600 3711 670 4865
rect 600 3655 607 3711
rect 663 3655 670 3711
rect 600 2501 670 3655
rect 600 2445 607 2501
rect 663 2445 670 2501
rect 600 1291 670 2445
rect 600 1235 607 1291
rect 663 1235 670 1291
rect 600 81 670 1235
rect 600 25 607 81
rect 663 25 670 81
rect 600 -16 670 25
rect 600 -72 607 -16
rect 663 -72 670 -16
rect 600 -77 670 -72
rect 800 4905 870 5070
rect 800 4849 807 4905
rect 863 4849 870 4905
rect 800 3695 870 4849
rect 800 3639 807 3695
rect 863 3639 870 3695
rect 800 2485 870 3639
rect 800 2429 807 2485
rect 863 2429 870 2485
rect 800 1275 870 2429
rect 800 1219 807 1275
rect 863 1219 870 1275
rect 800 65 870 1219
rect 800 9 807 65
rect 863 9 870 65
rect 800 -16 870 9
rect 800 -72 807 -16
rect 863 -72 870 -16
rect 800 -77 870 -72
rect 1000 4921 1070 5070
rect 1000 4865 1007 4921
rect 1063 4865 1070 4921
rect 1000 3711 1070 4865
rect 1000 3655 1007 3711
rect 1063 3655 1070 3711
rect 1000 2501 1070 3655
rect 1000 2445 1007 2501
rect 1063 2445 1070 2501
rect 1000 1291 1070 2445
rect 1000 1235 1007 1291
rect 1063 1235 1070 1291
rect 1000 81 1070 1235
rect 1000 25 1007 81
rect 1063 25 1070 81
rect 1000 -16 1070 25
rect 1000 -72 1007 -16
rect 1063 -72 1070 -16
rect 1000 -77 1070 -72
rect 1200 4905 1270 5070
rect 1200 4849 1207 4905
rect 1263 4849 1270 4905
rect 1200 3695 1270 4849
rect 1200 3639 1207 3695
rect 1263 3639 1270 3695
rect 1200 2485 1270 3639
rect 1200 2429 1207 2485
rect 1263 2429 1270 2485
rect 1200 1275 1270 2429
rect 1200 1219 1207 1275
rect 1263 1219 1270 1275
rect 1200 65 1270 1219
rect 1200 9 1207 65
rect 1263 9 1270 65
rect 1200 -16 1270 9
rect 1200 -72 1207 -16
rect 1263 -72 1270 -16
rect 1200 -77 1270 -72
rect 1400 4921 1470 5070
rect 1400 4865 1407 4921
rect 1463 4865 1470 4921
rect 1400 3711 1470 4865
rect 1400 3655 1407 3711
rect 1463 3655 1470 3711
rect 1400 2501 1470 3655
rect 1400 2445 1407 2501
rect 1463 2445 1470 2501
rect 1400 1291 1470 2445
rect 1400 1235 1407 1291
rect 1463 1235 1470 1291
rect 1400 81 1470 1235
rect 1400 25 1407 81
rect 1463 25 1470 81
rect 1400 -16 1470 25
rect 1400 -72 1407 -16
rect 1463 -72 1470 -16
rect 1400 -77 1470 -72
rect 1600 4905 1670 5070
rect 1600 4849 1607 4905
rect 1663 4849 1670 4905
rect 1600 3695 1670 4849
rect 1600 3639 1607 3695
rect 1663 3639 1670 3695
rect 1600 2485 1670 3639
rect 1600 2429 1607 2485
rect 1663 2429 1670 2485
rect 1600 1275 1670 2429
rect 1600 1219 1607 1275
rect 1663 1219 1670 1275
rect 1600 65 1670 1219
rect 1600 9 1607 65
rect 1663 9 1670 65
rect 1600 -16 1670 9
rect 1600 -72 1607 -16
rect 1663 -72 1670 -16
rect 1600 -77 1670 -72
rect 1800 4921 1870 5070
rect 1800 4865 1807 4921
rect 1863 4865 1870 4921
rect 1800 3711 1870 4865
rect 1800 3655 1807 3711
rect 1863 3655 1870 3711
rect 1800 2501 1870 3655
rect 1800 2445 1807 2501
rect 1863 2445 1870 2501
rect 1800 1291 1870 2445
rect 1800 1235 1807 1291
rect 1863 1235 1870 1291
rect 1800 81 1870 1235
rect 1800 25 1807 81
rect 1863 25 1870 81
rect 1800 -16 1870 25
rect 1800 -72 1807 -16
rect 1863 -72 1870 -16
rect 1800 -77 1870 -72
rect 2000 4905 2070 5070
rect 2000 4849 2007 4905
rect 2063 4849 2070 4905
rect 2000 3695 2070 4849
rect 2000 3639 2007 3695
rect 2063 3639 2070 3695
rect 2000 2485 2070 3639
rect 2000 2429 2007 2485
rect 2063 2429 2070 2485
rect 2000 1275 2070 2429
rect 2000 1219 2007 1275
rect 2063 1219 2070 1275
rect 2000 65 2070 1219
rect 2000 9 2007 65
rect 2063 9 2070 65
rect 2000 -16 2070 9
rect 2000 -72 2007 -16
rect 2063 -72 2070 -16
rect 2000 -77 2070 -72
rect 2200 4921 2270 5070
rect 2200 4865 2207 4921
rect 2263 4865 2270 4921
rect 2200 3711 2270 4865
rect 2200 3655 2207 3711
rect 2263 3655 2270 3711
rect 2200 2501 2270 3655
rect 2200 2445 2207 2501
rect 2263 2445 2270 2501
rect 2200 1291 2270 2445
rect 2200 1235 2207 1291
rect 2263 1235 2270 1291
rect 2200 81 2270 1235
rect 2200 25 2207 81
rect 2263 25 2270 81
rect 2200 -16 2270 25
rect 2200 -72 2207 -16
rect 2263 -72 2270 -16
rect 2200 -77 2270 -72
rect 2400 4905 2470 5070
rect 2400 4849 2407 4905
rect 2463 4849 2470 4905
rect 2400 3695 2470 4849
rect 2400 3639 2407 3695
rect 2463 3639 2470 3695
rect 2400 2485 2470 3639
rect 2400 2429 2407 2485
rect 2463 2429 2470 2485
rect 2400 1275 2470 2429
rect 2400 1219 2407 1275
rect 2463 1219 2470 1275
rect 2400 65 2470 1219
rect 2400 9 2407 65
rect 2463 9 2470 65
rect 2400 -16 2470 9
rect 2400 -72 2407 -16
rect 2463 -72 2470 -16
rect 2400 -77 2470 -72
rect 2600 4921 2670 5070
rect 2600 4865 2607 4921
rect 2663 4865 2670 4921
rect 2600 3711 2670 4865
rect 2600 3655 2607 3711
rect 2663 3655 2670 3711
rect 2600 2501 2670 3655
rect 2600 2445 2607 2501
rect 2663 2445 2670 2501
rect 2600 1291 2670 2445
rect 2600 1235 2607 1291
rect 2663 1235 2670 1291
rect 2600 81 2670 1235
rect 2600 25 2607 81
rect 2663 25 2670 81
rect 2600 -16 2670 25
rect 2600 -72 2607 -16
rect 2663 -72 2670 -16
rect 2600 -77 2670 -72
rect 2800 4905 2870 5070
rect 2800 4849 2807 4905
rect 2863 4849 2870 4905
rect 2800 3695 2870 4849
rect 2800 3639 2807 3695
rect 2863 3639 2870 3695
rect 2800 2485 2870 3639
rect 2800 2429 2807 2485
rect 2863 2429 2870 2485
rect 2800 1275 2870 2429
rect 2800 1219 2807 1275
rect 2863 1219 2870 1275
rect 2800 65 2870 1219
rect 2800 9 2807 65
rect 2863 9 2870 65
rect 2800 -16 2870 9
rect 2800 -72 2807 -16
rect 2863 -72 2870 -16
rect 2800 -77 2870 -72
rect 3000 4921 3070 5070
rect 3000 4865 3007 4921
rect 3063 4865 3070 4921
rect 3000 3711 3070 4865
rect 3000 3655 3007 3711
rect 3063 3655 3070 3711
rect 3000 2501 3070 3655
rect 3000 2445 3007 2501
rect 3063 2445 3070 2501
rect 3000 1291 3070 2445
rect 3000 1235 3007 1291
rect 3063 1235 3070 1291
rect 3000 81 3070 1235
rect 3000 25 3007 81
rect 3063 25 3070 81
rect 3000 -16 3070 25
rect 3000 -72 3007 -16
rect 3063 -72 3070 -16
rect 3000 -77 3070 -72
rect 3200 4905 3270 5070
rect 3200 4849 3207 4905
rect 3263 4849 3270 4905
rect 3200 3695 3270 4849
rect 3200 3639 3207 3695
rect 3263 3639 3270 3695
rect 3200 2485 3270 3639
rect 3200 2429 3207 2485
rect 3263 2429 3270 2485
rect 3200 1275 3270 2429
rect 3200 1219 3207 1275
rect 3263 1219 3270 1275
rect 3200 65 3270 1219
rect 3200 9 3207 65
rect 3263 9 3270 65
rect 3200 -16 3270 9
rect 3200 -72 3207 -16
rect 3263 -72 3270 -16
rect 3200 -77 3270 -72
rect 3400 4921 3470 5070
rect 3400 4865 3407 4921
rect 3463 4865 3470 4921
rect 3400 3711 3470 4865
rect 3400 3655 3407 3711
rect 3463 3655 3470 3711
rect 3400 2501 3470 3655
rect 3400 2445 3407 2501
rect 3463 2445 3470 2501
rect 3400 1291 3470 2445
rect 3400 1235 3407 1291
rect 3463 1235 3470 1291
rect 3400 81 3470 1235
rect 3400 25 3407 81
rect 3463 25 3470 81
rect 3400 -16 3470 25
rect 3400 -72 3407 -16
rect 3463 -72 3470 -16
rect 3400 -77 3470 -72
rect 3600 4905 3670 5070
rect 3600 4849 3607 4905
rect 3663 4849 3670 4905
rect 3600 3695 3670 4849
rect 3600 3639 3607 3695
rect 3663 3639 3670 3695
rect 3600 2485 3670 3639
rect 3600 2429 3607 2485
rect 3663 2429 3670 2485
rect 3600 1275 3670 2429
rect 3600 1219 3607 1275
rect 3663 1219 3670 1275
rect 3600 65 3670 1219
rect 3600 9 3607 65
rect 3663 9 3670 65
rect 3600 -16 3670 9
rect 3600 -72 3607 -16
rect 3663 -72 3670 -16
rect 3600 -77 3670 -72
rect 3800 4921 3870 5070
rect 3800 4865 3807 4921
rect 3863 4865 3870 4921
rect 3800 3711 3870 4865
rect 3800 3655 3807 3711
rect 3863 3655 3870 3711
rect 3800 2501 3870 3655
rect 3800 2445 3807 2501
rect 3863 2445 3870 2501
rect 3800 1291 3870 2445
rect 3800 1235 3807 1291
rect 3863 1235 3870 1291
rect 3800 81 3870 1235
rect 3800 25 3807 81
rect 3863 25 3870 81
rect 3800 -16 3870 25
rect 3800 -72 3807 -16
rect 3863 -72 3870 -16
rect 3800 -77 3870 -72
rect 4000 4905 4070 5070
rect 4000 4849 4007 4905
rect 4063 4849 4070 4905
rect 4000 3695 4070 4849
rect 4000 3639 4007 3695
rect 4063 3639 4070 3695
rect 4000 2485 4070 3639
rect 4000 2429 4007 2485
rect 4063 2429 4070 2485
rect 4000 1275 4070 2429
rect 4000 1219 4007 1275
rect 4063 1219 4070 1275
rect 4000 65 4070 1219
rect 4000 9 4007 65
rect 4063 9 4070 65
rect 4000 -16 4070 9
rect 4000 -72 4007 -16
rect 4063 -72 4070 -16
rect 4000 -77 4070 -72
rect 4200 4921 4270 5070
rect 4200 4865 4207 4921
rect 4263 4865 4270 4921
rect 4200 3711 4270 4865
rect 4200 3655 4207 3711
rect 4263 3655 4270 3711
rect 4200 2501 4270 3655
rect 4200 2445 4207 2501
rect 4263 2445 4270 2501
rect 4200 1291 4270 2445
rect 4200 1235 4207 1291
rect 4263 1235 4270 1291
rect 4200 81 4270 1235
rect 4200 25 4207 81
rect 4263 25 4270 81
rect 4200 -16 4270 25
rect 4200 -72 4207 -16
rect 4263 -72 4270 -16
rect 4200 -77 4270 -72
rect 4400 4905 4470 5070
rect 4400 4849 4407 4905
rect 4463 4849 4470 4905
rect 4400 3695 4470 4849
rect 4400 3639 4407 3695
rect 4463 3639 4470 3695
rect 4400 2485 4470 3639
rect 4400 2429 4407 2485
rect 4463 2429 4470 2485
rect 4400 1275 4470 2429
rect 4400 1219 4407 1275
rect 4463 1219 4470 1275
rect 4400 65 4470 1219
rect 4400 9 4407 65
rect 4463 9 4470 65
rect 4400 -16 4470 9
rect 4400 -72 4407 -16
rect 4463 -72 4470 -16
rect 4400 -77 4470 -72
rect 4600 4921 4670 5070
rect 4600 4865 4607 4921
rect 4663 4865 4670 4921
rect 4600 3711 4670 4865
rect 4600 3655 4607 3711
rect 4663 3655 4670 3711
rect 4600 2501 4670 3655
rect 4600 2445 4607 2501
rect 4663 2445 4670 2501
rect 4600 1291 4670 2445
rect 4600 1235 4607 1291
rect 4663 1235 4670 1291
rect 4600 81 4670 1235
rect 4600 25 4607 81
rect 4663 25 4670 81
rect 4600 -16 4670 25
rect 4600 -72 4607 -16
rect 4663 -72 4670 -16
rect 4600 -77 4670 -72
rect 4800 4905 4870 5070
rect 4800 4849 4807 4905
rect 4863 4849 4870 4905
rect 4800 3695 4870 4849
rect 4800 3639 4807 3695
rect 4863 3639 4870 3695
rect 4800 2485 4870 3639
rect 4800 2429 4807 2485
rect 4863 2429 4870 2485
rect 4800 1275 4870 2429
rect 4800 1219 4807 1275
rect 4863 1219 4870 1275
rect 4800 65 4870 1219
rect 4800 9 4807 65
rect 4863 9 4870 65
rect 4800 -16 4870 9
rect 4800 -72 4807 -16
rect 4863 -72 4870 -16
rect 4800 -77 4870 -72
rect 5000 4921 5070 5070
rect 5000 4865 5007 4921
rect 5063 4865 5070 4921
rect 5000 3711 5070 4865
rect 5000 3655 5007 3711
rect 5063 3655 5070 3711
rect 5000 2501 5070 3655
rect 5000 2445 5007 2501
rect 5063 2445 5070 2501
rect 5000 1291 5070 2445
rect 5000 1235 5007 1291
rect 5063 1235 5070 1291
rect 5000 81 5070 1235
rect 5000 25 5007 81
rect 5063 25 5070 81
rect 5000 -16 5070 25
rect 5000 -72 5007 -16
rect 5063 -72 5070 -16
rect 5000 -77 5070 -72
rect 5200 4905 5270 5070
rect 5200 4849 5207 4905
rect 5263 4849 5270 4905
rect 5200 3695 5270 4849
rect 5200 3639 5207 3695
rect 5263 3639 5270 3695
rect 5200 2485 5270 3639
rect 5200 2429 5207 2485
rect 5263 2429 5270 2485
rect 5200 1275 5270 2429
rect 5200 1219 5207 1275
rect 5263 1219 5270 1275
rect 5200 65 5270 1219
rect 5200 9 5207 65
rect 5263 9 5270 65
rect 5200 -16 5270 9
rect 5200 -72 5207 -16
rect 5263 -72 5270 -16
rect 5200 -77 5270 -72
rect 5400 4921 5470 5070
rect 5400 4865 5407 4921
rect 5463 4865 5470 4921
rect 5400 3711 5470 4865
rect 5400 3655 5407 3711
rect 5463 3655 5470 3711
rect 5400 2501 5470 3655
rect 5400 2445 5407 2501
rect 5463 2445 5470 2501
rect 5400 1291 5470 2445
rect 5400 1235 5407 1291
rect 5463 1235 5470 1291
rect 5400 81 5470 1235
rect 5400 25 5407 81
rect 5463 25 5470 81
rect 5400 -16 5470 25
rect 5400 -72 5407 -16
rect 5463 -72 5470 -16
rect 5400 -77 5470 -72
rect 5600 4905 5670 5070
rect 5600 4849 5607 4905
rect 5663 4849 5670 4905
rect 5600 3695 5670 4849
rect 5600 3639 5607 3695
rect 5663 3639 5670 3695
rect 5600 2485 5670 3639
rect 5600 2429 5607 2485
rect 5663 2429 5670 2485
rect 5600 1275 5670 2429
rect 5600 1219 5607 1275
rect 5663 1219 5670 1275
rect 5600 65 5670 1219
rect 5600 9 5607 65
rect 5663 9 5670 65
rect 5600 -16 5670 9
rect 5600 -72 5607 -16
rect 5663 -72 5670 -16
rect 5600 -77 5670 -72
rect 5800 4921 5870 5070
rect 5800 4865 5807 4921
rect 5863 4865 5870 4921
rect 5800 3711 5870 4865
rect 5800 3655 5807 3711
rect 5863 3655 5870 3711
rect 5800 2501 5870 3655
rect 5800 2445 5807 2501
rect 5863 2445 5870 2501
rect 5800 1291 5870 2445
rect 5800 1235 5807 1291
rect 5863 1235 5870 1291
rect 5800 81 5870 1235
rect 5800 25 5807 81
rect 5863 25 5870 81
rect 5800 -16 5870 25
rect 5800 -72 5807 -16
rect 5863 -72 5870 -16
rect 5800 -77 5870 -72
rect 6000 4905 6070 5070
rect 6000 4849 6007 4905
rect 6063 4849 6070 4905
rect 6000 3695 6070 4849
rect 6000 3639 6007 3695
rect 6063 3639 6070 3695
rect 6000 2485 6070 3639
rect 6000 2429 6007 2485
rect 6063 2429 6070 2485
rect 6000 1275 6070 2429
rect 6000 1219 6007 1275
rect 6063 1219 6070 1275
rect 6000 65 6070 1219
rect 6000 9 6007 65
rect 6063 9 6070 65
rect 6000 -16 6070 9
rect 6000 -72 6007 -16
rect 6063 -72 6070 -16
rect 6000 -77 6070 -72
rect 6200 4921 6270 5070
rect 6200 4865 6207 4921
rect 6263 4865 6270 4921
rect 6200 3711 6270 4865
rect 6200 3655 6207 3711
rect 6263 3655 6270 3711
rect 6200 2501 6270 3655
rect 6200 2445 6207 2501
rect 6263 2445 6270 2501
rect 6200 1291 6270 2445
rect 6200 1235 6207 1291
rect 6263 1235 6270 1291
rect 6200 81 6270 1235
rect 6200 25 6207 81
rect 6263 25 6270 81
rect 6200 -16 6270 25
rect 6200 -72 6207 -16
rect 6263 -72 6270 -16
rect 6200 -77 6270 -72
rect 6400 4905 6470 5070
rect 6400 4849 6407 4905
rect 6463 4849 6470 4905
rect 6400 3695 6470 4849
rect 6400 3639 6407 3695
rect 6463 3639 6470 3695
rect 6400 2485 6470 3639
rect 6400 2429 6407 2485
rect 6463 2429 6470 2485
rect 6400 1275 6470 2429
rect 6400 1219 6407 1275
rect 6463 1219 6470 1275
rect 6400 65 6470 1219
rect 6400 9 6407 65
rect 6463 9 6470 65
rect 6400 -16 6470 9
rect 6400 -72 6407 -16
rect 6463 -72 6470 -16
rect 6400 -77 6470 -72
rect 6600 4921 6670 5070
rect 6600 4865 6607 4921
rect 6663 4865 6670 4921
rect 6600 3711 6670 4865
rect 6600 3655 6607 3711
rect 6663 3655 6670 3711
rect 6600 2501 6670 3655
rect 6600 2445 6607 2501
rect 6663 2445 6670 2501
rect 6600 1291 6670 2445
rect 6600 1235 6607 1291
rect 6663 1235 6670 1291
rect 6600 81 6670 1235
rect 6600 25 6607 81
rect 6663 25 6670 81
rect 6600 -16 6670 25
rect 6600 -72 6607 -16
rect 6663 -72 6670 -16
rect 6600 -77 6670 -72
rect 6800 4905 6870 5070
rect 6800 4849 6807 4905
rect 6863 4849 6870 4905
rect 6800 3695 6870 4849
rect 6800 3639 6807 3695
rect 6863 3639 6870 3695
rect 6800 2485 6870 3639
rect 6800 2429 6807 2485
rect 6863 2429 6870 2485
rect 6800 1275 6870 2429
rect 6800 1219 6807 1275
rect 6863 1219 6870 1275
rect 6800 65 6870 1219
rect 6800 9 6807 65
rect 6863 9 6870 65
rect 6800 -16 6870 9
rect 6800 -72 6807 -16
rect 6863 -72 6870 -16
rect 6800 -77 6870 -72
rect 7000 4921 7070 5070
rect 7000 4865 7007 4921
rect 7063 4865 7070 4921
rect 7000 3711 7070 4865
rect 7000 3655 7007 3711
rect 7063 3655 7070 3711
rect 7000 2501 7070 3655
rect 7000 2445 7007 2501
rect 7063 2445 7070 2501
rect 7000 1291 7070 2445
rect 7000 1235 7007 1291
rect 7063 1235 7070 1291
rect 7000 81 7070 1235
rect 7000 25 7007 81
rect 7063 25 7070 81
rect 7000 -16 7070 25
rect 7000 -72 7007 -16
rect 7063 -72 7070 -16
rect 7000 -77 7070 -72
rect 7200 4905 7270 5070
rect 7200 4849 7207 4905
rect 7263 4849 7270 4905
rect 7200 3695 7270 4849
rect 7200 3639 7207 3695
rect 7263 3639 7270 3695
rect 7200 2485 7270 3639
rect 7200 2429 7207 2485
rect 7263 2429 7270 2485
rect 7200 1275 7270 2429
rect 7200 1219 7207 1275
rect 7263 1219 7270 1275
rect 7200 65 7270 1219
rect 7200 9 7207 65
rect 7263 9 7270 65
rect 7200 -16 7270 9
rect 7200 -72 7207 -16
rect 7263 -72 7270 -16
rect 7200 -77 7270 -72
rect 7400 4921 7470 5070
rect 7400 4865 7407 4921
rect 7463 4865 7470 4921
rect 7400 3711 7470 4865
rect 7400 3655 7407 3711
rect 7463 3655 7470 3711
rect 7400 2501 7470 3655
rect 7400 2445 7407 2501
rect 7463 2445 7470 2501
rect 7400 1291 7470 2445
rect 7400 1235 7407 1291
rect 7463 1235 7470 1291
rect 7400 81 7470 1235
rect 7400 25 7407 81
rect 7463 25 7470 81
rect 7400 -16 7470 25
rect 7400 -72 7407 -16
rect 7463 -72 7470 -16
rect 7400 -77 7470 -72
rect 7600 4905 7670 5070
rect 7600 4849 7607 4905
rect 7663 4849 7670 4905
rect 7600 3695 7670 4849
rect 7600 3639 7607 3695
rect 7663 3639 7670 3695
rect 7600 2485 7670 3639
rect 7600 2429 7607 2485
rect 7663 2429 7670 2485
rect 7600 1275 7670 2429
rect 7600 1219 7607 1275
rect 7663 1219 7670 1275
rect 7600 65 7670 1219
rect 7600 9 7607 65
rect 7663 9 7670 65
rect 7600 -16 7670 9
rect 7600 -72 7607 -16
rect 7663 -72 7670 -16
rect 7600 -77 7670 -72
rect 7800 4921 7870 5070
rect 7800 4865 7807 4921
rect 7863 4865 7870 4921
rect 7800 3711 7870 4865
rect 7800 3655 7807 3711
rect 7863 3655 7870 3711
rect 7800 2501 7870 3655
rect 7800 2445 7807 2501
rect 7863 2445 7870 2501
rect 7800 1291 7870 2445
rect 7800 1235 7807 1291
rect 7863 1235 7870 1291
rect 7800 81 7870 1235
rect 7800 25 7807 81
rect 7863 25 7870 81
rect 7800 -16 7870 25
rect 7800 -72 7807 -16
rect 7863 -72 7870 -16
rect 7800 -77 7870 -72
rect 8000 4905 8070 5070
rect 8000 4849 8007 4905
rect 8063 4849 8070 4905
rect 8000 3695 8070 4849
rect 8000 3639 8007 3695
rect 8063 3639 8070 3695
rect 8000 2485 8070 3639
rect 8000 2429 8007 2485
rect 8063 2429 8070 2485
rect 8000 1275 8070 2429
rect 8000 1219 8007 1275
rect 8063 1219 8070 1275
rect 8000 65 8070 1219
rect 8000 9 8007 65
rect 8063 9 8070 65
rect 8000 -16 8070 9
rect 8000 -72 8007 -16
rect 8063 -72 8070 -16
rect 8000 -77 8070 -72
rect 8200 4921 8270 5070
rect 8200 4865 8207 4921
rect 8263 4865 8270 4921
rect 8200 3711 8270 4865
rect 8200 3655 8207 3711
rect 8263 3655 8270 3711
rect 8200 2501 8270 3655
rect 8200 2445 8207 2501
rect 8263 2445 8270 2501
rect 8200 1291 8270 2445
rect 8200 1235 8207 1291
rect 8263 1235 8270 1291
rect 8200 81 8270 1235
rect 8200 25 8207 81
rect 8263 25 8270 81
rect 8200 -16 8270 25
rect 8200 -72 8207 -16
rect 8263 -72 8270 -16
rect 8200 -77 8270 -72
rect 8400 4905 8470 5070
rect 8400 4849 8407 4905
rect 8463 4849 8470 4905
rect 8400 3695 8470 4849
rect 8400 3639 8407 3695
rect 8463 3639 8470 3695
rect 8400 2485 8470 3639
rect 8400 2429 8407 2485
rect 8463 2429 8470 2485
rect 8400 1275 8470 2429
rect 8400 1219 8407 1275
rect 8463 1219 8470 1275
rect 8400 65 8470 1219
rect 8400 9 8407 65
rect 8463 9 8470 65
rect 8400 -16 8470 9
rect 8400 -72 8407 -16
rect 8463 -72 8470 -16
rect 8400 -77 8470 -72
rect 8600 4921 8670 5070
rect 8600 4865 8607 4921
rect 8663 4865 8670 4921
rect 8600 3711 8670 4865
rect 8600 3655 8607 3711
rect 8663 3655 8670 3711
rect 8600 2501 8670 3655
rect 8600 2445 8607 2501
rect 8663 2445 8670 2501
rect 8600 1291 8670 2445
rect 8600 1235 8607 1291
rect 8663 1235 8670 1291
rect 8600 81 8670 1235
rect 8600 25 8607 81
rect 8663 25 8670 81
rect 8600 -16 8670 25
rect 8600 -72 8607 -16
rect 8663 -72 8670 -16
rect 8600 -77 8670 -72
rect 8800 4905 8870 5070
rect 8800 4849 8807 4905
rect 8863 4849 8870 4905
rect 8800 3695 8870 4849
rect 8800 3639 8807 3695
rect 8863 3639 8870 3695
rect 8800 2485 8870 3639
rect 8800 2429 8807 2485
rect 8863 2429 8870 2485
rect 8800 1275 8870 2429
rect 8800 1219 8807 1275
rect 8863 1219 8870 1275
rect 8800 65 8870 1219
rect 8800 9 8807 65
rect 8863 9 8870 65
rect 8800 -16 8870 9
rect 8800 -72 8807 -16
rect 8863 -72 8870 -16
rect 8800 -77 8870 -72
rect 9000 4921 9070 5070
rect 9000 4865 9007 4921
rect 9063 4865 9070 4921
rect 9000 3711 9070 4865
rect 9000 3655 9007 3711
rect 9063 3655 9070 3711
rect 9000 2501 9070 3655
rect 9000 2445 9007 2501
rect 9063 2445 9070 2501
rect 9000 1291 9070 2445
rect 9000 1235 9007 1291
rect 9063 1235 9070 1291
rect 9000 81 9070 1235
rect 9000 25 9007 81
rect 9063 25 9070 81
rect 9000 -16 9070 25
rect 9000 -72 9007 -16
rect 9063 -72 9070 -16
rect 9000 -77 9070 -72
rect 9200 4905 9270 5070
rect 9200 4849 9207 4905
rect 9263 4849 9270 4905
rect 9200 3695 9270 4849
rect 9200 3639 9207 3695
rect 9263 3639 9270 3695
rect 9200 2485 9270 3639
rect 9200 2429 9207 2485
rect 9263 2429 9270 2485
rect 9200 1275 9270 2429
rect 9200 1219 9207 1275
rect 9263 1219 9270 1275
rect 9200 65 9270 1219
rect 9200 9 9207 65
rect 9263 9 9270 65
rect 9200 -16 9270 9
rect 9200 -72 9207 -16
rect 9263 -72 9270 -16
rect 9200 -77 9270 -72
rect 9400 4921 9470 5070
rect 9400 4865 9407 4921
rect 9463 4865 9470 4921
rect 9400 3711 9470 4865
rect 9400 3655 9407 3711
rect 9463 3655 9470 3711
rect 9400 2501 9470 3655
rect 9400 2445 9407 2501
rect 9463 2445 9470 2501
rect 9400 1291 9470 2445
rect 9400 1235 9407 1291
rect 9463 1235 9470 1291
rect 9400 81 9470 1235
rect 9400 25 9407 81
rect 9463 25 9470 81
rect 9400 -16 9470 25
rect 9400 -72 9407 -16
rect 9463 -72 9470 -16
rect 9400 -77 9470 -72
rect 9600 4905 9670 5070
rect 9600 4849 9607 4905
rect 9663 4849 9670 4905
rect 9600 3695 9670 4849
rect 9600 3639 9607 3695
rect 9663 3639 9670 3695
rect 9600 2485 9670 3639
rect 9600 2429 9607 2485
rect 9663 2429 9670 2485
rect 9600 1275 9670 2429
rect 9600 1219 9607 1275
rect 9663 1219 9670 1275
rect 9600 65 9670 1219
rect 9600 9 9607 65
rect 9663 9 9670 65
rect 9600 -16 9670 9
rect 9600 -72 9607 -16
rect 9663 -72 9670 -16
rect 9600 -77 9670 -72
rect 9800 4921 9870 5070
rect 9800 4865 9807 4921
rect 9863 4865 9870 4921
rect 9800 3711 9870 4865
rect 9800 3655 9807 3711
rect 9863 3655 9870 3711
rect 9800 2501 9870 3655
rect 9800 2445 9807 2501
rect 9863 2445 9870 2501
rect 9800 1291 9870 2445
rect 9800 1235 9807 1291
rect 9863 1235 9870 1291
rect 9800 81 9870 1235
rect 9800 25 9807 81
rect 9863 25 9870 81
rect 9800 -16 9870 25
rect 9800 -72 9807 -16
rect 9863 -72 9870 -16
rect 9800 -77 9870 -72
rect 10000 4905 10070 5070
rect 10000 4849 10007 4905
rect 10063 4849 10070 4905
rect 10000 3695 10070 4849
rect 10000 3639 10007 3695
rect 10063 3639 10070 3695
rect 10000 2485 10070 3639
rect 10000 2429 10007 2485
rect 10063 2429 10070 2485
rect 10000 1275 10070 2429
rect 10000 1219 10007 1275
rect 10063 1219 10070 1275
rect 10000 65 10070 1219
rect 10000 9 10007 65
rect 10063 9 10070 65
rect 10000 -16 10070 9
rect 10000 -72 10007 -16
rect 10063 -72 10070 -16
rect 10000 -77 10070 -72
rect 10200 4921 10270 5070
rect 10200 4865 10207 4921
rect 10263 4865 10270 4921
rect 10200 3711 10270 4865
rect 10200 3655 10207 3711
rect 10263 3655 10270 3711
rect 10200 2501 10270 3655
rect 10200 2445 10207 2501
rect 10263 2445 10270 2501
rect 10200 1291 10270 2445
rect 10200 1235 10207 1291
rect 10263 1235 10270 1291
rect 10200 81 10270 1235
rect 10200 25 10207 81
rect 10263 25 10270 81
rect 10200 -16 10270 25
rect 10200 -72 10207 -16
rect 10263 -72 10270 -16
rect 10200 -77 10270 -72
rect 10400 4905 10470 5070
rect 10400 4849 10407 4905
rect 10463 4849 10470 4905
rect 10400 3695 10470 4849
rect 10400 3639 10407 3695
rect 10463 3639 10470 3695
rect 10400 2485 10470 3639
rect 10400 2429 10407 2485
rect 10463 2429 10470 2485
rect 10400 1275 10470 2429
rect 10400 1219 10407 1275
rect 10463 1219 10470 1275
rect 10400 65 10470 1219
rect 10400 9 10407 65
rect 10463 9 10470 65
rect 10400 -16 10470 9
rect 10400 -72 10407 -16
rect 10463 -72 10470 -16
rect 10400 -77 10470 -72
rect 10600 4921 10670 5070
rect 10600 4865 10607 4921
rect 10663 4865 10670 4921
rect 10600 3711 10670 4865
rect 10600 3655 10607 3711
rect 10663 3655 10670 3711
rect 10600 2501 10670 3655
rect 10600 2445 10607 2501
rect 10663 2445 10670 2501
rect 10600 1291 10670 2445
rect 10600 1235 10607 1291
rect 10663 1235 10670 1291
rect 10600 81 10670 1235
rect 10600 25 10607 81
rect 10663 25 10670 81
rect 10600 -16 10670 25
rect 10600 -72 10607 -16
rect 10663 -72 10670 -16
rect 10600 -77 10670 -72
rect 10800 4905 10870 5070
rect 10800 4849 10807 4905
rect 10863 4849 10870 4905
rect 10800 3695 10870 4849
rect 10800 3639 10807 3695
rect 10863 3639 10870 3695
rect 10800 2485 10870 3639
rect 10800 2429 10807 2485
rect 10863 2429 10870 2485
rect 10800 1275 10870 2429
rect 10800 1219 10807 1275
rect 10863 1219 10870 1275
rect 10800 65 10870 1219
rect 10800 9 10807 65
rect 10863 9 10870 65
rect 10800 -16 10870 9
rect 10800 -72 10807 -16
rect 10863 -72 10870 -16
rect 10800 -77 10870 -72
rect 11000 4921 11070 5070
rect 11000 4865 11007 4921
rect 11063 4865 11070 4921
rect 11000 3711 11070 4865
rect 11000 3655 11007 3711
rect 11063 3655 11070 3711
rect 11000 2501 11070 3655
rect 11000 2445 11007 2501
rect 11063 2445 11070 2501
rect 11000 1291 11070 2445
rect 11000 1235 11007 1291
rect 11063 1235 11070 1291
rect 11000 81 11070 1235
rect 11000 25 11007 81
rect 11063 25 11070 81
rect 11000 -16 11070 25
rect 11000 -72 11007 -16
rect 11063 -72 11070 -16
rect 11000 -77 11070 -72
rect 11200 4905 11270 5070
rect 11200 4849 11207 4905
rect 11263 4849 11270 4905
rect 11200 3695 11270 4849
rect 11200 3639 11207 3695
rect 11263 3639 11270 3695
rect 11200 2485 11270 3639
rect 11200 2429 11207 2485
rect 11263 2429 11270 2485
rect 11200 1275 11270 2429
rect 11200 1219 11207 1275
rect 11263 1219 11270 1275
rect 11200 65 11270 1219
rect 11200 9 11207 65
rect 11263 9 11270 65
rect 11200 -16 11270 9
rect 11200 -72 11207 -16
rect 11263 -72 11270 -16
rect 11200 -77 11270 -72
rect 11400 4921 11470 5070
rect 11400 4865 11407 4921
rect 11463 4865 11470 4921
rect 11400 3711 11470 4865
rect 11400 3655 11407 3711
rect 11463 3655 11470 3711
rect 11400 2501 11470 3655
rect 11400 2445 11407 2501
rect 11463 2445 11470 2501
rect 11400 1291 11470 2445
rect 11400 1235 11407 1291
rect 11463 1235 11470 1291
rect 11400 81 11470 1235
rect 11400 25 11407 81
rect 11463 25 11470 81
rect 11400 -16 11470 25
rect 11400 -72 11407 -16
rect 11463 -72 11470 -16
rect 11400 -77 11470 -72
rect 11600 4905 11670 5070
rect 11600 4849 11607 4905
rect 11663 4849 11670 4905
rect 11600 3695 11670 4849
rect 11600 3639 11607 3695
rect 11663 3639 11670 3695
rect 11600 2485 11670 3639
rect 11600 2429 11607 2485
rect 11663 2429 11670 2485
rect 11600 1275 11670 2429
rect 11600 1219 11607 1275
rect 11663 1219 11670 1275
rect 11600 65 11670 1219
rect 11600 9 11607 65
rect 11663 9 11670 65
rect 11600 -16 11670 9
rect 11600 -72 11607 -16
rect 11663 -72 11670 -16
rect 11600 -77 11670 -72
rect 11800 4921 11870 5070
rect 11800 4865 11807 4921
rect 11863 4865 11870 4921
rect 11800 3711 11870 4865
rect 11800 3655 11807 3711
rect 11863 3655 11870 3711
rect 11800 2501 11870 3655
rect 11800 2445 11807 2501
rect 11863 2445 11870 2501
rect 11800 1291 11870 2445
rect 11800 1235 11807 1291
rect 11863 1235 11870 1291
rect 11800 81 11870 1235
rect 11800 25 11807 81
rect 11863 25 11870 81
rect 11800 -16 11870 25
rect 11800 -72 11807 -16
rect 11863 -72 11870 -16
rect 11800 -77 11870 -72
rect 12000 4905 12070 5070
rect 12000 4849 12007 4905
rect 12063 4849 12070 4905
rect 12000 3695 12070 4849
rect 12000 3639 12007 3695
rect 12063 3639 12070 3695
rect 12000 2485 12070 3639
rect 12000 2429 12007 2485
rect 12063 2429 12070 2485
rect 12000 1275 12070 2429
rect 12000 1219 12007 1275
rect 12063 1219 12070 1275
rect 12000 65 12070 1219
rect 12000 9 12007 65
rect 12063 9 12070 65
rect 12000 -16 12070 9
rect 12000 -72 12007 -16
rect 12063 -72 12070 -16
rect 12000 -77 12070 -72
rect 12200 4921 12270 5070
rect 12200 4865 12207 4921
rect 12263 4865 12270 4921
rect 12200 3711 12270 4865
rect 12200 3655 12207 3711
rect 12263 3655 12270 3711
rect 12200 2501 12270 3655
rect 12200 2445 12207 2501
rect 12263 2445 12270 2501
rect 12200 1291 12270 2445
rect 12200 1235 12207 1291
rect 12263 1235 12270 1291
rect 12200 81 12270 1235
rect 12200 25 12207 81
rect 12263 25 12270 81
rect 12200 -16 12270 25
rect 12200 -72 12207 -16
rect 12263 -72 12270 -16
rect 12200 -77 12270 -72
rect 12400 4905 12470 5070
rect 12400 4849 12407 4905
rect 12463 4849 12470 4905
rect 12400 3695 12470 4849
rect 12400 3639 12407 3695
rect 12463 3639 12470 3695
rect 12400 2485 12470 3639
rect 12400 2429 12407 2485
rect 12463 2429 12470 2485
rect 12400 1275 12470 2429
rect 12400 1219 12407 1275
rect 12463 1219 12470 1275
rect 12400 65 12470 1219
rect 12400 9 12407 65
rect 12463 9 12470 65
rect 12400 -16 12470 9
rect 12400 -72 12407 -16
rect 12463 -72 12470 -16
rect 12400 -77 12470 -72
rect 12600 4921 12670 5070
rect 12600 4865 12607 4921
rect 12663 4865 12670 4921
rect 12600 3711 12670 4865
rect 12600 3655 12607 3711
rect 12663 3655 12670 3711
rect 12600 2501 12670 3655
rect 12600 2445 12607 2501
rect 12663 2445 12670 2501
rect 12600 1291 12670 2445
rect 12600 1235 12607 1291
rect 12663 1235 12670 1291
rect 12600 81 12670 1235
rect 12600 25 12607 81
rect 12663 25 12670 81
rect 12600 -16 12670 25
rect 12600 -72 12607 -16
rect 12663 -72 12670 -16
rect 12600 -77 12670 -72
rect -138 -145 12808 -140
rect -138 -201 -133 -145
rect -77 -201 -53 -145
rect 3 -201 67 -145
rect 123 -201 147 -145
rect 203 -201 267 -145
rect 323 -201 347 -145
rect 403 -201 467 -145
rect 523 -201 547 -145
rect 603 -201 667 -145
rect 723 -201 747 -145
rect 803 -201 867 -145
rect 923 -201 947 -145
rect 1003 -201 1067 -145
rect 1123 -201 1147 -145
rect 1203 -201 1267 -145
rect 1323 -201 1347 -145
rect 1403 -201 1467 -145
rect 1523 -201 1547 -145
rect 1603 -201 1667 -145
rect 1723 -201 1747 -145
rect 1803 -201 1867 -145
rect 1923 -201 1947 -145
rect 2003 -201 2067 -145
rect 2123 -201 2147 -145
rect 2203 -201 2267 -145
rect 2323 -201 2347 -145
rect 2403 -201 2467 -145
rect 2523 -201 2547 -145
rect 2603 -201 2667 -145
rect 2723 -201 2747 -145
rect 2803 -201 2867 -145
rect 2923 -201 2947 -145
rect 3003 -201 3067 -145
rect 3123 -201 3147 -145
rect 3203 -201 3267 -145
rect 3323 -201 3347 -145
rect 3403 -201 3467 -145
rect 3523 -201 3547 -145
rect 3603 -201 3667 -145
rect 3723 -201 3747 -145
rect 3803 -201 3867 -145
rect 3923 -201 3947 -145
rect 4003 -201 4067 -145
rect 4123 -201 4147 -145
rect 4203 -201 4267 -145
rect 4323 -201 4347 -145
rect 4403 -201 4467 -145
rect 4523 -201 4547 -145
rect 4603 -201 4667 -145
rect 4723 -201 4747 -145
rect 4803 -201 4867 -145
rect 4923 -201 4947 -145
rect 5003 -201 5067 -145
rect 5123 -201 5147 -145
rect 5203 -201 5267 -145
rect 5323 -201 5347 -145
rect 5403 -201 5467 -145
rect 5523 -201 5547 -145
rect 5603 -201 5667 -145
rect 5723 -201 5747 -145
rect 5803 -201 5867 -145
rect 5923 -201 5947 -145
rect 6003 -201 6067 -145
rect 6123 -201 6147 -145
rect 6203 -201 6267 -145
rect 6323 -201 6347 -145
rect 6403 -201 6467 -145
rect 6523 -201 6547 -145
rect 6603 -201 6667 -145
rect 6723 -201 6747 -145
rect 6803 -201 6867 -145
rect 6923 -201 6947 -145
rect 7003 -201 7067 -145
rect 7123 -201 7147 -145
rect 7203 -201 7267 -145
rect 7323 -201 7347 -145
rect 7403 -201 7467 -145
rect 7523 -201 7547 -145
rect 7603 -201 7667 -145
rect 7723 -201 7747 -145
rect 7803 -201 7867 -145
rect 7923 -201 7947 -145
rect 8003 -201 8067 -145
rect 8123 -201 8147 -145
rect 8203 -201 8267 -145
rect 8323 -201 8347 -145
rect 8403 -201 8467 -145
rect 8523 -201 8547 -145
rect 8603 -201 8667 -145
rect 8723 -201 8747 -145
rect 8803 -201 8867 -145
rect 8923 -201 8947 -145
rect 9003 -201 9067 -145
rect 9123 -201 9147 -145
rect 9203 -201 9267 -145
rect 9323 -201 9347 -145
rect 9403 -201 9467 -145
rect 9523 -201 9547 -145
rect 9603 -201 9667 -145
rect 9723 -201 9747 -145
rect 9803 -201 9867 -145
rect 9923 -201 9947 -145
rect 10003 -201 10067 -145
rect 10123 -201 10147 -145
rect 10203 -201 10267 -145
rect 10323 -201 10347 -145
rect 10403 -201 10467 -145
rect 10523 -201 10547 -145
rect 10603 -201 10667 -145
rect 10723 -201 10747 -145
rect 10803 -201 10867 -145
rect 10923 -201 10947 -145
rect 11003 -201 11067 -145
rect 11123 -201 11147 -145
rect 11203 -201 11267 -145
rect 11323 -201 11347 -145
rect 11403 -201 11467 -145
rect 11523 -201 11547 -145
rect 11603 -201 11667 -145
rect 11723 -201 11747 -145
rect 11803 -201 11867 -145
rect 11923 -201 11947 -145
rect 12003 -201 12067 -145
rect 12123 -201 12147 -145
rect 12203 -201 12267 -145
rect 12323 -201 12347 -145
rect 12403 -201 12467 -145
rect 12523 -201 12547 -145
rect 12603 -201 12667 -145
rect 12723 -201 12747 -145
rect 12803 -201 12808 -145
rect -138 -240 12808 -201
rect 14521 -197 14702 -160
rect 14521 -253 14543 -197
rect 14599 -253 14623 -197
rect 14679 -253 14702 -197
rect -98 -348 12768 -324
rect -98 -404 -93 -348
rect -37 -404 107 -348
rect 163 -404 307 -348
rect 363 -404 507 -348
rect 563 -404 707 -348
rect 763 -404 907 -348
rect 963 -404 1107 -348
rect 1163 -404 1307 -348
rect 1363 -404 1507 -348
rect 1563 -404 1707 -348
rect 1763 -404 1907 -348
rect 1963 -404 2107 -348
rect 2163 -404 2307 -348
rect 2363 -404 2507 -348
rect 2563 -404 2707 -348
rect 2763 -404 2907 -348
rect 2963 -404 3107 -348
rect 3163 -404 3307 -348
rect 3363 -404 3507 -348
rect 3563 -404 3707 -348
rect 3763 -404 3907 -348
rect 3963 -404 4107 -348
rect 4163 -404 4307 -348
rect 4363 -404 4507 -348
rect 4563 -404 4707 -348
rect 4763 -404 4907 -348
rect 4963 -404 5107 -348
rect 5163 -404 5307 -348
rect 5363 -404 5507 -348
rect 5563 -404 5707 -348
rect 5763 -404 5907 -348
rect 5963 -404 6107 -348
rect 6163 -404 6307 -348
rect 6363 -404 6507 -348
rect 6563 -404 6707 -348
rect 6763 -404 6907 -348
rect 6963 -404 7107 -348
rect 7163 -404 7307 -348
rect 7363 -404 7507 -348
rect 7563 -404 7707 -348
rect 7763 -404 7907 -348
rect 7963 -404 8107 -348
rect 8163 -404 8307 -348
rect 8363 -404 8507 -348
rect 8563 -404 8707 -348
rect 8763 -404 8907 -348
rect 8963 -404 9107 -348
rect 9163 -404 9307 -348
rect 9363 -404 9507 -348
rect 9563 -404 9707 -348
rect 9763 -404 9907 -348
rect 9963 -404 10107 -348
rect 10163 -404 10307 -348
rect 10363 -404 10507 -348
rect 10563 -404 10707 -348
rect 10763 -404 10907 -348
rect 10963 -404 11107 -348
rect 11163 -404 11307 -348
rect 11363 -404 11507 -348
rect 11563 -404 11707 -348
rect 11763 -404 11907 -348
rect 11963 -404 12107 -348
rect 12163 -404 12307 -348
rect 12363 -404 12507 -348
rect 12563 -404 12707 -348
rect 12763 -404 12768 -348
rect -98 -428 12768 -404
rect -98 -484 -93 -428
rect -37 -484 107 -428
rect 163 -484 307 -428
rect 363 -484 507 -428
rect 563 -484 707 -428
rect 763 -484 907 -428
rect 963 -484 1107 -428
rect 1163 -484 1307 -428
rect 1363 -484 1507 -428
rect 1563 -484 1707 -428
rect 1763 -484 1907 -428
rect 1963 -484 2107 -428
rect 2163 -484 2307 -428
rect 2363 -484 2507 -428
rect 2563 -484 2707 -428
rect 2763 -484 2907 -428
rect 2963 -484 3107 -428
rect 3163 -484 3307 -428
rect 3363 -484 3507 -428
rect 3563 -484 3707 -428
rect 3763 -484 3907 -428
rect 3963 -484 4107 -428
rect 4163 -484 4307 -428
rect 4363 -484 4507 -428
rect 4563 -484 4707 -428
rect 4763 -484 4907 -428
rect 4963 -484 5107 -428
rect 5163 -484 5307 -428
rect 5363 -484 5507 -428
rect 5563 -484 5707 -428
rect 5763 -484 5907 -428
rect 5963 -484 6107 -428
rect 6163 -484 6307 -428
rect 6363 -484 6507 -428
rect 6563 -484 6707 -428
rect 6763 -484 6907 -428
rect 6963 -484 7107 -428
rect 7163 -484 7307 -428
rect 7363 -484 7507 -428
rect 7563 -484 7707 -428
rect 7763 -484 7907 -428
rect 7963 -484 8107 -428
rect 8163 -484 8307 -428
rect 8363 -484 8507 -428
rect 8563 -484 8707 -428
rect 8763 -484 8907 -428
rect 8963 -484 9107 -428
rect 9163 -484 9307 -428
rect 9363 -484 9507 -428
rect 9563 -484 9707 -428
rect 9763 -484 9907 -428
rect 9963 -484 10107 -428
rect 10163 -484 10307 -428
rect 10363 -484 10507 -428
rect 10563 -484 10707 -428
rect 10763 -484 10907 -428
rect 10963 -484 11107 -428
rect 11163 -484 11307 -428
rect 11363 -484 11507 -428
rect 11563 -484 11707 -428
rect 11763 -484 11907 -428
rect 11963 -484 12107 -428
rect 12163 -484 12307 -428
rect 12363 -484 12507 -428
rect 12563 -484 12707 -428
rect 12763 -484 12768 -428
rect -98 -508 12768 -484
rect 14521 -397 14702 -253
rect 14521 -453 14543 -397
rect 14599 -453 14623 -397
rect 14679 -453 14702 -397
rect 14521 -597 14702 -453
rect 14521 -653 14543 -597
rect 14599 -653 14623 -597
rect 14679 -653 14702 -597
rect 14521 -797 14702 -653
rect 14521 -853 14543 -797
rect 14599 -853 14623 -797
rect 14679 -853 14702 -797
rect 14521 -997 14702 -853
rect 14521 -1053 14543 -997
rect 14599 -1053 14623 -997
rect 14679 -1053 14702 -997
rect 14521 -1197 14702 -1053
rect 14521 -1253 14543 -1197
rect 14599 -1253 14623 -1197
rect 14679 -1253 14702 -1197
rect 14521 -1397 14702 -1253
rect 14521 -1453 14543 -1397
rect 14599 -1453 14623 -1397
rect 14679 -1453 14702 -1397
rect 14521 -1597 14702 -1453
rect 14521 -1653 14543 -1597
rect 14599 -1653 14623 -1597
rect 14679 -1653 14702 -1597
rect 14521 -1797 14702 -1653
rect 14521 -1853 14543 -1797
rect 14599 -1853 14623 -1797
rect 14679 -1853 14702 -1797
rect 14521 -1997 14702 -1853
rect 14521 -2053 14543 -1997
rect 14599 -2053 14623 -1997
rect 14679 -2053 14702 -1997
rect 14521 -2090 14702 -2053
rect 14800 -197 15141 -160
rect 14800 -253 14822 -197
rect 14878 -253 14902 -197
rect 14958 -253 14982 -197
rect 15038 -253 15062 -197
rect 15118 -253 15141 -197
rect 14800 -397 15141 -253
rect 14800 -453 14822 -397
rect 14878 -453 14902 -397
rect 14958 -453 14982 -397
rect 15038 -453 15062 -397
rect 15118 -453 15141 -397
rect 14800 -597 15141 -453
rect 14800 -653 14822 -597
rect 14878 -653 14902 -597
rect 14958 -653 14982 -597
rect 15038 -653 15062 -597
rect 15118 -653 15141 -597
rect 14800 -797 15141 -653
rect 14800 -853 14822 -797
rect 14878 -853 14902 -797
rect 14958 -853 14982 -797
rect 15038 -853 15062 -797
rect 15118 -853 15141 -797
rect 14800 -997 15141 -853
rect 14800 -1053 14822 -997
rect 14878 -1053 14902 -997
rect 14958 -1053 14982 -997
rect 15038 -1053 15062 -997
rect 15118 -1053 15141 -997
rect 14800 -1197 15141 -1053
rect 14800 -1253 14822 -1197
rect 14878 -1253 14902 -1197
rect 14958 -1253 14982 -1197
rect 15038 -1253 15062 -1197
rect 15118 -1253 15141 -1197
rect 14800 -1397 15141 -1253
rect 14800 -1453 14822 -1397
rect 14878 -1453 14902 -1397
rect 14958 -1453 14982 -1397
rect 15038 -1453 15062 -1397
rect 15118 -1453 15141 -1397
rect 14800 -1597 15141 -1453
rect 14800 -1653 14822 -1597
rect 14878 -1653 14902 -1597
rect 14958 -1653 14982 -1597
rect 15038 -1653 15062 -1597
rect 15118 -1653 15141 -1597
rect 14800 -1797 15141 -1653
rect 14800 -1853 14822 -1797
rect 14878 -1853 14902 -1797
rect 14958 -1853 14982 -1797
rect 15038 -1853 15062 -1797
rect 15118 -1853 15141 -1797
rect 14800 -1997 15141 -1853
rect 14800 -2053 14822 -1997
rect 14878 -2053 14902 -1997
rect 14958 -2053 14982 -1997
rect 15038 -2053 15062 -1997
rect 15118 -2053 15141 -1997
rect 14800 -2090 15141 -2053
rect 15201 -197 15542 -160
rect 15201 -253 15223 -197
rect 15279 -253 15303 -197
rect 15359 -253 15383 -197
rect 15439 -253 15463 -197
rect 15519 -253 15542 -197
rect 15201 -397 15542 -253
rect 15201 -453 15223 -397
rect 15279 -453 15303 -397
rect 15359 -453 15383 -397
rect 15439 -453 15463 -397
rect 15519 -453 15542 -397
rect 15201 -597 15542 -453
rect 15201 -653 15223 -597
rect 15279 -653 15303 -597
rect 15359 -653 15383 -597
rect 15439 -653 15463 -597
rect 15519 -653 15542 -597
rect 15201 -797 15542 -653
rect 15201 -853 15223 -797
rect 15279 -853 15303 -797
rect 15359 -853 15383 -797
rect 15439 -853 15463 -797
rect 15519 -853 15542 -797
rect 15201 -997 15542 -853
rect 15201 -1053 15223 -997
rect 15279 -1053 15303 -997
rect 15359 -1053 15383 -997
rect 15439 -1053 15463 -997
rect 15519 -1053 15542 -997
rect 15201 -1197 15542 -1053
rect 15201 -1253 15223 -1197
rect 15279 -1253 15303 -1197
rect 15359 -1253 15383 -1197
rect 15439 -1253 15463 -1197
rect 15519 -1253 15542 -1197
rect 15201 -1397 15542 -1253
rect 15201 -1453 15223 -1397
rect 15279 -1453 15303 -1397
rect 15359 -1453 15383 -1397
rect 15439 -1453 15463 -1397
rect 15519 -1453 15542 -1397
rect 15201 -1597 15542 -1453
rect 15201 -1653 15223 -1597
rect 15279 -1653 15303 -1597
rect 15359 -1653 15383 -1597
rect 15439 -1653 15463 -1597
rect 15519 -1653 15542 -1597
rect 15201 -1797 15542 -1653
rect 15201 -1853 15223 -1797
rect 15279 -1853 15303 -1797
rect 15359 -1853 15383 -1797
rect 15439 -1853 15463 -1797
rect 15519 -1853 15542 -1797
rect 15201 -1997 15542 -1853
rect 15201 -2053 15223 -1997
rect 15279 -2053 15303 -1997
rect 15359 -2053 15383 -1997
rect 15439 -2053 15463 -1997
rect 15519 -2053 15542 -1997
rect 15201 -2090 15542 -2053
rect 15640 -197 15821 -160
rect 15640 -253 15662 -197
rect 15718 -253 15742 -197
rect 15798 -253 15821 -197
rect 15640 -397 15821 -253
rect 15640 -453 15662 -397
rect 15718 -453 15742 -397
rect 15798 -453 15821 -397
rect 15640 -597 15821 -453
rect 15640 -653 15662 -597
rect 15718 -653 15742 -597
rect 15798 -653 15821 -597
rect 15640 -797 15821 -653
rect 15640 -853 15662 -797
rect 15718 -853 15742 -797
rect 15798 -853 15821 -797
rect 15640 -997 15821 -853
rect 15640 -1053 15662 -997
rect 15718 -1053 15742 -997
rect 15798 -1053 15821 -997
rect 15640 -1197 15821 -1053
rect 15640 -1253 15662 -1197
rect 15718 -1253 15742 -1197
rect 15798 -1253 15821 -1197
rect 15640 -1397 15821 -1253
rect 15640 -1453 15662 -1397
rect 15718 -1453 15742 -1397
rect 15798 -1453 15821 -1397
rect 15640 -1597 15821 -1453
rect 15640 -1653 15662 -1597
rect 15718 -1653 15742 -1597
rect 15798 -1653 15821 -1597
rect 15640 -1797 15821 -1653
rect 15640 -1853 15662 -1797
rect 15718 -1853 15742 -1797
rect 15798 -1853 15821 -1797
rect 15640 -1997 15821 -1853
rect 15640 -2053 15662 -1997
rect 15718 -2053 15742 -1997
rect 15798 -2053 15821 -1997
rect 15640 -2090 15821 -2053
<< properties >>
string GDS_END 5235316
string GDS_FILE ../gds/rom_4k_1_core.gds
string GDS_START 112
<< end >>
